
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i0_s5, io_i0_s6, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, 
        io_i1_s4, io_i1_s5, io_i1_s6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, 
        p_rand_4, p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, 
        p_rand_11, p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16, 
        p_rand_17, p_rand_18, p_rand_19, p_rand_20, p_rand_21, p_rand_22, 
        p_rand_23, p_rand_24, p_rand_25, p_rand_26, p_rand_27, p_rand_28, 
        p_rand_29, p_rand_30, p_rand_31, p_rand_32, p_rand_33, p_rand_34, 
        p_rand_35, p_rand_36, p_rand_37, p_rand_38, p_rand_39, p_rand_40, 
        p_rand_41, io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5, 
        io_o0_s6 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i0_s5, io_i0_s6, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4,
         io_i1_s5, io_i1_s6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4,
         p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10,
         p_rand_11, p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16,
         p_rand_17, p_rand_18, p_rand_19, p_rand_20, p_rand_21, p_rand_22,
         p_rand_23, p_rand_24, p_rand_25, p_rand_26, p_rand_27, p_rand_28,
         p_rand_29, p_rand_30, p_rand_31, p_rand_32, p_rand_33, p_rand_34,
         p_rand_35, p_rand_36, p_rand_37, p_rand_38, p_rand_39, p_rand_40,
         p_rand_41;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5, io_o0_s6;
  wire   n_hpc2_0_n161, n_hpc2_0_n160, n_hpc2_0_n159, n_hpc2_0_n158,
         n_hpc2_0_n157, n_hpc2_0_n156, n_hpc2_0_n155, n_hpc2_0_n154,
         n_hpc2_0_n153, n_hpc2_0_n152, n_hpc2_0_n151, n_hpc2_0_n150,
         n_hpc2_0_n149, n_hpc2_0_n148, n_hpc2_0_n147, n_hpc2_0_n146,
         n_hpc2_0_n145, n_hpc2_0_n144, n_hpc2_0_n143, n_hpc2_0_n142,
         n_hpc2_0_n141, n_hpc2_0_n140, n_hpc2_0_n139, n_hpc2_0_n138,
         n_hpc2_0_n137, n_hpc2_0_n136, n_hpc2_0_n135, n_hpc2_0_n134,
         n_hpc2_0_n133, n_hpc2_0_n132, n_hpc2_0_n131, n_hpc2_0_n130,
         n_hpc2_0_n129, n_hpc2_0_n128, n_hpc2_0_n127, n_hpc2_0_n126,
         n_hpc2_0_n125, n_hpc2_0_n124, n_hpc2_0_n123, n_hpc2_0_n122,
         n_hpc2_0_n121, n_hpc2_0_n120, n_hpc2_0_n119, n_hpc2_0_n118,
         n_hpc2_0_n117, n_hpc2_0_n116, n_hpc2_0_n115, n_hpc2_0_n114,
         n_hpc2_0_n113, n_hpc2_0_n112, n_hpc2_0_n111, n_hpc2_0_n110,
         n_hpc2_0_n109, n_hpc2_0_n108, n_hpc2_0_n107, n_hpc2_0_n106,
         n_hpc2_0_n105, n_hpc2_0_n104, n_hpc2_0_n103, n_hpc2_0_n102,
         n_hpc2_0_n101, n_hpc2_0_n100, n_hpc2_0_n99, n_hpc2_0_n98,
         n_hpc2_0_n97, n_hpc2_0_n96, n_hpc2_0_n95, n_hpc2_0_n94, n_hpc2_0_n93,
         n_hpc2_0_n92, n_hpc2_0_n91, n_hpc2_0_n90, n_hpc2_0_n89, n_hpc2_0_n88,
         n_hpc2_0_n87, n_hpc2_0_n86, n_hpc2_0_n85, n_hpc2_0_n84, n_hpc2_0_n83,
         n_hpc2_0_n82, n_hpc2_0_n81, n_hpc2_0_n80, n_hpc2_0_n79, n_hpc2_0_n78,
         n_hpc2_0_n77, n_hpc2_0_n76, n_hpc2_0_n75, n_hpc2_0_n74, n_hpc2_0_n73,
         n_hpc2_0_n72, n_hpc2_0_n71, n_hpc2_0_n70, n_hpc2_0_n69, n_hpc2_0_n68,
         n_hpc2_0_n67, n_hpc2_0_n66, n_hpc2_0_n65, n_hpc2_0_n64, n_hpc2_0_n63,
         n_hpc2_0_n62, n_hpc2_0_n61, n_hpc2_0_n60, n_hpc2_0_n59, n_hpc2_0_n58,
         n_hpc2_0_n57, n_hpc2_0_n56, n_hpc2_0_n55, n_hpc2_0_n54, n_hpc2_0_n53,
         n_hpc2_0_n52, n_hpc2_0_n51, n_hpc2_0_n50, n_hpc2_0_n49, n_hpc2_0_n48,
         n_hpc2_0_n47, n_hpc2_0_n46, n_hpc2_0_n45, n_hpc2_0_n44, n_hpc2_0_n43,
         n_hpc2_0_n42, n_hpc2_0_n41, n_hpc2_0_n40, n_hpc2_0_n39, n_hpc2_0_n38,
         n_hpc2_0_n37, n_hpc2_0_n36, n_hpc2_0_n35, n_hpc2_0_n34, n_hpc2_0_n33,
         n_hpc2_0_n32, n_hpc2_0_n31, n_hpc2_0_n30, n_hpc2_0_n29, n_hpc2_0_n28,
         n_hpc2_0_n27, n_hpc2_0_n26, n_hpc2_0_n25, n_hpc2_0_n24, n_hpc2_0_n23,
         n_hpc2_0_n22, n_hpc2_0_n21, n_hpc2_0_n20, n_hpc2_0_n19, n_hpc2_0_n18,
         n_hpc2_0_n17, n_hpc2_0_n16, n_hpc2_0_n15, n_hpc2_0_n14, n_hpc2_0_n13,
         n_hpc2_0_n12, n_hpc2_0_n11, n_hpc2_0_n10, n_hpc2_0_n9, n_hpc2_0_n8,
         n_hpc2_0_n7, n_hpc2_0_n6, n_hpc2_0_n5, n_hpc2_0_n4, n_hpc2_0_n3,
         n_hpc2_0_n2, n_hpc2_0_n1, n_hpc2_0_N55, n_hpc2_0_N54, n_hpc2_0_N53,
         n_hpc2_0_N52, n_hpc2_0_N51, n_hpc2_0_N50, n_hpc2_0_N49, n_hpc2_0_N48,
         n_hpc2_0_N47, n_hpc2_0_N46, n_hpc2_0_N45, n_hpc2_0_N44, n_hpc2_0_N43,
         n_hpc2_0_N42, n_hpc2_0_N41, n_hpc2_0_N40, n_hpc2_0_N39, n_hpc2_0_N38,
         n_hpc2_0_N37, n_hpc2_0_N36, n_hpc2_0_N35, n_hpc2_0_N34, n_hpc2_0_N33,
         n_hpc2_0_N32, n_hpc2_0_N31, n_hpc2_0_N30, n_hpc2_0_N29, n_hpc2_0_N28,
         n_hpc2_0_N27, n_hpc2_0_N26, n_hpc2_0_N25, n_hpc2_0_N24, n_hpc2_0_N23,
         n_hpc2_0_N22, n_hpc2_0_N21, n_hpc2_0_N20, n_hpc2_0_N19, n_hpc2_0_N18,
         n_hpc2_0_N17, n_hpc2_0_N16, n_hpc2_0_N15, n_hpc2_0_N14, n_hpc2_0_N13,
         n_hpc2_0_N12, n_hpc2_0_N11, n_hpc2_0_N10, n_hpc2_0_N9, n_hpc2_0_N8,
         n_hpc2_0_N7, n_hpc2_0_reg_pipeline_26, n_hpc2_0_reg_pipeline_25,
         n_hpc2_0_reg_pipeline_24, n_hpc2_0_reg_pipeline_23,
         n_hpc2_0_reg_pipeline_22, n_hpc2_0_reg_pipeline_21,
         n_hpc2_0_reg_pipeline_20, n_hpc2_0_reg_pipeline_19,
         n_hpc2_0_reg_pipeline_18, n_hpc2_0_reg_pipeline_17,
         n_hpc2_0_reg_pipeline_16, n_hpc2_0_reg_pipeline_15,
         n_hpc2_0_reg_pipeline_14, n_hpc2_0_reg_pipeline_13,
         n_hpc2_0_reg_pipeline_12, n_hpc2_0_reg_pipeline_11,
         n_hpc2_0_reg_pipeline_10, n_hpc2_0_reg_pipeline_9,
         n_hpc2_0_reg_pipeline_8, n_hpc2_0_reg_pipeline_7,
         n_hpc2_0_reg_pipeline_6, n_hpc2_0_reg_pipeline_5,
         n_hpc2_0_reg_pipeline_4, n_hpc2_0_reg_pipeline_3,
         n_hpc2_0_reg_pipeline_2, n_hpc2_0_reg_pipeline_1,
         n_hpc2_0_reg_pipeline_0, n_hpc2_0_reg_pipeline, n_hpc2_0_N6,
         n_hpc2_0_N5, n_hpc2_0_N4, n_hpc2_0_N3, n_hpc2_0_N2, n_hpc2_0_N1,
         n_hpc2_0_N0, n_hpc2_0__hpc1_z65, n_hpc2_0__hpc1_z55,
         n_hpc2_0__hpc1_z45, n_hpc2_0__hpc1_z35, n_hpc2_0__hpc1_z25,
         n_hpc2_0__hpc1_z15, n_hpc2_0__hpc1_z05;

  XOR2_X1 u_hpc2_0_U177 ( .A(io_i1_s0), .B(p_rand_5), .Z(n_hpc2_0_n118) );
  XOR2_X1 u_hpc2_0_U176 ( .A(p_rand_4), .B(p_rand_3), .Z(n_hpc2_0_n119) );
  XOR2_X1 u_hpc2_0_U175 ( .A(n_hpc2_0_n118), .B(n_hpc2_0_n119), .Z(
        n_hpc2_0_n115) );
  XOR2_X1 u_hpc2_0_U174 ( .A(p_rand_2), .B(p_rand_1), .Z(n_hpc2_0_n117) );
  XOR2_X1 u_hpc2_0_U173 ( .A(p_rand_0), .B(n_hpc2_0_n117), .Z(n_hpc2_0_n116)
         );
  XOR2_X1 u_hpc2_0_U172 ( .A(n_hpc2_0_n115), .B(n_hpc2_0_n116), .Z(n_hpc2_0_N0) );
  XOR2_X1 u_hpc2_0_U171 ( .A(io_i1_s1), .B(p_rand_9), .Z(n_hpc2_0_n113) );
  XOR2_X1 u_hpc2_0_U170 ( .A(p_rand_8), .B(p_rand_7), .Z(n_hpc2_0_n114) );
  XOR2_X1 u_hpc2_0_U169 ( .A(n_hpc2_0_n113), .B(n_hpc2_0_n114), .Z(
        n_hpc2_0_n110) );
  XOR2_X1 u_hpc2_0_U168 ( .A(p_rand_6), .B(p_rand_10), .Z(n_hpc2_0_n112) );
  XOR2_X1 u_hpc2_0_U167 ( .A(p_rand_0), .B(n_hpc2_0_n112), .Z(n_hpc2_0_n111)
         );
  XOR2_X1 u_hpc2_0_U166 ( .A(n_hpc2_0_n110), .B(n_hpc2_0_n111), .Z(n_hpc2_0_N1) );
  NAND2_X1 u_hpc2_0_U165 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_n109) );
  XNOR2_X1 u_hpc2_0_U164 ( .A(n_hpc2_0_reg_pipeline_2), .B(n_hpc2_0_n109), 
        .ZN(n_hpc2_0_N10) );
  NAND2_X1 u_hpc2_0_U163 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n6), .ZN(
        n_hpc2_0_n108) );
  XNOR2_X1 u_hpc2_0_U162 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n108), 
        .ZN(n_hpc2_0_N11) );
  NAND2_X1 u_hpc2_0_U161 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n5), .ZN(
        n_hpc2_0_n107) );
  XNOR2_X1 u_hpc2_0_U160 ( .A(n_hpc2_0_reg_pipeline_4), .B(n_hpc2_0_n107), 
        .ZN(n_hpc2_0_N12) );
  NAND2_X1 u_hpc2_0_U159 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n4), .ZN(
        n_hpc2_0_n106) );
  XNOR2_X1 u_hpc2_0_U158 ( .A(n_hpc2_0_reg_pipeline_5), .B(n_hpc2_0_n106), 
        .ZN(n_hpc2_0_N13) );
  NAND2_X1 u_hpc2_0_U157 ( .A1(n_hpc2_0_reg_pipeline_6), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n105) );
  XNOR2_X1 u_hpc2_0_U156 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n105), 
        .ZN(n_hpc2_0_N14) );
  AND2_X1 u_hpc2_0_U155 ( .A1(n_hpc2_0_n2), .A2(n_hpc2_0_reg_pipeline_6), .ZN(
        n_hpc2_0_N15) );
  NAND2_X1 u_hpc2_0_U154 ( .A1(n_hpc2_0_reg_pipeline_6), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n104) );
  XNOR2_X1 u_hpc2_0_U153 ( .A(n_hpc2_0_reg_pipeline_7), .B(n_hpc2_0_n104), 
        .ZN(n_hpc2_0_N16) );
  NAND2_X1 u_hpc2_0_U152 ( .A1(n_hpc2_0_reg_pipeline_6), .A2(n_hpc2_0_n7), 
        .ZN(n_hpc2_0_n103) );
  XNOR2_X1 u_hpc2_0_U151 ( .A(n_hpc2_0_reg_pipeline_8), .B(n_hpc2_0_n103), 
        .ZN(n_hpc2_0_N17) );
  NAND2_X1 u_hpc2_0_U150 ( .A1(n_hpc2_0_reg_pipeline_6), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n102) );
  XNOR2_X1 u_hpc2_0_U149 ( .A(n_hpc2_0_reg_pipeline_9), .B(n_hpc2_0_n102), 
        .ZN(n_hpc2_0_N18) );
  NAND2_X1 u_hpc2_0_U148 ( .A1(n_hpc2_0_reg_pipeline_6), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n101) );
  XNOR2_X1 u_hpc2_0_U147 ( .A(n_hpc2_0_reg_pipeline_10), .B(n_hpc2_0_n101), 
        .ZN(n_hpc2_0_N19) );
  XOR2_X1 u_hpc2_0_U146 ( .A(io_i1_s2), .B(p_rand_6), .Z(n_hpc2_0_n99) );
  XOR2_X1 u_hpc2_0_U145 ( .A(p_rand_14), .B(p_rand_13), .Z(n_hpc2_0_n100) );
  XOR2_X1 u_hpc2_0_U144 ( .A(n_hpc2_0_n99), .B(n_hpc2_0_n100), .Z(n_hpc2_0_n96) );
  XOR2_X1 u_hpc2_0_U143 ( .A(p_rand_12), .B(p_rand_11), .Z(n_hpc2_0_n98) );
  XOR2_X1 u_hpc2_0_U142 ( .A(p_rand_1), .B(n_hpc2_0_n98), .Z(n_hpc2_0_n97) );
  XOR2_X1 u_hpc2_0_U141 ( .A(n_hpc2_0_n96), .B(n_hpc2_0_n97), .Z(n_hpc2_0_N2)
         );
  NAND2_X1 u_hpc2_0_U140 ( .A1(n_hpc2_0_reg_pipeline_6), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n95) );
  XNOR2_X1 u_hpc2_0_U139 ( .A(n_hpc2_0_reg_pipeline_11), .B(n_hpc2_0_n95), 
        .ZN(n_hpc2_0_N20) );
  NAND2_X1 u_hpc2_0_U138 ( .A1(n_hpc2_0_reg_pipeline_12), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n94) );
  XNOR2_X1 u_hpc2_0_U137 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n94), .ZN(
        n_hpc2_0_N21) );
  NAND2_X1 u_hpc2_0_U136 ( .A1(n_hpc2_0_reg_pipeline_12), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n93) );
  XNOR2_X1 u_hpc2_0_U135 ( .A(n_hpc2_0_reg_pipeline_7), .B(n_hpc2_0_n93), .ZN(
        n_hpc2_0_N22) );
  AND2_X1 u_hpc2_0_U134 ( .A1(n_hpc2_0_n1), .A2(n_hpc2_0_reg_pipeline_12), 
        .ZN(n_hpc2_0_N23) );
  NAND2_X1 u_hpc2_0_U133 ( .A1(n_hpc2_0_reg_pipeline_12), .A2(n_hpc2_0_n7), 
        .ZN(n_hpc2_0_n92) );
  XNOR2_X1 u_hpc2_0_U132 ( .A(n_hpc2_0_reg_pipeline_13), .B(n_hpc2_0_n92), 
        .ZN(n_hpc2_0_N24) );
  NAND2_X1 u_hpc2_0_U131 ( .A1(n_hpc2_0_reg_pipeline_12), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n91) );
  XNOR2_X1 u_hpc2_0_U130 ( .A(n_hpc2_0_reg_pipeline_14), .B(n_hpc2_0_n91), 
        .ZN(n_hpc2_0_N25) );
  NAND2_X1 u_hpc2_0_U129 ( .A1(n_hpc2_0_reg_pipeline_12), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n90) );
  XNOR2_X1 u_hpc2_0_U128 ( .A(n_hpc2_0_reg_pipeline_15), .B(n_hpc2_0_n90), 
        .ZN(n_hpc2_0_N26) );
  NAND2_X1 u_hpc2_0_U127 ( .A1(n_hpc2_0_reg_pipeline_12), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n89) );
  XNOR2_X1 u_hpc2_0_U126 ( .A(n_hpc2_0_reg_pipeline_16), .B(n_hpc2_0_n89), 
        .ZN(n_hpc2_0_N27) );
  NAND2_X1 u_hpc2_0_U125 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n88) );
  XNOR2_X1 u_hpc2_0_U124 ( .A(n_hpc2_0_reg_pipeline_2), .B(n_hpc2_0_n88), .ZN(
        n_hpc2_0_N28) );
  NAND2_X1 u_hpc2_0_U123 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n87) );
  XNOR2_X1 u_hpc2_0_U122 ( .A(n_hpc2_0_reg_pipeline_8), .B(n_hpc2_0_n87), .ZN(
        n_hpc2_0_N29) );
  XOR2_X1 u_hpc2_0_U121 ( .A(io_i1_s3), .B(p_rand_7), .Z(n_hpc2_0_n85) );
  XOR2_X1 u_hpc2_0_U120 ( .A(p_rand_2), .B(p_rand_17), .Z(n_hpc2_0_n86) );
  XOR2_X1 u_hpc2_0_U119 ( .A(n_hpc2_0_n85), .B(n_hpc2_0_n86), .Z(n_hpc2_0_n82)
         );
  XOR2_X1 u_hpc2_0_U118 ( .A(p_rand_16), .B(p_rand_15), .Z(n_hpc2_0_n84) );
  XOR2_X1 u_hpc2_0_U117 ( .A(p_rand_11), .B(n_hpc2_0_n84), .Z(n_hpc2_0_n83) );
  XOR2_X1 u_hpc2_0_U116 ( .A(n_hpc2_0_n82), .B(n_hpc2_0_n83), .Z(n_hpc2_0_N3)
         );
  NAND2_X1 u_hpc2_0_U115 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n81) );
  XNOR2_X1 u_hpc2_0_U114 ( .A(n_hpc2_0_reg_pipeline_13), .B(n_hpc2_0_n81), 
        .ZN(n_hpc2_0_N30) );
  AND2_X1 u_hpc2_0_U113 ( .A1(n_hpc2_0_n7), .A2(n_hpc2_0_reg_pipeline_17), 
        .ZN(n_hpc2_0_N31) );
  NAND2_X1 u_hpc2_0_U112 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n80) );
  XNOR2_X1 u_hpc2_0_U111 ( .A(n_hpc2_0_reg_pipeline_18), .B(n_hpc2_0_n80), 
        .ZN(n_hpc2_0_N32) );
  NAND2_X1 u_hpc2_0_U110 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n79) );
  XNOR2_X1 u_hpc2_0_U109 ( .A(n_hpc2_0_reg_pipeline_19), .B(n_hpc2_0_n79), 
        .ZN(n_hpc2_0_N33) );
  NAND2_X1 u_hpc2_0_U108 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n78) );
  XNOR2_X1 u_hpc2_0_U107 ( .A(n_hpc2_0_reg_pipeline_20), .B(n_hpc2_0_n78), 
        .ZN(n_hpc2_0_N34) );
  NAND2_X1 u_hpc2_0_U106 ( .A1(n_hpc2_0_reg_pipeline_21), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n77) );
  XNOR2_X1 u_hpc2_0_U105 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n77), .ZN(
        n_hpc2_0_N35) );
  NAND2_X1 u_hpc2_0_U104 ( .A1(n_hpc2_0_reg_pipeline_21), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n76) );
  XNOR2_X1 u_hpc2_0_U103 ( .A(n_hpc2_0_reg_pipeline_9), .B(n_hpc2_0_n76), .ZN(
        n_hpc2_0_N36) );
  NAND2_X1 u_hpc2_0_U102 ( .A1(n_hpc2_0_reg_pipeline_21), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n75) );
  XNOR2_X1 u_hpc2_0_U101 ( .A(n_hpc2_0_reg_pipeline_14), .B(n_hpc2_0_n75), 
        .ZN(n_hpc2_0_N37) );
  NAND2_X1 u_hpc2_0_U100 ( .A1(n_hpc2_0_reg_pipeline_21), .A2(n_hpc2_0_n7), 
        .ZN(n_hpc2_0_n74) );
  XNOR2_X1 u_hpc2_0_U99 ( .A(n_hpc2_0_reg_pipeline_18), .B(n_hpc2_0_n74), .ZN(
        n_hpc2_0_N38) );
  AND2_X1 u_hpc2_0_U98 ( .A1(n_hpc2_0_n6), .A2(n_hpc2_0_reg_pipeline_21), .ZN(
        n_hpc2_0_N39) );
  XOR2_X1 u_hpc2_0_U97 ( .A(io_i1_s4), .B(p_rand_8), .Z(n_hpc2_0_n72) );
  XOR2_X1 u_hpc2_0_U96 ( .A(p_rand_3), .B(p_rand_19), .Z(n_hpc2_0_n73) );
  XOR2_X1 u_hpc2_0_U95 ( .A(n_hpc2_0_n72), .B(n_hpc2_0_n73), .Z(n_hpc2_0_n69)
         );
  XOR2_X1 u_hpc2_0_U94 ( .A(p_rand_18), .B(p_rand_15), .Z(n_hpc2_0_n71) );
  XOR2_X1 u_hpc2_0_U93 ( .A(p_rand_12), .B(n_hpc2_0_n71), .Z(n_hpc2_0_n70) );
  XOR2_X1 u_hpc2_0_U92 ( .A(n_hpc2_0_n69), .B(n_hpc2_0_n70), .Z(n_hpc2_0_N4)
         );
  NAND2_X1 u_hpc2_0_U91 ( .A1(n_hpc2_0_reg_pipeline_21), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n68) );
  XNOR2_X1 u_hpc2_0_U90 ( .A(n_hpc2_0_reg_pipeline_22), .B(n_hpc2_0_n68), .ZN(
        n_hpc2_0_N40) );
  NAND2_X1 u_hpc2_0_U89 ( .A1(n_hpc2_0_reg_pipeline_21), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n67) );
  XNOR2_X1 u_hpc2_0_U88 ( .A(n_hpc2_0_reg_pipeline_23), .B(n_hpc2_0_n67), .ZN(
        n_hpc2_0_N41) );
  NAND2_X1 u_hpc2_0_U87 ( .A1(n_hpc2_0_reg_pipeline_24), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n66) );
  XNOR2_X1 u_hpc2_0_U86 ( .A(n_hpc2_0_reg_pipeline_4), .B(n_hpc2_0_n66), .ZN(
        n_hpc2_0_N42) );
  NAND2_X1 u_hpc2_0_U85 ( .A1(n_hpc2_0_reg_pipeline_24), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n65) );
  XNOR2_X1 u_hpc2_0_U84 ( .A(n_hpc2_0_reg_pipeline_10), .B(n_hpc2_0_n65), .ZN(
        n_hpc2_0_N43) );
  NAND2_X1 u_hpc2_0_U83 ( .A1(n_hpc2_0_reg_pipeline_24), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n64) );
  XNOR2_X1 u_hpc2_0_U82 ( .A(n_hpc2_0_reg_pipeline_15), .B(n_hpc2_0_n64), .ZN(
        n_hpc2_0_N44) );
  NAND2_X1 u_hpc2_0_U81 ( .A1(n_hpc2_0_reg_pipeline_24), .A2(n_hpc2_0_n7), 
        .ZN(n_hpc2_0_n63) );
  XNOR2_X1 u_hpc2_0_U80 ( .A(n_hpc2_0_reg_pipeline_19), .B(n_hpc2_0_n63), .ZN(
        n_hpc2_0_N45) );
  NAND2_X1 u_hpc2_0_U79 ( .A1(n_hpc2_0_reg_pipeline_24), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n62) );
  XNOR2_X1 u_hpc2_0_U78 ( .A(n_hpc2_0_reg_pipeline_22), .B(n_hpc2_0_n62), .ZN(
        n_hpc2_0_N46) );
  AND2_X1 u_hpc2_0_U77 ( .A1(n_hpc2_0_n5), .A2(n_hpc2_0_reg_pipeline_24), .ZN(
        n_hpc2_0_N47) );
  NAND2_X1 u_hpc2_0_U76 ( .A1(n_hpc2_0_reg_pipeline_24), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n61) );
  XNOR2_X1 u_hpc2_0_U75 ( .A(n_hpc2_0_reg_pipeline_25), .B(n_hpc2_0_n61), .ZN(
        n_hpc2_0_N48) );
  NAND2_X1 u_hpc2_0_U74 ( .A1(n_hpc2_0_reg_pipeline_26), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n60) );
  XNOR2_X1 u_hpc2_0_U73 ( .A(n_hpc2_0_reg_pipeline_5), .B(n_hpc2_0_n60), .ZN(
        n_hpc2_0_N49) );
  XOR2_X1 u_hpc2_0_U72 ( .A(io_i1_s5), .B(p_rand_9), .Z(n_hpc2_0_n58) );
  XOR2_X1 u_hpc2_0_U71 ( .A(p_rand_4), .B(p_rand_20), .Z(n_hpc2_0_n59) );
  XOR2_X1 u_hpc2_0_U70 ( .A(n_hpc2_0_n58), .B(n_hpc2_0_n59), .Z(n_hpc2_0_n55)
         );
  XOR2_X1 u_hpc2_0_U69 ( .A(p_rand_18), .B(p_rand_16), .Z(n_hpc2_0_n57) );
  XOR2_X1 u_hpc2_0_U68 ( .A(p_rand_13), .B(n_hpc2_0_n57), .Z(n_hpc2_0_n56) );
  XOR2_X1 u_hpc2_0_U67 ( .A(n_hpc2_0_n55), .B(n_hpc2_0_n56), .Z(n_hpc2_0_N5)
         );
  NAND2_X1 u_hpc2_0_U66 ( .A1(n_hpc2_0_reg_pipeline_26), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n54) );
  XNOR2_X1 u_hpc2_0_U65 ( .A(n_hpc2_0_reg_pipeline_11), .B(n_hpc2_0_n54), .ZN(
        n_hpc2_0_N50) );
  NAND2_X1 u_hpc2_0_U64 ( .A1(n_hpc2_0_reg_pipeline_26), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n53) );
  XNOR2_X1 u_hpc2_0_U63 ( .A(n_hpc2_0_reg_pipeline_16), .B(n_hpc2_0_n53), .ZN(
        n_hpc2_0_N51) );
  NAND2_X1 u_hpc2_0_U62 ( .A1(n_hpc2_0_reg_pipeline_26), .A2(n_hpc2_0_n7), 
        .ZN(n_hpc2_0_n52) );
  XNOR2_X1 u_hpc2_0_U61 ( .A(n_hpc2_0_reg_pipeline_20), .B(n_hpc2_0_n52), .ZN(
        n_hpc2_0_N52) );
  NAND2_X1 u_hpc2_0_U60 ( .A1(n_hpc2_0_reg_pipeline_26), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n51) );
  XNOR2_X1 u_hpc2_0_U59 ( .A(n_hpc2_0_reg_pipeline_23), .B(n_hpc2_0_n51), .ZN(
        n_hpc2_0_N53) );
  NAND2_X1 u_hpc2_0_U58 ( .A1(n_hpc2_0_reg_pipeline_26), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n50) );
  XNOR2_X1 u_hpc2_0_U57 ( .A(n_hpc2_0_reg_pipeline_25), .B(n_hpc2_0_n50), .ZN(
        n_hpc2_0_N54) );
  AND2_X1 u_hpc2_0_U56 ( .A1(n_hpc2_0_n4), .A2(n_hpc2_0_reg_pipeline_26), .ZN(
        n_hpc2_0_N55) );
  XOR2_X1 u_hpc2_0_U55 ( .A(io_i1_s6), .B(p_rand_5), .Z(n_hpc2_0_n48) );
  XOR2_X1 u_hpc2_0_U54 ( .A(p_rand_20), .B(p_rand_19), .Z(n_hpc2_0_n49) );
  XOR2_X1 u_hpc2_0_U53 ( .A(n_hpc2_0_n48), .B(n_hpc2_0_n49), .Z(n_hpc2_0_n45)
         );
  XOR2_X1 u_hpc2_0_U52 ( .A(p_rand_17), .B(p_rand_14), .Z(n_hpc2_0_n47) );
  XOR2_X1 u_hpc2_0_U51 ( .A(p_rand_10), .B(n_hpc2_0_n47), .Z(n_hpc2_0_n46) );
  XOR2_X1 u_hpc2_0_U50 ( .A(n_hpc2_0_n45), .B(n_hpc2_0_n46), .Z(n_hpc2_0_N6)
         );
  AND2_X1 u_hpc2_0_U49 ( .A1(n_hpc2_0_n3), .A2(n_hpc2_0_reg_pipeline), .ZN(
        n_hpc2_0_N7) );
  NAND2_X1 u_hpc2_0_U48 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n44) );
  XNOR2_X1 u_hpc2_0_U47 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n44), .ZN(
        n_hpc2_0_N8) );
  NAND2_X1 u_hpc2_0_U46 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n43) );
  XNOR2_X1 u_hpc2_0_U45 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n43), .ZN(
        n_hpc2_0_N9) );
  XOR2_X1 u_hpc2_0_U44 ( .A(n_hpc2_0__hpc1_z05), .B(n_hpc2_0_n158), .Z(
        n_hpc2_0_n41) );
  XOR2_X1 u_hpc2_0_U43 ( .A(n_hpc2_0_n156), .B(n_hpc2_0_n157), .Z(n_hpc2_0_n42) );
  XOR2_X1 u_hpc2_0_U42 ( .A(n_hpc2_0_n41), .B(n_hpc2_0_n42), .Z(n_hpc2_0_n38)
         );
  XOR2_X1 u_hpc2_0_U41 ( .A(n_hpc2_0_n159), .B(n_hpc2_0_n160), .Z(n_hpc2_0_n40) );
  XOR2_X1 u_hpc2_0_U40 ( .A(n_hpc2_0_n161), .B(n_hpc2_0_n40), .Z(n_hpc2_0_n39)
         );
  XOR2_X1 u_hpc2_0_U39 ( .A(n_hpc2_0_n38), .B(n_hpc2_0_n39), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U38 ( .A(n_hpc2_0__hpc1_z15), .B(n_hpc2_0_n152), .Z(
        n_hpc2_0_n36) );
  XOR2_X1 u_hpc2_0_U37 ( .A(n_hpc2_0_n150), .B(n_hpc2_0_n151), .Z(n_hpc2_0_n37) );
  XOR2_X1 u_hpc2_0_U36 ( .A(n_hpc2_0_n36), .B(n_hpc2_0_n37), .Z(n_hpc2_0_n33)
         );
  XOR2_X1 u_hpc2_0_U35 ( .A(n_hpc2_0_n153), .B(n_hpc2_0_n154), .Z(n_hpc2_0_n35) );
  XOR2_X1 u_hpc2_0_U34 ( .A(n_hpc2_0_n155), .B(n_hpc2_0_n35), .Z(n_hpc2_0_n34)
         );
  XOR2_X1 u_hpc2_0_U33 ( .A(n_hpc2_0_n33), .B(n_hpc2_0_n34), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U32 ( .A(n_hpc2_0__hpc1_z25), .B(n_hpc2_0_n146), .Z(
        n_hpc2_0_n31) );
  XOR2_X1 u_hpc2_0_U31 ( .A(n_hpc2_0_n144), .B(n_hpc2_0_n145), .Z(n_hpc2_0_n32) );
  XOR2_X1 u_hpc2_0_U30 ( .A(n_hpc2_0_n31), .B(n_hpc2_0_n32), .Z(n_hpc2_0_n28)
         );
  XOR2_X1 u_hpc2_0_U29 ( .A(n_hpc2_0_n147), .B(n_hpc2_0_n148), .Z(n_hpc2_0_n30) );
  XOR2_X1 u_hpc2_0_U28 ( .A(n_hpc2_0_n149), .B(n_hpc2_0_n30), .Z(n_hpc2_0_n29)
         );
  XOR2_X1 u_hpc2_0_U27 ( .A(n_hpc2_0_n28), .B(n_hpc2_0_n29), .Z(io_o0_s2) );
  XOR2_X1 u_hpc2_0_U26 ( .A(n_hpc2_0__hpc1_z35), .B(n_hpc2_0_n140), .Z(
        n_hpc2_0_n26) );
  XOR2_X1 u_hpc2_0_U25 ( .A(n_hpc2_0_n138), .B(n_hpc2_0_n139), .Z(n_hpc2_0_n27) );
  XOR2_X1 u_hpc2_0_U24 ( .A(n_hpc2_0_n26), .B(n_hpc2_0_n27), .Z(n_hpc2_0_n23)
         );
  XOR2_X1 u_hpc2_0_U23 ( .A(n_hpc2_0_n141), .B(n_hpc2_0_n142), .Z(n_hpc2_0_n25) );
  XOR2_X1 u_hpc2_0_U22 ( .A(n_hpc2_0_n143), .B(n_hpc2_0_n25), .Z(n_hpc2_0_n24)
         );
  XOR2_X1 u_hpc2_0_U21 ( .A(n_hpc2_0_n23), .B(n_hpc2_0_n24), .Z(io_o0_s3) );
  XOR2_X1 u_hpc2_0_U20 ( .A(n_hpc2_0__hpc1_z45), .B(n_hpc2_0_n134), .Z(
        n_hpc2_0_n21) );
  XOR2_X1 u_hpc2_0_U19 ( .A(n_hpc2_0_n132), .B(n_hpc2_0_n133), .Z(n_hpc2_0_n22) );
  XOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0_n21), .B(n_hpc2_0_n22), .Z(n_hpc2_0_n18)
         );
  XOR2_X1 u_hpc2_0_U17 ( .A(n_hpc2_0_n135), .B(n_hpc2_0_n136), .Z(n_hpc2_0_n20) );
  XOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_n137), .B(n_hpc2_0_n20), .Z(n_hpc2_0_n19)
         );
  XOR2_X1 u_hpc2_0_U15 ( .A(n_hpc2_0_n18), .B(n_hpc2_0_n19), .Z(io_o0_s4) );
  XOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0__hpc1_z55), .B(n_hpc2_0_n128), .Z(
        n_hpc2_0_n16) );
  XOR2_X1 u_hpc2_0_U13 ( .A(n_hpc2_0_n126), .B(n_hpc2_0_n127), .Z(n_hpc2_0_n17) );
  XOR2_X1 u_hpc2_0_U12 ( .A(n_hpc2_0_n16), .B(n_hpc2_0_n17), .Z(n_hpc2_0_n13)
         );
  XOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_n129), .B(n_hpc2_0_n130), .Z(n_hpc2_0_n15) );
  XOR2_X1 u_hpc2_0_U10 ( .A(n_hpc2_0_n131), .B(n_hpc2_0_n15), .Z(n_hpc2_0_n14)
         );
  XOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_n13), .B(n_hpc2_0_n14), .Z(io_o0_s5) );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0__hpc1_z65), .B(n_hpc2_0_n122), .Z(
        n_hpc2_0_n11) );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0_n120), .B(n_hpc2_0_n121), .Z(n_hpc2_0_n12)
         );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0_n11), .B(n_hpc2_0_n12), .Z(n_hpc2_0_n8) );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0_n123), .B(n_hpc2_0_n124), .Z(n_hpc2_0_n10)
         );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0_n125), .B(n_hpc2_0_n10), .Z(n_hpc2_0_n9)
         );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n8), .B(n_hpc2_0_n9), .Z(io_o0_s6) );
  DFF_X1 u_hpc2_0__hpc1_z56_reg ( .D(n_hpc2_0_N48), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n129) );
  DFF_X1 u_hpc2_0__hpc1_z55_reg ( .D(n_hpc2_0_N47), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z55), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z54_reg ( .D(n_hpc2_0_N46), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n131) );
  DFF_X1 u_hpc2_0__hpc1_z53_reg ( .D(n_hpc2_0_N45), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n130) );
  DFF_X1 u_hpc2_0__hpc1_z52_reg ( .D(n_hpc2_0_N44), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n128) );
  DFF_X1 u_hpc2_0__hpc1_z51_reg ( .D(n_hpc2_0_N43), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n127) );
  DFF_X1 u_hpc2_0__hpc1_z50_reg ( .D(n_hpc2_0_N42), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n126) );
  DFF_X1 u_hpc2_0__hpc1_z46_reg ( .D(n_hpc2_0_N41), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n135) );
  DFF_X1 u_hpc2_0__hpc1_z45_reg ( .D(n_hpc2_0_N40), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z45), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z44_reg ( .D(n_hpc2_0_N39), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n137) );
  DFF_X1 u_hpc2_0__hpc1_z43_reg ( .D(n_hpc2_0_N38), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n136) );
  DFF_X1 u_hpc2_0__hpc1_z42_reg ( .D(n_hpc2_0_N37), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n134) );
  DFF_X1 u_hpc2_0__hpc1_z41_reg ( .D(n_hpc2_0_N36), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n133) );
  DFF_X1 u_hpc2_0__hpc1_z40_reg ( .D(n_hpc2_0_N35), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n132) );
  DFF_X1 u_hpc2_0__hpc1_z36_reg ( .D(n_hpc2_0_N34), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n141) );
  DFF_X1 u_hpc2_0__hpc1_z35_reg ( .D(n_hpc2_0_N33), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z35), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z34_reg ( .D(n_hpc2_0_N32), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n143) );
  DFF_X1 u_hpc2_0__hpc1_z33_reg ( .D(n_hpc2_0_N31), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n142) );
  DFF_X1 u_hpc2_0__hpc1_z32_reg ( .D(n_hpc2_0_N30), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n140) );
  DFF_X1 u_hpc2_0__hpc1_z31_reg ( .D(n_hpc2_0_N29), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n139) );
  DFF_X1 u_hpc2_0__hpc1_z30_reg ( .D(n_hpc2_0_N28), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n138) );
  DFF_X1 u_hpc2_0__hpc1_z26_reg ( .D(n_hpc2_0_N27), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n147) );
  DFF_X1 u_hpc2_0__hpc1_z25_reg ( .D(n_hpc2_0_N26), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z25), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z24_reg ( .D(n_hpc2_0_N25), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n149) );
  DFF_X1 u_hpc2_0__hpc1_z23_reg ( .D(n_hpc2_0_N24), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n148) );
  DFF_X1 u_hpc2_0__hpc1_z22_reg ( .D(n_hpc2_0_N23), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n146) );
  DFF_X1 u_hpc2_0__hpc1_z21_reg ( .D(n_hpc2_0_N22), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n145) );
  DFF_X1 u_hpc2_0__hpc1_z20_reg ( .D(n_hpc2_0_N21), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n144) );
  DFF_X1 u_hpc2_0__hpc1_z16_reg ( .D(n_hpc2_0_N20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n153) );
  DFF_X1 u_hpc2_0__hpc1_z15_reg ( .D(n_hpc2_0_N19), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z15), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z14_reg ( .D(n_hpc2_0_N18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n155) );
  DFF_X1 u_hpc2_0__hpc1_z13_reg ( .D(n_hpc2_0_N17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n154) );
  DFF_X1 u_hpc2_0__hpc1_z12_reg ( .D(n_hpc2_0_N16), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n152) );
  DFF_X1 u_hpc2_0__hpc1_z11_reg ( .D(n_hpc2_0_N15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n151) );
  DFF_X1 u_hpc2_0__hpc1_z10_reg ( .D(n_hpc2_0_N14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n150) );
  DFF_X1 u_hpc2_0__hpc1_z06_reg ( .D(n_hpc2_0_N13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n159) );
  DFF_X1 u_hpc2_0__hpc1_z05_reg ( .D(n_hpc2_0_N12), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z05), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z04_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n161) );
  DFF_X1 u_hpc2_0__hpc1_z03_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n160) );
  DFF_X1 u_hpc2_0__hpc1_z02_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n158) );
  DFF_X1 u_hpc2_0__hpc1_z01_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n157) );
  DFF_X1 u_hpc2_0__hpc1_z00_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n156) );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(p_rand_23), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_2), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(io_i0_s0), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z65_reg ( .D(n_hpc2_0_N54), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z65), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_25_reg ( .D(p_rand_41), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_25), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(p_rand_22), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_1), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_6_reg ( .D(io_i0_s1), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_6), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z61_reg ( .D(n_hpc2_0_N50), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n121) );
  DFF_X1 u_hpc2_0_reg_pipeline_11_reg ( .D(p_rand_31), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_11), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z66_reg ( .D(n_hpc2_0_N55), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n123) );
  DFF_X1 u_hpc2_0__hpc1_ref_v6_reg ( .D(n_hpc2_0_N6), .CK(clock_0), .Q(
        n_hpc2_0_n4), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_13_reg ( .D(p_rand_32), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_13), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z63_reg ( .D(n_hpc2_0_N52), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n124) );
  DFF_X1 u_hpc2_0__hpc1_ref_v3_reg ( .D(n_hpc2_0_N3), .CK(clock_0), .Q(
        n_hpc2_0_n7), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_15_reg ( .D(p_rand_34), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_15), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v1_reg ( .D(n_hpc2_0_N1), .CK(clock_0), .Q(
        n_hpc2_0_n2), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_17_reg ( .D(io_i0_s3), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_17), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_19_reg ( .D(p_rand_37), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_19), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z60_reg ( .D(n_hpc2_0_N49), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n120) );
  DFF_X1 u_hpc2_0__hpc1_ref_v0_reg ( .D(n_hpc2_0_N0), .CK(clock_0), .Q(
        n_hpc2_0_n3), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_18_reg ( .D(p_rand_36), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_18), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z64_reg ( .D(n_hpc2_0_N53), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n125) );
  DFF_X1 u_hpc2_0_reg_pipeline_24_reg ( .D(io_i0_s5), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_24), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z62_reg ( .D(n_hpc2_0_N51), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n122) );
  DFF_X1 u_hpc2_0_reg_pipeline_16_reg ( .D(p_rand_35), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_16), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_5_reg ( .D(p_rand_26), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_5), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_23_reg ( .D(p_rand_40), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_23), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_14_reg ( .D(p_rand_33), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_14), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_9_reg ( .D(p_rand_29), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_9), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(p_rand_25), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_4), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_22_reg ( .D(p_rand_39), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_22), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_12_reg ( .D(io_i0_s2), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_12), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v4_reg ( .D(n_hpc2_0_N4), .CK(clock_0), .Q(
        n_hpc2_0_n6), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_8_reg ( .D(p_rand_28), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_8), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(p_rand_24), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_3), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_21_reg ( .D(io_i0_s4), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_21), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_10_reg ( .D(p_rand_30), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_10), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v2_reg ( .D(n_hpc2_0_N2), .CK(clock_0), .Q(
        n_hpc2_0_n1), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v5_reg ( .D(n_hpc2_0_N5), .CK(clock_0), .Q(
        n_hpc2_0_n5), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_7_reg ( .D(p_rand_27), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_7), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_26_reg ( .D(io_i0_s6), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_26), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_20_reg ( .D(p_rand_38), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_20), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(p_rand_21), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_0), .QN() );
endmodule

