
module AesSbox_keyAdd ( clock, reset, io_state, io_key, io_out );
  input [7:0] io_state;
  input [7:0] io_key;
  output [7:0] io_out;
  input clock, reset;
  wire   sbox_io_o0, sbox_io_o1, sbox_io_o2, sbox_io_o3, sbox_io_o4,
         sbox_io_o5, sbox_io_o6, sbox_io_o7, sbox_n127, sbox_n126, sbox_n125,
         sbox_n124, sbox_n123, sbox_n122, sbox_n121, sbox_n120, sbox_n119,
         sbox_n118, sbox_n117, sbox_n116, sbox_n115, sbox_n114, sbox_n113,
         sbox_n112, sbox_n111, sbox_n110, sbox_n109, sbox_n108, sbox_n107,
         sbox_n106, sbox_n105, sbox_n104, sbox_n103, sbox_n102, sbox_n101,
         sbox_n100, sbox_n99, sbox_n98, sbox_n97, sbox_n96, sbox_n95, sbox_n94,
         sbox_n93, sbox_n92, sbox_n91, sbox_n90, sbox_n89, sbox_n88, sbox_n87,
         sbox_n86, sbox_n85, sbox_n84, sbox_n83, sbox_n82, sbox_n81, sbox_n80,
         sbox_n79, sbox_n78, sbox_n77, sbox_n76, sbox_n75, sbox_n74, sbox_n73,
         sbox_n72, sbox_n71, sbox_n70, sbox_n69, sbox_n68, sbox_n67, sbox_n66,
         sbox_n65, sbox_n64, sbox_n63, sbox_n62, sbox_n61, sbox_n60, sbox_n59,
         sbox_n58, sbox_n57, sbox_n56, sbox_n55, sbox_n54, sbox_n53, sbox_n52,
         sbox_n51, sbox_n50, sbox_n49, sbox_n48, sbox_n47, sbox_n46, sbox_n45,
         sbox_n44, sbox_n43, sbox_n42, sbox_n41, sbox_n40, sbox_n39, sbox_n38,
         sbox_n37, sbox_n36, sbox_n35, sbox_n34, sbox_n33, sbox_n32, sbox_n31,
         sbox_n30, sbox_n29, sbox_n28, sbox_n27, sbox_n26, sbox_n25, sbox_n24,
         sbox_n23, sbox_n22, sbox_n21, sbox_n20, sbox_n19, sbox_n18, sbox_n17,
         sbox_n16, sbox_n15, sbox_n14, sbox_n13, sbox_n12, sbox_n11, sbox_n10,
         sbox_n9, sbox_n8, sbox_n7, sbox_n6, sbox_n5, sbox_n4, sbox_n3,
         sbox_n2, sbox_n1;

  XOR2_X1 U9 ( .A(sbox_io_o7), .B(io_key[7]), .Z(io_out[7]) );
  XOR2_X1 U10 ( .A(sbox_io_o6), .B(io_key[6]), .Z(io_out[6]) );
  XOR2_X1 U11 ( .A(sbox_io_o5), .B(io_key[5]), .Z(io_out[5]) );
  XOR2_X1 U12 ( .A(sbox_io_o4), .B(io_key[4]), .Z(io_out[4]) );
  XOR2_X1 U13 ( .A(sbox_io_o3), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 U14 ( .A(sbox_io_o2), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 U15 ( .A(sbox_io_o1), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 U16 ( .A(sbox_io_o0), .B(io_key[0]), .Z(io_out[0]) );
  XOR2_X1 sbox_U135 ( .A(io_state[0]), .B(io_state[3]), .Z(sbox_n72) );
  XOR2_X1 sbox_U134 ( .A(io_state[2]), .B(io_state[5]), .Z(sbox_n108) );
  XOR2_X1 sbox_U133 ( .A(sbox_n72), .B(sbox_n108), .Z(sbox_n78) );
  XOR2_X1 sbox_U132 ( .A(io_state[1]), .B(io_state[5]), .Z(sbox_n125) );
  XOR2_X1 sbox_U131 ( .A(io_state[6]), .B(io_state[4]), .Z(sbox_n124) );
  INV_X1 sbox_U130 ( .A(sbox_n124), .ZN(sbox_n109) );
  XNOR2_X1 sbox_U129 ( .A(sbox_n109), .B(sbox_n125), .ZN(sbox_n77) );
  NAND2_X1 sbox_U128 ( .A1(sbox_n77), .A2(sbox_n72), .ZN(sbox_n116) );
  XOR2_X1 sbox_U127 ( .A(io_state[3]), .B(io_state[5]), .Z(sbox_n74) );
  INV_X1 sbox_U126 ( .A(sbox_n74), .ZN(sbox_n123) );
  XNOR2_X1 sbox_U125 ( .A(sbox_n108), .B(sbox_n72), .ZN(sbox_n127) );
  NOR2_X1 sbox_U124 ( .A1(sbox_n123), .A2(sbox_n127), .ZN(sbox_n126) );
  XNOR2_X1 sbox_U123 ( .A(sbox_n116), .B(sbox_n126), .ZN(sbox_n101) );
  XNOR2_X1 sbox_U122 ( .A(sbox_n125), .B(sbox_n101), .ZN(sbox_n119) );
  XOR2_X1 sbox_U121 ( .A(sbox_n124), .B(sbox_n72), .Z(sbox_n62) );
  XOR2_X1 sbox_U120 ( .A(io_state[0]), .B(io_state[6]), .Z(sbox_n48) );
  XNOR2_X1 sbox_U119 ( .A(sbox_n123), .B(sbox_n48), .ZN(sbox_n64) );
  NAND2_X1 sbox_U118 ( .A1(sbox_n64), .A2(sbox_n62), .ZN(sbox_n114) );
  XOR2_X1 sbox_U117 ( .A(io_state[1]), .B(io_state[2]), .Z(sbox_n118) );
  XOR2_X1 sbox_U116 ( .A(io_state[7]), .B(sbox_n118), .Z(sbox_n68) );
  XOR2_X1 sbox_U115 ( .A(sbox_n68), .B(io_state[6]), .Z(sbox_n14) );
  XOR2_X1 sbox_U114 ( .A(io_state[0]), .B(io_state[5]), .Z(sbox_n43) );
  XNOR2_X1 sbox_U113 ( .A(sbox_n14), .B(sbox_n43), .ZN(sbox_n67) );
  XNOR2_X1 sbox_U112 ( .A(io_state[7]), .B(sbox_n62), .ZN(sbox_n59) );
  NOR2_X1 sbox_U111 ( .A1(sbox_n67), .A2(sbox_n59), .ZN(sbox_n122) );
  XOR2_X1 sbox_U110 ( .A(sbox_n114), .B(sbox_n122), .Z(sbox_n121) );
  XNOR2_X1 sbox_U109 ( .A(sbox_n62), .B(sbox_n121), .ZN(sbox_n120) );
  XNOR2_X1 sbox_U108 ( .A(sbox_n119), .B(sbox_n120), .ZN(sbox_n95) );
  INV_X1 sbox_U107 ( .A(sbox_n43), .ZN(sbox_n112) );
  XNOR2_X1 sbox_U106 ( .A(sbox_n118), .B(sbox_n62), .ZN(sbox_n45) );
  NOR2_X1 sbox_U105 ( .A1(sbox_n112), .A2(sbox_n45), .ZN(sbox_n117) );
  XOR2_X1 sbox_U104 ( .A(sbox_n116), .B(sbox_n117), .Z(sbox_n105) );
  XNOR2_X1 sbox_U103 ( .A(sbox_n105), .B(sbox_n45), .ZN(sbox_n110) );
  XOR2_X1 sbox_U102 ( .A(sbox_n68), .B(io_state[3]), .Z(sbox_n25) );
  AND2_X1 sbox_U101 ( .A1(sbox_n25), .A2(io_state[7]), .ZN(sbox_n115) );
  XNOR2_X1 sbox_U100 ( .A(sbox_n114), .B(sbox_n115), .ZN(sbox_n113) );
  XNOR2_X1 sbox_U99 ( .A(sbox_n112), .B(sbox_n113), .ZN(sbox_n111) );
  XNOR2_X1 sbox_U98 ( .A(sbox_n110), .B(sbox_n111), .ZN(sbox_n88) );
  INV_X1 sbox_U97 ( .A(sbox_n88), .ZN(sbox_n80) );
  XNOR2_X1 sbox_U96 ( .A(sbox_n95), .B(sbox_n80), .ZN(sbox_n82) );
  AND2_X1 sbox_U95 ( .A1(sbox_n95), .A2(sbox_n82), .ZN(sbox_n102) );
  XNOR2_X1 sbox_U94 ( .A(sbox_n108), .B(sbox_n109), .ZN(sbox_n75) );
  AND2_X1 sbox_U93 ( .A1(sbox_n75), .A2(sbox_n48), .ZN(sbox_n99) );
  XNOR2_X1 sbox_U92 ( .A(sbox_n25), .B(sbox_n72), .ZN(sbox_n50) );
  XNOR2_X1 sbox_U91 ( .A(sbox_n68), .B(sbox_n75), .ZN(sbox_n33) );
  NOR2_X1 sbox_U90 ( .A1(sbox_n50), .A2(sbox_n33), .ZN(sbox_n107) );
  XOR2_X1 sbox_U89 ( .A(sbox_n99), .B(sbox_n107), .Z(sbox_n106) );
  XOR2_X1 sbox_U88 ( .A(sbox_n105), .B(sbox_n106), .Z(sbox_n103) );
  XOR2_X1 sbox_U87 ( .A(sbox_n50), .B(sbox_n33), .Z(sbox_n104) );
  XNOR2_X1 sbox_U86 ( .A(sbox_n103), .B(sbox_n104), .ZN(sbox_n84) );
  NAND2_X1 sbox_U85 ( .A1(sbox_n102), .A2(sbox_n84), .ZN(sbox_n94) );
  XNOR2_X1 sbox_U84 ( .A(sbox_n75), .B(sbox_n101), .ZN(sbox_n96) );
  AND2_X1 sbox_U83 ( .A1(sbox_n68), .A2(sbox_n14), .ZN(sbox_n100) );
  XOR2_X1 sbox_U82 ( .A(sbox_n99), .B(sbox_n100), .Z(sbox_n98) );
  XOR2_X1 sbox_U81 ( .A(sbox_n48), .B(sbox_n98), .Z(sbox_n97) );
  XNOR2_X1 sbox_U80 ( .A(sbox_n96), .B(sbox_n97), .ZN(sbox_n92) );
  NAND2_X1 sbox_U79 ( .A1(sbox_n92), .A2(sbox_n95), .ZN(sbox_n83) );
  XNOR2_X1 sbox_U78 ( .A(sbox_n94), .B(sbox_n83), .ZN(sbox_n93) );
  XNOR2_X1 sbox_U77 ( .A(sbox_n93), .B(sbox_n82), .ZN(sbox_n13) );
  AND2_X1 sbox_U76 ( .A1(sbox_n88), .A2(sbox_n92), .ZN(sbox_n91) );
  XOR2_X1 sbox_U75 ( .A(sbox_n84), .B(sbox_n92), .Z(sbox_n87) );
  NAND2_X1 sbox_U74 ( .A1(sbox_n91), .A2(sbox_n87), .ZN(sbox_n90) );
  XNOR2_X1 sbox_U73 ( .A(sbox_n90), .B(sbox_n83), .ZN(sbox_n89) );
  XNOR2_X1 sbox_U72 ( .A(sbox_n89), .B(sbox_n87), .ZN(sbox_n65) );
  INV_X1 sbox_U71 ( .A(sbox_n65), .ZN(sbox_n60) );
  XNOR2_X1 sbox_U70 ( .A(sbox_n13), .B(sbox_n60), .ZN(sbox_n42) );
  INV_X1 sbox_U69 ( .A(sbox_n42), .ZN(sbox_n46) );
  XNOR2_X1 sbox_U68 ( .A(sbox_n83), .B(sbox_n88), .ZN(sbox_n86) );
  NAND2_X1 sbox_U67 ( .A1(sbox_n86), .A2(sbox_n87), .ZN(sbox_n85) );
  XNOR2_X1 sbox_U66 ( .A(sbox_n85), .B(sbox_n84), .ZN(sbox_n24) );
  INV_X1 sbox_U65 ( .A(sbox_n24), .ZN(sbox_n66) );
  XNOR2_X1 sbox_U64 ( .A(sbox_n83), .B(sbox_n84), .ZN(sbox_n81) );
  NAND2_X1 sbox_U63 ( .A1(sbox_n81), .A2(sbox_n82), .ZN(sbox_n79) );
  XOR2_X1 sbox_U62 ( .A(sbox_n79), .B(sbox_n80), .Z(sbox_n51) );
  XNOR2_X1 sbox_U61 ( .A(sbox_n66), .B(sbox_n51), .ZN(sbox_n71) );
  XNOR2_X1 sbox_U60 ( .A(sbox_n46), .B(sbox_n71), .ZN(sbox_n73) );
  NAND2_X1 sbox_U59 ( .A1(sbox_n78), .A2(sbox_n73), .ZN(sbox_n22) );
  NAND2_X1 sbox_U58 ( .A1(sbox_n77), .A2(sbox_n71), .ZN(sbox_n40) );
  XOR2_X1 sbox_U57 ( .A(sbox_n22), .B(sbox_n40), .Z(sbox_n56) );
  INV_X1 sbox_U56 ( .A(sbox_n13), .ZN(sbox_n76) );
  XNOR2_X1 sbox_U55 ( .A(sbox_n76), .B(sbox_n51), .ZN(sbox_n47) );
  NAND2_X1 sbox_U54 ( .A1(sbox_n47), .A2(sbox_n75), .ZN(sbox_n69) );
  NAND2_X1 sbox_U53 ( .A1(sbox_n73), .A2(sbox_n74), .ZN(sbox_n70) );
  AND2_X1 sbox_U52 ( .A1(sbox_n71), .A2(sbox_n72), .ZN(sbox_n41) );
  XNOR2_X1 sbox_U51 ( .A(sbox_n70), .B(sbox_n41), .ZN(sbox_n16) );
  XOR2_X1 sbox_U50 ( .A(sbox_n69), .B(sbox_n16), .Z(sbox_n6) );
  NAND2_X1 sbox_U49 ( .A1(sbox_n13), .A2(sbox_n68), .ZN(sbox_n15) );
  NOR2_X1 sbox_U48 ( .A1(sbox_n60), .A2(sbox_n67), .ZN(sbox_n55) );
  XOR2_X1 sbox_U47 ( .A(sbox_n15), .B(sbox_n55), .Z(sbox_n28) );
  XOR2_X1 sbox_U46 ( .A(sbox_n6), .B(sbox_n28), .Z(sbox_n35) );
  XNOR2_X1 sbox_U45 ( .A(sbox_n65), .B(sbox_n66), .ZN(sbox_n61) );
  AND2_X1 sbox_U44 ( .A1(sbox_n61), .A2(sbox_n64), .ZN(sbox_n57) );
  XNOR2_X1 sbox_U43 ( .A(sbox_n35), .B(sbox_n57), .ZN(sbox_n63) );
  XNOR2_X1 sbox_U42 ( .A(sbox_n56), .B(sbox_n63), .ZN(sbox_io_o0) );
  NAND2_X1 sbox_U41 ( .A1(sbox_n61), .A2(sbox_n62), .ZN(sbox_n52) );
  NOR2_X1 sbox_U40 ( .A1(sbox_n59), .A2(sbox_n60), .ZN(sbox_n58) );
  XOR2_X1 sbox_U39 ( .A(sbox_n57), .B(sbox_n58), .Z(sbox_n29) );
  XNOR2_X1 sbox_U38 ( .A(sbox_n52), .B(sbox_n29), .ZN(sbox_n34) );
  XNOR2_X1 sbox_U37 ( .A(sbox_n34), .B(sbox_n56), .ZN(sbox_n53) );
  XOR2_X1 sbox_U36 ( .A(sbox_n55), .B(sbox_n16), .Z(sbox_n54) );
  XOR2_X1 sbox_U35 ( .A(sbox_n53), .B(sbox_n54), .Z(sbox_io_o1) );
  AND2_X1 sbox_U34 ( .A1(io_state[7]), .A2(sbox_n24), .ZN(sbox_n31) );
  XNOR2_X1 sbox_U33 ( .A(sbox_n52), .B(sbox_n31), .ZN(sbox_n4) );
  INV_X1 sbox_U32 ( .A(sbox_n51), .ZN(sbox_n32) );
  NOR2_X1 sbox_U31 ( .A1(sbox_n50), .A2(sbox_n32), .ZN(sbox_n49) );
  XOR2_X1 sbox_U30 ( .A(sbox_n4), .B(sbox_n49), .Z(sbox_n20) );
  NAND2_X1 sbox_U29 ( .A1(sbox_n47), .A2(sbox_n48), .ZN(sbox_n7) );
  NOR2_X1 sbox_U28 ( .A1(sbox_n45), .A2(sbox_n46), .ZN(sbox_n44) );
  XNOR2_X1 sbox_U27 ( .A(sbox_n7), .B(sbox_n44), .ZN(sbox_n23) );
  XNOR2_X1 sbox_U26 ( .A(sbox_n20), .B(sbox_n23), .ZN(sbox_n36) );
  NAND2_X1 sbox_U25 ( .A1(sbox_n42), .A2(sbox_n43), .ZN(sbox_n38) );
  XOR2_X1 sbox_U24 ( .A(sbox_n40), .B(sbox_n41), .Z(sbox_n39) );
  XOR2_X1 sbox_U23 ( .A(sbox_n38), .B(sbox_n39), .Z(sbox_n37) );
  XOR2_X1 sbox_U22 ( .A(sbox_n36), .B(sbox_n37), .Z(sbox_io_o2) );
  INV_X1 sbox_U21 ( .A(sbox_n35), .ZN(sbox_n19) );
  XNOR2_X1 sbox_U20 ( .A(sbox_n19), .B(sbox_n34), .ZN(sbox_io_o3) );
  NOR2_X1 sbox_U19 ( .A1(sbox_n32), .A2(sbox_n33), .ZN(sbox_n12) );
  XOR2_X1 sbox_U18 ( .A(sbox_n31), .B(sbox_n12), .Z(sbox_n30) );
  XOR2_X1 sbox_U17 ( .A(sbox_n16), .B(sbox_n30), .Z(sbox_n26) );
  XNOR2_X1 sbox_U16 ( .A(sbox_n28), .B(sbox_n29), .ZN(sbox_n27) );
  XOR2_X1 sbox_U15 ( .A(sbox_n26), .B(sbox_n27), .Z(sbox_io_o4) );
  NAND2_X1 sbox_U14 ( .A1(sbox_n24), .A2(sbox_n25), .ZN(sbox_n21) );
  XOR2_X1 sbox_U13 ( .A(sbox_n22), .B(sbox_n23), .Z(sbox_n10) );
  XOR2_X1 sbox_U12 ( .A(sbox_n21), .B(sbox_n10), .Z(sbox_n17) );
  XNOR2_X1 sbox_U11 ( .A(sbox_n19), .B(sbox_n20), .ZN(sbox_n18) );
  XOR2_X1 sbox_U10 ( .A(sbox_n17), .B(sbox_n18), .Z(sbox_io_o5) );
  XOR2_X1 sbox_U9 ( .A(sbox_n15), .B(sbox_n16), .Z(sbox_n8) );
  NAND2_X1 sbox_U8 ( .A1(sbox_n13), .A2(sbox_n14), .ZN(sbox_n11) );
  XNOR2_X1 sbox_U7 ( .A(sbox_n11), .B(sbox_n12), .ZN(sbox_n5) );
  XNOR2_X1 sbox_U6 ( .A(sbox_n5), .B(sbox_n10), .ZN(sbox_n9) );
  XOR2_X1 sbox_U5 ( .A(sbox_n8), .B(sbox_n9), .Z(sbox_io_o6) );
  XNOR2_X1 sbox_U4 ( .A(sbox_n6), .B(sbox_n7), .ZN(sbox_n1) );
  INV_X1 sbox_U3 ( .A(sbox_n5), .ZN(sbox_n3) );
  XNOR2_X1 sbox_U2 ( .A(sbox_n3), .B(sbox_n4), .ZN(sbox_n2) );
  XOR2_X1 sbox_U1 ( .A(sbox_n1), .B(sbox_n2), .Z(sbox_io_o7) );
endmodule

