
module PresentSbox_keyAdd_detection_noFlag ( clock, reset, io_state, io_key, 
        io_out );
  input [3:0] io_state;
  input [3:0] io_key;
  output [3:0] io_out;
  input clock, reset;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         PresentSbox_keyAdd_sbox_io_o3, PresentSbox_keyAdd_sbox_io_o2,
         PresentSbox_keyAdd_sbox_io_o1, PresentSbox_keyAdd_sbox_io_o0,
         PresentSbox_keyAdd_sbox_n18, PresentSbox_keyAdd_sbox_n17,
         PresentSbox_keyAdd_sbox_n16, PresentSbox_keyAdd_sbox_n15,
         PresentSbox_keyAdd_sbox_n14, PresentSbox_keyAdd_sbox_n13,
         PresentSbox_keyAdd_sbox_n12, PresentSbox_keyAdd_sbox_n11,
         PresentSbox_keyAdd_sbox_n10, PresentSbox_keyAdd_sbox_n9,
         PresentSbox_keyAdd_sbox_n8, PresentSbox_keyAdd_sbox_n7,
         PresentSbox_keyAdd_sbox_n6, PresentSbox_keyAdd_sbox_n5,
         PresentSbox_keyAdd_sbox_n4, PresentSbox_keyAdd_sbox_n3,
         PresentSbox_keyAdd_sbox_n2, PresentSbox_keyAdd_sbox_n1,
         PresentSbox_keyAdd_1_sbox_io_o3, PresentSbox_keyAdd_1_sbox_io_o2,
         PresentSbox_keyAdd_1_sbox_io_o1, PresentSbox_keyAdd_1_sbox_io_o0,
         PresentSbox_keyAdd_1_sbox_n18, PresentSbox_keyAdd_1_sbox_n17,
         PresentSbox_keyAdd_1_sbox_n16, PresentSbox_keyAdd_1_sbox_n15,
         PresentSbox_keyAdd_1_sbox_n14, PresentSbox_keyAdd_1_sbox_n13,
         PresentSbox_keyAdd_1_sbox_n12, PresentSbox_keyAdd_1_sbox_n11,
         PresentSbox_keyAdd_1_sbox_n10, PresentSbox_keyAdd_1_sbox_n9,
         PresentSbox_keyAdd_1_sbox_n8, PresentSbox_keyAdd_1_sbox_n7,
         PresentSbox_keyAdd_1_sbox_n6, PresentSbox_keyAdd_1_sbox_n5,
         PresentSbox_keyAdd_1_sbox_n4, PresentSbox_keyAdd_1_sbox_n3,
         PresentSbox_keyAdd_1_sbox_n2, PresentSbox_keyAdd_1_sbox_n1;
  wire   [3:0] output_sbox_0;
  wire   [3:0] output_sbox_1;
  wire io_state0, io_state1, io_state2, io_state3;

  BUF_X1 B00 ( .A(io_state[0]), .Z(io_state0) );
  BUF_X1 B01 ( .A(io_state[1]), .Z(io_state1) );
  BUF_X1 B02 ( .A(io_state[2]), .Z(io_state2) );
  BUF_X1 B03 ( .A(io_state[3]), .Z(io_state3) );

  NOR2_X1 det_U16 ( .A1(n12), .A2(n13), .ZN(io_out[3]) );
  INV_X1 det_U17 ( .A(output_sbox_0[3]), .ZN(n12) );
  NOR2_X1 det_U18 ( .A1(n14), .A2(n13), .ZN(io_out[2]) );
  INV_X1 det_U19 ( .A(output_sbox_0[2]), .ZN(n14) );
  NOR2_X1 det_U20 ( .A1(n15), .A2(n13), .ZN(io_out[1]) );
  INV_X1 det_U21 ( .A(output_sbox_0[1]), .ZN(n15) );
  NOR2_X1 det_U22 ( .A1(n16), .A2(n13), .ZN(io_out[0]) );
  NAND2_X1 det_U23 ( .A1(n17), .A2(n18), .ZN(n13) );
  NOR2_X1 det_U24 ( .A1(n19), .A2(n20), .ZN(n18) );
  XOR2_X1 det_U25 ( .A(output_sbox_1[1]), .B(output_sbox_0[1]), .Z(n20) );
  XOR2_X1 det_U26 ( .A(output_sbox_1[0]), .B(output_sbox_0[0]), .Z(n19) );
  NOR2_X1 det_U27 ( .A1(n21), .A2(n22), .ZN(n17) );
  XOR2_X1 det_U28 ( .A(output_sbox_1[3]), .B(output_sbox_0[3]), .Z(n22) );
  XOR2_X1 det_U29 ( .A(output_sbox_1[2]), .B(output_sbox_0[2]), .Z(n21) );
  INV_X1 det_U30 ( .A(output_sbox_0[0]), .ZN(n16) );
  XOR2_X1 PresentSbox_keyAdd_U4 ( .A(PresentSbox_keyAdd_sbox_io_o0), .B(
        io_key[0]), .Z(output_sbox_0[0]) );
  XOR2_X1 PresentSbox_keyAdd_U3 ( .A(PresentSbox_keyAdd_sbox_io_o1), .B(
        io_key[1]), .Z(output_sbox_0[1]) );
  XOR2_X1 PresentSbox_keyAdd_U2 ( .A(PresentSbox_keyAdd_sbox_io_o2), .B(
        io_key[2]), .Z(output_sbox_0[2]) );
  XOR2_X1 PresentSbox_keyAdd_U1 ( .A(PresentSbox_keyAdd_sbox_io_o3), .B(
        io_key[3]), .Z(output_sbox_0[3]) );
  INV_X1 PresentSbox_keyAdd_sbox_U022 ( .A(io_state[1]), .ZN(
        PresentSbox_keyAdd_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U021 ( .A1(PresentSbox_keyAdd_sbox_n18), .A2(
        io_state[2]), .ZN(PresentSbox_keyAdd_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_sbox_U020 ( .A1(io_state[2]), .A2(
        PresentSbox_keyAdd_sbox_n18), .ZN(PresentSbox_keyAdd_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_sbox_U019 ( .A1(PresentSbox_keyAdd_sbox_n1), .A2(
        PresentSbox_keyAdd_sbox_n17), .ZN(PresentSbox_keyAdd_sbox_n13) );
  INV_X1 PresentSbox_keyAdd_sbox_U018 ( .A(io_state[3]), .ZN(
        PresentSbox_keyAdd_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U017 ( .A(PresentSbox_keyAdd_sbox_n13), .B(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n15) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U016 ( .A1(PresentSbox_keyAdd_sbox_n13), .A2(
        io_state[0]), .ZN(PresentSbox_keyAdd_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_sbox_U015 ( .A1(PresentSbox_keyAdd_sbox_n11), .A2(
        PresentSbox_keyAdd_sbox_n1), .ZN(PresentSbox_keyAdd_sbox_n14) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U014 ( .A(io_state[0]), .B(io_state[2]), 
        .ZN(PresentSbox_keyAdd_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U013 ( .A(PresentSbox_keyAdd_sbox_n14), .B(
        PresentSbox_keyAdd_sbox_n4), .Z(PresentSbox_keyAdd_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_sbox_U012 ( .A1(PresentSbox_keyAdd_sbox_n15), 
        .A2(PresentSbox_keyAdd_sbox_n16), .ZN(PresentSbox_keyAdd_sbox_n3) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U011 ( .A(PresentSbox_keyAdd_sbox_n14), .B(
        io_state[3]), .ZN(PresentSbox_keyAdd_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U010 ( .A(PresentSbox_keyAdd_sbox_n3), .B(
        PresentSbox_keyAdd_sbox_n6), .Z(PresentSbox_keyAdd_sbox_io_o0) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U009 ( .A(io_state[0]), .B(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U008 ( .A(PresentSbox_keyAdd_sbox_n13), .B(
        PresentSbox_keyAdd_sbox_n2), .Z(PresentSbox_keyAdd_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U007 ( .A1(PresentSbox_keyAdd_sbox_n11), .A2(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n10) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U006 ( .A(PresentSbox_keyAdd_sbox_n4), .B(
        PresentSbox_keyAdd_sbox_n10), .Z(PresentSbox_keyAdd_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_sbox_U005 ( .A1(PresentSbox_keyAdd_sbox_n8), .A2(
        PresentSbox_keyAdd_sbox_n9), .ZN(PresentSbox_keyAdd_sbox_n7) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U004 ( .A(PresentSbox_keyAdd_sbox_n7), .B(
        io_state[2]), .Z(PresentSbox_keyAdd_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U003 ( .A(PresentSbox_keyAdd_sbox_n5), .B(
        PresentSbox_keyAdd_sbox_n6), .Z(PresentSbox_keyAdd_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U002 ( .A(PresentSbox_keyAdd_sbox_n3), .B(
        PresentSbox_keyAdd_sbox_n4), .Z(PresentSbox_keyAdd_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U001 ( .A(PresentSbox_keyAdd_sbox_n1), .B(
        PresentSbox_keyAdd_sbox_n2), .Z(PresentSbox_keyAdd_sbox_io_o3) );
  XOR2_X1 PresentSbox_keyAdd_1_U4 ( .A(PresentSbox_keyAdd_1_sbox_io_o0), .B(
        io_key[0]), .Z(output_sbox_1[0]) );
  XOR2_X1 PresentSbox_keyAdd_1_U3 ( .A(PresentSbox_keyAdd_1_sbox_io_o1), .B(
        io_key[1]), .Z(output_sbox_1[1]) );
  XOR2_X1 PresentSbox_keyAdd_1_U2 ( .A(PresentSbox_keyAdd_1_sbox_io_o2), .B(
        io_key[2]), .Z(output_sbox_1[2]) );
  XOR2_X1 PresentSbox_keyAdd_1_U1 ( .A(PresentSbox_keyAdd_1_sbox_io_o3), .B(
        io_key[3]), .Z(output_sbox_1[3]) );
  INV_X1 PresentSbox_keyAdd_1_sbox_U022 ( .A(io_state1), .ZN(
        PresentSbox_keyAdd_1_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U021 ( .A1(PresentSbox_keyAdd_1_sbox_n18), 
        .A2(io_state2), .ZN(PresentSbox_keyAdd_1_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_1_sbox_U020 ( .A1(io_state2), .A2(
        PresentSbox_keyAdd_1_sbox_n18), .ZN(PresentSbox_keyAdd_1_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U019 ( .A1(PresentSbox_keyAdd_1_sbox_n1), 
        .A2(PresentSbox_keyAdd_1_sbox_n17), .ZN(PresentSbox_keyAdd_1_sbox_n13)
         );
  INV_X1 PresentSbox_keyAdd_1_sbox_U018 ( .A(io_state3), .ZN(
        PresentSbox_keyAdd_1_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U017 ( .A(PresentSbox_keyAdd_1_sbox_n13), 
        .B(PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n15)
         );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U016 ( .A1(PresentSbox_keyAdd_1_sbox_n13), 
        .A2(io_state0), .ZN(PresentSbox_keyAdd_1_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U015 ( .A1(PresentSbox_keyAdd_1_sbox_n11), 
        .A2(PresentSbox_keyAdd_1_sbox_n1), .ZN(PresentSbox_keyAdd_1_sbox_n14)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U014 ( .A(io_state0), .B(io_state2), 
        .ZN(PresentSbox_keyAdd_1_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U013 ( .A(PresentSbox_keyAdd_1_sbox_n14), 
        .B(PresentSbox_keyAdd_1_sbox_n4), .Z(PresentSbox_keyAdd_1_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U012 ( .A1(PresentSbox_keyAdd_1_sbox_n15), 
        .A2(PresentSbox_keyAdd_1_sbox_n16), .ZN(PresentSbox_keyAdd_1_sbox_n3)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U011 ( .A(PresentSbox_keyAdd_1_sbox_n14), 
        .B(io_state3), .ZN(PresentSbox_keyAdd_1_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U010 ( .A(PresentSbox_keyAdd_1_sbox_n3), 
        .B(PresentSbox_keyAdd_1_sbox_n6), .Z(PresentSbox_keyAdd_1_sbox_io_o0)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U009 ( .A(io_state0), .B(
        PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U008 ( .A(PresentSbox_keyAdd_1_sbox_n13), 
        .B(PresentSbox_keyAdd_1_sbox_n2), .Z(PresentSbox_keyAdd_1_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U007 ( .A1(PresentSbox_keyAdd_1_sbox_n11), 
        .A2(PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n10)
         );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U006 ( .A(PresentSbox_keyAdd_1_sbox_n4), .B(
        PresentSbox_keyAdd_1_sbox_n10), .Z(PresentSbox_keyAdd_1_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U005 ( .A1(PresentSbox_keyAdd_1_sbox_n8), 
        .A2(PresentSbox_keyAdd_1_sbox_n9), .ZN(PresentSbox_keyAdd_1_sbox_n7)
         );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U004 ( .A(PresentSbox_keyAdd_1_sbox_n7), .B(
        io_state2), .Z(PresentSbox_keyAdd_1_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U003 ( .A(PresentSbox_keyAdd_1_sbox_n5), .B(
        PresentSbox_keyAdd_1_sbox_n6), .Z(PresentSbox_keyAdd_1_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U002 ( .A(PresentSbox_keyAdd_1_sbox_n3), .B(
        PresentSbox_keyAdd_1_sbox_n4), .Z(PresentSbox_keyAdd_1_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U001 ( .A(PresentSbox_keyAdd_1_sbox_n1), .B(
        PresentSbox_keyAdd_1_sbox_n2), .Z(PresentSbox_keyAdd_1_sbox_io_o3) );
endmodule

