
module Shared_Chi5_SifaTest ( port_a_in, port_b_in, port_c_in, port_d_in, 
        port_e_in, port_rand, port_det_out );
  input [1:0] port_a_in;
  input [1:0] port_b_in;
  input [1:0] port_c_in;
  input [1:0] port_d_in;
  input [1:0] port_e_in;
  input [0:0] port_rand;
  output [1:0] port_det_out;
  wire   chi5_1_port_e_out_1_, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         chi5_0_st0_t0_n2, chi5_0_st0_t0_n1, chi5_0_st0_t2_n1,
         chi5_0_st0_t1_n2, chi5_0_st0_t1_n1, chi5_0_st0_t3_n1,
         chi5_0_st1_t0_n2, chi5_0_st1_t0_n1, chi5_0_st1_t2_n1,
         chi5_0_st1_t1_n2, chi5_0_st1_t1_n1, chi5_0_st1_t3_n1,
         chi5_0_st2_t0_n2, chi5_0_st2_t0_n1, chi5_0_st2_t2_n1,
         chi5_0_st2_t1_n2, chi5_0_st2_t1_n1, chi5_0_st2_t3_n1,
         chi5_0_st3_t0_n2, chi5_0_st3_t0_n1, chi5_0_st3_t2_n1,
         chi5_0_st3_t1_n2, chi5_0_st3_t1_n1, chi5_0_st3_t3_n1,
         chi5_0_st4_t0_n2, chi5_0_st4_t0_n1, chi5_0_st4_t2_n1,
         chi5_0_st4_t1_n2, chi5_0_st4_t1_n1, chi5_0_st4_t3_n1,
         chi5_1_port_e_out_0_, chi5_1_st0_t0_n2, chi5_1_st0_t0_n1,
         chi5_1_st0_t2_n1, chi5_1_st0_t1_n2, chi5_1_st0_t1_n1,
         chi5_1_st0_t3_n1, chi5_1_st1_t0_n2, chi5_1_st1_t0_n1,
         chi5_1_st1_t2_n1, chi5_1_st1_t1_n2, chi5_1_st1_t1_n1,
         chi5_1_st1_t3_n1, chi5_1_st2_t0_n2, chi5_1_st2_t0_n1,
         chi5_1_st2_t2_n1, chi5_1_st2_t1_n2, chi5_1_st2_t1_n1,
         chi5_1_st2_t3_n1, chi5_1_st3_t0_n2, chi5_1_st3_t0_n1,
         chi5_1_st3_t2_n1, chi5_1_st3_t1_n2, chi5_1_st3_t1_n1,
         chi5_1_st3_t3_n1, chi5_1_st4_t0_n2, chi5_1_st4_t0_n1,
         chi5_1_st4_t2_n1, chi5_1_st4_t1_n2, chi5_1_st4_t1_n1,
         chi5_1_st4_t3_n1;
  wire   [1:0] chi5_0_port_a_out;
  wire   [1:0] chi5_0_port_b_out;
  wire   [1:0] chi5_0_port_c_out;
  wire   [1:0] chi5_0_port_d_out;
  wire   [1:0] chi5_0_port_e_out;
  wire   [1:0] chi5_1_port_a_out;
  wire   [1:0] chi5_1_port_b_out;
  wire   [1:0] chi5_1_port_c_out;
  wire   [1:0] chi5_1_port_d_out;
  wire   [1:0] chi5_0__zz_port_d_out_1;
  wire   [1:0] chi5_0_st0_a_temp;
  wire   [1:0] chi5_0_st1_a_temp;
  wire   [1:0] chi5_0_st2_a_temp;
  wire   [1:0] chi5_0_st3_a_temp;
  wire   [1:0] chi5_0_st4_a_temp;
  wire   [1:0] chi5_1__zz_port_d_out_1;
  wire   [1:0] chi5_1_st0_a_temp;
  wire   [1:0] chi5_1_st1_a_temp;
  wire   [1:0] chi5_1_st2_a_temp;
  wire   [1:0] chi5_1_st3_a_temp;
  wire   [1:0] chi5_1_st4_a_temp;
  wire port_a_in0, port_a_in1;

  BUF_X1 B00 ( .A(port_a_in[0]), .Z(port_a_in0) );
  BUF_X1 B01 ( .A(port_a_in[1]), .Z(port_a_in1) );

  NOR2_X1 U19 ( .A1(n17), .A2(n18), .ZN(port_det_out[1]) );
  NAND2_X1 U20 ( .A1(n19), .A2(n20), .ZN(n18) );
  XNOR2_X1 U21 ( .A(chi5_1_port_a_out[1]), .B(chi5_0_port_a_out[1]), .ZN(n20)
         );
  XNOR2_X1 U22 ( .A(chi5_1_port_b_out[1]), .B(chi5_0_port_b_out[1]), .ZN(n19)
         );
  NAND2_X1 U23 ( .A1(n21), .A2(n22), .ZN(n17) );
  XNOR2_X1 U24 ( .A(chi5_1_port_d_out[1]), .B(chi5_0_port_d_out[1]), .ZN(n22)
         );
  NOR2_X1 U25 ( .A1(n23), .A2(n24), .ZN(n21) );
  XOR2_X1 U26 ( .A(chi5_1_port_c_out[1]), .B(chi5_0_port_c_out[1]), .Z(n24) );
  XOR2_X1 U27 ( .A(chi5_1_port_e_out_1_), .B(chi5_0_port_e_out[1]), .Z(n23) );
  NOR2_X1 U28 ( .A1(n25), .A2(n26), .ZN(port_det_out[0]) );
  NAND2_X1 U29 ( .A1(n27), .A2(n28), .ZN(n26) );
  XNOR2_X1 U30 ( .A(chi5_1_port_b_out[0]), .B(chi5_0_port_b_out[0]), .ZN(n28)
         );
  NOR2_X1 U31 ( .A1(n29), .A2(n30), .ZN(n27) );
  NOR2_X1 U32 ( .A1(chi5_0_port_d_out[0]), .A2(n31), .ZN(n30) );
  NOR2_X1 U33 ( .A1(chi5_0_port_e_out[0]), .A2(n32), .ZN(n29) );
  INV_X1 U34 ( .A(chi5_0_port_d_out[0]), .ZN(n32) );
  NAND2_X1 U35 ( .A1(n33), .A2(n34), .ZN(n25) );
  XNOR2_X1 U36 ( .A(chi5_1_port_c_out[0]), .B(chi5_0_port_c_out[0]), .ZN(n34)
         );
  NOR2_X1 U37 ( .A1(n35), .A2(n36), .ZN(n33) );
  XOR2_X1 U38 ( .A(chi5_1_port_a_out[0]), .B(chi5_0_port_a_out[0]), .Z(n36) );
  AND2_X1 U39 ( .A1(n31), .A2(chi5_0_port_e_out[0]), .ZN(n35) );
  INV_X1 U40 ( .A(chi5_1_port_d_out[0]), .ZN(n31) );
  XOR2_X1 chi5_0_U2 ( .A(port_d_in[0]), .B(chi5_0__zz_port_d_out_1[0]), .Z(
        chi5_0_port_d_out[0]) );
  XOR2_X1 chi5_0_U1 ( .A(port_d_in[1]), .B(chi5_0__zz_port_d_out_1[1]), .Z(
        chi5_0_port_d_out[1]) );
  INV_X1 chi5_0_st0_t0_U3 ( .A(port_a_in1), .ZN(chi5_0_st0_t0_n2) );
  NOR2_X1 chi5_0_st0_t0_U2 ( .A1(port_e_in[0]), .A2(chi5_0_st0_t0_n2), .ZN(
        chi5_0_st0_t0_n1) );
  XOR2_X1 chi5_0_st0_t0_U1 ( .A(port_rand[0]), .B(chi5_0_st0_t0_n1), .Z(
        chi5_0_st0_a_temp[0]) );
  NAND2_X1 chi5_0_st0_t2_U2 ( .A1(port_a_in1), .A2(port_e_in[1]), .ZN(
        chi5_0_st0_t2_n1) );
  XNOR2_X1 chi5_0_st0_t2_U1 ( .A(port_rand[0]), .B(chi5_0_st0_t2_n1), .ZN(
        chi5_0_st0_a_temp[1]) );
  INV_X1 chi5_0_st0_t1_U3 ( .A(port_a_in0), .ZN(chi5_0_st0_t1_n2) );
  NOR2_X1 chi5_0_st0_t1_U2 ( .A1(port_e_in[0]), .A2(chi5_0_st0_t1_n2), .ZN(
        chi5_0_st0_t1_n1) );
  XOR2_X1 chi5_0_st0_t1_U1 ( .A(chi5_0_st0_a_temp[0]), .B(chi5_0_st0_t1_n1), 
        .Z(chi5_0__zz_port_d_out_1[0]) );
  NAND2_X1 chi5_0_st0_t3_U2 ( .A1(port_a_in0), .A2(port_e_in[1]), .ZN(
        chi5_0_st0_t3_n1) );
  XNOR2_X1 chi5_0_st0_t3_U1 ( .A(chi5_0_st0_a_temp[1]), .B(chi5_0_st0_t3_n1), 
        .ZN(chi5_0__zz_port_d_out_1[1]) );
  INV_X1 chi5_0_st1_t0_U3 ( .A(port_c_in[1]), .ZN(chi5_0_st1_t0_n2) );
  NOR2_X1 chi5_0_st1_t0_U2 ( .A1(port_b_in[0]), .A2(chi5_0_st1_t0_n2), .ZN(
        chi5_0_st1_t0_n1) );
  XOR2_X1 chi5_0_st1_t0_U1 ( .A(port_a_in0), .B(chi5_0_st1_t0_n1), .Z(
        chi5_0_st1_a_temp[0]) );
  NAND2_X1 chi5_0_st1_t2_U2 ( .A1(port_c_in[1]), .A2(port_b_in[1]), .ZN(
        chi5_0_st1_t2_n1) );
  XNOR2_X1 chi5_0_st1_t2_U1 ( .A(port_a_in1), .B(chi5_0_st1_t2_n1), .ZN(
        chi5_0_st1_a_temp[1]) );
  INV_X1 chi5_0_st1_t1_U3 ( .A(port_c_in[0]), .ZN(chi5_0_st1_t1_n2) );
  NOR2_X1 chi5_0_st1_t1_U2 ( .A1(port_b_in[0]), .A2(chi5_0_st1_t1_n2), .ZN(
        chi5_0_st1_t1_n1) );
  XOR2_X1 chi5_0_st1_t1_U1 ( .A(chi5_0_st1_a_temp[0]), .B(chi5_0_st1_t1_n1), 
        .Z(chi5_0_port_a_out[0]) );
  NAND2_X1 chi5_0_st1_t3_U2 ( .A1(port_c_in[0]), .A2(port_b_in[1]), .ZN(
        chi5_0_st1_t3_n1) );
  XNOR2_X1 chi5_0_st1_t3_U1 ( .A(chi5_0_st1_a_temp[1]), .B(chi5_0_st1_t3_n1), 
        .ZN(chi5_0_port_a_out[1]) );
  INV_X1 chi5_0_st2_t0_U3 ( .A(port_e_in[1]), .ZN(chi5_0_st2_t0_n2) );
  NOR2_X1 chi5_0_st2_t0_U2 ( .A1(port_d_in[0]), .A2(chi5_0_st2_t0_n2), .ZN(
        chi5_0_st2_t0_n1) );
  XOR2_X1 chi5_0_st2_t0_U1 ( .A(port_c_in[0]), .B(chi5_0_st2_t0_n1), .Z(
        chi5_0_st2_a_temp[0]) );
  NAND2_X1 chi5_0_st2_t2_U2 ( .A1(port_e_in[1]), .A2(port_d_in[1]), .ZN(
        chi5_0_st2_t2_n1) );
  XNOR2_X1 chi5_0_st2_t2_U1 ( .A(port_c_in[1]), .B(chi5_0_st2_t2_n1), .ZN(
        chi5_0_st2_a_temp[1]) );
  INV_X1 chi5_0_st2_t1_U3 ( .A(port_e_in[0]), .ZN(chi5_0_st2_t1_n2) );
  NOR2_X1 chi5_0_st2_t1_U2 ( .A1(port_d_in[0]), .A2(chi5_0_st2_t1_n2), .ZN(
        chi5_0_st2_t1_n1) );
  XOR2_X1 chi5_0_st2_t1_U1 ( .A(chi5_0_st2_a_temp[0]), .B(chi5_0_st2_t1_n1), 
        .Z(chi5_0_port_c_out[0]) );
  NAND2_X1 chi5_0_st2_t3_U2 ( .A1(port_e_in[0]), .A2(port_d_in[1]), .ZN(
        chi5_0_st2_t3_n1) );
  XNOR2_X1 chi5_0_st2_t3_U1 ( .A(chi5_0_st2_a_temp[1]), .B(chi5_0_st2_t3_n1), 
        .ZN(chi5_0_port_c_out[1]) );
  INV_X1 chi5_0_st3_t0_U3 ( .A(port_b_in[1]), .ZN(chi5_0_st3_t0_n2) );
  NOR2_X1 chi5_0_st3_t0_U2 ( .A1(port_a_in0), .A2(chi5_0_st3_t0_n2), .ZN(
        chi5_0_st3_t0_n1) );
  XOR2_X1 chi5_0_st3_t0_U1 ( .A(port_e_in[0]), .B(chi5_0_st3_t0_n1), .Z(
        chi5_0_st3_a_temp[0]) );
  NAND2_X1 chi5_0_st3_t2_U2 ( .A1(port_b_in[1]), .A2(port_a_in1), .ZN(
        chi5_0_st3_t2_n1) );
  XNOR2_X1 chi5_0_st3_t2_U1 ( .A(port_e_in[1]), .B(chi5_0_st3_t2_n1), .ZN(
        chi5_0_st3_a_temp[1]) );
  INV_X1 chi5_0_st3_t1_U3 ( .A(port_b_in[0]), .ZN(chi5_0_st3_t1_n2) );
  NOR2_X1 chi5_0_st3_t1_U2 ( .A1(port_a_in0), .A2(chi5_0_st3_t1_n2), .ZN(
        chi5_0_st3_t1_n1) );
  XOR2_X1 chi5_0_st3_t1_U1 ( .A(chi5_0_st3_a_temp[0]), .B(chi5_0_st3_t1_n1), 
        .Z(chi5_0_port_e_out[0]) );
  NAND2_X1 chi5_0_st3_t3_U2 ( .A1(port_b_in[0]), .A2(port_a_in1), .ZN(
        chi5_0_st3_t3_n1) );
  XNOR2_X1 chi5_0_st3_t3_U1 ( .A(chi5_0_st3_a_temp[1]), .B(chi5_0_st3_t3_n1), 
        .ZN(chi5_0_port_e_out[1]) );
  INV_X1 chi5_0_st4_t0_U3 ( .A(port_d_in[1]), .ZN(chi5_0_st4_t0_n2) );
  NOR2_X1 chi5_0_st4_t0_U2 ( .A1(port_c_in[0]), .A2(chi5_0_st4_t0_n2), .ZN(
        chi5_0_st4_t0_n1) );
  XOR2_X1 chi5_0_st4_t0_U1 ( .A(port_b_in[0]), .B(chi5_0_st4_t0_n1), .Z(
        chi5_0_st4_a_temp[0]) );
  NAND2_X1 chi5_0_st4_t2_U2 ( .A1(port_d_in[1]), .A2(port_c_in[1]), .ZN(
        chi5_0_st4_t2_n1) );
  XNOR2_X1 chi5_0_st4_t2_U1 ( .A(port_b_in[1]), .B(chi5_0_st4_t2_n1), .ZN(
        chi5_0_st4_a_temp[1]) );
  INV_X1 chi5_0_st4_t1_U3 ( .A(port_d_in[0]), .ZN(chi5_0_st4_t1_n2) );
  NOR2_X1 chi5_0_st4_t1_U2 ( .A1(port_c_in[0]), .A2(chi5_0_st4_t1_n2), .ZN(
        chi5_0_st4_t1_n1) );
  XOR2_X1 chi5_0_st4_t1_U1 ( .A(chi5_0_st4_a_temp[0]), .B(chi5_0_st4_t1_n1), 
        .Z(chi5_0_port_b_out[0]) );
  NAND2_X1 chi5_0_st4_t3_U2 ( .A1(port_d_in[0]), .A2(port_c_in[1]), .ZN(
        chi5_0_st4_t3_n1) );
  XNOR2_X1 chi5_0_st4_t3_U1 ( .A(chi5_0_st4_a_temp[1]), .B(chi5_0_st4_t3_n1), 
        .ZN(chi5_0_port_b_out[1]) );
  XOR2_X1 chi5_1_U2 ( .A(port_d_in[0]), .B(chi5_1__zz_port_d_out_1[0]), .Z(
        chi5_1_port_d_out[0]) );
  XOR2_X1 chi5_1_U1 ( .A(port_d_in[1]), .B(chi5_1__zz_port_d_out_1[1]), .Z(
        chi5_1_port_d_out[1]) );
  INV_X1 chi5_1_st0_t0_U3 ( .A(port_a_in[1]), .ZN(chi5_1_st0_t0_n2) );
  NOR2_X1 chi5_1_st0_t0_U2 ( .A1(port_e_in[0]), .A2(chi5_1_st0_t0_n2), .ZN(
        chi5_1_st0_t0_n1) );
  XOR2_X1 chi5_1_st0_t0_U1 ( .A(port_rand[0]), .B(chi5_1_st0_t0_n1), .Z(
        chi5_1_st0_a_temp[0]) );
  NAND2_X1 chi5_1_st0_t2_U2 ( .A1(port_a_in[1]), .A2(port_e_in[1]), .ZN(
        chi5_1_st0_t2_n1) );
  XNOR2_X1 chi5_1_st0_t2_U1 ( .A(port_rand[0]), .B(chi5_1_st0_t2_n1), .ZN(
        chi5_1_st0_a_temp[1]) );
  INV_X1 chi5_1_st0_t1_U3 ( .A(port_a_in[0]), .ZN(chi5_1_st0_t1_n2) );
  NOR2_X1 chi5_1_st0_t1_U2 ( .A1(port_e_in[0]), .A2(chi5_1_st0_t1_n2), .ZN(
        chi5_1_st0_t1_n1) );
  XOR2_X1 chi5_1_st0_t1_U1 ( .A(chi5_1_st0_a_temp[0]), .B(chi5_1_st0_t1_n1), 
        .Z(chi5_1__zz_port_d_out_1[0]) );
  NAND2_X1 chi5_1_st0_t3_U2 ( .A1(port_a_in[0]), .A2(port_e_in[1]), .ZN(
        chi5_1_st0_t3_n1) );
  XNOR2_X1 chi5_1_st0_t3_U1 ( .A(chi5_1_st0_a_temp[1]), .B(chi5_1_st0_t3_n1), 
        .ZN(chi5_1__zz_port_d_out_1[1]) );
  INV_X1 chi5_1_st1_t0_U3 ( .A(port_c_in[1]), .ZN(chi5_1_st1_t0_n2) );
  NOR2_X1 chi5_1_st1_t0_U2 ( .A1(port_b_in[0]), .A2(chi5_1_st1_t0_n2), .ZN(
        chi5_1_st1_t0_n1) );
  XOR2_X1 chi5_1_st1_t0_U1 ( .A(port_a_in[0]), .B(chi5_1_st1_t0_n1), .Z(
        chi5_1_st1_a_temp[0]) );
  NAND2_X1 chi5_1_st1_t2_U2 ( .A1(port_c_in[1]), .A2(port_b_in[1]), .ZN(
        chi5_1_st1_t2_n1) );
  XNOR2_X1 chi5_1_st1_t2_U1 ( .A(port_a_in[1]), .B(chi5_1_st1_t2_n1), .ZN(
        chi5_1_st1_a_temp[1]) );
  INV_X1 chi5_1_st1_t1_U3 ( .A(port_c_in[0]), .ZN(chi5_1_st1_t1_n2) );
  NOR2_X1 chi5_1_st1_t1_U2 ( .A1(port_b_in[0]), .A2(chi5_1_st1_t1_n2), .ZN(
        chi5_1_st1_t1_n1) );
  XOR2_X1 chi5_1_st1_t1_U1 ( .A(chi5_1_st1_a_temp[0]), .B(chi5_1_st1_t1_n1), 
        .Z(chi5_1_port_a_out[0]) );
  NAND2_X1 chi5_1_st1_t3_U2 ( .A1(port_c_in[0]), .A2(port_b_in[1]), .ZN(
        chi5_1_st1_t3_n1) );
  XNOR2_X1 chi5_1_st1_t3_U1 ( .A(chi5_1_st1_a_temp[1]), .B(chi5_1_st1_t3_n1), 
        .ZN(chi5_1_port_a_out[1]) );
  INV_X1 chi5_1_st2_t0_U3 ( .A(port_e_in[1]), .ZN(chi5_1_st2_t0_n2) );
  NOR2_X1 chi5_1_st2_t0_U2 ( .A1(port_d_in[0]), .A2(chi5_1_st2_t0_n2), .ZN(
        chi5_1_st2_t0_n1) );
  XOR2_X1 chi5_1_st2_t0_U1 ( .A(port_c_in[0]), .B(chi5_1_st2_t0_n1), .Z(
        chi5_1_st2_a_temp[0]) );
  NAND2_X1 chi5_1_st2_t2_U2 ( .A1(port_e_in[1]), .A2(port_d_in[1]), .ZN(
        chi5_1_st2_t2_n1) );
  XNOR2_X1 chi5_1_st2_t2_U1 ( .A(port_c_in[1]), .B(chi5_1_st2_t2_n1), .ZN(
        chi5_1_st2_a_temp[1]) );
  INV_X1 chi5_1_st2_t1_U3 ( .A(port_e_in[0]), .ZN(chi5_1_st2_t1_n2) );
  NOR2_X1 chi5_1_st2_t1_U2 ( .A1(port_d_in[0]), .A2(chi5_1_st2_t1_n2), .ZN(
        chi5_1_st2_t1_n1) );
  XOR2_X1 chi5_1_st2_t1_U1 ( .A(chi5_1_st2_a_temp[0]), .B(chi5_1_st2_t1_n1), 
        .Z(chi5_1_port_c_out[0]) );
  NAND2_X1 chi5_1_st2_t3_U2 ( .A1(port_e_in[0]), .A2(port_d_in[1]), .ZN(
        chi5_1_st2_t3_n1) );
  XNOR2_X1 chi5_1_st2_t3_U1 ( .A(chi5_1_st2_a_temp[1]), .B(chi5_1_st2_t3_n1), 
        .ZN(chi5_1_port_c_out[1]) );
  INV_X1 chi5_1_st3_t0_U3 ( .A(port_b_in[1]), .ZN(chi5_1_st3_t0_n2) );
  NOR2_X1 chi5_1_st3_t0_U2 ( .A1(port_a_in[0]), .A2(chi5_1_st3_t0_n2), .ZN(
        chi5_1_st3_t0_n1) );
  XOR2_X1 chi5_1_st3_t0_U1 ( .A(port_e_in[0]), .B(chi5_1_st3_t0_n1), .Z(
        chi5_1_st3_a_temp[0]) );
  NAND2_X1 chi5_1_st3_t2_U2 ( .A1(port_b_in[1]), .A2(port_a_in[1]), .ZN(
        chi5_1_st3_t2_n1) );
  XNOR2_X1 chi5_1_st3_t2_U1 ( .A(port_e_in[1]), .B(chi5_1_st3_t2_n1), .ZN(
        chi5_1_st3_a_temp[1]) );
  INV_X1 chi5_1_st3_t1_U3 ( .A(port_b_in[0]), .ZN(chi5_1_st3_t1_n2) );
  NOR2_X1 chi5_1_st3_t1_U2 ( .A1(port_a_in[0]), .A2(chi5_1_st3_t1_n2), .ZN(
        chi5_1_st3_t1_n1) );
  XOR2_X1 chi5_1_st3_t1_U1 ( .A(chi5_1_st3_a_temp[0]), .B(chi5_1_st3_t1_n1), 
        .Z(chi5_1_port_e_out_0_) );
  NAND2_X1 chi5_1_st3_t3_U2 ( .A1(port_b_in[0]), .A2(port_a_in[1]), .ZN(
        chi5_1_st3_t3_n1) );
  XNOR2_X1 chi5_1_st3_t3_U1 ( .A(chi5_1_st3_a_temp[1]), .B(chi5_1_st3_t3_n1), 
        .ZN(chi5_1_port_e_out_1_) );
  INV_X1 chi5_1_st4_t0_U3 ( .A(port_d_in[1]), .ZN(chi5_1_st4_t0_n2) );
  NOR2_X1 chi5_1_st4_t0_U2 ( .A1(port_c_in[0]), .A2(chi5_1_st4_t0_n2), .ZN(
        chi5_1_st4_t0_n1) );
  XOR2_X1 chi5_1_st4_t0_U1 ( .A(port_b_in[0]), .B(chi5_1_st4_t0_n1), .Z(
        chi5_1_st4_a_temp[0]) );
  NAND2_X1 chi5_1_st4_t2_U2 ( .A1(port_d_in[1]), .A2(port_c_in[1]), .ZN(
        chi5_1_st4_t2_n1) );
  XNOR2_X1 chi5_1_st4_t2_U1 ( .A(port_b_in[1]), .B(chi5_1_st4_t2_n1), .ZN(
        chi5_1_st4_a_temp[1]) );
  INV_X1 chi5_1_st4_t1_U3 ( .A(port_d_in[0]), .ZN(chi5_1_st4_t1_n2) );
  NOR2_X1 chi5_1_st4_t1_U2 ( .A1(port_c_in[0]), .A2(chi5_1_st4_t1_n2), .ZN(
        chi5_1_st4_t1_n1) );
  XOR2_X1 chi5_1_st4_t1_U1 ( .A(chi5_1_st4_a_temp[0]), .B(chi5_1_st4_t1_n1), 
        .Z(chi5_1_port_b_out[0]) );
  NAND2_X1 chi5_1_st4_t3_U2 ( .A1(port_d_in[0]), .A2(port_c_in[1]), .ZN(
        chi5_1_st4_t3_n1) );
  XNOR2_X1 chi5_1_st4_t3_U1 ( .A(chi5_1_st4_a_temp[1]), .B(chi5_1_st4_t3_n1), 
        .ZN(chi5_1_port_b_out[1]) );
endmodule

