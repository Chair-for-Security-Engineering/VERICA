
module CINI3 ( port_a_0, port_a_1, port_a_2, port_a_3, port_b_0, port_b_1, 
        port_b_2, port_b_3, port_c_0, port_c_1, port_c_2, port_c_3, 
        port_rand_ref, port_rand_mul, clk, reset );
  input [4:0] port_a_0;
  input [4:0] port_a_1;
  input [4:0] port_a_2;
  input [4:0] port_a_3;
  input [4:0] port_b_0;
  input [4:0] port_b_1;
  input [4:0] port_b_2;
  input [4:0] port_b_3;
  output [4:0] port_c_0;
  output [4:0] port_c_1;
  output [4:0] port_c_2;
  output [4:0] port_c_3;
  input [5:0] port_rand_ref;
  input [5:0] port_rand_mul;
  input clk, reset;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, ref_1_n40, ref_1_n39,
         ref_1_n38, ref_1_n37, ref_1_n36, ref_1_n35, ref_1_n34, ref_1_n33,
         ref_1_n32, ref_1_n31, ref_1_n30, ref_1_n29, ref_1_n28, ref_1_n27,
         ref_1_n26, ref_1_n25, ref_1_n24, ref_1_n23, ref_1_n22, ref_1_n21,
         ref_1_n20, ref_1_n19, ref_1_n18, ref_1_n17, ref_1_n16, ref_1_n15,
         ref_1_n14, ref_1_n13, ref_1_n12, ref_1_n11, ref_1_n10, ref_1_n9,
         ref_1_n8, ref_1_n7, ref_1_n6, ref_1_n5, ref_1_n4, ref_1_n3, ref_1_n2,
         ref_1_n1, ref_1_maj_159_port_o, ref_1_maj_158_port_o,
         ref_1_maj_157_port_o, ref_1_maj_156_port_o, ref_1_maj_155_port_o,
         ref_1_maj_154_port_o, ref_1_maj_153_port_o, ref_1_maj_152_port_o,
         ref_1_maj_151_port_o, ref_1_maj_150_port_o, ref_1_maj_149_port_o,
         ref_1_maj_148_port_o, ref_1_maj_147_port_o, ref_1_maj_146_port_o,
         ref_1_maj_145_port_o, ref_1_maj_144_port_o, ref_1_maj_143_port_o,
         ref_1_maj_142_port_o, ref_1_maj_141_port_o, ref_1_maj_140_port_o,
         ref_1_maj_139_port_o, ref_1_maj_138_port_o, ref_1_maj_137_port_o,
         ref_1_maj_136_port_o, ref_1_maj_135_port_o, ref_1_maj_134_port_o,
         ref_1_maj_133_port_o, ref_1_maj_132_port_o, ref_1_maj_131_port_o,
         ref_1_maj_130_port_o, ref_1_maj_129_port_o, ref_1_maj_128_port_o,
         ref_1_maj_127_port_o, ref_1_maj_126_port_o, ref_1_maj_125_port_o,
         ref_1_maj_124_port_o, ref_1_maj_123_port_o, ref_1_maj_122_port_o,
         ref_1_maj_121_port_o, ref_1_maj_120_port_o, ref_1_maj_119_port_o,
         ref_1_maj_118_port_o, ref_1_maj_117_port_o, ref_1_maj_116_port_o,
         ref_1_maj_115_port_o, ref_1_maj_114_port_o, ref_1_maj_113_port_o,
         ref_1_maj_112_port_o, ref_1_maj_111_port_o, ref_1_maj_110_port_o,
         ref_1_maj_109_port_o, ref_1_maj_108_port_o, ref_1_maj_107_port_o,
         ref_1_maj_106_port_o, ref_1_maj_105_port_o, ref_1_maj_104_port_o,
         ref_1_maj_103_port_o, ref_1_maj_102_port_o, ref_1_maj_101_port_o,
         ref_1_maj_100_port_o, ref_1_maj_99_port_o, ref_1_maj_98_port_o,
         ref_1_maj_97_port_o, ref_1_maj_96_port_o, ref_1_maj_95_port_o,
         ref_1_maj_94_port_o, ref_1_maj_93_port_o, ref_1_maj_92_port_o,
         ref_1_refreshed_3_0_, ref_1_refreshed_3_1_, ref_1_refreshed_3_2_,
         ref_1_refreshed_3_3_, ref_1_refreshed_3_4_, ref_1_maj_91_port_o,
         ref_1_maj_90_port_o, ref_1_maj_89_port_o, ref_1_maj_88_port_o,
         ref_1_refreshed_2_0_, ref_1_refreshed_2_1_, ref_1_refreshed_2_2_,
         ref_1_refreshed_2_3_, ref_1_refreshed_2_4_, ref_1_maj_87_port_o,
         ref_1_maj_86_port_o, ref_1_maj_85_port_o, ref_1_maj_84_port_o,
         ref_1_refreshed_1_0_, ref_1_refreshed_1_1_, ref_1_refreshed_1_2_,
         ref_1_refreshed_1_3_, ref_1_refreshed_1_4_, ref_1_maj_83_port_o,
         ref_1_maj_82_port_o, ref_1_maj_81_port_o, ref_1_maj_80_port_o,
         ref_1_refreshed_0_0_, ref_1_refreshed_0_1_, ref_1_refreshed_0_2_,
         ref_1_refreshed_0_3_, ref_1_refreshed_0_4_,
         ref_1_simpleXor_118_port_z, ref_1_simpleXor_117_port_z,
         ref_1_simpleXor_115_port_z, ref_1_simpleXor_114_port_z,
         ref_1_simpleXor_112_port_z, ref_1_simpleXor_111_port_z,
         ref_1_simpleXor_109_port_z, ref_1_simpleXor_108_port_z,
         ref_1_simpleXor_106_port_z, ref_1_simpleXor_105_port_z,
         ref_1_simpleXor_103_port_z, ref_1_simpleXor_102_port_z,
         ref_1_simpleXor_100_port_z, ref_1_simpleXor_99_port_z,
         ref_1_simpleXor_97_port_z, ref_1_simpleXor_96_port_z,
         ref_1_simpleXor_94_port_z, ref_1_simpleXor_93_port_z,
         ref_1_simpleXor_91_port_z, ref_1_simpleXor_90_port_z,
         ref_1_simpleXor_88_port_z, ref_1_simpleXor_87_port_z,
         ref_1_simpleXor_85_port_z, ref_1_simpleXor_84_port_z,
         ref_1_simpleXor_82_port_z, ref_1_simpleXor_81_port_z,
         ref_1_simpleXor_79_port_z, ref_1_simpleXor_78_port_z,
         ref_1_simpleXor_76_port_z, ref_1_simpleXor_75_port_z,
         ref_1_simpleXor_73_port_z, ref_1_simpleXor_72_port_z,
         ref_1_simpleXor_70_port_z, ref_1_simpleXor_69_port_z,
         ref_1_simpleXor_67_port_z, ref_1_simpleXor_66_port_z,
         ref_1_simpleXor_64_port_z, ref_1_simpleXor_63_port_z,
         ref_1_simpleXor_61_port_z, ref_1_simpleXor_60_port_z,
         ref_1_maj_80_n13, ref_1_maj_80_n12, ref_1_maj_80_n11,
         ref_1_maj_80_n10, ref_1_maj_80_n9, ref_1_maj_80_n8, ref_1_maj_80_n7,
         ref_1_maj_80_n6, ref_1_maj_80_n5, ref_1_maj_80_n4, ref_1_maj_80_n3,
         ref_1_maj_80_n2, ref_1_maj_80_n1, ref_1_maj_81_n26, ref_1_maj_81_n25,
         ref_1_maj_81_n24, ref_1_maj_81_n23, ref_1_maj_81_n22,
         ref_1_maj_81_n21, ref_1_maj_81_n20, ref_1_maj_81_n19,
         ref_1_maj_81_n18, ref_1_maj_81_n17, ref_1_maj_81_n16,
         ref_1_maj_81_n15, ref_1_maj_81_n14, ref_1_maj_82_n26,
         ref_1_maj_82_n25, ref_1_maj_82_n24, ref_1_maj_82_n23,
         ref_1_maj_82_n22, ref_1_maj_82_n21, ref_1_maj_82_n20,
         ref_1_maj_82_n19, ref_1_maj_82_n18, ref_1_maj_82_n17,
         ref_1_maj_82_n16, ref_1_maj_82_n15, ref_1_maj_82_n14,
         ref_1_maj_83_n26, ref_1_maj_83_n25, ref_1_maj_83_n24,
         ref_1_maj_83_n23, ref_1_maj_83_n22, ref_1_maj_83_n21,
         ref_1_maj_83_n20, ref_1_maj_83_n19, ref_1_maj_83_n18,
         ref_1_maj_83_n17, ref_1_maj_83_n16, ref_1_maj_83_n15,
         ref_1_maj_83_n14, ref_1_maj_84_n26, ref_1_maj_84_n25,
         ref_1_maj_84_n24, ref_1_maj_84_n23, ref_1_maj_84_n22,
         ref_1_maj_84_n21, ref_1_maj_84_n20, ref_1_maj_84_n19,
         ref_1_maj_84_n18, ref_1_maj_84_n17, ref_1_maj_84_n16,
         ref_1_maj_84_n15, ref_1_maj_84_n14, ref_1_maj_85_n26,
         ref_1_maj_85_n25, ref_1_maj_85_n24, ref_1_maj_85_n23,
         ref_1_maj_85_n22, ref_1_maj_85_n21, ref_1_maj_85_n20,
         ref_1_maj_85_n19, ref_1_maj_85_n18, ref_1_maj_85_n17,
         ref_1_maj_85_n16, ref_1_maj_85_n15, ref_1_maj_85_n14,
         ref_1_maj_86_n26, ref_1_maj_86_n25, ref_1_maj_86_n24,
         ref_1_maj_86_n23, ref_1_maj_86_n22, ref_1_maj_86_n21,
         ref_1_maj_86_n20, ref_1_maj_86_n19, ref_1_maj_86_n18,
         ref_1_maj_86_n17, ref_1_maj_86_n16, ref_1_maj_86_n15,
         ref_1_maj_86_n14, ref_1_maj_87_n26, ref_1_maj_87_n25,
         ref_1_maj_87_n24, ref_1_maj_87_n23, ref_1_maj_87_n22,
         ref_1_maj_87_n21, ref_1_maj_87_n20, ref_1_maj_87_n19,
         ref_1_maj_87_n18, ref_1_maj_87_n17, ref_1_maj_87_n16,
         ref_1_maj_87_n15, ref_1_maj_87_n14, ref_1_maj_88_n26,
         ref_1_maj_88_n25, ref_1_maj_88_n24, ref_1_maj_88_n23,
         ref_1_maj_88_n22, ref_1_maj_88_n21, ref_1_maj_88_n20,
         ref_1_maj_88_n19, ref_1_maj_88_n18, ref_1_maj_88_n17,
         ref_1_maj_88_n16, ref_1_maj_88_n15, ref_1_maj_88_n14,
         ref_1_maj_89_n26, ref_1_maj_89_n25, ref_1_maj_89_n24,
         ref_1_maj_89_n23, ref_1_maj_89_n22, ref_1_maj_89_n21,
         ref_1_maj_89_n20, ref_1_maj_89_n19, ref_1_maj_89_n18,
         ref_1_maj_89_n17, ref_1_maj_89_n16, ref_1_maj_89_n15,
         ref_1_maj_89_n14, ref_1_maj_90_n26, ref_1_maj_90_n25,
         ref_1_maj_90_n24, ref_1_maj_90_n23, ref_1_maj_90_n22,
         ref_1_maj_90_n21, ref_1_maj_90_n20, ref_1_maj_90_n19,
         ref_1_maj_90_n18, ref_1_maj_90_n17, ref_1_maj_90_n16,
         ref_1_maj_90_n15, ref_1_maj_90_n14, ref_1_maj_91_n26,
         ref_1_maj_91_n25, ref_1_maj_91_n24, ref_1_maj_91_n23,
         ref_1_maj_91_n22, ref_1_maj_91_n21, ref_1_maj_91_n20,
         ref_1_maj_91_n19, ref_1_maj_91_n18, ref_1_maj_91_n17,
         ref_1_maj_91_n16, ref_1_maj_91_n15, ref_1_maj_91_n14,
         ref_1_maj_92_n26, ref_1_maj_92_n25, ref_1_maj_92_n24,
         ref_1_maj_92_n23, ref_1_maj_92_n22, ref_1_maj_92_n21,
         ref_1_maj_92_n20, ref_1_maj_92_n19, ref_1_maj_92_n18,
         ref_1_maj_92_n17, ref_1_maj_92_n16, ref_1_maj_92_n15,
         ref_1_maj_92_n14, ref_1_maj_93_n26, ref_1_maj_93_n25,
         ref_1_maj_93_n24, ref_1_maj_93_n23, ref_1_maj_93_n22,
         ref_1_maj_93_n21, ref_1_maj_93_n20, ref_1_maj_93_n19,
         ref_1_maj_93_n18, ref_1_maj_93_n17, ref_1_maj_93_n16,
         ref_1_maj_93_n15, ref_1_maj_93_n14, ref_1_maj_94_n26,
         ref_1_maj_94_n25, ref_1_maj_94_n24, ref_1_maj_94_n23,
         ref_1_maj_94_n22, ref_1_maj_94_n21, ref_1_maj_94_n20,
         ref_1_maj_94_n19, ref_1_maj_94_n18, ref_1_maj_94_n17,
         ref_1_maj_94_n16, ref_1_maj_94_n15, ref_1_maj_94_n14,
         ref_1_maj_95_n26, ref_1_maj_95_n25, ref_1_maj_95_n24,
         ref_1_maj_95_n23, ref_1_maj_95_n22, ref_1_maj_95_n21,
         ref_1_maj_95_n20, ref_1_maj_95_n19, ref_1_maj_95_n18,
         ref_1_maj_95_n17, ref_1_maj_95_n16, ref_1_maj_95_n15,
         ref_1_maj_95_n14, ref_1_maj_96_n26, ref_1_maj_96_n25,
         ref_1_maj_96_n24, ref_1_maj_96_n23, ref_1_maj_96_n22,
         ref_1_maj_96_n21, ref_1_maj_96_n20, ref_1_maj_96_n19,
         ref_1_maj_96_n18, ref_1_maj_96_n17, ref_1_maj_96_n16,
         ref_1_maj_96_n15, ref_1_maj_96_n14, ref_1_maj_97_n26,
         ref_1_maj_97_n25, ref_1_maj_97_n24, ref_1_maj_97_n23,
         ref_1_maj_97_n22, ref_1_maj_97_n21, ref_1_maj_97_n20,
         ref_1_maj_97_n19, ref_1_maj_97_n18, ref_1_maj_97_n17,
         ref_1_maj_97_n16, ref_1_maj_97_n15, ref_1_maj_97_n14,
         ref_1_maj_98_n26, ref_1_maj_98_n25, ref_1_maj_98_n24,
         ref_1_maj_98_n23, ref_1_maj_98_n22, ref_1_maj_98_n21,
         ref_1_maj_98_n20, ref_1_maj_98_n19, ref_1_maj_98_n18,
         ref_1_maj_98_n17, ref_1_maj_98_n16, ref_1_maj_98_n15,
         ref_1_maj_98_n14, ref_1_maj_99_n26, ref_1_maj_99_n25,
         ref_1_maj_99_n24, ref_1_maj_99_n23, ref_1_maj_99_n22,
         ref_1_maj_99_n21, ref_1_maj_99_n20, ref_1_maj_99_n19,
         ref_1_maj_99_n18, ref_1_maj_99_n17, ref_1_maj_99_n16,
         ref_1_maj_99_n15, ref_1_maj_99_n14, ref_1_maj_100_n26,
         ref_1_maj_100_n25, ref_1_maj_100_n24, ref_1_maj_100_n23,
         ref_1_maj_100_n22, ref_1_maj_100_n21, ref_1_maj_100_n20,
         ref_1_maj_100_n19, ref_1_maj_100_n18, ref_1_maj_100_n17,
         ref_1_maj_100_n16, ref_1_maj_100_n15, ref_1_maj_100_n14,
         ref_1_maj_101_n26, ref_1_maj_101_n25, ref_1_maj_101_n24,
         ref_1_maj_101_n23, ref_1_maj_101_n22, ref_1_maj_101_n21,
         ref_1_maj_101_n20, ref_1_maj_101_n19, ref_1_maj_101_n18,
         ref_1_maj_101_n17, ref_1_maj_101_n16, ref_1_maj_101_n15,
         ref_1_maj_101_n14, ref_1_maj_102_n26, ref_1_maj_102_n25,
         ref_1_maj_102_n24, ref_1_maj_102_n23, ref_1_maj_102_n22,
         ref_1_maj_102_n21, ref_1_maj_102_n20, ref_1_maj_102_n19,
         ref_1_maj_102_n18, ref_1_maj_102_n17, ref_1_maj_102_n16,
         ref_1_maj_102_n15, ref_1_maj_102_n14, ref_1_maj_103_n26,
         ref_1_maj_103_n25, ref_1_maj_103_n24, ref_1_maj_103_n23,
         ref_1_maj_103_n22, ref_1_maj_103_n21, ref_1_maj_103_n20,
         ref_1_maj_103_n19, ref_1_maj_103_n18, ref_1_maj_103_n17,
         ref_1_maj_103_n16, ref_1_maj_103_n15, ref_1_maj_103_n14,
         ref_1_maj_104_n26, ref_1_maj_104_n25, ref_1_maj_104_n24,
         ref_1_maj_104_n23, ref_1_maj_104_n22, ref_1_maj_104_n21,
         ref_1_maj_104_n20, ref_1_maj_104_n19, ref_1_maj_104_n18,
         ref_1_maj_104_n17, ref_1_maj_104_n16, ref_1_maj_104_n15,
         ref_1_maj_104_n14, ref_1_maj_105_n26, ref_1_maj_105_n25,
         ref_1_maj_105_n24, ref_1_maj_105_n23, ref_1_maj_105_n22,
         ref_1_maj_105_n21, ref_1_maj_105_n20, ref_1_maj_105_n19,
         ref_1_maj_105_n18, ref_1_maj_105_n17, ref_1_maj_105_n16,
         ref_1_maj_105_n15, ref_1_maj_105_n14, ref_1_maj_106_n26,
         ref_1_maj_106_n25, ref_1_maj_106_n24, ref_1_maj_106_n23,
         ref_1_maj_106_n22, ref_1_maj_106_n21, ref_1_maj_106_n20,
         ref_1_maj_106_n19, ref_1_maj_106_n18, ref_1_maj_106_n17,
         ref_1_maj_106_n16, ref_1_maj_106_n15, ref_1_maj_106_n14,
         ref_1_maj_107_n26, ref_1_maj_107_n25, ref_1_maj_107_n24,
         ref_1_maj_107_n23, ref_1_maj_107_n22, ref_1_maj_107_n21,
         ref_1_maj_107_n20, ref_1_maj_107_n19, ref_1_maj_107_n18,
         ref_1_maj_107_n17, ref_1_maj_107_n16, ref_1_maj_107_n15,
         ref_1_maj_107_n14, ref_1_maj_108_n26, ref_1_maj_108_n25,
         ref_1_maj_108_n24, ref_1_maj_108_n23, ref_1_maj_108_n22,
         ref_1_maj_108_n21, ref_1_maj_108_n20, ref_1_maj_108_n19,
         ref_1_maj_108_n18, ref_1_maj_108_n17, ref_1_maj_108_n16,
         ref_1_maj_108_n15, ref_1_maj_108_n14, ref_1_maj_109_n26,
         ref_1_maj_109_n25, ref_1_maj_109_n24, ref_1_maj_109_n23,
         ref_1_maj_109_n22, ref_1_maj_109_n21, ref_1_maj_109_n20,
         ref_1_maj_109_n19, ref_1_maj_109_n18, ref_1_maj_109_n17,
         ref_1_maj_109_n16, ref_1_maj_109_n15, ref_1_maj_109_n14,
         ref_1_maj_110_n26, ref_1_maj_110_n25, ref_1_maj_110_n24,
         ref_1_maj_110_n23, ref_1_maj_110_n22, ref_1_maj_110_n21,
         ref_1_maj_110_n20, ref_1_maj_110_n19, ref_1_maj_110_n18,
         ref_1_maj_110_n17, ref_1_maj_110_n16, ref_1_maj_110_n15,
         ref_1_maj_110_n14, ref_1_maj_111_n26, ref_1_maj_111_n25,
         ref_1_maj_111_n24, ref_1_maj_111_n23, ref_1_maj_111_n22,
         ref_1_maj_111_n21, ref_1_maj_111_n20, ref_1_maj_111_n19,
         ref_1_maj_111_n18, ref_1_maj_111_n17, ref_1_maj_111_n16,
         ref_1_maj_111_n15, ref_1_maj_111_n14, ref_1_maj_112_n26,
         ref_1_maj_112_n25, ref_1_maj_112_n24, ref_1_maj_112_n23,
         ref_1_maj_112_n22, ref_1_maj_112_n21, ref_1_maj_112_n20,
         ref_1_maj_112_n19, ref_1_maj_112_n18, ref_1_maj_112_n17,
         ref_1_maj_112_n16, ref_1_maj_112_n15, ref_1_maj_112_n14,
         ref_1_maj_113_n26, ref_1_maj_113_n25, ref_1_maj_113_n24,
         ref_1_maj_113_n23, ref_1_maj_113_n22, ref_1_maj_113_n21,
         ref_1_maj_113_n20, ref_1_maj_113_n19, ref_1_maj_113_n18,
         ref_1_maj_113_n17, ref_1_maj_113_n16, ref_1_maj_113_n15,
         ref_1_maj_113_n14, ref_1_maj_114_n26, ref_1_maj_114_n25,
         ref_1_maj_114_n24, ref_1_maj_114_n23, ref_1_maj_114_n22,
         ref_1_maj_114_n21, ref_1_maj_114_n20, ref_1_maj_114_n19,
         ref_1_maj_114_n18, ref_1_maj_114_n17, ref_1_maj_114_n16,
         ref_1_maj_114_n15, ref_1_maj_114_n14, ref_1_maj_115_n26,
         ref_1_maj_115_n25, ref_1_maj_115_n24, ref_1_maj_115_n23,
         ref_1_maj_115_n22, ref_1_maj_115_n21, ref_1_maj_115_n20,
         ref_1_maj_115_n19, ref_1_maj_115_n18, ref_1_maj_115_n17,
         ref_1_maj_115_n16, ref_1_maj_115_n15, ref_1_maj_115_n14,
         ref_1_maj_116_n26, ref_1_maj_116_n25, ref_1_maj_116_n24,
         ref_1_maj_116_n23, ref_1_maj_116_n22, ref_1_maj_116_n21,
         ref_1_maj_116_n20, ref_1_maj_116_n19, ref_1_maj_116_n18,
         ref_1_maj_116_n17, ref_1_maj_116_n16, ref_1_maj_116_n15,
         ref_1_maj_116_n14, ref_1_maj_117_n26, ref_1_maj_117_n25,
         ref_1_maj_117_n24, ref_1_maj_117_n23, ref_1_maj_117_n22,
         ref_1_maj_117_n21, ref_1_maj_117_n20, ref_1_maj_117_n19,
         ref_1_maj_117_n18, ref_1_maj_117_n17, ref_1_maj_117_n16,
         ref_1_maj_117_n15, ref_1_maj_117_n14, ref_1_maj_118_n26,
         ref_1_maj_118_n25, ref_1_maj_118_n24, ref_1_maj_118_n23,
         ref_1_maj_118_n22, ref_1_maj_118_n21, ref_1_maj_118_n20,
         ref_1_maj_118_n19, ref_1_maj_118_n18, ref_1_maj_118_n17,
         ref_1_maj_118_n16, ref_1_maj_118_n15, ref_1_maj_118_n14,
         ref_1_maj_119_n26, ref_1_maj_119_n25, ref_1_maj_119_n24,
         ref_1_maj_119_n23, ref_1_maj_119_n22, ref_1_maj_119_n21,
         ref_1_maj_119_n20, ref_1_maj_119_n19, ref_1_maj_119_n18,
         ref_1_maj_119_n17, ref_1_maj_119_n16, ref_1_maj_119_n15,
         ref_1_maj_119_n14, ref_1_maj_120_n26, ref_1_maj_120_n25,
         ref_1_maj_120_n24, ref_1_maj_120_n23, ref_1_maj_120_n22,
         ref_1_maj_120_n21, ref_1_maj_120_n20, ref_1_maj_120_n19,
         ref_1_maj_120_n18, ref_1_maj_120_n17, ref_1_maj_120_n16,
         ref_1_maj_120_n15, ref_1_maj_120_n14, ref_1_maj_121_n26,
         ref_1_maj_121_n25, ref_1_maj_121_n24, ref_1_maj_121_n23,
         ref_1_maj_121_n22, ref_1_maj_121_n21, ref_1_maj_121_n20,
         ref_1_maj_121_n19, ref_1_maj_121_n18, ref_1_maj_121_n17,
         ref_1_maj_121_n16, ref_1_maj_121_n15, ref_1_maj_121_n14,
         ref_1_maj_122_n26, ref_1_maj_122_n25, ref_1_maj_122_n24,
         ref_1_maj_122_n23, ref_1_maj_122_n22, ref_1_maj_122_n21,
         ref_1_maj_122_n20, ref_1_maj_122_n19, ref_1_maj_122_n18,
         ref_1_maj_122_n17, ref_1_maj_122_n16, ref_1_maj_122_n15,
         ref_1_maj_122_n14, ref_1_maj_123_n26, ref_1_maj_123_n25,
         ref_1_maj_123_n24, ref_1_maj_123_n23, ref_1_maj_123_n22,
         ref_1_maj_123_n21, ref_1_maj_123_n20, ref_1_maj_123_n19,
         ref_1_maj_123_n18, ref_1_maj_123_n17, ref_1_maj_123_n16,
         ref_1_maj_123_n15, ref_1_maj_123_n14, ref_1_maj_124_n26,
         ref_1_maj_124_n25, ref_1_maj_124_n24, ref_1_maj_124_n23,
         ref_1_maj_124_n22, ref_1_maj_124_n21, ref_1_maj_124_n20,
         ref_1_maj_124_n19, ref_1_maj_124_n18, ref_1_maj_124_n17,
         ref_1_maj_124_n16, ref_1_maj_124_n15, ref_1_maj_124_n14,
         ref_1_maj_125_n26, ref_1_maj_125_n25, ref_1_maj_125_n24,
         ref_1_maj_125_n23, ref_1_maj_125_n22, ref_1_maj_125_n21,
         ref_1_maj_125_n20, ref_1_maj_125_n19, ref_1_maj_125_n18,
         ref_1_maj_125_n17, ref_1_maj_125_n16, ref_1_maj_125_n15,
         ref_1_maj_125_n14, ref_1_maj_126_n26, ref_1_maj_126_n25,
         ref_1_maj_126_n24, ref_1_maj_126_n23, ref_1_maj_126_n22,
         ref_1_maj_126_n21, ref_1_maj_126_n20, ref_1_maj_126_n19,
         ref_1_maj_126_n18, ref_1_maj_126_n17, ref_1_maj_126_n16,
         ref_1_maj_126_n15, ref_1_maj_126_n14, ref_1_maj_127_n26,
         ref_1_maj_127_n25, ref_1_maj_127_n24, ref_1_maj_127_n23,
         ref_1_maj_127_n22, ref_1_maj_127_n21, ref_1_maj_127_n20,
         ref_1_maj_127_n19, ref_1_maj_127_n18, ref_1_maj_127_n17,
         ref_1_maj_127_n16, ref_1_maj_127_n15, ref_1_maj_127_n14,
         ref_1_maj_128_n26, ref_1_maj_128_n25, ref_1_maj_128_n24,
         ref_1_maj_128_n23, ref_1_maj_128_n22, ref_1_maj_128_n21,
         ref_1_maj_128_n20, ref_1_maj_128_n19, ref_1_maj_128_n18,
         ref_1_maj_128_n17, ref_1_maj_128_n16, ref_1_maj_128_n15,
         ref_1_maj_128_n14, ref_1_maj_129_n26, ref_1_maj_129_n25,
         ref_1_maj_129_n24, ref_1_maj_129_n23, ref_1_maj_129_n22,
         ref_1_maj_129_n21, ref_1_maj_129_n20, ref_1_maj_129_n19,
         ref_1_maj_129_n18, ref_1_maj_129_n17, ref_1_maj_129_n16,
         ref_1_maj_129_n15, ref_1_maj_129_n14, ref_1_maj_130_n26,
         ref_1_maj_130_n25, ref_1_maj_130_n24, ref_1_maj_130_n23,
         ref_1_maj_130_n22, ref_1_maj_130_n21, ref_1_maj_130_n20,
         ref_1_maj_130_n19, ref_1_maj_130_n18, ref_1_maj_130_n17,
         ref_1_maj_130_n16, ref_1_maj_130_n15, ref_1_maj_130_n14,
         ref_1_maj_131_n26, ref_1_maj_131_n25, ref_1_maj_131_n24,
         ref_1_maj_131_n23, ref_1_maj_131_n22, ref_1_maj_131_n21,
         ref_1_maj_131_n20, ref_1_maj_131_n19, ref_1_maj_131_n18,
         ref_1_maj_131_n17, ref_1_maj_131_n16, ref_1_maj_131_n15,
         ref_1_maj_131_n14, ref_1_maj_132_n26, ref_1_maj_132_n25,
         ref_1_maj_132_n24, ref_1_maj_132_n23, ref_1_maj_132_n22,
         ref_1_maj_132_n21, ref_1_maj_132_n20, ref_1_maj_132_n19,
         ref_1_maj_132_n18, ref_1_maj_132_n17, ref_1_maj_132_n16,
         ref_1_maj_132_n15, ref_1_maj_132_n14, ref_1_maj_133_n26,
         ref_1_maj_133_n25, ref_1_maj_133_n24, ref_1_maj_133_n23,
         ref_1_maj_133_n22, ref_1_maj_133_n21, ref_1_maj_133_n20,
         ref_1_maj_133_n19, ref_1_maj_133_n18, ref_1_maj_133_n17,
         ref_1_maj_133_n16, ref_1_maj_133_n15, ref_1_maj_133_n14,
         ref_1_maj_134_n26, ref_1_maj_134_n25, ref_1_maj_134_n24,
         ref_1_maj_134_n23, ref_1_maj_134_n22, ref_1_maj_134_n21,
         ref_1_maj_134_n20, ref_1_maj_134_n19, ref_1_maj_134_n18,
         ref_1_maj_134_n17, ref_1_maj_134_n16, ref_1_maj_134_n15,
         ref_1_maj_134_n14, ref_1_maj_135_n26, ref_1_maj_135_n25,
         ref_1_maj_135_n24, ref_1_maj_135_n23, ref_1_maj_135_n22,
         ref_1_maj_135_n21, ref_1_maj_135_n20, ref_1_maj_135_n19,
         ref_1_maj_135_n18, ref_1_maj_135_n17, ref_1_maj_135_n16,
         ref_1_maj_135_n15, ref_1_maj_135_n14, ref_1_maj_136_n26,
         ref_1_maj_136_n25, ref_1_maj_136_n24, ref_1_maj_136_n23,
         ref_1_maj_136_n22, ref_1_maj_136_n21, ref_1_maj_136_n20,
         ref_1_maj_136_n19, ref_1_maj_136_n18, ref_1_maj_136_n17,
         ref_1_maj_136_n16, ref_1_maj_136_n15, ref_1_maj_136_n14,
         ref_1_maj_137_n26, ref_1_maj_137_n25, ref_1_maj_137_n24,
         ref_1_maj_137_n23, ref_1_maj_137_n22, ref_1_maj_137_n21,
         ref_1_maj_137_n20, ref_1_maj_137_n19, ref_1_maj_137_n18,
         ref_1_maj_137_n17, ref_1_maj_137_n16, ref_1_maj_137_n15,
         ref_1_maj_137_n14, ref_1_maj_138_n26, ref_1_maj_138_n25,
         ref_1_maj_138_n24, ref_1_maj_138_n23, ref_1_maj_138_n22,
         ref_1_maj_138_n21, ref_1_maj_138_n20, ref_1_maj_138_n19,
         ref_1_maj_138_n18, ref_1_maj_138_n17, ref_1_maj_138_n16,
         ref_1_maj_138_n15, ref_1_maj_138_n14, ref_1_maj_139_n26,
         ref_1_maj_139_n25, ref_1_maj_139_n24, ref_1_maj_139_n23,
         ref_1_maj_139_n22, ref_1_maj_139_n21, ref_1_maj_139_n20,
         ref_1_maj_139_n19, ref_1_maj_139_n18, ref_1_maj_139_n17,
         ref_1_maj_139_n16, ref_1_maj_139_n15, ref_1_maj_139_n14,
         ref_1_maj_140_n26, ref_1_maj_140_n25, ref_1_maj_140_n24,
         ref_1_maj_140_n23, ref_1_maj_140_n22, ref_1_maj_140_n21,
         ref_1_maj_140_n20, ref_1_maj_140_n19, ref_1_maj_140_n18,
         ref_1_maj_140_n17, ref_1_maj_140_n16, ref_1_maj_140_n15,
         ref_1_maj_140_n14, ref_1_maj_141_n26, ref_1_maj_141_n25,
         ref_1_maj_141_n24, ref_1_maj_141_n23, ref_1_maj_141_n22,
         ref_1_maj_141_n21, ref_1_maj_141_n20, ref_1_maj_141_n19,
         ref_1_maj_141_n18, ref_1_maj_141_n17, ref_1_maj_141_n16,
         ref_1_maj_141_n15, ref_1_maj_141_n14, ref_1_maj_142_n26,
         ref_1_maj_142_n25, ref_1_maj_142_n24, ref_1_maj_142_n23,
         ref_1_maj_142_n22, ref_1_maj_142_n21, ref_1_maj_142_n20,
         ref_1_maj_142_n19, ref_1_maj_142_n18, ref_1_maj_142_n17,
         ref_1_maj_142_n16, ref_1_maj_142_n15, ref_1_maj_142_n14,
         ref_1_maj_143_n26, ref_1_maj_143_n25, ref_1_maj_143_n24,
         ref_1_maj_143_n23, ref_1_maj_143_n22, ref_1_maj_143_n21,
         ref_1_maj_143_n20, ref_1_maj_143_n19, ref_1_maj_143_n18,
         ref_1_maj_143_n17, ref_1_maj_143_n16, ref_1_maj_143_n15,
         ref_1_maj_143_n14, ref_1_maj_144_n26, ref_1_maj_144_n25,
         ref_1_maj_144_n24, ref_1_maj_144_n23, ref_1_maj_144_n22,
         ref_1_maj_144_n21, ref_1_maj_144_n20, ref_1_maj_144_n19,
         ref_1_maj_144_n18, ref_1_maj_144_n17, ref_1_maj_144_n16,
         ref_1_maj_144_n15, ref_1_maj_144_n14, ref_1_maj_145_n26,
         ref_1_maj_145_n25, ref_1_maj_145_n24, ref_1_maj_145_n23,
         ref_1_maj_145_n22, ref_1_maj_145_n21, ref_1_maj_145_n20,
         ref_1_maj_145_n19, ref_1_maj_145_n18, ref_1_maj_145_n17,
         ref_1_maj_145_n16, ref_1_maj_145_n15, ref_1_maj_145_n14,
         ref_1_maj_146_n26, ref_1_maj_146_n25, ref_1_maj_146_n24,
         ref_1_maj_146_n23, ref_1_maj_146_n22, ref_1_maj_146_n21,
         ref_1_maj_146_n20, ref_1_maj_146_n19, ref_1_maj_146_n18,
         ref_1_maj_146_n17, ref_1_maj_146_n16, ref_1_maj_146_n15,
         ref_1_maj_146_n14, ref_1_maj_147_n26, ref_1_maj_147_n25,
         ref_1_maj_147_n24, ref_1_maj_147_n23, ref_1_maj_147_n22,
         ref_1_maj_147_n21, ref_1_maj_147_n20, ref_1_maj_147_n19,
         ref_1_maj_147_n18, ref_1_maj_147_n17, ref_1_maj_147_n16,
         ref_1_maj_147_n15, ref_1_maj_147_n14, ref_1_maj_148_n26,
         ref_1_maj_148_n25, ref_1_maj_148_n24, ref_1_maj_148_n23,
         ref_1_maj_148_n22, ref_1_maj_148_n21, ref_1_maj_148_n20,
         ref_1_maj_148_n19, ref_1_maj_148_n18, ref_1_maj_148_n17,
         ref_1_maj_148_n16, ref_1_maj_148_n15, ref_1_maj_148_n14,
         ref_1_maj_149_n26, ref_1_maj_149_n25, ref_1_maj_149_n24,
         ref_1_maj_149_n23, ref_1_maj_149_n22, ref_1_maj_149_n21,
         ref_1_maj_149_n20, ref_1_maj_149_n19, ref_1_maj_149_n18,
         ref_1_maj_149_n17, ref_1_maj_149_n16, ref_1_maj_149_n15,
         ref_1_maj_149_n14, ref_1_maj_150_n26, ref_1_maj_150_n25,
         ref_1_maj_150_n24, ref_1_maj_150_n23, ref_1_maj_150_n22,
         ref_1_maj_150_n21, ref_1_maj_150_n20, ref_1_maj_150_n19,
         ref_1_maj_150_n18, ref_1_maj_150_n17, ref_1_maj_150_n16,
         ref_1_maj_150_n15, ref_1_maj_150_n14, ref_1_maj_151_n26,
         ref_1_maj_151_n25, ref_1_maj_151_n24, ref_1_maj_151_n23,
         ref_1_maj_151_n22, ref_1_maj_151_n21, ref_1_maj_151_n20,
         ref_1_maj_151_n19, ref_1_maj_151_n18, ref_1_maj_151_n17,
         ref_1_maj_151_n16, ref_1_maj_151_n15, ref_1_maj_151_n14,
         ref_1_maj_152_n26, ref_1_maj_152_n25, ref_1_maj_152_n24,
         ref_1_maj_152_n23, ref_1_maj_152_n22, ref_1_maj_152_n21,
         ref_1_maj_152_n20, ref_1_maj_152_n19, ref_1_maj_152_n18,
         ref_1_maj_152_n17, ref_1_maj_152_n16, ref_1_maj_152_n15,
         ref_1_maj_152_n14, ref_1_maj_153_n26, ref_1_maj_153_n25,
         ref_1_maj_153_n24, ref_1_maj_153_n23, ref_1_maj_153_n22,
         ref_1_maj_153_n21, ref_1_maj_153_n20, ref_1_maj_153_n19,
         ref_1_maj_153_n18, ref_1_maj_153_n17, ref_1_maj_153_n16,
         ref_1_maj_153_n15, ref_1_maj_153_n14, ref_1_maj_154_n26,
         ref_1_maj_154_n25, ref_1_maj_154_n24, ref_1_maj_154_n23,
         ref_1_maj_154_n22, ref_1_maj_154_n21, ref_1_maj_154_n20,
         ref_1_maj_154_n19, ref_1_maj_154_n18, ref_1_maj_154_n17,
         ref_1_maj_154_n16, ref_1_maj_154_n15, ref_1_maj_154_n14,
         ref_1_maj_155_n26, ref_1_maj_155_n25, ref_1_maj_155_n24,
         ref_1_maj_155_n23, ref_1_maj_155_n22, ref_1_maj_155_n21,
         ref_1_maj_155_n20, ref_1_maj_155_n19, ref_1_maj_155_n18,
         ref_1_maj_155_n17, ref_1_maj_155_n16, ref_1_maj_155_n15,
         ref_1_maj_155_n14, ref_1_maj_156_n26, ref_1_maj_156_n25,
         ref_1_maj_156_n24, ref_1_maj_156_n23, ref_1_maj_156_n22,
         ref_1_maj_156_n21, ref_1_maj_156_n20, ref_1_maj_156_n19,
         ref_1_maj_156_n18, ref_1_maj_156_n17, ref_1_maj_156_n16,
         ref_1_maj_156_n15, ref_1_maj_156_n14, ref_1_maj_157_n26,
         ref_1_maj_157_n25, ref_1_maj_157_n24, ref_1_maj_157_n23,
         ref_1_maj_157_n22, ref_1_maj_157_n21, ref_1_maj_157_n20,
         ref_1_maj_157_n19, ref_1_maj_157_n18, ref_1_maj_157_n17,
         ref_1_maj_157_n16, ref_1_maj_157_n15, ref_1_maj_157_n14,
         ref_1_maj_158_n26, ref_1_maj_158_n25, ref_1_maj_158_n24,
         ref_1_maj_158_n23, ref_1_maj_158_n22, ref_1_maj_158_n21,
         ref_1_maj_158_n20, ref_1_maj_158_n19, ref_1_maj_158_n18,
         ref_1_maj_158_n17, ref_1_maj_158_n16, ref_1_maj_158_n15,
         ref_1_maj_158_n14, ref_1_maj_159_n26, ref_1_maj_159_n25,
         ref_1_maj_159_n24, ref_1_maj_159_n23, ref_1_maj_159_n22,
         ref_1_maj_159_n21, ref_1_maj_159_n20, ref_1_maj_159_n19,
         ref_1_maj_159_n18, ref_1_maj_159_n17, ref_1_maj_159_n16,
         ref_1_maj_159_n15, ref_1_maj_159_n14;
  wire   [4:0] ref_1_port_o_0_0;
  wire   [4:0] ref_1_port_o_0_1;
  wire   [4:0] ref_1_port_o_0_2;
  wire   [4:0] ref_1_port_o_0_3;
  wire   [4:0] ref_1_port_o_1_0;
  wire   [4:0] ref_1_port_o_1_1;
  wire   [4:0] ref_1_port_o_1_2;
  wire   [4:0] ref_1_port_o_1_3;
  wire   [4:0] ref_1_port_o_2_0;
  wire   [4:0] ref_1_port_o_2_1;
  wire   [4:0] ref_1_port_o_2_2;
  wire   [4:0] ref_1_port_o_2_3;
  wire   [4:0] ref_1_port_o_3_0;
  wire   [4:0] ref_1_port_o_3_1;
  wire   [4:0] ref_1_port_o_3_2;
  wire   [4:0] ref_1_port_o_3_3;
  wire   [4:0] temp_0_0;
  wire   [4:0] mult_ab_0_1;
  wire   [4:0] mult_ab_0_2;
  wire   [4:0] mult_ab_0_3;
  wire   [4:0] temp_0_1;
  wire   [4:0] mult_ab_1_0;
  wire   [4:0] mult_ab_1_2;
  wire   [4:0] mult_ab_1_3;
  wire   [4:0] temp_0_2;
  wire   [4:0] mult_ab_2_0;
  wire   [4:0] mult_ab_2_1;
  wire   [4:0] mult_ab_2_3;
  wire   [4:0] temp_0_3;
  wire   [4:0] mult_ab_3_0;
  wire   [4:0] mult_ab_3_1;
  wire   [4:0] mult_ab_3_2;

  DFF_X1 mult_ab_0_0_reg_4_ ( .D(N64), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 mult_ab_0_0_reg_3_ ( .D(N48), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 mult_ab_0_0_reg_2_ ( .D(N32), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 mult_ab_0_0_reg_1_ ( .D(N16), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 mult_ab_0_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 mult_ab_3_3_reg_4_ ( .D(N79), .CK(clk), .Q(temp_0_3[4]), .QN() );
  DFF_X1 mult_ab_3_3_reg_3_ ( .D(N63), .CK(clk), .Q(temp_0_3[3]), .QN() );
  DFF_X1 mult_ab_3_3_reg_2_ ( .D(N47), .CK(clk), .Q(temp_0_3[2]), .QN() );
  DFF_X1 mult_ab_3_3_reg_1_ ( .D(N31), .CK(clk), .Q(temp_0_3[1]), .QN() );
  DFF_X1 mult_ab_3_3_reg_0_ ( .D(N15), .CK(clk), .Q(temp_0_3[0]), .QN() );
  DFF_X1 mult_ab_0_1_reg_4_ ( .D(N65), .CK(clk), .Q(mult_ab_0_1[4]), .QN() );
  DFF_X1 mult_ab_0_1_reg_3_ ( .D(N49), .CK(clk), .Q(mult_ab_0_1[3]), .QN() );
  DFF_X1 mult_ab_0_1_reg_2_ ( .D(N33), .CK(clk), .Q(mult_ab_0_1[2]), .QN() );
  DFF_X1 mult_ab_0_1_reg_1_ ( .D(N17), .CK(clk), .Q(mult_ab_0_1[1]), .QN() );
  DFF_X1 mult_ab_0_1_reg_0_ ( .D(N1), .CK(clk), .Q(mult_ab_0_1[0]), .QN() );
  DFF_X1 mult_ab_0_2_reg_4_ ( .D(N66), .CK(clk), .Q(mult_ab_0_2[4]), .QN() );
  DFF_X1 mult_ab_0_2_reg_3_ ( .D(N50), .CK(clk), .Q(mult_ab_0_2[3]), .QN() );
  DFF_X1 mult_ab_0_2_reg_2_ ( .D(N34), .CK(clk), .Q(mult_ab_0_2[2]), .QN() );
  DFF_X1 mult_ab_0_2_reg_1_ ( .D(N18), .CK(clk), .Q(mult_ab_0_2[1]), .QN() );
  DFF_X1 mult_ab_0_2_reg_0_ ( .D(N2), .CK(clk), .Q(mult_ab_0_2[0]), .QN() );
  DFF_X1 mult_ab_2_3_reg_4_ ( .D(N75), .CK(clk), .Q(mult_ab_2_3[4]), .QN() );
  DFF_X1 mult_ab_2_3_reg_3_ ( .D(N59), .CK(clk), .Q(mult_ab_2_3[3]), .QN() );
  DFF_X1 mult_ab_2_3_reg_2_ ( .D(N43), .CK(clk), .Q(mult_ab_2_3[2]), .QN() );
  DFF_X1 mult_ab_2_3_reg_1_ ( .D(N27), .CK(clk), .Q(mult_ab_2_3[1]), .QN() );
  DFF_X1 mult_ab_2_3_reg_0_ ( .D(N11), .CK(clk), .Q(mult_ab_2_3[0]), .QN() );
  DFF_X1 mult_ab_1_3_reg_4_ ( .D(N71), .CK(clk), .Q(mult_ab_1_3[4]), .QN() );
  DFF_X1 mult_ab_1_3_reg_3_ ( .D(N55), .CK(clk), .Q(mult_ab_1_3[3]), .QN() );
  DFF_X1 mult_ab_1_3_reg_2_ ( .D(N39), .CK(clk), .Q(mult_ab_1_3[2]), .QN() );
  DFF_X1 mult_ab_1_3_reg_1_ ( .D(N23), .CK(clk), .Q(mult_ab_1_3[1]), .QN() );
  DFF_X1 mult_ab_1_3_reg_0_ ( .D(N7), .CK(clk), .Q(mult_ab_1_3[0]), .QN() );
  DFF_X1 mult_ab_0_3_reg_4_ ( .D(N67), .CK(clk), .Q(mult_ab_0_3[4]), .QN() );
  DFF_X1 mult_ab_0_3_reg_3_ ( .D(N51), .CK(clk), .Q(mult_ab_0_3[3]), .QN() );
  DFF_X1 mult_ab_0_3_reg_2_ ( .D(N35), .CK(clk), .Q(mult_ab_0_3[2]), .QN() );
  DFF_X1 mult_ab_0_3_reg_1_ ( .D(N19), .CK(clk), .Q(mult_ab_0_3[1]), .QN() );
  DFF_X1 mult_ab_0_3_reg_0_ ( .D(N3), .CK(clk), .Q(mult_ab_0_3[0]), .QN() );
  DFF_X1 mult_ab_3_1_reg_4_ ( .D(N77), .CK(clk), .Q(mult_ab_3_1[4]), .QN() );
  DFF_X1 mult_ab_3_1_reg_3_ ( .D(N61), .CK(clk), .Q(mult_ab_3_1[3]), .QN() );
  DFF_X1 mult_ab_3_1_reg_2_ ( .D(N45), .CK(clk), .Q(mult_ab_3_1[2]), .QN() );
  DFF_X1 mult_ab_3_1_reg_1_ ( .D(N29), .CK(clk), .Q(mult_ab_3_1[1]), .QN() );
  DFF_X1 mult_ab_3_1_reg_0_ ( .D(N13), .CK(clk), .Q(mult_ab_3_1[0]), .QN() );
  DFF_X1 mult_ab_1_1_reg_4_ ( .D(N69), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 mult_ab_1_1_reg_3_ ( .D(N53), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 mult_ab_1_1_reg_2_ ( .D(N37), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 mult_ab_1_1_reg_1_ ( .D(N21), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 mult_ab_1_1_reg_0_ ( .D(N5), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 mult_ab_3_0_reg_4_ ( .D(N76), .CK(clk), .Q(mult_ab_3_0[4]), .QN() );
  DFF_X1 mult_ab_3_0_reg_3_ ( .D(N60), .CK(clk), .Q(mult_ab_3_0[3]), .QN() );
  DFF_X1 mult_ab_3_0_reg_2_ ( .D(N44), .CK(clk), .Q(mult_ab_3_0[2]), .QN() );
  DFF_X1 mult_ab_3_0_reg_1_ ( .D(N28), .CK(clk), .Q(mult_ab_3_0[1]), .QN() );
  DFF_X1 mult_ab_3_0_reg_0_ ( .D(N12), .CK(clk), .Q(mult_ab_3_0[0]), .QN() );
  DFF_X1 mult_ab_2_2_reg_4_ ( .D(N74), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 mult_ab_2_2_reg_3_ ( .D(N58), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 mult_ab_2_2_reg_2_ ( .D(N42), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 mult_ab_2_2_reg_1_ ( .D(N26), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 mult_ab_2_2_reg_0_ ( .D(N10), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 mult_ab_3_2_reg_4_ ( .D(N78), .CK(clk), .Q(mult_ab_3_2[4]), .QN() );
  DFF_X1 mult_ab_3_2_reg_3_ ( .D(N62), .CK(clk), .Q(mult_ab_3_2[3]), .QN() );
  DFF_X1 mult_ab_3_2_reg_2_ ( .D(N46), .CK(clk), .Q(mult_ab_3_2[2]), .QN() );
  DFF_X1 mult_ab_3_2_reg_1_ ( .D(N30), .CK(clk), .Q(mult_ab_3_2[1]), .QN() );
  DFF_X1 mult_ab_3_2_reg_0_ ( .D(N14), .CK(clk), .Q(mult_ab_3_2[0]), .QN() );
  DFF_X1 mult_ab_1_2_reg_4_ ( .D(N70), .CK(clk), .Q(mult_ab_1_2[4]), .QN() );
  DFF_X1 mult_ab_1_2_reg_3_ ( .D(N54), .CK(clk), .Q(mult_ab_1_2[3]), .QN() );
  DFF_X1 mult_ab_1_2_reg_2_ ( .D(N38), .CK(clk), .Q(mult_ab_1_2[2]), .QN() );
  DFF_X1 mult_ab_1_2_reg_1_ ( .D(N22), .CK(clk), .Q(mult_ab_1_2[1]), .QN() );
  DFF_X1 mult_ab_1_2_reg_0_ ( .D(N6), .CK(clk), .Q(mult_ab_1_2[0]), .QN() );
  DFF_X1 mult_ab_2_0_reg_4_ ( .D(N72), .CK(clk), .Q(mult_ab_2_0[4]), .QN() );
  DFF_X1 mult_ab_2_0_reg_3_ ( .D(N56), .CK(clk), .Q(mult_ab_2_0[3]), .QN() );
  DFF_X1 mult_ab_2_0_reg_2_ ( .D(N40), .CK(clk), .Q(mult_ab_2_0[2]), .QN() );
  DFF_X1 mult_ab_2_0_reg_1_ ( .D(N24), .CK(clk), .Q(mult_ab_2_0[1]), .QN() );
  DFF_X1 mult_ab_2_0_reg_0_ ( .D(N8), .CK(clk), .Q(mult_ab_2_0[0]), .QN() );
  DFF_X1 mult_ab_2_1_reg_4_ ( .D(N73), .CK(clk), .Q(mult_ab_2_1[4]), .QN() );
  DFF_X1 mult_ab_2_1_reg_3_ ( .D(N57), .CK(clk), .Q(mult_ab_2_1[3]), .QN() );
  DFF_X1 mult_ab_2_1_reg_2_ ( .D(N41), .CK(clk), .Q(mult_ab_2_1[2]), .QN() );
  DFF_X1 mult_ab_2_1_reg_1_ ( .D(N25), .CK(clk), .Q(mult_ab_2_1[1]), .QN() );
  DFF_X1 mult_ab_2_1_reg_0_ ( .D(N9), .CK(clk), .Q(mult_ab_2_1[0]), .QN() );
  DFF_X1 mult_ab_1_0_reg_4_ ( .D(N68), .CK(clk), .Q(mult_ab_1_0[4]), .QN() );
  DFF_X1 mult_ab_1_0_reg_3_ ( .D(N52), .CK(clk), .Q(mult_ab_1_0[3]), .QN() );
  DFF_X1 mult_ab_1_0_reg_2_ ( .D(N36), .CK(clk), .Q(mult_ab_1_0[2]), .QN() );
  DFF_X1 mult_ab_1_0_reg_1_ ( .D(N20), .CK(clk), .Q(mult_ab_1_0[1]), .QN() );
  DFF_X1 mult_ab_1_0_reg_0_ ( .D(N4), .CK(clk), .Q(mult_ab_1_0[0]), .QN() );
  XNOR2_X1 U203 ( .A(port_rand_mul[0]), .B(n75), .ZN(N4) );
  NAND2_X1 U204 ( .A1(ref_1_port_o_1_0[0]), .A2(port_a_1[0]), .ZN(n75) );
  XNOR2_X1 U205 ( .A(port_rand_mul[0]), .B(n91), .ZN(N20) );
  NAND2_X1 U206 ( .A1(ref_1_port_o_1_0[1]), .A2(port_a_1[1]), .ZN(n91) );
  XNOR2_X1 U207 ( .A(port_rand_mul[0]), .B(n78), .ZN(N36) );
  NAND2_X1 U208 ( .A1(ref_1_port_o_1_0[2]), .A2(port_a_1[2]), .ZN(n78) );
  XNOR2_X1 U209 ( .A(port_rand_mul[0]), .B(n65), .ZN(N52) );
  NAND2_X1 U210 ( .A1(ref_1_port_o_1_0[3]), .A2(port_a_1[3]), .ZN(n65) );
  XNOR2_X1 U211 ( .A(port_rand_mul[0]), .B(n52), .ZN(N68) );
  NAND2_X1 U212 ( .A1(ref_1_port_o_1_0[4]), .A2(port_a_1[4]), .ZN(n52) );
  XNOR2_X1 U213 ( .A(port_rand_mul[3]), .B(n41), .ZN(N9) );
  NAND2_X1 U214 ( .A1(ref_1_port_o_2_1[0]), .A2(port_a_2[0]), .ZN(n41) );
  XNOR2_X1 U215 ( .A(port_rand_mul[3]), .B(n87), .ZN(N25) );
  NAND2_X1 U216 ( .A1(ref_1_port_o_2_1[1]), .A2(port_a_2[1]), .ZN(n87) );
  XNOR2_X1 U217 ( .A(port_rand_mul[3]), .B(n73), .ZN(N41) );
  NAND2_X1 U218 ( .A1(ref_1_port_o_2_1[2]), .A2(port_a_2[2]), .ZN(n73) );
  XNOR2_X1 U219 ( .A(port_rand_mul[3]), .B(n61), .ZN(N57) );
  NAND2_X1 U220 ( .A1(ref_1_port_o_2_1[3]), .A2(port_a_2[3]), .ZN(n61) );
  XNOR2_X1 U221 ( .A(port_rand_mul[3]), .B(n47), .ZN(N73) );
  NAND2_X1 U222 ( .A1(ref_1_port_o_2_1[4]), .A2(port_a_2[4]), .ZN(n47) );
  XNOR2_X1 U223 ( .A(port_rand_mul[1]), .B(n42), .ZN(N8) );
  NAND2_X1 U224 ( .A1(ref_1_port_o_2_0[0]), .A2(port_a_2[0]), .ZN(n42) );
  XNOR2_X1 U225 ( .A(port_rand_mul[1]), .B(n88), .ZN(N24) );
  NAND2_X1 U226 ( .A1(ref_1_port_o_2_0[1]), .A2(port_a_2[1]), .ZN(n88) );
  XNOR2_X1 U227 ( .A(port_rand_mul[1]), .B(n74), .ZN(N40) );
  NAND2_X1 U228 ( .A1(ref_1_port_o_2_0[2]), .A2(port_a_2[2]), .ZN(n74) );
  XNOR2_X1 U229 ( .A(port_rand_mul[1]), .B(n62), .ZN(N56) );
  NAND2_X1 U230 ( .A1(ref_1_port_o_2_0[3]), .A2(port_a_2[3]), .ZN(n62) );
  XNOR2_X1 U231 ( .A(port_rand_mul[1]), .B(n48), .ZN(N72) );
  NAND2_X1 U232 ( .A1(ref_1_port_o_2_0[4]), .A2(port_a_2[4]), .ZN(n48) );
  XNOR2_X1 U233 ( .A(port_rand_mul[3]), .B(n59), .ZN(N6) );
  NAND2_X1 U234 ( .A1(ref_1_port_o_1_2[0]), .A2(port_a_1[0]), .ZN(n59) );
  XNOR2_X1 U235 ( .A(port_rand_mul[3]), .B(n90), .ZN(N22) );
  NAND2_X1 U236 ( .A1(ref_1_port_o_1_2[1]), .A2(port_a_1[1]), .ZN(n90) );
  XNOR2_X1 U237 ( .A(port_rand_mul[3]), .B(n77), .ZN(N38) );
  NAND2_X1 U238 ( .A1(ref_1_port_o_1_2[2]), .A2(port_a_1[2]), .ZN(n77) );
  XNOR2_X1 U239 ( .A(port_rand_mul[3]), .B(n64), .ZN(N54) );
  NAND2_X1 U240 ( .A1(ref_1_port_o_1_2[3]), .A2(port_a_1[3]), .ZN(n64) );
  XNOR2_X1 U241 ( .A(port_rand_mul[3]), .B(n50), .ZN(N70) );
  NAND2_X1 U242 ( .A1(ref_1_port_o_1_2[4]), .A2(port_a_1[4]), .ZN(n50) );
  XNOR2_X1 U243 ( .A(port_rand_mul[5]), .B(n96), .ZN(N14) );
  NAND2_X1 U244 ( .A1(ref_1_port_o_3_2[0]), .A2(port_a_3[0]), .ZN(n96) );
  XNOR2_X1 U245 ( .A(port_rand_mul[5]), .B(n82), .ZN(N30) );
  NAND2_X1 U246 ( .A1(ref_1_port_o_3_2[1]), .A2(port_a_3[1]), .ZN(n82) );
  XNOR2_X1 U247 ( .A(port_rand_mul[5]), .B(n69), .ZN(N46) );
  NAND2_X1 U248 ( .A1(ref_1_port_o_3_2[2]), .A2(port_a_3[2]), .ZN(n69) );
  XNOR2_X1 U249 ( .A(port_rand_mul[5]), .B(n56), .ZN(N62) );
  NAND2_X1 U250 ( .A1(ref_1_port_o_3_2[3]), .A2(port_a_3[3]), .ZN(n56) );
  XNOR2_X1 U251 ( .A(port_rand_mul[5]), .B(n43), .ZN(N78) );
  NAND2_X1 U252 ( .A1(ref_1_port_o_3_2[4]), .A2(port_a_3[4]), .ZN(n43) );
  XNOR2_X1 U253 ( .A(port_rand_mul[2]), .B(n98), .ZN(N12) );
  NAND2_X1 U254 ( .A1(ref_1_port_o_3_0[0]), .A2(port_a_3[0]), .ZN(n98) );
  XNOR2_X1 U255 ( .A(port_rand_mul[2]), .B(n85), .ZN(N28) );
  NAND2_X1 U256 ( .A1(ref_1_port_o_3_0[1]), .A2(port_a_3[1]), .ZN(n85) );
  XNOR2_X1 U257 ( .A(port_rand_mul[2]), .B(n71), .ZN(N44) );
  NAND2_X1 U258 ( .A1(ref_1_port_o_3_0[2]), .A2(port_a_3[2]), .ZN(n71) );
  XNOR2_X1 U259 ( .A(port_rand_mul[2]), .B(n58), .ZN(N60) );
  NAND2_X1 U260 ( .A1(ref_1_port_o_3_0[3]), .A2(port_a_3[3]), .ZN(n58) );
  XNOR2_X1 U261 ( .A(port_rand_mul[2]), .B(n45), .ZN(N76) );
  NAND2_X1 U262 ( .A1(ref_1_port_o_3_0[4]), .A2(port_a_3[4]), .ZN(n45) );
  XNOR2_X1 U263 ( .A(port_rand_mul[4]), .B(n97), .ZN(N13) );
  NAND2_X1 U264 ( .A1(ref_1_port_o_3_1[0]), .A2(port_a_3[0]), .ZN(n97) );
  XNOR2_X1 U265 ( .A(port_rand_mul[4]), .B(n84), .ZN(N29) );
  NAND2_X1 U266 ( .A1(ref_1_port_o_3_1[1]), .A2(port_a_3[1]), .ZN(n84) );
  XNOR2_X1 U267 ( .A(port_rand_mul[4]), .B(n70), .ZN(N45) );
  NAND2_X1 U268 ( .A1(ref_1_port_o_3_1[2]), .A2(port_a_3[2]), .ZN(n70) );
  XNOR2_X1 U269 ( .A(port_rand_mul[4]), .B(n57), .ZN(N61) );
  NAND2_X1 U270 ( .A1(ref_1_port_o_3_1[3]), .A2(port_a_3[3]), .ZN(n57) );
  XNOR2_X1 U271 ( .A(port_rand_mul[4]), .B(n44), .ZN(N77) );
  NAND2_X1 U272 ( .A1(ref_1_port_o_3_1[4]), .A2(port_a_3[4]), .ZN(n44) );
  XNOR2_X1 U273 ( .A(port_rand_mul[2]), .B(n83), .ZN(N3) );
  NAND2_X1 U274 ( .A1(ref_1_port_o_0_3[0]), .A2(port_a_0[0]), .ZN(n83) );
  XNOR2_X1 U275 ( .A(port_rand_mul[2]), .B(n93), .ZN(N19) );
  NAND2_X1 U276 ( .A1(ref_1_port_o_0_3[1]), .A2(port_a_0[1]), .ZN(n93) );
  XNOR2_X1 U277 ( .A(port_rand_mul[2]), .B(n79), .ZN(N35) );
  NAND2_X1 U278 ( .A1(ref_1_port_o_0_3[2]), .A2(port_a_0[2]), .ZN(n79) );
  XNOR2_X1 U279 ( .A(port_rand_mul[2]), .B(n66), .ZN(N51) );
  NAND2_X1 U280 ( .A1(ref_1_port_o_0_3[3]), .A2(port_a_0[3]), .ZN(n66) );
  XNOR2_X1 U281 ( .A(port_rand_mul[2]), .B(n53), .ZN(N67) );
  NAND2_X1 U282 ( .A1(ref_1_port_o_0_3[4]), .A2(port_a_0[4]), .ZN(n53) );
  XNOR2_X1 U283 ( .A(port_rand_mul[4]), .B(n51), .ZN(N7) );
  NAND2_X1 U284 ( .A1(ref_1_port_o_1_3[0]), .A2(port_a_1[0]), .ZN(n51) );
  XNOR2_X1 U285 ( .A(port_rand_mul[4]), .B(n89), .ZN(N23) );
  NAND2_X1 U286 ( .A1(ref_1_port_o_1_3[1]), .A2(port_a_1[1]), .ZN(n89) );
  XNOR2_X1 U287 ( .A(port_rand_mul[4]), .B(n76), .ZN(N39) );
  NAND2_X1 U288 ( .A1(ref_1_port_o_1_3[2]), .A2(port_a_1[2]), .ZN(n76) );
  XNOR2_X1 U289 ( .A(port_rand_mul[4]), .B(n63), .ZN(N55) );
  NAND2_X1 U290 ( .A1(ref_1_port_o_1_3[3]), .A2(port_a_1[3]), .ZN(n63) );
  XNOR2_X1 U291 ( .A(port_rand_mul[4]), .B(n49), .ZN(N71) );
  NAND2_X1 U292 ( .A1(ref_1_port_o_1_3[4]), .A2(port_a_1[4]), .ZN(n49) );
  XNOR2_X1 U293 ( .A(port_rand_mul[5]), .B(n99), .ZN(N11) );
  NAND2_X1 U294 ( .A1(ref_1_port_o_2_3[0]), .A2(port_a_2[0]), .ZN(n99) );
  XNOR2_X1 U295 ( .A(port_rand_mul[5]), .B(n86), .ZN(N27) );
  NAND2_X1 U296 ( .A1(ref_1_port_o_2_3[1]), .A2(port_a_2[1]), .ZN(n86) );
  XNOR2_X1 U297 ( .A(port_rand_mul[5]), .B(n72), .ZN(N43) );
  NAND2_X1 U298 ( .A1(ref_1_port_o_2_3[2]), .A2(port_a_2[2]), .ZN(n72) );
  XNOR2_X1 U299 ( .A(port_rand_mul[5]), .B(n60), .ZN(N59) );
  NAND2_X1 U300 ( .A1(ref_1_port_o_2_3[3]), .A2(port_a_2[3]), .ZN(n60) );
  XNOR2_X1 U301 ( .A(port_rand_mul[5]), .B(n46), .ZN(N75) );
  NAND2_X1 U302 ( .A1(ref_1_port_o_2_3[4]), .A2(port_a_2[4]), .ZN(n46) );
  XNOR2_X1 U303 ( .A(port_rand_mul[1]), .B(n92), .ZN(N2) );
  NAND2_X1 U304 ( .A1(ref_1_port_o_0_2[0]), .A2(port_a_0[0]), .ZN(n92) );
  XNOR2_X1 U305 ( .A(port_rand_mul[1]), .B(n94), .ZN(N18) );
  NAND2_X1 U306 ( .A1(ref_1_port_o_0_2[1]), .A2(port_a_0[1]), .ZN(n94) );
  XNOR2_X1 U307 ( .A(port_rand_mul[1]), .B(n80), .ZN(N34) );
  NAND2_X1 U308 ( .A1(ref_1_port_o_0_2[2]), .A2(port_a_0[2]), .ZN(n80) );
  XNOR2_X1 U309 ( .A(port_rand_mul[1]), .B(n67), .ZN(N50) );
  NAND2_X1 U310 ( .A1(ref_1_port_o_0_2[3]), .A2(port_a_0[3]), .ZN(n67) );
  XNOR2_X1 U311 ( .A(port_rand_mul[1]), .B(n54), .ZN(N66) );
  NAND2_X1 U312 ( .A1(ref_1_port_o_0_2[4]), .A2(port_a_0[4]), .ZN(n54) );
  XNOR2_X1 U313 ( .A(port_rand_mul[0]), .B(n100), .ZN(N1) );
  NAND2_X1 U314 ( .A1(ref_1_port_o_0_1[0]), .A2(port_a_0[0]), .ZN(n100) );
  XNOR2_X1 U315 ( .A(port_rand_mul[0]), .B(n95), .ZN(N17) );
  NAND2_X1 U316 ( .A1(ref_1_port_o_0_1[1]), .A2(port_a_0[1]), .ZN(n95) );
  XNOR2_X1 U317 ( .A(port_rand_mul[0]), .B(n81), .ZN(N33) );
  NAND2_X1 U318 ( .A1(ref_1_port_o_0_1[2]), .A2(port_a_0[2]), .ZN(n81) );
  XNOR2_X1 U319 ( .A(port_rand_mul[0]), .B(n68), .ZN(N49) );
  NAND2_X1 U320 ( .A1(ref_1_port_o_0_1[3]), .A2(port_a_0[3]), .ZN(n68) );
  XNOR2_X1 U321 ( .A(port_rand_mul[0]), .B(n55), .ZN(N65) );
  NAND2_X1 U322 ( .A1(ref_1_port_o_0_1[4]), .A2(port_a_0[4]), .ZN(n55) );
  AND2_X1 U323 ( .A1(ref_1_port_o_2_2[0]), .A2(port_a_2[0]), .ZN(N10) );
  AND2_X1 U324 ( .A1(ref_1_port_o_2_2[1]), .A2(port_a_2[1]), .ZN(N26) );
  AND2_X1 U325 ( .A1(ref_1_port_o_2_2[2]), .A2(port_a_2[2]), .ZN(N42) );
  AND2_X1 U326 ( .A1(ref_1_port_o_2_2[3]), .A2(port_a_2[3]), .ZN(N58) );
  AND2_X1 U327 ( .A1(ref_1_port_o_2_2[4]), .A2(port_a_2[4]), .ZN(N74) );
  AND2_X1 U328 ( .A1(ref_1_port_o_1_1[0]), .A2(port_a_1[0]), .ZN(N5) );
  AND2_X1 U329 ( .A1(ref_1_port_o_1_1[1]), .A2(port_a_1[1]), .ZN(N21) );
  AND2_X1 U330 ( .A1(ref_1_port_o_1_1[2]), .A2(port_a_1[2]), .ZN(N37) );
  AND2_X1 U331 ( .A1(ref_1_port_o_1_1[3]), .A2(port_a_1[3]), .ZN(N53) );
  AND2_X1 U332 ( .A1(ref_1_port_o_1_1[4]), .A2(port_a_1[4]), .ZN(N69) );
  AND2_X1 U333 ( .A1(ref_1_port_o_3_3[0]), .A2(port_a_3[0]), .ZN(N15) );
  AND2_X1 U334 ( .A1(ref_1_port_o_3_3[1]), .A2(port_a_3[1]), .ZN(N31) );
  AND2_X1 U335 ( .A1(ref_1_port_o_3_3[2]), .A2(port_a_3[2]), .ZN(N47) );
  AND2_X1 U336 ( .A1(ref_1_port_o_3_3[3]), .A2(port_a_3[3]), .ZN(N63) );
  AND2_X1 U337 ( .A1(ref_1_port_o_3_3[4]), .A2(port_a_3[4]), .ZN(N79) );
  AND2_X1 U338 ( .A1(ref_1_port_o_0_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U339 ( .A1(ref_1_port_o_0_0[1]), .A2(port_a_0[1]), .ZN(N16) );
  AND2_X1 U340 ( .A1(ref_1_port_o_0_0[2]), .A2(port_a_0[2]), .ZN(N32) );
  AND2_X1 U341 ( .A1(ref_1_port_o_0_0[3]), .A2(port_a_0[3]), .ZN(N48) );
  AND2_X1 U342 ( .A1(ref_1_port_o_0_0[4]), .A2(port_a_0[4]), .ZN(N64) );
  XOR2_X1 U343 ( .A(n9), .B(n10), .Z(port_c_3[0]) );
  XNOR2_X1 U344 ( .A(temp_0_3[0]), .B(mult_ab_3_2[0]), .ZN(n9) );
  XNOR2_X1 U345 ( .A(mult_ab_3_1[0]), .B(mult_ab_3_0[0]), .ZN(n10) );
  XOR2_X1 U346 ( .A(n7), .B(n8), .Z(port_c_3[1]) );
  XNOR2_X1 U347 ( .A(temp_0_3[1]), .B(mult_ab_3_2[1]), .ZN(n7) );
  XNOR2_X1 U348 ( .A(mult_ab_3_1[1]), .B(mult_ab_3_0[1]), .ZN(n8) );
  XOR2_X1 U349 ( .A(n5), .B(n6), .Z(port_c_3[2]) );
  XNOR2_X1 U350 ( .A(temp_0_3[2]), .B(mult_ab_3_2[2]), .ZN(n5) );
  XNOR2_X1 U351 ( .A(mult_ab_3_1[2]), .B(mult_ab_3_0[2]), .ZN(n6) );
  XOR2_X1 U352 ( .A(n3), .B(n4), .Z(port_c_3[3]) );
  XNOR2_X1 U353 ( .A(temp_0_3[3]), .B(mult_ab_3_2[3]), .ZN(n3) );
  XNOR2_X1 U354 ( .A(mult_ab_3_1[3]), .B(mult_ab_3_0[3]), .ZN(n4) );
  XOR2_X1 U355 ( .A(n1), .B(n2), .Z(port_c_3[4]) );
  XNOR2_X1 U356 ( .A(temp_0_3[4]), .B(mult_ab_3_2[4]), .ZN(n1) );
  XNOR2_X1 U357 ( .A(mult_ab_3_1[4]), .B(mult_ab_3_0[4]), .ZN(n2) );
  XOR2_X1 U358 ( .A(n19), .B(n20), .Z(port_c_2[0]) );
  XNOR2_X1 U359 ( .A(temp_0_2[0]), .B(mult_ab_2_3[0]), .ZN(n19) );
  XNOR2_X1 U360 ( .A(mult_ab_2_1[0]), .B(mult_ab_2_0[0]), .ZN(n20) );
  XOR2_X1 U361 ( .A(n17), .B(n18), .Z(port_c_2[1]) );
  XNOR2_X1 U362 ( .A(temp_0_2[1]), .B(mult_ab_2_3[1]), .ZN(n17) );
  XNOR2_X1 U363 ( .A(mult_ab_2_1[1]), .B(mult_ab_2_0[1]), .ZN(n18) );
  XOR2_X1 U364 ( .A(n15), .B(n16), .Z(port_c_2[2]) );
  XNOR2_X1 U365 ( .A(temp_0_2[2]), .B(mult_ab_2_3[2]), .ZN(n15) );
  XNOR2_X1 U366 ( .A(mult_ab_2_1[2]), .B(mult_ab_2_0[2]), .ZN(n16) );
  XOR2_X1 U367 ( .A(n13), .B(n14), .Z(port_c_2[3]) );
  XNOR2_X1 U368 ( .A(temp_0_2[3]), .B(mult_ab_2_3[3]), .ZN(n13) );
  XNOR2_X1 U369 ( .A(mult_ab_2_1[3]), .B(mult_ab_2_0[3]), .ZN(n14) );
  XOR2_X1 U370 ( .A(n11), .B(n12), .Z(port_c_2[4]) );
  XNOR2_X1 U371 ( .A(temp_0_2[4]), .B(mult_ab_2_3[4]), .ZN(n11) );
  XNOR2_X1 U372 ( .A(mult_ab_2_1[4]), .B(mult_ab_2_0[4]), .ZN(n12) );
  XOR2_X1 U373 ( .A(n29), .B(n30), .Z(port_c_1[0]) );
  XNOR2_X1 U374 ( .A(temp_0_1[0]), .B(mult_ab_1_3[0]), .ZN(n29) );
  XNOR2_X1 U375 ( .A(mult_ab_1_2[0]), .B(mult_ab_1_0[0]), .ZN(n30) );
  XOR2_X1 U376 ( .A(n27), .B(n28), .Z(port_c_1[1]) );
  XNOR2_X1 U377 ( .A(temp_0_1[1]), .B(mult_ab_1_3[1]), .ZN(n27) );
  XNOR2_X1 U378 ( .A(mult_ab_1_2[1]), .B(mult_ab_1_0[1]), .ZN(n28) );
  XOR2_X1 U379 ( .A(n25), .B(n26), .Z(port_c_1[2]) );
  XNOR2_X1 U380 ( .A(temp_0_1[2]), .B(mult_ab_1_3[2]), .ZN(n25) );
  XNOR2_X1 U381 ( .A(mult_ab_1_2[2]), .B(mult_ab_1_0[2]), .ZN(n26) );
  XOR2_X1 U382 ( .A(n23), .B(n24), .Z(port_c_1[3]) );
  XNOR2_X1 U383 ( .A(temp_0_1[3]), .B(mult_ab_1_3[3]), .ZN(n23) );
  XNOR2_X1 U384 ( .A(mult_ab_1_2[3]), .B(mult_ab_1_0[3]), .ZN(n24) );
  XOR2_X1 U385 ( .A(n21), .B(n22), .Z(port_c_1[4]) );
  XNOR2_X1 U386 ( .A(temp_0_1[4]), .B(mult_ab_1_3[4]), .ZN(n21) );
  XNOR2_X1 U387 ( .A(mult_ab_1_2[4]), .B(mult_ab_1_0[4]), .ZN(n22) );
  XOR2_X1 U388 ( .A(n39), .B(n40), .Z(port_c_0[0]) );
  XNOR2_X1 U389 ( .A(temp_0_0[0]), .B(mult_ab_0_3[0]), .ZN(n39) );
  XNOR2_X1 U390 ( .A(mult_ab_0_2[0]), .B(mult_ab_0_1[0]), .ZN(n40) );
  XOR2_X1 U391 ( .A(n37), .B(n38), .Z(port_c_0[1]) );
  XNOR2_X1 U392 ( .A(temp_0_0[1]), .B(mult_ab_0_3[1]), .ZN(n37) );
  XNOR2_X1 U393 ( .A(mult_ab_0_2[1]), .B(mult_ab_0_1[1]), .ZN(n38) );
  XOR2_X1 U394 ( .A(n35), .B(n36), .Z(port_c_0[2]) );
  XNOR2_X1 U395 ( .A(temp_0_0[2]), .B(mult_ab_0_3[2]), .ZN(n35) );
  XNOR2_X1 U396 ( .A(mult_ab_0_2[2]), .B(mult_ab_0_1[2]), .ZN(n36) );
  XOR2_X1 U397 ( .A(n33), .B(n34), .Z(port_c_0[3]) );
  XNOR2_X1 U398 ( .A(temp_0_0[3]), .B(mult_ab_0_3[3]), .ZN(n33) );
  XNOR2_X1 U399 ( .A(mult_ab_0_2[3]), .B(mult_ab_0_1[3]), .ZN(n34) );
  XOR2_X1 U400 ( .A(n31), .B(n32), .Z(port_c_0[4]) );
  XNOR2_X1 U401 ( .A(temp_0_0[4]), .B(mult_ab_0_3[4]), .ZN(n31) );
  XNOR2_X1 U402 ( .A(mult_ab_0_2[4]), .B(mult_ab_0_1[4]), .ZN(n32) );
  BUF_X1 ref_1_U42 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n40) );
  BUF_X1 ref_1_U41 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n39) );
  BUF_X1 ref_1_U40 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n38) );
  BUF_X1 ref_1_U39 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n37) );
  BUF_X1 ref_1_U38 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n36) );
  BUF_X1 ref_1_U37 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n35) );
  BUF_X1 ref_1_U36 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n34) );
  BUF_X1 ref_1_U35 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n33) );
  BUF_X1 ref_1_U34 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n32) );
  BUF_X1 ref_1_U33 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n31) );
  BUF_X1 ref_1_U32 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n30) );
  BUF_X1 ref_1_U31 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n29) );
  BUF_X1 ref_1_U30 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n28) );
  BUF_X1 ref_1_U29 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n27) );
  BUF_X1 ref_1_U28 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n26) );
  BUF_X1 ref_1_U27 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n25) );
  BUF_X1 ref_1_U26 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n24) );
  BUF_X1 ref_1_U25 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n23) );
  BUF_X1 ref_1_U24 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n22) );
  BUF_X1 ref_1_U23 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n21) );
  BUF_X1 ref_1_U22 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n20) );
  BUF_X1 ref_1_U21 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n19) );
  BUF_X1 ref_1_U20 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n18) );
  BUF_X1 ref_1_U19 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n17) );
  BUF_X1 ref_1_U18 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n16) );
  BUF_X1 ref_1_U17 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n15) );
  BUF_X1 ref_1_U16 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n14) );
  BUF_X1 ref_1_U15 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n13) );
  BUF_X1 ref_1_U14 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n12) );
  BUF_X1 ref_1_U13 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n11) );
  BUF_X1 ref_1_U12 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n10) );
  BUF_X1 ref_1_U11 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n9) );
  BUF_X1 ref_1_U10 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n8) );
  BUF_X1 ref_1_U9 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n7) );
  BUF_X1 ref_1_U8 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n6) );
  BUF_X1 ref_1_U7 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n5) );
  BUF_X1 ref_1_U6 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n4) );
  BUF_X1 ref_1_U5 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n3) );
  BUF_X1 ref_1_U4 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n2) );
  BUF_X1 ref_1_U3 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n1) );
  DFF_X1 ref_1_reg_out_3_3_reg_0_ ( .D(ref_1_maj_95_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_1_ ( .D(ref_1_maj_111_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_2_ ( .D(ref_1_maj_127_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_3_ ( .D(ref_1_maj_143_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_4_ ( .D(ref_1_maj_159_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_0_ ( .D(ref_1_maj_94_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_1_ ( .D(ref_1_maj_110_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_2_ ( .D(ref_1_maj_126_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_3_ ( .D(ref_1_maj_142_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_4_ ( .D(ref_1_maj_158_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_0_ ( .D(ref_1_maj_93_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_1_ ( .D(ref_1_maj_109_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_2_ ( .D(ref_1_maj_125_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_3_ ( .D(ref_1_maj_141_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_4_ ( .D(ref_1_maj_157_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_0_ ( .D(ref_1_maj_92_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_1_ ( .D(ref_1_maj_108_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_2_ ( .D(ref_1_maj_124_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_3_ ( .D(ref_1_maj_140_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_4_ ( .D(ref_1_maj_156_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_0_ ( .D(ref_1_maj_91_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_1_ ( .D(ref_1_maj_107_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_2_ ( .D(ref_1_maj_123_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_3_ ( .D(ref_1_maj_139_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_4_ ( .D(ref_1_maj_155_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_0_ ( .D(ref_1_maj_90_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_1_ ( .D(ref_1_maj_106_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_2_ ( .D(ref_1_maj_122_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_3_ ( .D(ref_1_maj_138_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_4_ ( .D(ref_1_maj_154_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_0_ ( .D(ref_1_maj_89_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_1_ ( .D(ref_1_maj_105_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_2_ ( .D(ref_1_maj_121_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_3_ ( .D(ref_1_maj_137_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_4_ ( .D(ref_1_maj_153_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_0_ ( .D(ref_1_maj_88_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_1_ ( .D(ref_1_maj_104_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_2_ ( .D(ref_1_maj_120_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_3_ ( .D(ref_1_maj_136_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_4_ ( .D(ref_1_maj_152_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_0_ ( .D(ref_1_maj_87_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_1_ ( .D(ref_1_maj_103_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_2_ ( .D(ref_1_maj_119_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_3_ ( .D(ref_1_maj_135_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_4_ ( .D(ref_1_maj_151_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_0_ ( .D(ref_1_maj_86_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_1_ ( .D(ref_1_maj_102_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_2_ ( .D(ref_1_maj_118_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_3_ ( .D(ref_1_maj_134_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_4_ ( .D(ref_1_maj_150_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_0_ ( .D(ref_1_maj_85_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_1_ ( .D(ref_1_maj_101_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_2_ ( .D(ref_1_maj_117_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_3_ ( .D(ref_1_maj_133_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_4_ ( .D(ref_1_maj_149_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_0_ ( .D(ref_1_maj_84_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_1_ ( .D(ref_1_maj_100_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_2_ ( .D(ref_1_maj_116_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_3_ ( .D(ref_1_maj_132_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_4_ ( .D(ref_1_maj_148_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_0_ ( .D(ref_1_maj_83_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_1_ ( .D(ref_1_maj_99_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_2_ ( .D(ref_1_maj_115_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_3_ ( .D(ref_1_maj_131_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_4_ ( .D(ref_1_maj_147_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_0_ ( .D(ref_1_maj_82_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_1_ ( .D(ref_1_maj_98_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_2_ ( .D(ref_1_maj_114_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_3_ ( .D(ref_1_maj_130_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_4_ ( .D(ref_1_maj_146_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_0_ ( .D(ref_1_maj_81_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_1_ ( .D(ref_1_maj_97_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_2_ ( .D(ref_1_maj_113_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_3_ ( .D(ref_1_maj_129_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_4_ ( .D(ref_1_maj_145_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_0_ ( .D(ref_1_maj_80_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_1_ ( .D(ref_1_maj_96_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_2_ ( .D(ref_1_maj_112_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_3_ ( .D(ref_1_maj_128_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_4_ ( .D(ref_1_maj_144_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[4]), .QN() );
  XOR2_X1 ref_1_simpleXor_60_U1 ( .A(port_rand_ref[0]), .B(port_b_0[0]), .Z(
        ref_1_simpleXor_60_port_z) );
  XOR2_X1 ref_1_simpleXor_61_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_60_port_z), .Z(ref_1_simpleXor_61_port_z) );
  XOR2_X1 ref_1_simpleXor_62_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_61_port_z), .Z(ref_1_refreshed_0_0_) );
  XOR2_X1 ref_1_simpleXor_63_U1 ( .A(port_rand_ref[0]), .B(port_b_1[0]), .Z(
        ref_1_simpleXor_63_port_z) );
  XOR2_X1 ref_1_simpleXor_64_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_63_port_z), .Z(ref_1_simpleXor_64_port_z) );
  XOR2_X1 ref_1_simpleXor_65_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_64_port_z), .Z(ref_1_refreshed_1_0_) );
  XOR2_X1 ref_1_simpleXor_66_U1 ( .A(port_rand_ref[1]), .B(port_b_2[0]), .Z(
        ref_1_simpleXor_66_port_z) );
  XOR2_X1 ref_1_simpleXor_67_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_66_port_z), .Z(ref_1_simpleXor_67_port_z) );
  XOR2_X1 ref_1_simpleXor_68_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_67_port_z), .Z(ref_1_refreshed_2_0_) );
  XOR2_X1 ref_1_simpleXor_69_U1 ( .A(port_rand_ref[2]), .B(port_b_3[0]), .Z(
        ref_1_simpleXor_69_port_z) );
  XOR2_X1 ref_1_simpleXor_70_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_69_port_z), .Z(ref_1_simpleXor_70_port_z) );
  XOR2_X1 ref_1_simpleXor_71_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_70_port_z), .Z(ref_1_refreshed_3_0_) );
  XOR2_X1 ref_1_simpleXor_72_U1 ( .A(port_rand_ref[0]), .B(port_b_0[1]), .Z(
        ref_1_simpleXor_72_port_z) );
  XOR2_X1 ref_1_simpleXor_73_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_72_port_z), .Z(ref_1_simpleXor_73_port_z) );
  XOR2_X1 ref_1_simpleXor_74_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_73_port_z), .Z(ref_1_refreshed_0_1_) );
  XOR2_X1 ref_1_simpleXor_75_U1 ( .A(port_rand_ref[0]), .B(port_b_1[1]), .Z(
        ref_1_simpleXor_75_port_z) );
  XOR2_X1 ref_1_simpleXor_76_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_75_port_z), .Z(ref_1_simpleXor_76_port_z) );
  XOR2_X1 ref_1_simpleXor_77_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_76_port_z), .Z(ref_1_refreshed_1_1_) );
  XOR2_X1 ref_1_simpleXor_78_U1 ( .A(port_rand_ref[1]), .B(port_b_2[1]), .Z(
        ref_1_simpleXor_78_port_z) );
  XOR2_X1 ref_1_simpleXor_79_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_78_port_z), .Z(ref_1_simpleXor_79_port_z) );
  XOR2_X1 ref_1_simpleXor_80_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_79_port_z), .Z(ref_1_refreshed_2_1_) );
  XOR2_X1 ref_1_simpleXor_81_U1 ( .A(port_rand_ref[2]), .B(port_b_3[1]), .Z(
        ref_1_simpleXor_81_port_z) );
  XOR2_X1 ref_1_simpleXor_82_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_81_port_z), .Z(ref_1_simpleXor_82_port_z) );
  XOR2_X1 ref_1_simpleXor_83_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_82_port_z), .Z(ref_1_refreshed_3_1_) );
  XOR2_X1 ref_1_simpleXor_84_U1 ( .A(port_rand_ref[0]), .B(port_b_0[2]), .Z(
        ref_1_simpleXor_84_port_z) );
  XOR2_X1 ref_1_simpleXor_85_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_84_port_z), .Z(ref_1_simpleXor_85_port_z) );
  XOR2_X1 ref_1_simpleXor_86_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_85_port_z), .Z(ref_1_refreshed_0_2_) );
  XOR2_X1 ref_1_simpleXor_87_U1 ( .A(port_rand_ref[0]), .B(port_b_1[2]), .Z(
        ref_1_simpleXor_87_port_z) );
  XOR2_X1 ref_1_simpleXor_88_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_87_port_z), .Z(ref_1_simpleXor_88_port_z) );
  XOR2_X1 ref_1_simpleXor_89_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_88_port_z), .Z(ref_1_refreshed_1_2_) );
  XOR2_X1 ref_1_simpleXor_90_U1 ( .A(port_rand_ref[1]), .B(port_b_2[2]), .Z(
        ref_1_simpleXor_90_port_z) );
  XOR2_X1 ref_1_simpleXor_91_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_90_port_z), .Z(ref_1_simpleXor_91_port_z) );
  XOR2_X1 ref_1_simpleXor_92_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_91_port_z), .Z(ref_1_refreshed_2_2_) );
  XOR2_X1 ref_1_simpleXor_93_U1 ( .A(port_rand_ref[2]), .B(port_b_3[2]), .Z(
        ref_1_simpleXor_93_port_z) );
  XOR2_X1 ref_1_simpleXor_94_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_93_port_z), .Z(ref_1_simpleXor_94_port_z) );
  XOR2_X1 ref_1_simpleXor_95_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_94_port_z), .Z(ref_1_refreshed_3_2_) );
  XOR2_X1 ref_1_simpleXor_96_U1 ( .A(port_rand_ref[0]), .B(port_b_0[3]), .Z(
        ref_1_simpleXor_96_port_z) );
  XOR2_X1 ref_1_simpleXor_97_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_96_port_z), .Z(ref_1_simpleXor_97_port_z) );
  XOR2_X1 ref_1_simpleXor_98_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_97_port_z), .Z(ref_1_refreshed_0_3_) );
  XOR2_X1 ref_1_simpleXor_99_U1 ( .A(port_rand_ref[0]), .B(port_b_1[3]), .Z(
        ref_1_simpleXor_99_port_z) );
  XOR2_X1 ref_1_simpleXor_100_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_99_port_z), .Z(ref_1_simpleXor_100_port_z) );
  XOR2_X1 ref_1_simpleXor_101_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_100_port_z), .Z(ref_1_refreshed_1_3_) );
  XOR2_X1 ref_1_simpleXor_102_U1 ( .A(port_rand_ref[1]), .B(port_b_2[3]), .Z(
        ref_1_simpleXor_102_port_z) );
  XOR2_X1 ref_1_simpleXor_103_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_102_port_z), .Z(ref_1_simpleXor_103_port_z) );
  XOR2_X1 ref_1_simpleXor_104_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_103_port_z), .Z(ref_1_refreshed_2_3_) );
  XOR2_X1 ref_1_simpleXor_105_U1 ( .A(port_rand_ref[2]), .B(port_b_3[3]), .Z(
        ref_1_simpleXor_105_port_z) );
  XOR2_X1 ref_1_simpleXor_106_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_105_port_z), .Z(ref_1_simpleXor_106_port_z) );
  XOR2_X1 ref_1_simpleXor_107_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_106_port_z), .Z(ref_1_refreshed_3_3_) );
  XOR2_X1 ref_1_simpleXor_108_U1 ( .A(port_rand_ref[0]), .B(port_b_0[4]), .Z(
        ref_1_simpleXor_108_port_z) );
  XOR2_X1 ref_1_simpleXor_109_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_108_port_z), .Z(ref_1_simpleXor_109_port_z) );
  XOR2_X1 ref_1_simpleXor_110_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_109_port_z), .Z(ref_1_refreshed_0_4_) );
  XOR2_X1 ref_1_simpleXor_111_U1 ( .A(port_rand_ref[0]), .B(port_b_1[4]), .Z(
        ref_1_simpleXor_111_port_z) );
  XOR2_X1 ref_1_simpleXor_112_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_111_port_z), .Z(ref_1_simpleXor_112_port_z) );
  XOR2_X1 ref_1_simpleXor_113_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_112_port_z), .Z(ref_1_refreshed_1_4_) );
  XOR2_X1 ref_1_simpleXor_114_U1 ( .A(port_rand_ref[1]), .B(port_b_2[4]), .Z(
        ref_1_simpleXor_114_port_z) );
  XOR2_X1 ref_1_simpleXor_115_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_114_port_z), .Z(ref_1_simpleXor_115_port_z) );
  XOR2_X1 ref_1_simpleXor_116_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_115_port_z), .Z(ref_1_refreshed_2_4_) );
  XOR2_X1 ref_1_simpleXor_117_U1 ( .A(port_rand_ref[2]), .B(port_b_3[4]), .Z(
        ref_1_simpleXor_117_port_z) );
  XOR2_X1 ref_1_simpleXor_118_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_117_port_z), .Z(ref_1_simpleXor_118_port_z) );
  XOR2_X1 ref_1_simpleXor_119_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_118_port_z), .Z(ref_1_refreshed_3_4_) );
  NAND2_X1 ref_1_maj_80_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_80_n9) );
  NAND2_X1 ref_1_maj_80_U14 ( .A1(ref_1_maj_80_n6), .A2(ref_1_maj_80_n5), .ZN(
        ref_1_maj_80_n10) );
  NAND2_X1 ref_1_maj_80_U13 ( .A1(ref_1_maj_80_n9), .A2(ref_1_maj_80_n10), 
        .ZN(ref_1_maj_80_n8) );
  NAND2_X1 ref_1_maj_80_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_80_n11), .ZN(
        ref_1_maj_80_n13) );
  NAND2_X1 ref_1_maj_80_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_80_n12) );
  NAND2_X1 ref_1_maj_80_U10 ( .A1(ref_1_maj_80_n12), .A2(ref_1_maj_80_n13), 
        .ZN(ref_1_maj_80_n7) );
  XOR2_X1 ref_1_maj_80_U9 ( .A(ref_1_n36), .B(ref_1_maj_80_n11), .Z(
        ref_1_maj_80_n6) );
  XOR2_X1 ref_1_maj_80_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_80_n5)
         );
  XOR2_X1 ref_1_maj_80_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_80_n11)
         );
  OR2_X1 ref_1_maj_80_U6 ( .A1(ref_1_maj_80_n7), .A2(ref_1_maj_80_n8), .ZN(
        ref_1_maj_80_n3) );
  NAND2_X1 ref_1_maj_80_U5 ( .A1(ref_1_maj_80_n3), .A2(ref_1_maj_80_n4), .ZN(
        ref_1_maj_80_n2) );
  NAND2_X1 ref_1_maj_80_U4 ( .A1(ref_1_maj_80_n7), .A2(ref_1_maj_80_n8), .ZN(
        ref_1_maj_80_n1) );
  NAND2_X1 ref_1_maj_80_U3 ( .A1(ref_1_maj_80_n1), .A2(ref_1_maj_80_n2), .ZN(
        ref_1_maj_80_port_o) );
  XOR2_X1 ref_1_maj_80_U2 ( .A(ref_1_maj_80_n5), .B(ref_1_maj_80_n6), .Z(
        ref_1_maj_80_n4) );
  NAND2_X1 ref_1_maj_81_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_81_n18) );
  NAND2_X1 ref_1_maj_81_U14 ( .A1(ref_1_maj_81_n21), .A2(ref_1_maj_81_n22), 
        .ZN(ref_1_maj_81_n17) );
  NAND2_X1 ref_1_maj_81_U13 ( .A1(ref_1_maj_81_n18), .A2(ref_1_maj_81_n17), 
        .ZN(ref_1_maj_81_n19) );
  NAND2_X1 ref_1_maj_81_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_81_n16), .ZN(
        ref_1_maj_81_n14) );
  NAND2_X1 ref_1_maj_81_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_81_n15) );
  NAND2_X1 ref_1_maj_81_U10 ( .A1(ref_1_maj_81_n15), .A2(ref_1_maj_81_n14), 
        .ZN(ref_1_maj_81_n20) );
  XOR2_X1 ref_1_maj_81_U9 ( .A(ref_1_n36), .B(ref_1_maj_81_n16), .Z(
        ref_1_maj_81_n21) );
  XOR2_X1 ref_1_maj_81_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_81_n22)
         );
  XOR2_X1 ref_1_maj_81_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_81_n16)
         );
  OR2_X1 ref_1_maj_81_U6 ( .A1(ref_1_maj_81_n20), .A2(ref_1_maj_81_n19), .ZN(
        ref_1_maj_81_n24) );
  NAND2_X1 ref_1_maj_81_U5 ( .A1(ref_1_maj_81_n24), .A2(ref_1_maj_81_n23), 
        .ZN(ref_1_maj_81_n25) );
  NAND2_X1 ref_1_maj_81_U4 ( .A1(ref_1_maj_81_n20), .A2(ref_1_maj_81_n19), 
        .ZN(ref_1_maj_81_n26) );
  NAND2_X1 ref_1_maj_81_U3 ( .A1(ref_1_maj_81_n26), .A2(ref_1_maj_81_n25), 
        .ZN(ref_1_maj_81_port_o) );
  XOR2_X1 ref_1_maj_81_U2 ( .A(ref_1_maj_81_n22), .B(ref_1_maj_81_n21), .Z(
        ref_1_maj_81_n23) );
  NAND2_X1 ref_1_maj_82_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_82_n18) );
  NAND2_X1 ref_1_maj_82_U14 ( .A1(ref_1_maj_82_n21), .A2(ref_1_maj_82_n22), 
        .ZN(ref_1_maj_82_n17) );
  NAND2_X1 ref_1_maj_82_U13 ( .A1(ref_1_maj_82_n18), .A2(ref_1_maj_82_n17), 
        .ZN(ref_1_maj_82_n19) );
  NAND2_X1 ref_1_maj_82_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_82_n16), 
        .ZN(ref_1_maj_82_n14) );
  NAND2_X1 ref_1_maj_82_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_82_n15) );
  NAND2_X1 ref_1_maj_82_U10 ( .A1(ref_1_maj_82_n15), .A2(ref_1_maj_82_n14), 
        .ZN(ref_1_maj_82_n20) );
  XOR2_X1 ref_1_maj_82_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_82_n16), 
        .Z(ref_1_maj_82_n21) );
  XOR2_X1 ref_1_maj_82_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_82_n22) );
  XOR2_X1 ref_1_maj_82_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), 
        .Z(ref_1_maj_82_n16) );
  OR2_X1 ref_1_maj_82_U6 ( .A1(ref_1_maj_82_n20), .A2(ref_1_maj_82_n19), .ZN(
        ref_1_maj_82_n24) );
  NAND2_X1 ref_1_maj_82_U5 ( .A1(ref_1_maj_82_n24), .A2(ref_1_maj_82_n23), 
        .ZN(ref_1_maj_82_n25) );
  NAND2_X1 ref_1_maj_82_U4 ( .A1(ref_1_maj_82_n20), .A2(ref_1_maj_82_n19), 
        .ZN(ref_1_maj_82_n26) );
  NAND2_X1 ref_1_maj_82_U3 ( .A1(ref_1_maj_82_n26), .A2(ref_1_maj_82_n25), 
        .ZN(ref_1_maj_82_port_o) );
  XOR2_X1 ref_1_maj_82_U2 ( .A(ref_1_maj_82_n22), .B(ref_1_maj_82_n21), .Z(
        ref_1_maj_82_n23) );
  NAND2_X1 ref_1_maj_83_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_83_n18) );
  NAND2_X1 ref_1_maj_83_U14 ( .A1(ref_1_maj_83_n21), .A2(ref_1_maj_83_n22), 
        .ZN(ref_1_maj_83_n17) );
  NAND2_X1 ref_1_maj_83_U13 ( .A1(ref_1_maj_83_n18), .A2(ref_1_maj_83_n17), 
        .ZN(ref_1_maj_83_n19) );
  NAND2_X1 ref_1_maj_83_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_83_n16), 
        .ZN(ref_1_maj_83_n14) );
  NAND2_X1 ref_1_maj_83_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_83_n15) );
  NAND2_X1 ref_1_maj_83_U10 ( .A1(ref_1_maj_83_n15), .A2(ref_1_maj_83_n14), 
        .ZN(ref_1_maj_83_n20) );
  XOR2_X1 ref_1_maj_83_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_83_n16), 
        .Z(ref_1_maj_83_n21) );
  XOR2_X1 ref_1_maj_83_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_83_n22) );
  XOR2_X1 ref_1_maj_83_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), 
        .Z(ref_1_maj_83_n16) );
  OR2_X1 ref_1_maj_83_U6 ( .A1(ref_1_maj_83_n20), .A2(ref_1_maj_83_n19), .ZN(
        ref_1_maj_83_n24) );
  NAND2_X1 ref_1_maj_83_U5 ( .A1(ref_1_maj_83_n24), .A2(ref_1_maj_83_n23), 
        .ZN(ref_1_maj_83_n25) );
  NAND2_X1 ref_1_maj_83_U4 ( .A1(ref_1_maj_83_n20), .A2(ref_1_maj_83_n19), 
        .ZN(ref_1_maj_83_n26) );
  NAND2_X1 ref_1_maj_83_U3 ( .A1(ref_1_maj_83_n26), .A2(ref_1_maj_83_n25), 
        .ZN(ref_1_maj_83_port_o) );
  XOR2_X1 ref_1_maj_83_U2 ( .A(ref_1_maj_83_n22), .B(ref_1_maj_83_n21), .Z(
        ref_1_maj_83_n23) );
  NAND2_X1 ref_1_maj_84_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_84_n18) );
  NAND2_X1 ref_1_maj_84_U14 ( .A1(ref_1_maj_84_n21), .A2(ref_1_maj_84_n22), 
        .ZN(ref_1_maj_84_n17) );
  NAND2_X1 ref_1_maj_84_U13 ( .A1(ref_1_maj_84_n18), .A2(ref_1_maj_84_n17), 
        .ZN(ref_1_maj_84_n19) );
  NAND2_X1 ref_1_maj_84_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_84_n16), .ZN(
        ref_1_maj_84_n14) );
  NAND2_X1 ref_1_maj_84_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_84_n15) );
  NAND2_X1 ref_1_maj_84_U10 ( .A1(ref_1_maj_84_n15), .A2(ref_1_maj_84_n14), 
        .ZN(ref_1_maj_84_n20) );
  XOR2_X1 ref_1_maj_84_U9 ( .A(ref_1_n26), .B(ref_1_maj_84_n16), .Z(
        ref_1_maj_84_n21) );
  XOR2_X1 ref_1_maj_84_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_84_n22)
         );
  XOR2_X1 ref_1_maj_84_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(ref_1_maj_84_n16)
         );
  OR2_X1 ref_1_maj_84_U6 ( .A1(ref_1_maj_84_n20), .A2(ref_1_maj_84_n19), .ZN(
        ref_1_maj_84_n24) );
  NAND2_X1 ref_1_maj_84_U5 ( .A1(ref_1_maj_84_n24), .A2(ref_1_maj_84_n23), 
        .ZN(ref_1_maj_84_n25) );
  NAND2_X1 ref_1_maj_84_U4 ( .A1(ref_1_maj_84_n20), .A2(ref_1_maj_84_n19), 
        .ZN(ref_1_maj_84_n26) );
  NAND2_X1 ref_1_maj_84_U3 ( .A1(ref_1_maj_84_n26), .A2(ref_1_maj_84_n25), 
        .ZN(ref_1_maj_84_port_o) );
  XOR2_X1 ref_1_maj_84_U2 ( .A(ref_1_maj_84_n22), .B(ref_1_maj_84_n21), .Z(
        ref_1_maj_84_n23) );
  NAND2_X1 ref_1_maj_85_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_85_n18) );
  NAND2_X1 ref_1_maj_85_U14 ( .A1(ref_1_maj_85_n21), .A2(ref_1_maj_85_n22), 
        .ZN(ref_1_maj_85_n17) );
  NAND2_X1 ref_1_maj_85_U13 ( .A1(ref_1_maj_85_n18), .A2(ref_1_maj_85_n17), 
        .ZN(ref_1_maj_85_n19) );
  NAND2_X1 ref_1_maj_85_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_85_n16), 
        .ZN(ref_1_maj_85_n14) );
  NAND2_X1 ref_1_maj_85_U11 ( .A1(ref_1_refreshed_1_0_), .A2(
        ref_1_refreshed_1_1_), .ZN(ref_1_maj_85_n15) );
  NAND2_X1 ref_1_maj_85_U10 ( .A1(ref_1_maj_85_n15), .A2(ref_1_maj_85_n14), 
        .ZN(ref_1_maj_85_n20) );
  XOR2_X1 ref_1_maj_85_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_85_n16), 
        .Z(ref_1_maj_85_n21) );
  XOR2_X1 ref_1_maj_85_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_85_n22) );
  XOR2_X1 ref_1_maj_85_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_refreshed_1_1_), 
        .Z(ref_1_maj_85_n16) );
  OR2_X1 ref_1_maj_85_U6 ( .A1(ref_1_maj_85_n20), .A2(ref_1_maj_85_n19), .ZN(
        ref_1_maj_85_n24) );
  NAND2_X1 ref_1_maj_85_U5 ( .A1(ref_1_maj_85_n24), .A2(ref_1_maj_85_n23), 
        .ZN(ref_1_maj_85_n25) );
  NAND2_X1 ref_1_maj_85_U4 ( .A1(ref_1_maj_85_n20), .A2(ref_1_maj_85_n19), 
        .ZN(ref_1_maj_85_n26) );
  NAND2_X1 ref_1_maj_85_U3 ( .A1(ref_1_maj_85_n26), .A2(ref_1_maj_85_n25), 
        .ZN(ref_1_maj_85_port_o) );
  XOR2_X1 ref_1_maj_85_U2 ( .A(ref_1_maj_85_n22), .B(ref_1_maj_85_n21), .Z(
        ref_1_maj_85_n23) );
  NAND2_X1 ref_1_maj_86_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_86_n18) );
  NAND2_X1 ref_1_maj_86_U14 ( .A1(ref_1_maj_86_n21), .A2(ref_1_maj_86_n22), 
        .ZN(ref_1_maj_86_n17) );
  NAND2_X1 ref_1_maj_86_U13 ( .A1(ref_1_maj_86_n18), .A2(ref_1_maj_86_n17), 
        .ZN(ref_1_maj_86_n19) );
  NAND2_X1 ref_1_maj_86_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_86_n16), 
        .ZN(ref_1_maj_86_n14) );
  NAND2_X1 ref_1_maj_86_U11 ( .A1(ref_1_refreshed_1_0_), .A2(
        ref_1_refreshed_1_1_), .ZN(ref_1_maj_86_n15) );
  NAND2_X1 ref_1_maj_86_U10 ( .A1(ref_1_maj_86_n15), .A2(ref_1_maj_86_n14), 
        .ZN(ref_1_maj_86_n20) );
  XOR2_X1 ref_1_maj_86_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_86_n16), 
        .Z(ref_1_maj_86_n21) );
  XOR2_X1 ref_1_maj_86_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_86_n22) );
  XOR2_X1 ref_1_maj_86_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_refreshed_1_1_), 
        .Z(ref_1_maj_86_n16) );
  OR2_X1 ref_1_maj_86_U6 ( .A1(ref_1_maj_86_n20), .A2(ref_1_maj_86_n19), .ZN(
        ref_1_maj_86_n24) );
  NAND2_X1 ref_1_maj_86_U5 ( .A1(ref_1_maj_86_n24), .A2(ref_1_maj_86_n23), 
        .ZN(ref_1_maj_86_n25) );
  NAND2_X1 ref_1_maj_86_U4 ( .A1(ref_1_maj_86_n20), .A2(ref_1_maj_86_n19), 
        .ZN(ref_1_maj_86_n26) );
  NAND2_X1 ref_1_maj_86_U3 ( .A1(ref_1_maj_86_n26), .A2(ref_1_maj_86_n25), 
        .ZN(ref_1_maj_86_port_o) );
  XOR2_X1 ref_1_maj_86_U2 ( .A(ref_1_maj_86_n22), .B(ref_1_maj_86_n21), .Z(
        ref_1_maj_86_n23) );
  NAND2_X1 ref_1_maj_87_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_87_n18) );
  NAND2_X1 ref_1_maj_87_U14 ( .A1(ref_1_maj_87_n21), .A2(ref_1_maj_87_n22), 
        .ZN(ref_1_maj_87_n17) );
  NAND2_X1 ref_1_maj_87_U13 ( .A1(ref_1_maj_87_n18), .A2(ref_1_maj_87_n17), 
        .ZN(ref_1_maj_87_n19) );
  NAND2_X1 ref_1_maj_87_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_87_n16), 
        .ZN(ref_1_maj_87_n14) );
  NAND2_X1 ref_1_maj_87_U11 ( .A1(ref_1_refreshed_1_0_), .A2(
        ref_1_refreshed_1_1_), .ZN(ref_1_maj_87_n15) );
  NAND2_X1 ref_1_maj_87_U10 ( .A1(ref_1_maj_87_n15), .A2(ref_1_maj_87_n14), 
        .ZN(ref_1_maj_87_n20) );
  XOR2_X1 ref_1_maj_87_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_87_n16), 
        .Z(ref_1_maj_87_n21) );
  XOR2_X1 ref_1_maj_87_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_87_n22) );
  XOR2_X1 ref_1_maj_87_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_refreshed_1_1_), 
        .Z(ref_1_maj_87_n16) );
  OR2_X1 ref_1_maj_87_U6 ( .A1(ref_1_maj_87_n20), .A2(ref_1_maj_87_n19), .ZN(
        ref_1_maj_87_n24) );
  NAND2_X1 ref_1_maj_87_U5 ( .A1(ref_1_maj_87_n24), .A2(ref_1_maj_87_n23), 
        .ZN(ref_1_maj_87_n25) );
  NAND2_X1 ref_1_maj_87_U4 ( .A1(ref_1_maj_87_n20), .A2(ref_1_maj_87_n19), 
        .ZN(ref_1_maj_87_n26) );
  NAND2_X1 ref_1_maj_87_U3 ( .A1(ref_1_maj_87_n26), .A2(ref_1_maj_87_n25), 
        .ZN(ref_1_maj_87_port_o) );
  XOR2_X1 ref_1_maj_87_U2 ( .A(ref_1_maj_87_n22), .B(ref_1_maj_87_n21), .Z(
        ref_1_maj_87_n23) );
  NAND2_X1 ref_1_maj_88_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_88_n18) );
  NAND2_X1 ref_1_maj_88_U14 ( .A1(ref_1_maj_88_n21), .A2(ref_1_maj_88_n22), 
        .ZN(ref_1_maj_88_n17) );
  NAND2_X1 ref_1_maj_88_U13 ( .A1(ref_1_maj_88_n18), .A2(ref_1_maj_88_n17), 
        .ZN(ref_1_maj_88_n19) );
  NAND2_X1 ref_1_maj_88_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_88_n16), .ZN(
        ref_1_maj_88_n14) );
  NAND2_X1 ref_1_maj_88_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_88_n15) );
  NAND2_X1 ref_1_maj_88_U10 ( .A1(ref_1_maj_88_n15), .A2(ref_1_maj_88_n14), 
        .ZN(ref_1_maj_88_n20) );
  XOR2_X1 ref_1_maj_88_U9 ( .A(ref_1_n16), .B(ref_1_maj_88_n16), .Z(
        ref_1_maj_88_n21) );
  XOR2_X1 ref_1_maj_88_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_88_n22)
         );
  XOR2_X1 ref_1_maj_88_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(ref_1_maj_88_n16)
         );
  OR2_X1 ref_1_maj_88_U6 ( .A1(ref_1_maj_88_n20), .A2(ref_1_maj_88_n19), .ZN(
        ref_1_maj_88_n24) );
  NAND2_X1 ref_1_maj_88_U5 ( .A1(ref_1_maj_88_n24), .A2(ref_1_maj_88_n23), 
        .ZN(ref_1_maj_88_n25) );
  NAND2_X1 ref_1_maj_88_U4 ( .A1(ref_1_maj_88_n20), .A2(ref_1_maj_88_n19), 
        .ZN(ref_1_maj_88_n26) );
  NAND2_X1 ref_1_maj_88_U3 ( .A1(ref_1_maj_88_n26), .A2(ref_1_maj_88_n25), 
        .ZN(ref_1_maj_88_port_o) );
  XOR2_X1 ref_1_maj_88_U2 ( .A(ref_1_maj_88_n22), .B(ref_1_maj_88_n21), .Z(
        ref_1_maj_88_n23) );
  NAND2_X1 ref_1_maj_89_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_89_n18) );
  NAND2_X1 ref_1_maj_89_U14 ( .A1(ref_1_maj_89_n21), .A2(ref_1_maj_89_n22), 
        .ZN(ref_1_maj_89_n17) );
  NAND2_X1 ref_1_maj_89_U13 ( .A1(ref_1_maj_89_n18), .A2(ref_1_maj_89_n17), 
        .ZN(ref_1_maj_89_n19) );
  NAND2_X1 ref_1_maj_89_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_89_n16), 
        .ZN(ref_1_maj_89_n14) );
  NAND2_X1 ref_1_maj_89_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_89_n15) );
  NAND2_X1 ref_1_maj_89_U10 ( .A1(ref_1_maj_89_n15), .A2(ref_1_maj_89_n14), 
        .ZN(ref_1_maj_89_n20) );
  XOR2_X1 ref_1_maj_89_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_89_n16), 
        .Z(ref_1_maj_89_n21) );
  XOR2_X1 ref_1_maj_89_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_89_n22) );
  XOR2_X1 ref_1_maj_89_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), 
        .Z(ref_1_maj_89_n16) );
  OR2_X1 ref_1_maj_89_U6 ( .A1(ref_1_maj_89_n20), .A2(ref_1_maj_89_n19), .ZN(
        ref_1_maj_89_n24) );
  NAND2_X1 ref_1_maj_89_U5 ( .A1(ref_1_maj_89_n24), .A2(ref_1_maj_89_n23), 
        .ZN(ref_1_maj_89_n25) );
  NAND2_X1 ref_1_maj_89_U4 ( .A1(ref_1_maj_89_n20), .A2(ref_1_maj_89_n19), 
        .ZN(ref_1_maj_89_n26) );
  NAND2_X1 ref_1_maj_89_U3 ( .A1(ref_1_maj_89_n26), .A2(ref_1_maj_89_n25), 
        .ZN(ref_1_maj_89_port_o) );
  XOR2_X1 ref_1_maj_89_U2 ( .A(ref_1_maj_89_n22), .B(ref_1_maj_89_n21), .Z(
        ref_1_maj_89_n23) );
  NAND2_X1 ref_1_maj_90_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_90_n18) );
  NAND2_X1 ref_1_maj_90_U14 ( .A1(ref_1_maj_90_n21), .A2(ref_1_maj_90_n22), 
        .ZN(ref_1_maj_90_n17) );
  NAND2_X1 ref_1_maj_90_U13 ( .A1(ref_1_maj_90_n18), .A2(ref_1_maj_90_n17), 
        .ZN(ref_1_maj_90_n19) );
  NAND2_X1 ref_1_maj_90_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_90_n16), 
        .ZN(ref_1_maj_90_n14) );
  NAND2_X1 ref_1_maj_90_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_90_n15) );
  NAND2_X1 ref_1_maj_90_U10 ( .A1(ref_1_maj_90_n15), .A2(ref_1_maj_90_n14), 
        .ZN(ref_1_maj_90_n20) );
  XOR2_X1 ref_1_maj_90_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_90_n16), 
        .Z(ref_1_maj_90_n21) );
  XOR2_X1 ref_1_maj_90_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_90_n22) );
  XOR2_X1 ref_1_maj_90_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), 
        .Z(ref_1_maj_90_n16) );
  OR2_X1 ref_1_maj_90_U6 ( .A1(ref_1_maj_90_n20), .A2(ref_1_maj_90_n19), .ZN(
        ref_1_maj_90_n24) );
  NAND2_X1 ref_1_maj_90_U5 ( .A1(ref_1_maj_90_n24), .A2(ref_1_maj_90_n23), 
        .ZN(ref_1_maj_90_n25) );
  NAND2_X1 ref_1_maj_90_U4 ( .A1(ref_1_maj_90_n20), .A2(ref_1_maj_90_n19), 
        .ZN(ref_1_maj_90_n26) );
  NAND2_X1 ref_1_maj_90_U3 ( .A1(ref_1_maj_90_n26), .A2(ref_1_maj_90_n25), 
        .ZN(ref_1_maj_90_port_o) );
  XOR2_X1 ref_1_maj_90_U2 ( .A(ref_1_maj_90_n22), .B(ref_1_maj_90_n21), .Z(
        ref_1_maj_90_n23) );
  NAND2_X1 ref_1_maj_91_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_91_n18) );
  NAND2_X1 ref_1_maj_91_U14 ( .A1(ref_1_maj_91_n21), .A2(ref_1_maj_91_n22), 
        .ZN(ref_1_maj_91_n17) );
  NAND2_X1 ref_1_maj_91_U13 ( .A1(ref_1_maj_91_n18), .A2(ref_1_maj_91_n17), 
        .ZN(ref_1_maj_91_n19) );
  NAND2_X1 ref_1_maj_91_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_91_n16), 
        .ZN(ref_1_maj_91_n14) );
  NAND2_X1 ref_1_maj_91_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_91_n15) );
  NAND2_X1 ref_1_maj_91_U10 ( .A1(ref_1_maj_91_n15), .A2(ref_1_maj_91_n14), 
        .ZN(ref_1_maj_91_n20) );
  XOR2_X1 ref_1_maj_91_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_91_n16), 
        .Z(ref_1_maj_91_n21) );
  XOR2_X1 ref_1_maj_91_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_91_n22) );
  XOR2_X1 ref_1_maj_91_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), 
        .Z(ref_1_maj_91_n16) );
  OR2_X1 ref_1_maj_91_U6 ( .A1(ref_1_maj_91_n20), .A2(ref_1_maj_91_n19), .ZN(
        ref_1_maj_91_n24) );
  NAND2_X1 ref_1_maj_91_U5 ( .A1(ref_1_maj_91_n24), .A2(ref_1_maj_91_n23), 
        .ZN(ref_1_maj_91_n25) );
  NAND2_X1 ref_1_maj_91_U4 ( .A1(ref_1_maj_91_n20), .A2(ref_1_maj_91_n19), 
        .ZN(ref_1_maj_91_n26) );
  NAND2_X1 ref_1_maj_91_U3 ( .A1(ref_1_maj_91_n26), .A2(ref_1_maj_91_n25), 
        .ZN(ref_1_maj_91_port_o) );
  XOR2_X1 ref_1_maj_91_U2 ( .A(ref_1_maj_91_n22), .B(ref_1_maj_91_n21), .Z(
        ref_1_maj_91_n23) );
  NAND2_X1 ref_1_maj_92_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_92_n18) );
  NAND2_X1 ref_1_maj_92_U14 ( .A1(ref_1_maj_92_n21), .A2(ref_1_maj_92_n22), 
        .ZN(ref_1_maj_92_n17) );
  NAND2_X1 ref_1_maj_92_U13 ( .A1(ref_1_maj_92_n18), .A2(ref_1_maj_92_n17), 
        .ZN(ref_1_maj_92_n19) );
  NAND2_X1 ref_1_maj_92_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_92_n16), .ZN(
        ref_1_maj_92_n14) );
  NAND2_X1 ref_1_maj_92_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_92_n15) );
  NAND2_X1 ref_1_maj_92_U10 ( .A1(ref_1_maj_92_n15), .A2(ref_1_maj_92_n14), 
        .ZN(ref_1_maj_92_n20) );
  XOR2_X1 ref_1_maj_92_U9 ( .A(ref_1_n6), .B(ref_1_maj_92_n16), .Z(
        ref_1_maj_92_n21) );
  XOR2_X1 ref_1_maj_92_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_92_n22)
         );
  XOR2_X1 ref_1_maj_92_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_92_n16)
         );
  OR2_X1 ref_1_maj_92_U6 ( .A1(ref_1_maj_92_n20), .A2(ref_1_maj_92_n19), .ZN(
        ref_1_maj_92_n24) );
  NAND2_X1 ref_1_maj_92_U5 ( .A1(ref_1_maj_92_n24), .A2(ref_1_maj_92_n23), 
        .ZN(ref_1_maj_92_n25) );
  NAND2_X1 ref_1_maj_92_U4 ( .A1(ref_1_maj_92_n20), .A2(ref_1_maj_92_n19), 
        .ZN(ref_1_maj_92_n26) );
  NAND2_X1 ref_1_maj_92_U3 ( .A1(ref_1_maj_92_n26), .A2(ref_1_maj_92_n25), 
        .ZN(ref_1_maj_92_port_o) );
  XOR2_X1 ref_1_maj_92_U2 ( .A(ref_1_maj_92_n22), .B(ref_1_maj_92_n21), .Z(
        ref_1_maj_92_n23) );
  NAND2_X1 ref_1_maj_93_U15 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_93_n18) );
  NAND2_X1 ref_1_maj_93_U14 ( .A1(ref_1_maj_93_n21), .A2(ref_1_maj_93_n22), 
        .ZN(ref_1_maj_93_n17) );
  NAND2_X1 ref_1_maj_93_U13 ( .A1(ref_1_maj_93_n18), .A2(ref_1_maj_93_n17), 
        .ZN(ref_1_maj_93_n19) );
  NAND2_X1 ref_1_maj_93_U12 ( .A1(ref_1_refreshed_3_2_), .A2(ref_1_maj_93_n16), 
        .ZN(ref_1_maj_93_n14) );
  NAND2_X1 ref_1_maj_93_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_93_n15) );
  NAND2_X1 ref_1_maj_93_U10 ( .A1(ref_1_maj_93_n15), .A2(ref_1_maj_93_n14), 
        .ZN(ref_1_maj_93_n20) );
  XOR2_X1 ref_1_maj_93_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_93_n16), 
        .Z(ref_1_maj_93_n21) );
  XOR2_X1 ref_1_maj_93_U8 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), 
        .Z(ref_1_maj_93_n22) );
  XOR2_X1 ref_1_maj_93_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), 
        .Z(ref_1_maj_93_n16) );
  OR2_X1 ref_1_maj_93_U6 ( .A1(ref_1_maj_93_n20), .A2(ref_1_maj_93_n19), .ZN(
        ref_1_maj_93_n24) );
  NAND2_X1 ref_1_maj_93_U5 ( .A1(ref_1_maj_93_n24), .A2(ref_1_maj_93_n23), 
        .ZN(ref_1_maj_93_n25) );
  NAND2_X1 ref_1_maj_93_U4 ( .A1(ref_1_maj_93_n20), .A2(ref_1_maj_93_n19), 
        .ZN(ref_1_maj_93_n26) );
  NAND2_X1 ref_1_maj_93_U3 ( .A1(ref_1_maj_93_n26), .A2(ref_1_maj_93_n25), 
        .ZN(ref_1_maj_93_port_o) );
  XOR2_X1 ref_1_maj_93_U2 ( .A(ref_1_maj_93_n22), .B(ref_1_maj_93_n21), .Z(
        ref_1_maj_93_n23) );
  NAND2_X1 ref_1_maj_94_U15 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_94_n18) );
  NAND2_X1 ref_1_maj_94_U14 ( .A1(ref_1_maj_94_n21), .A2(ref_1_maj_94_n22), 
        .ZN(ref_1_maj_94_n17) );
  NAND2_X1 ref_1_maj_94_U13 ( .A1(ref_1_maj_94_n18), .A2(ref_1_maj_94_n17), 
        .ZN(ref_1_maj_94_n19) );
  NAND2_X1 ref_1_maj_94_U12 ( .A1(ref_1_refreshed_3_2_), .A2(ref_1_maj_94_n16), 
        .ZN(ref_1_maj_94_n14) );
  NAND2_X1 ref_1_maj_94_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_94_n15) );
  NAND2_X1 ref_1_maj_94_U10 ( .A1(ref_1_maj_94_n15), .A2(ref_1_maj_94_n14), 
        .ZN(ref_1_maj_94_n20) );
  XOR2_X1 ref_1_maj_94_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_94_n16), 
        .Z(ref_1_maj_94_n21) );
  XOR2_X1 ref_1_maj_94_U8 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), 
        .Z(ref_1_maj_94_n22) );
  XOR2_X1 ref_1_maj_94_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), 
        .Z(ref_1_maj_94_n16) );
  OR2_X1 ref_1_maj_94_U6 ( .A1(ref_1_maj_94_n20), .A2(ref_1_maj_94_n19), .ZN(
        ref_1_maj_94_n24) );
  NAND2_X1 ref_1_maj_94_U5 ( .A1(ref_1_maj_94_n24), .A2(ref_1_maj_94_n23), 
        .ZN(ref_1_maj_94_n25) );
  NAND2_X1 ref_1_maj_94_U4 ( .A1(ref_1_maj_94_n20), .A2(ref_1_maj_94_n19), 
        .ZN(ref_1_maj_94_n26) );
  NAND2_X1 ref_1_maj_94_U3 ( .A1(ref_1_maj_94_n26), .A2(ref_1_maj_94_n25), 
        .ZN(ref_1_maj_94_port_o) );
  XOR2_X1 ref_1_maj_94_U2 ( .A(ref_1_maj_94_n22), .B(ref_1_maj_94_n21), .Z(
        ref_1_maj_94_n23) );
  NAND2_X1 ref_1_maj_95_U15 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_95_n18) );
  NAND2_X1 ref_1_maj_95_U14 ( .A1(ref_1_maj_95_n21), .A2(ref_1_maj_95_n22), 
        .ZN(ref_1_maj_95_n17) );
  NAND2_X1 ref_1_maj_95_U13 ( .A1(ref_1_maj_95_n18), .A2(ref_1_maj_95_n17), 
        .ZN(ref_1_maj_95_n19) );
  NAND2_X1 ref_1_maj_95_U12 ( .A1(ref_1_refreshed_3_2_), .A2(ref_1_maj_95_n16), 
        .ZN(ref_1_maj_95_n14) );
  NAND2_X1 ref_1_maj_95_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_95_n15) );
  NAND2_X1 ref_1_maj_95_U10 ( .A1(ref_1_maj_95_n15), .A2(ref_1_maj_95_n14), 
        .ZN(ref_1_maj_95_n20) );
  XOR2_X1 ref_1_maj_95_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_95_n16), 
        .Z(ref_1_maj_95_n21) );
  XOR2_X1 ref_1_maj_95_U8 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), 
        .Z(ref_1_maj_95_n22) );
  XOR2_X1 ref_1_maj_95_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), 
        .Z(ref_1_maj_95_n16) );
  OR2_X1 ref_1_maj_95_U6 ( .A1(ref_1_maj_95_n20), .A2(ref_1_maj_95_n19), .ZN(
        ref_1_maj_95_n24) );
  NAND2_X1 ref_1_maj_95_U5 ( .A1(ref_1_maj_95_n24), .A2(ref_1_maj_95_n23), 
        .ZN(ref_1_maj_95_n25) );
  NAND2_X1 ref_1_maj_95_U4 ( .A1(ref_1_maj_95_n20), .A2(ref_1_maj_95_n19), 
        .ZN(ref_1_maj_95_n26) );
  NAND2_X1 ref_1_maj_95_U3 ( .A1(ref_1_maj_95_n26), .A2(ref_1_maj_95_n25), 
        .ZN(ref_1_maj_95_port_o) );
  XOR2_X1 ref_1_maj_95_U2 ( .A(ref_1_maj_95_n22), .B(ref_1_maj_95_n21), .Z(
        ref_1_maj_95_n23) );
  NAND2_X1 ref_1_maj_96_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_96_n18) );
  NAND2_X1 ref_1_maj_96_U14 ( .A1(ref_1_maj_96_n21), .A2(ref_1_maj_96_n22), 
        .ZN(ref_1_maj_96_n17) );
  NAND2_X1 ref_1_maj_96_U13 ( .A1(ref_1_maj_96_n18), .A2(ref_1_maj_96_n17), 
        .ZN(ref_1_maj_96_n19) );
  NAND2_X1 ref_1_maj_96_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_96_n16), 
        .ZN(ref_1_maj_96_n14) );
  NAND2_X1 ref_1_maj_96_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_96_n15) );
  NAND2_X1 ref_1_maj_96_U10 ( .A1(ref_1_maj_96_n15), .A2(ref_1_maj_96_n14), 
        .ZN(ref_1_maj_96_n20) );
  XOR2_X1 ref_1_maj_96_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_96_n16), 
        .Z(ref_1_maj_96_n21) );
  XOR2_X1 ref_1_maj_96_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_96_n22) );
  XOR2_X1 ref_1_maj_96_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), 
        .Z(ref_1_maj_96_n16) );
  OR2_X1 ref_1_maj_96_U6 ( .A1(ref_1_maj_96_n20), .A2(ref_1_maj_96_n19), .ZN(
        ref_1_maj_96_n24) );
  NAND2_X1 ref_1_maj_96_U5 ( .A1(ref_1_maj_96_n24), .A2(ref_1_maj_96_n23), 
        .ZN(ref_1_maj_96_n25) );
  NAND2_X1 ref_1_maj_96_U4 ( .A1(ref_1_maj_96_n20), .A2(ref_1_maj_96_n19), 
        .ZN(ref_1_maj_96_n26) );
  NAND2_X1 ref_1_maj_96_U3 ( .A1(ref_1_maj_96_n26), .A2(ref_1_maj_96_n25), 
        .ZN(ref_1_maj_96_port_o) );
  XOR2_X1 ref_1_maj_96_U2 ( .A(ref_1_maj_96_n22), .B(ref_1_maj_96_n21), .Z(
        ref_1_maj_96_n23) );
  NAND2_X1 ref_1_maj_97_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_97_n18) );
  NAND2_X1 ref_1_maj_97_U14 ( .A1(ref_1_maj_97_n21), .A2(ref_1_maj_97_n22), 
        .ZN(ref_1_maj_97_n17) );
  NAND2_X1 ref_1_maj_97_U13 ( .A1(ref_1_maj_97_n18), .A2(ref_1_maj_97_n17), 
        .ZN(ref_1_maj_97_n19) );
  NAND2_X1 ref_1_maj_97_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_97_n16), .ZN(
        ref_1_maj_97_n14) );
  NAND2_X1 ref_1_maj_97_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_97_n15) );
  NAND2_X1 ref_1_maj_97_U10 ( .A1(ref_1_maj_97_n15), .A2(ref_1_maj_97_n14), 
        .ZN(ref_1_maj_97_n20) );
  XOR2_X1 ref_1_maj_97_U9 ( .A(ref_1_n35), .B(ref_1_maj_97_n16), .Z(
        ref_1_maj_97_n21) );
  XOR2_X1 ref_1_maj_97_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(ref_1_maj_97_n22)
         );
  XOR2_X1 ref_1_maj_97_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(ref_1_maj_97_n16)
         );
  OR2_X1 ref_1_maj_97_U6 ( .A1(ref_1_maj_97_n20), .A2(ref_1_maj_97_n19), .ZN(
        ref_1_maj_97_n24) );
  NAND2_X1 ref_1_maj_97_U5 ( .A1(ref_1_maj_97_n24), .A2(ref_1_maj_97_n23), 
        .ZN(ref_1_maj_97_n25) );
  NAND2_X1 ref_1_maj_97_U4 ( .A1(ref_1_maj_97_n20), .A2(ref_1_maj_97_n19), 
        .ZN(ref_1_maj_97_n26) );
  NAND2_X1 ref_1_maj_97_U3 ( .A1(ref_1_maj_97_n26), .A2(ref_1_maj_97_n25), 
        .ZN(ref_1_maj_97_port_o) );
  XOR2_X1 ref_1_maj_97_U2 ( .A(ref_1_maj_97_n22), .B(ref_1_maj_97_n21), .Z(
        ref_1_maj_97_n23) );
  NAND2_X1 ref_1_maj_98_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_98_n18) );
  NAND2_X1 ref_1_maj_98_U14 ( .A1(ref_1_maj_98_n21), .A2(ref_1_maj_98_n22), 
        .ZN(ref_1_maj_98_n17) );
  NAND2_X1 ref_1_maj_98_U13 ( .A1(ref_1_maj_98_n18), .A2(ref_1_maj_98_n17), 
        .ZN(ref_1_maj_98_n19) );
  NAND2_X1 ref_1_maj_98_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_98_n16), .ZN(
        ref_1_maj_98_n14) );
  NAND2_X1 ref_1_maj_98_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_98_n15) );
  NAND2_X1 ref_1_maj_98_U10 ( .A1(ref_1_maj_98_n15), .A2(ref_1_maj_98_n14), 
        .ZN(ref_1_maj_98_n20) );
  XOR2_X1 ref_1_maj_98_U9 ( .A(ref_1_n36), .B(ref_1_maj_98_n16), .Z(
        ref_1_maj_98_n21) );
  XOR2_X1 ref_1_maj_98_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_98_n22)
         );
  XOR2_X1 ref_1_maj_98_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_98_n16)
         );
  OR2_X1 ref_1_maj_98_U6 ( .A1(ref_1_maj_98_n20), .A2(ref_1_maj_98_n19), .ZN(
        ref_1_maj_98_n24) );
  NAND2_X1 ref_1_maj_98_U5 ( .A1(ref_1_maj_98_n24), .A2(ref_1_maj_98_n23), 
        .ZN(ref_1_maj_98_n25) );
  NAND2_X1 ref_1_maj_98_U4 ( .A1(ref_1_maj_98_n20), .A2(ref_1_maj_98_n19), 
        .ZN(ref_1_maj_98_n26) );
  NAND2_X1 ref_1_maj_98_U3 ( .A1(ref_1_maj_98_n26), .A2(ref_1_maj_98_n25), 
        .ZN(ref_1_maj_98_port_o) );
  XOR2_X1 ref_1_maj_98_U2 ( .A(ref_1_maj_98_n22), .B(ref_1_maj_98_n21), .Z(
        ref_1_maj_98_n23) );
  NAND2_X1 ref_1_maj_99_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_99_n18) );
  NAND2_X1 ref_1_maj_99_U14 ( .A1(ref_1_maj_99_n21), .A2(ref_1_maj_99_n22), 
        .ZN(ref_1_maj_99_n17) );
  NAND2_X1 ref_1_maj_99_U13 ( .A1(ref_1_maj_99_n18), .A2(ref_1_maj_99_n17), 
        .ZN(ref_1_maj_99_n19) );
  NAND2_X1 ref_1_maj_99_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_99_n16), .ZN(
        ref_1_maj_99_n14) );
  NAND2_X1 ref_1_maj_99_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_99_n15) );
  NAND2_X1 ref_1_maj_99_U10 ( .A1(ref_1_maj_99_n15), .A2(ref_1_maj_99_n14), 
        .ZN(ref_1_maj_99_n20) );
  XOR2_X1 ref_1_maj_99_U9 ( .A(ref_1_n36), .B(ref_1_maj_99_n16), .Z(
        ref_1_maj_99_n21) );
  XOR2_X1 ref_1_maj_99_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_99_n22)
         );
  XOR2_X1 ref_1_maj_99_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_99_n16)
         );
  OR2_X1 ref_1_maj_99_U6 ( .A1(ref_1_maj_99_n20), .A2(ref_1_maj_99_n19), .ZN(
        ref_1_maj_99_n24) );
  NAND2_X1 ref_1_maj_99_U5 ( .A1(ref_1_maj_99_n24), .A2(ref_1_maj_99_n23), 
        .ZN(ref_1_maj_99_n25) );
  NAND2_X1 ref_1_maj_99_U4 ( .A1(ref_1_maj_99_n20), .A2(ref_1_maj_99_n19), 
        .ZN(ref_1_maj_99_n26) );
  NAND2_X1 ref_1_maj_99_U3 ( .A1(ref_1_maj_99_n26), .A2(ref_1_maj_99_n25), 
        .ZN(ref_1_maj_99_port_o) );
  XOR2_X1 ref_1_maj_99_U2 ( .A(ref_1_maj_99_n22), .B(ref_1_maj_99_n21), .Z(
        ref_1_maj_99_n23) );
  NAND2_X1 ref_1_maj_100_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_100_n18) );
  NAND2_X1 ref_1_maj_100_U14 ( .A1(ref_1_maj_100_n21), .A2(ref_1_maj_100_n22), 
        .ZN(ref_1_maj_100_n17) );
  NAND2_X1 ref_1_maj_100_U13 ( .A1(ref_1_maj_100_n18), .A2(ref_1_maj_100_n17), 
        .ZN(ref_1_maj_100_n19) );
  NAND2_X1 ref_1_maj_100_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_100_n16), .ZN(
        ref_1_maj_100_n14) );
  NAND2_X1 ref_1_maj_100_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_100_n15) );
  NAND2_X1 ref_1_maj_100_U10 ( .A1(ref_1_maj_100_n15), .A2(ref_1_maj_100_n14), 
        .ZN(ref_1_maj_100_n20) );
  XOR2_X1 ref_1_maj_100_U9 ( .A(ref_1_n25), .B(ref_1_maj_100_n16), .Z(
        ref_1_maj_100_n21) );
  XOR2_X1 ref_1_maj_100_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_100_n22) );
  XOR2_X1 ref_1_maj_100_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_100_n16) );
  OR2_X1 ref_1_maj_100_U6 ( .A1(ref_1_maj_100_n20), .A2(ref_1_maj_100_n19), 
        .ZN(ref_1_maj_100_n24) );
  NAND2_X1 ref_1_maj_100_U5 ( .A1(ref_1_maj_100_n24), .A2(ref_1_maj_100_n23), 
        .ZN(ref_1_maj_100_n25) );
  NAND2_X1 ref_1_maj_100_U4 ( .A1(ref_1_maj_100_n20), .A2(ref_1_maj_100_n19), 
        .ZN(ref_1_maj_100_n26) );
  NAND2_X1 ref_1_maj_100_U3 ( .A1(ref_1_maj_100_n26), .A2(ref_1_maj_100_n25), 
        .ZN(ref_1_maj_100_port_o) );
  XOR2_X1 ref_1_maj_100_U2 ( .A(ref_1_maj_100_n22), .B(ref_1_maj_100_n21), .Z(
        ref_1_maj_100_n23) );
  NAND2_X1 ref_1_maj_101_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_101_n18) );
  NAND2_X1 ref_1_maj_101_U14 ( .A1(ref_1_maj_101_n21), .A2(ref_1_maj_101_n22), 
        .ZN(ref_1_maj_101_n17) );
  NAND2_X1 ref_1_maj_101_U13 ( .A1(ref_1_maj_101_n18), .A2(ref_1_maj_101_n17), 
        .ZN(ref_1_maj_101_n19) );
  NAND2_X1 ref_1_maj_101_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_101_n16), .ZN(
        ref_1_maj_101_n14) );
  NAND2_X1 ref_1_maj_101_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_101_n15) );
  NAND2_X1 ref_1_maj_101_U10 ( .A1(ref_1_maj_101_n15), .A2(ref_1_maj_101_n14), 
        .ZN(ref_1_maj_101_n20) );
  XOR2_X1 ref_1_maj_101_U9 ( .A(ref_1_n26), .B(ref_1_maj_101_n16), .Z(
        ref_1_maj_101_n21) );
  XOR2_X1 ref_1_maj_101_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_101_n22) );
  XOR2_X1 ref_1_maj_101_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_101_n16) );
  OR2_X1 ref_1_maj_101_U6 ( .A1(ref_1_maj_101_n20), .A2(ref_1_maj_101_n19), 
        .ZN(ref_1_maj_101_n24) );
  NAND2_X1 ref_1_maj_101_U5 ( .A1(ref_1_maj_101_n24), .A2(ref_1_maj_101_n23), 
        .ZN(ref_1_maj_101_n25) );
  NAND2_X1 ref_1_maj_101_U4 ( .A1(ref_1_maj_101_n20), .A2(ref_1_maj_101_n19), 
        .ZN(ref_1_maj_101_n26) );
  NAND2_X1 ref_1_maj_101_U3 ( .A1(ref_1_maj_101_n26), .A2(ref_1_maj_101_n25), 
        .ZN(ref_1_maj_101_port_o) );
  XOR2_X1 ref_1_maj_101_U2 ( .A(ref_1_maj_101_n22), .B(ref_1_maj_101_n21), .Z(
        ref_1_maj_101_n23) );
  NAND2_X1 ref_1_maj_102_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_102_n18) );
  NAND2_X1 ref_1_maj_102_U14 ( .A1(ref_1_maj_102_n21), .A2(ref_1_maj_102_n22), 
        .ZN(ref_1_maj_102_n17) );
  NAND2_X1 ref_1_maj_102_U13 ( .A1(ref_1_maj_102_n18), .A2(ref_1_maj_102_n17), 
        .ZN(ref_1_maj_102_n19) );
  NAND2_X1 ref_1_maj_102_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_102_n16), .ZN(
        ref_1_maj_102_n14) );
  NAND2_X1 ref_1_maj_102_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_102_n15) );
  NAND2_X1 ref_1_maj_102_U10 ( .A1(ref_1_maj_102_n15), .A2(ref_1_maj_102_n14), 
        .ZN(ref_1_maj_102_n20) );
  XOR2_X1 ref_1_maj_102_U9 ( .A(ref_1_n26), .B(ref_1_maj_102_n16), .Z(
        ref_1_maj_102_n21) );
  XOR2_X1 ref_1_maj_102_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_102_n22) );
  XOR2_X1 ref_1_maj_102_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_102_n16) );
  OR2_X1 ref_1_maj_102_U6 ( .A1(ref_1_maj_102_n20), .A2(ref_1_maj_102_n19), 
        .ZN(ref_1_maj_102_n24) );
  NAND2_X1 ref_1_maj_102_U5 ( .A1(ref_1_maj_102_n24), .A2(ref_1_maj_102_n23), 
        .ZN(ref_1_maj_102_n25) );
  NAND2_X1 ref_1_maj_102_U4 ( .A1(ref_1_maj_102_n20), .A2(ref_1_maj_102_n19), 
        .ZN(ref_1_maj_102_n26) );
  NAND2_X1 ref_1_maj_102_U3 ( .A1(ref_1_maj_102_n26), .A2(ref_1_maj_102_n25), 
        .ZN(ref_1_maj_102_port_o) );
  XOR2_X1 ref_1_maj_102_U2 ( .A(ref_1_maj_102_n22), .B(ref_1_maj_102_n21), .Z(
        ref_1_maj_102_n23) );
  NAND2_X1 ref_1_maj_103_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_103_n18) );
  NAND2_X1 ref_1_maj_103_U14 ( .A1(ref_1_maj_103_n21), .A2(ref_1_maj_103_n22), 
        .ZN(ref_1_maj_103_n17) );
  NAND2_X1 ref_1_maj_103_U13 ( .A1(ref_1_maj_103_n18), .A2(ref_1_maj_103_n17), 
        .ZN(ref_1_maj_103_n19) );
  NAND2_X1 ref_1_maj_103_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_103_n16), .ZN(
        ref_1_maj_103_n14) );
  NAND2_X1 ref_1_maj_103_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_103_n15) );
  NAND2_X1 ref_1_maj_103_U10 ( .A1(ref_1_maj_103_n15), .A2(ref_1_maj_103_n14), 
        .ZN(ref_1_maj_103_n20) );
  XOR2_X1 ref_1_maj_103_U9 ( .A(ref_1_n25), .B(ref_1_maj_103_n16), .Z(
        ref_1_maj_103_n21) );
  XOR2_X1 ref_1_maj_103_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_103_n22) );
  XOR2_X1 ref_1_maj_103_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_103_n16) );
  OR2_X1 ref_1_maj_103_U6 ( .A1(ref_1_maj_103_n20), .A2(ref_1_maj_103_n19), 
        .ZN(ref_1_maj_103_n24) );
  NAND2_X1 ref_1_maj_103_U5 ( .A1(ref_1_maj_103_n24), .A2(ref_1_maj_103_n23), 
        .ZN(ref_1_maj_103_n25) );
  NAND2_X1 ref_1_maj_103_U4 ( .A1(ref_1_maj_103_n20), .A2(ref_1_maj_103_n19), 
        .ZN(ref_1_maj_103_n26) );
  NAND2_X1 ref_1_maj_103_U3 ( .A1(ref_1_maj_103_n26), .A2(ref_1_maj_103_n25), 
        .ZN(ref_1_maj_103_port_o) );
  XOR2_X1 ref_1_maj_103_U2 ( .A(ref_1_maj_103_n22), .B(ref_1_maj_103_n21), .Z(
        ref_1_maj_103_n23) );
  NAND2_X1 ref_1_maj_104_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_104_n18) );
  NAND2_X1 ref_1_maj_104_U14 ( .A1(ref_1_maj_104_n21), .A2(ref_1_maj_104_n22), 
        .ZN(ref_1_maj_104_n17) );
  NAND2_X1 ref_1_maj_104_U13 ( .A1(ref_1_maj_104_n18), .A2(ref_1_maj_104_n17), 
        .ZN(ref_1_maj_104_n19) );
  NAND2_X1 ref_1_maj_104_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_104_n16), .ZN(
        ref_1_maj_104_n14) );
  NAND2_X1 ref_1_maj_104_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_104_n15) );
  NAND2_X1 ref_1_maj_104_U10 ( .A1(ref_1_maj_104_n15), .A2(ref_1_maj_104_n14), 
        .ZN(ref_1_maj_104_n20) );
  XOR2_X1 ref_1_maj_104_U9 ( .A(ref_1_n15), .B(ref_1_maj_104_n16), .Z(
        ref_1_maj_104_n21) );
  XOR2_X1 ref_1_maj_104_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_104_n22) );
  XOR2_X1 ref_1_maj_104_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_104_n16) );
  OR2_X1 ref_1_maj_104_U6 ( .A1(ref_1_maj_104_n20), .A2(ref_1_maj_104_n19), 
        .ZN(ref_1_maj_104_n24) );
  NAND2_X1 ref_1_maj_104_U5 ( .A1(ref_1_maj_104_n24), .A2(ref_1_maj_104_n23), 
        .ZN(ref_1_maj_104_n25) );
  NAND2_X1 ref_1_maj_104_U4 ( .A1(ref_1_maj_104_n20), .A2(ref_1_maj_104_n19), 
        .ZN(ref_1_maj_104_n26) );
  NAND2_X1 ref_1_maj_104_U3 ( .A1(ref_1_maj_104_n26), .A2(ref_1_maj_104_n25), 
        .ZN(ref_1_maj_104_port_o) );
  XOR2_X1 ref_1_maj_104_U2 ( .A(ref_1_maj_104_n22), .B(ref_1_maj_104_n21), .Z(
        ref_1_maj_104_n23) );
  NAND2_X1 ref_1_maj_105_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_105_n18) );
  NAND2_X1 ref_1_maj_105_U14 ( .A1(ref_1_maj_105_n21), .A2(ref_1_maj_105_n22), 
        .ZN(ref_1_maj_105_n17) );
  NAND2_X1 ref_1_maj_105_U13 ( .A1(ref_1_maj_105_n18), .A2(ref_1_maj_105_n17), 
        .ZN(ref_1_maj_105_n19) );
  NAND2_X1 ref_1_maj_105_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_105_n16), .ZN(
        ref_1_maj_105_n14) );
  NAND2_X1 ref_1_maj_105_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_105_n15) );
  NAND2_X1 ref_1_maj_105_U10 ( .A1(ref_1_maj_105_n15), .A2(ref_1_maj_105_n14), 
        .ZN(ref_1_maj_105_n20) );
  XOR2_X1 ref_1_maj_105_U9 ( .A(ref_1_n16), .B(ref_1_maj_105_n16), .Z(
        ref_1_maj_105_n21) );
  XOR2_X1 ref_1_maj_105_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_105_n22) );
  XOR2_X1 ref_1_maj_105_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_105_n16) );
  OR2_X1 ref_1_maj_105_U6 ( .A1(ref_1_maj_105_n20), .A2(ref_1_maj_105_n19), 
        .ZN(ref_1_maj_105_n24) );
  NAND2_X1 ref_1_maj_105_U5 ( .A1(ref_1_maj_105_n24), .A2(ref_1_maj_105_n23), 
        .ZN(ref_1_maj_105_n25) );
  NAND2_X1 ref_1_maj_105_U4 ( .A1(ref_1_maj_105_n20), .A2(ref_1_maj_105_n19), 
        .ZN(ref_1_maj_105_n26) );
  NAND2_X1 ref_1_maj_105_U3 ( .A1(ref_1_maj_105_n26), .A2(ref_1_maj_105_n25), 
        .ZN(ref_1_maj_105_port_o) );
  XOR2_X1 ref_1_maj_105_U2 ( .A(ref_1_maj_105_n22), .B(ref_1_maj_105_n21), .Z(
        ref_1_maj_105_n23) );
  NAND2_X1 ref_1_maj_106_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_106_n18) );
  NAND2_X1 ref_1_maj_106_U14 ( .A1(ref_1_maj_106_n21), .A2(ref_1_maj_106_n22), 
        .ZN(ref_1_maj_106_n17) );
  NAND2_X1 ref_1_maj_106_U13 ( .A1(ref_1_maj_106_n18), .A2(ref_1_maj_106_n17), 
        .ZN(ref_1_maj_106_n19) );
  NAND2_X1 ref_1_maj_106_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_106_n16), .ZN(
        ref_1_maj_106_n14) );
  NAND2_X1 ref_1_maj_106_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_106_n15) );
  NAND2_X1 ref_1_maj_106_U10 ( .A1(ref_1_maj_106_n15), .A2(ref_1_maj_106_n14), 
        .ZN(ref_1_maj_106_n20) );
  XOR2_X1 ref_1_maj_106_U9 ( .A(ref_1_n16), .B(ref_1_maj_106_n16), .Z(
        ref_1_maj_106_n21) );
  XOR2_X1 ref_1_maj_106_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_106_n22) );
  XOR2_X1 ref_1_maj_106_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_106_n16) );
  OR2_X1 ref_1_maj_106_U6 ( .A1(ref_1_maj_106_n20), .A2(ref_1_maj_106_n19), 
        .ZN(ref_1_maj_106_n24) );
  NAND2_X1 ref_1_maj_106_U5 ( .A1(ref_1_maj_106_n24), .A2(ref_1_maj_106_n23), 
        .ZN(ref_1_maj_106_n25) );
  NAND2_X1 ref_1_maj_106_U4 ( .A1(ref_1_maj_106_n20), .A2(ref_1_maj_106_n19), 
        .ZN(ref_1_maj_106_n26) );
  NAND2_X1 ref_1_maj_106_U3 ( .A1(ref_1_maj_106_n26), .A2(ref_1_maj_106_n25), 
        .ZN(ref_1_maj_106_port_o) );
  XOR2_X1 ref_1_maj_106_U2 ( .A(ref_1_maj_106_n22), .B(ref_1_maj_106_n21), .Z(
        ref_1_maj_106_n23) );
  NAND2_X1 ref_1_maj_107_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_107_n18) );
  NAND2_X1 ref_1_maj_107_U14 ( .A1(ref_1_maj_107_n21), .A2(ref_1_maj_107_n22), 
        .ZN(ref_1_maj_107_n17) );
  NAND2_X1 ref_1_maj_107_U13 ( .A1(ref_1_maj_107_n18), .A2(ref_1_maj_107_n17), 
        .ZN(ref_1_maj_107_n19) );
  NAND2_X1 ref_1_maj_107_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_107_n16), .ZN(
        ref_1_maj_107_n14) );
  NAND2_X1 ref_1_maj_107_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_107_n15) );
  NAND2_X1 ref_1_maj_107_U10 ( .A1(ref_1_maj_107_n15), .A2(ref_1_maj_107_n14), 
        .ZN(ref_1_maj_107_n20) );
  XOR2_X1 ref_1_maj_107_U9 ( .A(ref_1_n15), .B(ref_1_maj_107_n16), .Z(
        ref_1_maj_107_n21) );
  XOR2_X1 ref_1_maj_107_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_107_n22) );
  XOR2_X1 ref_1_maj_107_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_107_n16) );
  OR2_X1 ref_1_maj_107_U6 ( .A1(ref_1_maj_107_n20), .A2(ref_1_maj_107_n19), 
        .ZN(ref_1_maj_107_n24) );
  NAND2_X1 ref_1_maj_107_U5 ( .A1(ref_1_maj_107_n24), .A2(ref_1_maj_107_n23), 
        .ZN(ref_1_maj_107_n25) );
  NAND2_X1 ref_1_maj_107_U4 ( .A1(ref_1_maj_107_n20), .A2(ref_1_maj_107_n19), 
        .ZN(ref_1_maj_107_n26) );
  NAND2_X1 ref_1_maj_107_U3 ( .A1(ref_1_maj_107_n26), .A2(ref_1_maj_107_n25), 
        .ZN(ref_1_maj_107_port_o) );
  XOR2_X1 ref_1_maj_107_U2 ( .A(ref_1_maj_107_n22), .B(ref_1_maj_107_n21), .Z(
        ref_1_maj_107_n23) );
  NAND2_X1 ref_1_maj_108_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_108_n18) );
  NAND2_X1 ref_1_maj_108_U14 ( .A1(ref_1_maj_108_n21), .A2(ref_1_maj_108_n22), 
        .ZN(ref_1_maj_108_n17) );
  NAND2_X1 ref_1_maj_108_U13 ( .A1(ref_1_maj_108_n18), .A2(ref_1_maj_108_n17), 
        .ZN(ref_1_maj_108_n19) );
  NAND2_X1 ref_1_maj_108_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_108_n16), .ZN(
        ref_1_maj_108_n14) );
  NAND2_X1 ref_1_maj_108_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_108_n15) );
  NAND2_X1 ref_1_maj_108_U10 ( .A1(ref_1_maj_108_n15), .A2(ref_1_maj_108_n14), 
        .ZN(ref_1_maj_108_n20) );
  XOR2_X1 ref_1_maj_108_U9 ( .A(ref_1_n5), .B(ref_1_maj_108_n16), .Z(
        ref_1_maj_108_n21) );
  XOR2_X1 ref_1_maj_108_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_108_n22)
         );
  XOR2_X1 ref_1_maj_108_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_108_n16)
         );
  OR2_X1 ref_1_maj_108_U6 ( .A1(ref_1_maj_108_n20), .A2(ref_1_maj_108_n19), 
        .ZN(ref_1_maj_108_n24) );
  NAND2_X1 ref_1_maj_108_U5 ( .A1(ref_1_maj_108_n24), .A2(ref_1_maj_108_n23), 
        .ZN(ref_1_maj_108_n25) );
  NAND2_X1 ref_1_maj_108_U4 ( .A1(ref_1_maj_108_n20), .A2(ref_1_maj_108_n19), 
        .ZN(ref_1_maj_108_n26) );
  NAND2_X1 ref_1_maj_108_U3 ( .A1(ref_1_maj_108_n26), .A2(ref_1_maj_108_n25), 
        .ZN(ref_1_maj_108_port_o) );
  XOR2_X1 ref_1_maj_108_U2 ( .A(ref_1_maj_108_n22), .B(ref_1_maj_108_n21), .Z(
        ref_1_maj_108_n23) );
  NAND2_X1 ref_1_maj_109_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_109_n18) );
  NAND2_X1 ref_1_maj_109_U14 ( .A1(ref_1_maj_109_n21), .A2(ref_1_maj_109_n22), 
        .ZN(ref_1_maj_109_n17) );
  NAND2_X1 ref_1_maj_109_U13 ( .A1(ref_1_maj_109_n18), .A2(ref_1_maj_109_n17), 
        .ZN(ref_1_maj_109_n19) );
  NAND2_X1 ref_1_maj_109_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_109_n16), .ZN(
        ref_1_maj_109_n14) );
  NAND2_X1 ref_1_maj_109_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_109_n15) );
  NAND2_X1 ref_1_maj_109_U10 ( .A1(ref_1_maj_109_n15), .A2(ref_1_maj_109_n14), 
        .ZN(ref_1_maj_109_n20) );
  XOR2_X1 ref_1_maj_109_U9 ( .A(ref_1_n6), .B(ref_1_maj_109_n16), .Z(
        ref_1_maj_109_n21) );
  XOR2_X1 ref_1_maj_109_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_109_n22) );
  XOR2_X1 ref_1_maj_109_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_109_n16)
         );
  OR2_X1 ref_1_maj_109_U6 ( .A1(ref_1_maj_109_n20), .A2(ref_1_maj_109_n19), 
        .ZN(ref_1_maj_109_n24) );
  NAND2_X1 ref_1_maj_109_U5 ( .A1(ref_1_maj_109_n24), .A2(ref_1_maj_109_n23), 
        .ZN(ref_1_maj_109_n25) );
  NAND2_X1 ref_1_maj_109_U4 ( .A1(ref_1_maj_109_n20), .A2(ref_1_maj_109_n19), 
        .ZN(ref_1_maj_109_n26) );
  NAND2_X1 ref_1_maj_109_U3 ( .A1(ref_1_maj_109_n26), .A2(ref_1_maj_109_n25), 
        .ZN(ref_1_maj_109_port_o) );
  XOR2_X1 ref_1_maj_109_U2 ( .A(ref_1_maj_109_n22), .B(ref_1_maj_109_n21), .Z(
        ref_1_maj_109_n23) );
  NAND2_X1 ref_1_maj_110_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_110_n18) );
  NAND2_X1 ref_1_maj_110_U14 ( .A1(ref_1_maj_110_n21), .A2(ref_1_maj_110_n22), 
        .ZN(ref_1_maj_110_n17) );
  NAND2_X1 ref_1_maj_110_U13 ( .A1(ref_1_maj_110_n18), .A2(ref_1_maj_110_n17), 
        .ZN(ref_1_maj_110_n19) );
  NAND2_X1 ref_1_maj_110_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_110_n16), .ZN(
        ref_1_maj_110_n14) );
  NAND2_X1 ref_1_maj_110_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_110_n15) );
  NAND2_X1 ref_1_maj_110_U10 ( .A1(ref_1_maj_110_n15), .A2(ref_1_maj_110_n14), 
        .ZN(ref_1_maj_110_n20) );
  XOR2_X1 ref_1_maj_110_U9 ( .A(ref_1_n6), .B(ref_1_maj_110_n16), .Z(
        ref_1_maj_110_n21) );
  XOR2_X1 ref_1_maj_110_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_110_n22) );
  XOR2_X1 ref_1_maj_110_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_110_n16)
         );
  OR2_X1 ref_1_maj_110_U6 ( .A1(ref_1_maj_110_n20), .A2(ref_1_maj_110_n19), 
        .ZN(ref_1_maj_110_n24) );
  NAND2_X1 ref_1_maj_110_U5 ( .A1(ref_1_maj_110_n24), .A2(ref_1_maj_110_n23), 
        .ZN(ref_1_maj_110_n25) );
  NAND2_X1 ref_1_maj_110_U4 ( .A1(ref_1_maj_110_n20), .A2(ref_1_maj_110_n19), 
        .ZN(ref_1_maj_110_n26) );
  NAND2_X1 ref_1_maj_110_U3 ( .A1(ref_1_maj_110_n26), .A2(ref_1_maj_110_n25), 
        .ZN(ref_1_maj_110_port_o) );
  XOR2_X1 ref_1_maj_110_U2 ( .A(ref_1_maj_110_n22), .B(ref_1_maj_110_n21), .Z(
        ref_1_maj_110_n23) );
  NAND2_X1 ref_1_maj_111_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_111_n18) );
  NAND2_X1 ref_1_maj_111_U14 ( .A1(ref_1_maj_111_n21), .A2(ref_1_maj_111_n22), 
        .ZN(ref_1_maj_111_n17) );
  NAND2_X1 ref_1_maj_111_U13 ( .A1(ref_1_maj_111_n18), .A2(ref_1_maj_111_n17), 
        .ZN(ref_1_maj_111_n19) );
  NAND2_X1 ref_1_maj_111_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_111_n16), .ZN(
        ref_1_maj_111_n14) );
  NAND2_X1 ref_1_maj_111_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_111_n15) );
  NAND2_X1 ref_1_maj_111_U10 ( .A1(ref_1_maj_111_n15), .A2(ref_1_maj_111_n14), 
        .ZN(ref_1_maj_111_n20) );
  XOR2_X1 ref_1_maj_111_U9 ( .A(ref_1_n5), .B(ref_1_maj_111_n16), .Z(
        ref_1_maj_111_n21) );
  XOR2_X1 ref_1_maj_111_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_111_n22)
         );
  XOR2_X1 ref_1_maj_111_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_111_n16)
         );
  OR2_X1 ref_1_maj_111_U6 ( .A1(ref_1_maj_111_n20), .A2(ref_1_maj_111_n19), 
        .ZN(ref_1_maj_111_n24) );
  NAND2_X1 ref_1_maj_111_U5 ( .A1(ref_1_maj_111_n24), .A2(ref_1_maj_111_n23), 
        .ZN(ref_1_maj_111_n25) );
  NAND2_X1 ref_1_maj_111_U4 ( .A1(ref_1_maj_111_n20), .A2(ref_1_maj_111_n19), 
        .ZN(ref_1_maj_111_n26) );
  NAND2_X1 ref_1_maj_111_U3 ( .A1(ref_1_maj_111_n26), .A2(ref_1_maj_111_n25), 
        .ZN(ref_1_maj_111_port_o) );
  XOR2_X1 ref_1_maj_111_U2 ( .A(ref_1_maj_111_n22), .B(ref_1_maj_111_n21), .Z(
        ref_1_maj_111_n23) );
  NAND2_X1 ref_1_maj_112_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_112_n18) );
  NAND2_X1 ref_1_maj_112_U14 ( .A1(ref_1_maj_112_n21), .A2(ref_1_maj_112_n22), 
        .ZN(ref_1_maj_112_n17) );
  NAND2_X1 ref_1_maj_112_U13 ( .A1(ref_1_maj_112_n18), .A2(ref_1_maj_112_n17), 
        .ZN(ref_1_maj_112_n19) );
  NAND2_X1 ref_1_maj_112_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_112_n16), .ZN(
        ref_1_maj_112_n14) );
  NAND2_X1 ref_1_maj_112_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_112_n15) );
  NAND2_X1 ref_1_maj_112_U10 ( .A1(ref_1_maj_112_n15), .A2(ref_1_maj_112_n14), 
        .ZN(ref_1_maj_112_n20) );
  XOR2_X1 ref_1_maj_112_U9 ( .A(ref_1_n35), .B(ref_1_maj_112_n16), .Z(
        ref_1_maj_112_n21) );
  XOR2_X1 ref_1_maj_112_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_112_n22) );
  XOR2_X1 ref_1_maj_112_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_112_n16) );
  OR2_X1 ref_1_maj_112_U6 ( .A1(ref_1_maj_112_n20), .A2(ref_1_maj_112_n19), 
        .ZN(ref_1_maj_112_n24) );
  NAND2_X1 ref_1_maj_112_U5 ( .A1(ref_1_maj_112_n24), .A2(ref_1_maj_112_n23), 
        .ZN(ref_1_maj_112_n25) );
  NAND2_X1 ref_1_maj_112_U4 ( .A1(ref_1_maj_112_n20), .A2(ref_1_maj_112_n19), 
        .ZN(ref_1_maj_112_n26) );
  NAND2_X1 ref_1_maj_112_U3 ( .A1(ref_1_maj_112_n26), .A2(ref_1_maj_112_n25), 
        .ZN(ref_1_maj_112_port_o) );
  XOR2_X1 ref_1_maj_112_U2 ( .A(ref_1_maj_112_n22), .B(ref_1_maj_112_n21), .Z(
        ref_1_maj_112_n23) );
  NAND2_X1 ref_1_maj_113_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_113_n18) );
  NAND2_X1 ref_1_maj_113_U14 ( .A1(ref_1_maj_113_n21), .A2(ref_1_maj_113_n22), 
        .ZN(ref_1_maj_113_n17) );
  NAND2_X1 ref_1_maj_113_U13 ( .A1(ref_1_maj_113_n18), .A2(ref_1_maj_113_n17), 
        .ZN(ref_1_maj_113_n19) );
  NAND2_X1 ref_1_maj_113_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_113_n16), .ZN(
        ref_1_maj_113_n14) );
  NAND2_X1 ref_1_maj_113_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_113_n15) );
  NAND2_X1 ref_1_maj_113_U10 ( .A1(ref_1_maj_113_n15), .A2(ref_1_maj_113_n14), 
        .ZN(ref_1_maj_113_n20) );
  XOR2_X1 ref_1_maj_113_U9 ( .A(ref_1_n36), .B(ref_1_maj_113_n16), .Z(
        ref_1_maj_113_n21) );
  XOR2_X1 ref_1_maj_113_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_113_n22) );
  XOR2_X1 ref_1_maj_113_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_113_n16) );
  OR2_X1 ref_1_maj_113_U6 ( .A1(ref_1_maj_113_n20), .A2(ref_1_maj_113_n19), 
        .ZN(ref_1_maj_113_n24) );
  NAND2_X1 ref_1_maj_113_U5 ( .A1(ref_1_maj_113_n24), .A2(ref_1_maj_113_n23), 
        .ZN(ref_1_maj_113_n25) );
  NAND2_X1 ref_1_maj_113_U4 ( .A1(ref_1_maj_113_n20), .A2(ref_1_maj_113_n19), 
        .ZN(ref_1_maj_113_n26) );
  NAND2_X1 ref_1_maj_113_U3 ( .A1(ref_1_maj_113_n26), .A2(ref_1_maj_113_n25), 
        .ZN(ref_1_maj_113_port_o) );
  XOR2_X1 ref_1_maj_113_U2 ( .A(ref_1_maj_113_n22), .B(ref_1_maj_113_n21), .Z(
        ref_1_maj_113_n23) );
  NAND2_X1 ref_1_maj_114_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_114_n18) );
  NAND2_X1 ref_1_maj_114_U14 ( .A1(ref_1_maj_114_n21), .A2(ref_1_maj_114_n22), 
        .ZN(ref_1_maj_114_n17) );
  NAND2_X1 ref_1_maj_114_U13 ( .A1(ref_1_maj_114_n18), .A2(ref_1_maj_114_n17), 
        .ZN(ref_1_maj_114_n19) );
  NAND2_X1 ref_1_maj_114_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_114_n16), .ZN(
        ref_1_maj_114_n14) );
  NAND2_X1 ref_1_maj_114_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_114_n15) );
  NAND2_X1 ref_1_maj_114_U10 ( .A1(ref_1_maj_114_n15), .A2(ref_1_maj_114_n14), 
        .ZN(ref_1_maj_114_n20) );
  XOR2_X1 ref_1_maj_114_U9 ( .A(ref_1_n35), .B(ref_1_maj_114_n16), .Z(
        ref_1_maj_114_n21) );
  XOR2_X1 ref_1_maj_114_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_114_n22) );
  XOR2_X1 ref_1_maj_114_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_114_n16) );
  OR2_X1 ref_1_maj_114_U6 ( .A1(ref_1_maj_114_n20), .A2(ref_1_maj_114_n19), 
        .ZN(ref_1_maj_114_n24) );
  NAND2_X1 ref_1_maj_114_U5 ( .A1(ref_1_maj_114_n24), .A2(ref_1_maj_114_n23), 
        .ZN(ref_1_maj_114_n25) );
  NAND2_X1 ref_1_maj_114_U4 ( .A1(ref_1_maj_114_n20), .A2(ref_1_maj_114_n19), 
        .ZN(ref_1_maj_114_n26) );
  NAND2_X1 ref_1_maj_114_U3 ( .A1(ref_1_maj_114_n26), .A2(ref_1_maj_114_n25), 
        .ZN(ref_1_maj_114_port_o) );
  XOR2_X1 ref_1_maj_114_U2 ( .A(ref_1_maj_114_n22), .B(ref_1_maj_114_n21), .Z(
        ref_1_maj_114_n23) );
  NAND2_X1 ref_1_maj_115_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_115_n18) );
  NAND2_X1 ref_1_maj_115_U14 ( .A1(ref_1_maj_115_n21), .A2(ref_1_maj_115_n22), 
        .ZN(ref_1_maj_115_n17) );
  NAND2_X1 ref_1_maj_115_U13 ( .A1(ref_1_maj_115_n18), .A2(ref_1_maj_115_n17), 
        .ZN(ref_1_maj_115_n19) );
  NAND2_X1 ref_1_maj_115_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_115_n16), .ZN(
        ref_1_maj_115_n14) );
  NAND2_X1 ref_1_maj_115_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_115_n15) );
  NAND2_X1 ref_1_maj_115_U10 ( .A1(ref_1_maj_115_n15), .A2(ref_1_maj_115_n14), 
        .ZN(ref_1_maj_115_n20) );
  XOR2_X1 ref_1_maj_115_U9 ( .A(ref_1_n36), .B(ref_1_maj_115_n16), .Z(
        ref_1_maj_115_n21) );
  XOR2_X1 ref_1_maj_115_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_115_n22) );
  XOR2_X1 ref_1_maj_115_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_115_n16) );
  OR2_X1 ref_1_maj_115_U6 ( .A1(ref_1_maj_115_n20), .A2(ref_1_maj_115_n19), 
        .ZN(ref_1_maj_115_n24) );
  NAND2_X1 ref_1_maj_115_U5 ( .A1(ref_1_maj_115_n24), .A2(ref_1_maj_115_n23), 
        .ZN(ref_1_maj_115_n25) );
  NAND2_X1 ref_1_maj_115_U4 ( .A1(ref_1_maj_115_n20), .A2(ref_1_maj_115_n19), 
        .ZN(ref_1_maj_115_n26) );
  NAND2_X1 ref_1_maj_115_U3 ( .A1(ref_1_maj_115_n26), .A2(ref_1_maj_115_n25), 
        .ZN(ref_1_maj_115_port_o) );
  XOR2_X1 ref_1_maj_115_U2 ( .A(ref_1_maj_115_n22), .B(ref_1_maj_115_n21), .Z(
        ref_1_maj_115_n23) );
  NAND2_X1 ref_1_maj_116_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_116_n18) );
  NAND2_X1 ref_1_maj_116_U14 ( .A1(ref_1_maj_116_n21), .A2(ref_1_maj_116_n22), 
        .ZN(ref_1_maj_116_n17) );
  NAND2_X1 ref_1_maj_116_U13 ( .A1(ref_1_maj_116_n18), .A2(ref_1_maj_116_n17), 
        .ZN(ref_1_maj_116_n19) );
  NAND2_X1 ref_1_maj_116_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_116_n16), .ZN(
        ref_1_maj_116_n14) );
  NAND2_X1 ref_1_maj_116_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_116_n15) );
  NAND2_X1 ref_1_maj_116_U10 ( .A1(ref_1_maj_116_n15), .A2(ref_1_maj_116_n14), 
        .ZN(ref_1_maj_116_n20) );
  XOR2_X1 ref_1_maj_116_U9 ( .A(ref_1_n26), .B(ref_1_maj_116_n16), .Z(
        ref_1_maj_116_n21) );
  XOR2_X1 ref_1_maj_116_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_116_n22) );
  XOR2_X1 ref_1_maj_116_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_116_n16) );
  OR2_X1 ref_1_maj_116_U6 ( .A1(ref_1_maj_116_n20), .A2(ref_1_maj_116_n19), 
        .ZN(ref_1_maj_116_n24) );
  NAND2_X1 ref_1_maj_116_U5 ( .A1(ref_1_maj_116_n24), .A2(ref_1_maj_116_n23), 
        .ZN(ref_1_maj_116_n25) );
  NAND2_X1 ref_1_maj_116_U4 ( .A1(ref_1_maj_116_n20), .A2(ref_1_maj_116_n19), 
        .ZN(ref_1_maj_116_n26) );
  NAND2_X1 ref_1_maj_116_U3 ( .A1(ref_1_maj_116_n26), .A2(ref_1_maj_116_n25), 
        .ZN(ref_1_maj_116_port_o) );
  XOR2_X1 ref_1_maj_116_U2 ( .A(ref_1_maj_116_n22), .B(ref_1_maj_116_n21), .Z(
        ref_1_maj_116_n23) );
  NAND2_X1 ref_1_maj_117_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_117_n18) );
  NAND2_X1 ref_1_maj_117_U14 ( .A1(ref_1_maj_117_n21), .A2(ref_1_maj_117_n22), 
        .ZN(ref_1_maj_117_n17) );
  NAND2_X1 ref_1_maj_117_U13 ( .A1(ref_1_maj_117_n18), .A2(ref_1_maj_117_n17), 
        .ZN(ref_1_maj_117_n19) );
  NAND2_X1 ref_1_maj_117_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_117_n16), .ZN(
        ref_1_maj_117_n14) );
  NAND2_X1 ref_1_maj_117_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_117_n15) );
  NAND2_X1 ref_1_maj_117_U10 ( .A1(ref_1_maj_117_n15), .A2(ref_1_maj_117_n14), 
        .ZN(ref_1_maj_117_n20) );
  XOR2_X1 ref_1_maj_117_U9 ( .A(ref_1_n25), .B(ref_1_maj_117_n16), .Z(
        ref_1_maj_117_n21) );
  XOR2_X1 ref_1_maj_117_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_117_n22) );
  XOR2_X1 ref_1_maj_117_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_117_n16) );
  OR2_X1 ref_1_maj_117_U6 ( .A1(ref_1_maj_117_n20), .A2(ref_1_maj_117_n19), 
        .ZN(ref_1_maj_117_n24) );
  NAND2_X1 ref_1_maj_117_U5 ( .A1(ref_1_maj_117_n24), .A2(ref_1_maj_117_n23), 
        .ZN(ref_1_maj_117_n25) );
  NAND2_X1 ref_1_maj_117_U4 ( .A1(ref_1_maj_117_n20), .A2(ref_1_maj_117_n19), 
        .ZN(ref_1_maj_117_n26) );
  NAND2_X1 ref_1_maj_117_U3 ( .A1(ref_1_maj_117_n26), .A2(ref_1_maj_117_n25), 
        .ZN(ref_1_maj_117_port_o) );
  XOR2_X1 ref_1_maj_117_U2 ( .A(ref_1_maj_117_n22), .B(ref_1_maj_117_n21), .Z(
        ref_1_maj_117_n23) );
  NAND2_X1 ref_1_maj_118_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_118_n18) );
  NAND2_X1 ref_1_maj_118_U14 ( .A1(ref_1_maj_118_n21), .A2(ref_1_maj_118_n22), 
        .ZN(ref_1_maj_118_n17) );
  NAND2_X1 ref_1_maj_118_U13 ( .A1(ref_1_maj_118_n18), .A2(ref_1_maj_118_n17), 
        .ZN(ref_1_maj_118_n19) );
  NAND2_X1 ref_1_maj_118_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_118_n16), .ZN(
        ref_1_maj_118_n14) );
  NAND2_X1 ref_1_maj_118_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_118_n15) );
  NAND2_X1 ref_1_maj_118_U10 ( .A1(ref_1_maj_118_n15), .A2(ref_1_maj_118_n14), 
        .ZN(ref_1_maj_118_n20) );
  XOR2_X1 ref_1_maj_118_U9 ( .A(ref_1_n26), .B(ref_1_maj_118_n16), .Z(
        ref_1_maj_118_n21) );
  XOR2_X1 ref_1_maj_118_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_118_n22) );
  XOR2_X1 ref_1_maj_118_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_118_n16) );
  OR2_X1 ref_1_maj_118_U6 ( .A1(ref_1_maj_118_n20), .A2(ref_1_maj_118_n19), 
        .ZN(ref_1_maj_118_n24) );
  NAND2_X1 ref_1_maj_118_U5 ( .A1(ref_1_maj_118_n24), .A2(ref_1_maj_118_n23), 
        .ZN(ref_1_maj_118_n25) );
  NAND2_X1 ref_1_maj_118_U4 ( .A1(ref_1_maj_118_n20), .A2(ref_1_maj_118_n19), 
        .ZN(ref_1_maj_118_n26) );
  NAND2_X1 ref_1_maj_118_U3 ( .A1(ref_1_maj_118_n26), .A2(ref_1_maj_118_n25), 
        .ZN(ref_1_maj_118_port_o) );
  XOR2_X1 ref_1_maj_118_U2 ( .A(ref_1_maj_118_n22), .B(ref_1_maj_118_n21), .Z(
        ref_1_maj_118_n23) );
  NAND2_X1 ref_1_maj_119_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_119_n18) );
  NAND2_X1 ref_1_maj_119_U14 ( .A1(ref_1_maj_119_n21), .A2(ref_1_maj_119_n22), 
        .ZN(ref_1_maj_119_n17) );
  NAND2_X1 ref_1_maj_119_U13 ( .A1(ref_1_maj_119_n18), .A2(ref_1_maj_119_n17), 
        .ZN(ref_1_maj_119_n19) );
  NAND2_X1 ref_1_maj_119_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_119_n16), .ZN(
        ref_1_maj_119_n14) );
  NAND2_X1 ref_1_maj_119_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_119_n15) );
  NAND2_X1 ref_1_maj_119_U10 ( .A1(ref_1_maj_119_n15), .A2(ref_1_maj_119_n14), 
        .ZN(ref_1_maj_119_n20) );
  XOR2_X1 ref_1_maj_119_U9 ( .A(ref_1_n25), .B(ref_1_maj_119_n16), .Z(
        ref_1_maj_119_n21) );
  XOR2_X1 ref_1_maj_119_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_119_n22) );
  XOR2_X1 ref_1_maj_119_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_119_n16) );
  OR2_X1 ref_1_maj_119_U6 ( .A1(ref_1_maj_119_n20), .A2(ref_1_maj_119_n19), 
        .ZN(ref_1_maj_119_n24) );
  NAND2_X1 ref_1_maj_119_U5 ( .A1(ref_1_maj_119_n24), .A2(ref_1_maj_119_n23), 
        .ZN(ref_1_maj_119_n25) );
  NAND2_X1 ref_1_maj_119_U4 ( .A1(ref_1_maj_119_n20), .A2(ref_1_maj_119_n19), 
        .ZN(ref_1_maj_119_n26) );
  NAND2_X1 ref_1_maj_119_U3 ( .A1(ref_1_maj_119_n26), .A2(ref_1_maj_119_n25), 
        .ZN(ref_1_maj_119_port_o) );
  XOR2_X1 ref_1_maj_119_U2 ( .A(ref_1_maj_119_n22), .B(ref_1_maj_119_n21), .Z(
        ref_1_maj_119_n23) );
  NAND2_X1 ref_1_maj_120_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_120_n18) );
  NAND2_X1 ref_1_maj_120_U14 ( .A1(ref_1_maj_120_n21), .A2(ref_1_maj_120_n22), 
        .ZN(ref_1_maj_120_n17) );
  NAND2_X1 ref_1_maj_120_U13 ( .A1(ref_1_maj_120_n18), .A2(ref_1_maj_120_n17), 
        .ZN(ref_1_maj_120_n19) );
  NAND2_X1 ref_1_maj_120_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_120_n16), .ZN(
        ref_1_maj_120_n14) );
  NAND2_X1 ref_1_maj_120_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_120_n15) );
  NAND2_X1 ref_1_maj_120_U10 ( .A1(ref_1_maj_120_n15), .A2(ref_1_maj_120_n14), 
        .ZN(ref_1_maj_120_n20) );
  XOR2_X1 ref_1_maj_120_U9 ( .A(ref_1_n16), .B(ref_1_maj_120_n16), .Z(
        ref_1_maj_120_n21) );
  XOR2_X1 ref_1_maj_120_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_120_n22) );
  XOR2_X1 ref_1_maj_120_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_120_n16) );
  OR2_X1 ref_1_maj_120_U6 ( .A1(ref_1_maj_120_n20), .A2(ref_1_maj_120_n19), 
        .ZN(ref_1_maj_120_n24) );
  NAND2_X1 ref_1_maj_120_U5 ( .A1(ref_1_maj_120_n24), .A2(ref_1_maj_120_n23), 
        .ZN(ref_1_maj_120_n25) );
  NAND2_X1 ref_1_maj_120_U4 ( .A1(ref_1_maj_120_n20), .A2(ref_1_maj_120_n19), 
        .ZN(ref_1_maj_120_n26) );
  NAND2_X1 ref_1_maj_120_U3 ( .A1(ref_1_maj_120_n26), .A2(ref_1_maj_120_n25), 
        .ZN(ref_1_maj_120_port_o) );
  XOR2_X1 ref_1_maj_120_U2 ( .A(ref_1_maj_120_n22), .B(ref_1_maj_120_n21), .Z(
        ref_1_maj_120_n23) );
  NAND2_X1 ref_1_maj_121_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_121_n18) );
  NAND2_X1 ref_1_maj_121_U14 ( .A1(ref_1_maj_121_n21), .A2(ref_1_maj_121_n22), 
        .ZN(ref_1_maj_121_n17) );
  NAND2_X1 ref_1_maj_121_U13 ( .A1(ref_1_maj_121_n18), .A2(ref_1_maj_121_n17), 
        .ZN(ref_1_maj_121_n19) );
  NAND2_X1 ref_1_maj_121_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_121_n16), .ZN(
        ref_1_maj_121_n14) );
  NAND2_X1 ref_1_maj_121_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_121_n15) );
  NAND2_X1 ref_1_maj_121_U10 ( .A1(ref_1_maj_121_n15), .A2(ref_1_maj_121_n14), 
        .ZN(ref_1_maj_121_n20) );
  XOR2_X1 ref_1_maj_121_U9 ( .A(ref_1_n15), .B(ref_1_maj_121_n16), .Z(
        ref_1_maj_121_n21) );
  XOR2_X1 ref_1_maj_121_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_121_n22) );
  XOR2_X1 ref_1_maj_121_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_121_n16) );
  OR2_X1 ref_1_maj_121_U6 ( .A1(ref_1_maj_121_n20), .A2(ref_1_maj_121_n19), 
        .ZN(ref_1_maj_121_n24) );
  NAND2_X1 ref_1_maj_121_U5 ( .A1(ref_1_maj_121_n24), .A2(ref_1_maj_121_n23), 
        .ZN(ref_1_maj_121_n25) );
  NAND2_X1 ref_1_maj_121_U4 ( .A1(ref_1_maj_121_n20), .A2(ref_1_maj_121_n19), 
        .ZN(ref_1_maj_121_n26) );
  NAND2_X1 ref_1_maj_121_U3 ( .A1(ref_1_maj_121_n26), .A2(ref_1_maj_121_n25), 
        .ZN(ref_1_maj_121_port_o) );
  XOR2_X1 ref_1_maj_121_U2 ( .A(ref_1_maj_121_n22), .B(ref_1_maj_121_n21), .Z(
        ref_1_maj_121_n23) );
  NAND2_X1 ref_1_maj_122_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_122_n18) );
  NAND2_X1 ref_1_maj_122_U14 ( .A1(ref_1_maj_122_n21), .A2(ref_1_maj_122_n22), 
        .ZN(ref_1_maj_122_n17) );
  NAND2_X1 ref_1_maj_122_U13 ( .A1(ref_1_maj_122_n18), .A2(ref_1_maj_122_n17), 
        .ZN(ref_1_maj_122_n19) );
  NAND2_X1 ref_1_maj_122_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_122_n16), .ZN(
        ref_1_maj_122_n14) );
  NAND2_X1 ref_1_maj_122_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_122_n15) );
  NAND2_X1 ref_1_maj_122_U10 ( .A1(ref_1_maj_122_n15), .A2(ref_1_maj_122_n14), 
        .ZN(ref_1_maj_122_n20) );
  XOR2_X1 ref_1_maj_122_U9 ( .A(ref_1_n16), .B(ref_1_maj_122_n16), .Z(
        ref_1_maj_122_n21) );
  XOR2_X1 ref_1_maj_122_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_122_n22) );
  XOR2_X1 ref_1_maj_122_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_122_n16) );
  OR2_X1 ref_1_maj_122_U6 ( .A1(ref_1_maj_122_n20), .A2(ref_1_maj_122_n19), 
        .ZN(ref_1_maj_122_n24) );
  NAND2_X1 ref_1_maj_122_U5 ( .A1(ref_1_maj_122_n24), .A2(ref_1_maj_122_n23), 
        .ZN(ref_1_maj_122_n25) );
  NAND2_X1 ref_1_maj_122_U4 ( .A1(ref_1_maj_122_n20), .A2(ref_1_maj_122_n19), 
        .ZN(ref_1_maj_122_n26) );
  NAND2_X1 ref_1_maj_122_U3 ( .A1(ref_1_maj_122_n26), .A2(ref_1_maj_122_n25), 
        .ZN(ref_1_maj_122_port_o) );
  XOR2_X1 ref_1_maj_122_U2 ( .A(ref_1_maj_122_n22), .B(ref_1_maj_122_n21), .Z(
        ref_1_maj_122_n23) );
  NAND2_X1 ref_1_maj_123_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_123_n18) );
  NAND2_X1 ref_1_maj_123_U14 ( .A1(ref_1_maj_123_n21), .A2(ref_1_maj_123_n22), 
        .ZN(ref_1_maj_123_n17) );
  NAND2_X1 ref_1_maj_123_U13 ( .A1(ref_1_maj_123_n18), .A2(ref_1_maj_123_n17), 
        .ZN(ref_1_maj_123_n19) );
  NAND2_X1 ref_1_maj_123_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_123_n16), .ZN(
        ref_1_maj_123_n14) );
  NAND2_X1 ref_1_maj_123_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_123_n15) );
  NAND2_X1 ref_1_maj_123_U10 ( .A1(ref_1_maj_123_n15), .A2(ref_1_maj_123_n14), 
        .ZN(ref_1_maj_123_n20) );
  XOR2_X1 ref_1_maj_123_U9 ( .A(ref_1_n15), .B(ref_1_maj_123_n16), .Z(
        ref_1_maj_123_n21) );
  XOR2_X1 ref_1_maj_123_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_123_n22) );
  XOR2_X1 ref_1_maj_123_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_123_n16) );
  OR2_X1 ref_1_maj_123_U6 ( .A1(ref_1_maj_123_n20), .A2(ref_1_maj_123_n19), 
        .ZN(ref_1_maj_123_n24) );
  NAND2_X1 ref_1_maj_123_U5 ( .A1(ref_1_maj_123_n24), .A2(ref_1_maj_123_n23), 
        .ZN(ref_1_maj_123_n25) );
  NAND2_X1 ref_1_maj_123_U4 ( .A1(ref_1_maj_123_n20), .A2(ref_1_maj_123_n19), 
        .ZN(ref_1_maj_123_n26) );
  NAND2_X1 ref_1_maj_123_U3 ( .A1(ref_1_maj_123_n26), .A2(ref_1_maj_123_n25), 
        .ZN(ref_1_maj_123_port_o) );
  XOR2_X1 ref_1_maj_123_U2 ( .A(ref_1_maj_123_n22), .B(ref_1_maj_123_n21), .Z(
        ref_1_maj_123_n23) );
  NAND2_X1 ref_1_maj_124_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_124_n18) );
  NAND2_X1 ref_1_maj_124_U14 ( .A1(ref_1_maj_124_n21), .A2(ref_1_maj_124_n22), 
        .ZN(ref_1_maj_124_n17) );
  NAND2_X1 ref_1_maj_124_U13 ( .A1(ref_1_maj_124_n18), .A2(ref_1_maj_124_n17), 
        .ZN(ref_1_maj_124_n19) );
  NAND2_X1 ref_1_maj_124_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_124_n16), .ZN(
        ref_1_maj_124_n14) );
  NAND2_X1 ref_1_maj_124_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_124_n15) );
  NAND2_X1 ref_1_maj_124_U10 ( .A1(ref_1_maj_124_n15), .A2(ref_1_maj_124_n14), 
        .ZN(ref_1_maj_124_n20) );
  XOR2_X1 ref_1_maj_124_U9 ( .A(ref_1_n6), .B(ref_1_maj_124_n16), .Z(
        ref_1_maj_124_n21) );
  XOR2_X1 ref_1_maj_124_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_124_n22) );
  XOR2_X1 ref_1_maj_124_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_124_n16)
         );
  OR2_X1 ref_1_maj_124_U6 ( .A1(ref_1_maj_124_n20), .A2(ref_1_maj_124_n19), 
        .ZN(ref_1_maj_124_n24) );
  NAND2_X1 ref_1_maj_124_U5 ( .A1(ref_1_maj_124_n24), .A2(ref_1_maj_124_n23), 
        .ZN(ref_1_maj_124_n25) );
  NAND2_X1 ref_1_maj_124_U4 ( .A1(ref_1_maj_124_n20), .A2(ref_1_maj_124_n19), 
        .ZN(ref_1_maj_124_n26) );
  NAND2_X1 ref_1_maj_124_U3 ( .A1(ref_1_maj_124_n26), .A2(ref_1_maj_124_n25), 
        .ZN(ref_1_maj_124_port_o) );
  XOR2_X1 ref_1_maj_124_U2 ( .A(ref_1_maj_124_n22), .B(ref_1_maj_124_n21), .Z(
        ref_1_maj_124_n23) );
  NAND2_X1 ref_1_maj_125_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_125_n18) );
  NAND2_X1 ref_1_maj_125_U14 ( .A1(ref_1_maj_125_n21), .A2(ref_1_maj_125_n22), 
        .ZN(ref_1_maj_125_n17) );
  NAND2_X1 ref_1_maj_125_U13 ( .A1(ref_1_maj_125_n18), .A2(ref_1_maj_125_n17), 
        .ZN(ref_1_maj_125_n19) );
  NAND2_X1 ref_1_maj_125_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_125_n16), .ZN(
        ref_1_maj_125_n14) );
  NAND2_X1 ref_1_maj_125_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_125_n15) );
  NAND2_X1 ref_1_maj_125_U10 ( .A1(ref_1_maj_125_n15), .A2(ref_1_maj_125_n14), 
        .ZN(ref_1_maj_125_n20) );
  XOR2_X1 ref_1_maj_125_U9 ( .A(ref_1_n5), .B(ref_1_maj_125_n16), .Z(
        ref_1_maj_125_n21) );
  XOR2_X1 ref_1_maj_125_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_125_n22)
         );
  XOR2_X1 ref_1_maj_125_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_125_n16)
         );
  OR2_X1 ref_1_maj_125_U6 ( .A1(ref_1_maj_125_n20), .A2(ref_1_maj_125_n19), 
        .ZN(ref_1_maj_125_n24) );
  NAND2_X1 ref_1_maj_125_U5 ( .A1(ref_1_maj_125_n24), .A2(ref_1_maj_125_n23), 
        .ZN(ref_1_maj_125_n25) );
  NAND2_X1 ref_1_maj_125_U4 ( .A1(ref_1_maj_125_n20), .A2(ref_1_maj_125_n19), 
        .ZN(ref_1_maj_125_n26) );
  NAND2_X1 ref_1_maj_125_U3 ( .A1(ref_1_maj_125_n26), .A2(ref_1_maj_125_n25), 
        .ZN(ref_1_maj_125_port_o) );
  XOR2_X1 ref_1_maj_125_U2 ( .A(ref_1_maj_125_n22), .B(ref_1_maj_125_n21), .Z(
        ref_1_maj_125_n23) );
  NAND2_X1 ref_1_maj_126_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_126_n18) );
  NAND2_X1 ref_1_maj_126_U14 ( .A1(ref_1_maj_126_n21), .A2(ref_1_maj_126_n22), 
        .ZN(ref_1_maj_126_n17) );
  NAND2_X1 ref_1_maj_126_U13 ( .A1(ref_1_maj_126_n18), .A2(ref_1_maj_126_n17), 
        .ZN(ref_1_maj_126_n19) );
  NAND2_X1 ref_1_maj_126_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_126_n16), .ZN(
        ref_1_maj_126_n14) );
  NAND2_X1 ref_1_maj_126_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_126_n15) );
  NAND2_X1 ref_1_maj_126_U10 ( .A1(ref_1_maj_126_n15), .A2(ref_1_maj_126_n14), 
        .ZN(ref_1_maj_126_n20) );
  XOR2_X1 ref_1_maj_126_U9 ( .A(ref_1_n6), .B(ref_1_maj_126_n16), .Z(
        ref_1_maj_126_n21) );
  XOR2_X1 ref_1_maj_126_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_126_n22) );
  XOR2_X1 ref_1_maj_126_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_126_n16)
         );
  OR2_X1 ref_1_maj_126_U6 ( .A1(ref_1_maj_126_n20), .A2(ref_1_maj_126_n19), 
        .ZN(ref_1_maj_126_n24) );
  NAND2_X1 ref_1_maj_126_U5 ( .A1(ref_1_maj_126_n24), .A2(ref_1_maj_126_n23), 
        .ZN(ref_1_maj_126_n25) );
  NAND2_X1 ref_1_maj_126_U4 ( .A1(ref_1_maj_126_n20), .A2(ref_1_maj_126_n19), 
        .ZN(ref_1_maj_126_n26) );
  NAND2_X1 ref_1_maj_126_U3 ( .A1(ref_1_maj_126_n26), .A2(ref_1_maj_126_n25), 
        .ZN(ref_1_maj_126_port_o) );
  XOR2_X1 ref_1_maj_126_U2 ( .A(ref_1_maj_126_n22), .B(ref_1_maj_126_n21), .Z(
        ref_1_maj_126_n23) );
  NAND2_X1 ref_1_maj_127_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_127_n18) );
  NAND2_X1 ref_1_maj_127_U14 ( .A1(ref_1_maj_127_n21), .A2(ref_1_maj_127_n22), 
        .ZN(ref_1_maj_127_n17) );
  NAND2_X1 ref_1_maj_127_U13 ( .A1(ref_1_maj_127_n18), .A2(ref_1_maj_127_n17), 
        .ZN(ref_1_maj_127_n19) );
  NAND2_X1 ref_1_maj_127_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_127_n16), .ZN(
        ref_1_maj_127_n14) );
  NAND2_X1 ref_1_maj_127_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_127_n15) );
  NAND2_X1 ref_1_maj_127_U10 ( .A1(ref_1_maj_127_n15), .A2(ref_1_maj_127_n14), 
        .ZN(ref_1_maj_127_n20) );
  XOR2_X1 ref_1_maj_127_U9 ( .A(ref_1_n5), .B(ref_1_maj_127_n16), .Z(
        ref_1_maj_127_n21) );
  XOR2_X1 ref_1_maj_127_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_127_n22)
         );
  XOR2_X1 ref_1_maj_127_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_127_n16)
         );
  OR2_X1 ref_1_maj_127_U6 ( .A1(ref_1_maj_127_n20), .A2(ref_1_maj_127_n19), 
        .ZN(ref_1_maj_127_n24) );
  NAND2_X1 ref_1_maj_127_U5 ( .A1(ref_1_maj_127_n24), .A2(ref_1_maj_127_n23), 
        .ZN(ref_1_maj_127_n25) );
  NAND2_X1 ref_1_maj_127_U4 ( .A1(ref_1_maj_127_n20), .A2(ref_1_maj_127_n19), 
        .ZN(ref_1_maj_127_n26) );
  NAND2_X1 ref_1_maj_127_U3 ( .A1(ref_1_maj_127_n26), .A2(ref_1_maj_127_n25), 
        .ZN(ref_1_maj_127_port_o) );
  XOR2_X1 ref_1_maj_127_U2 ( .A(ref_1_maj_127_n22), .B(ref_1_maj_127_n21), .Z(
        ref_1_maj_127_n23) );
  NAND2_X1 ref_1_maj_128_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_128_n18) );
  NAND2_X1 ref_1_maj_128_U14 ( .A1(ref_1_maj_128_n21), .A2(ref_1_maj_128_n22), 
        .ZN(ref_1_maj_128_n17) );
  NAND2_X1 ref_1_maj_128_U13 ( .A1(ref_1_maj_128_n18), .A2(ref_1_maj_128_n17), 
        .ZN(ref_1_maj_128_n19) );
  NAND2_X1 ref_1_maj_128_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_128_n16), .ZN(
        ref_1_maj_128_n14) );
  NAND2_X1 ref_1_maj_128_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_128_n15) );
  NAND2_X1 ref_1_maj_128_U10 ( .A1(ref_1_maj_128_n15), .A2(ref_1_maj_128_n14), 
        .ZN(ref_1_maj_128_n20) );
  XOR2_X1 ref_1_maj_128_U9 ( .A(ref_1_n35), .B(ref_1_maj_128_n16), .Z(
        ref_1_maj_128_n21) );
  XOR2_X1 ref_1_maj_128_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_128_n22) );
  XOR2_X1 ref_1_maj_128_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_128_n16) );
  OR2_X1 ref_1_maj_128_U6 ( .A1(ref_1_maj_128_n20), .A2(ref_1_maj_128_n19), 
        .ZN(ref_1_maj_128_n24) );
  NAND2_X1 ref_1_maj_128_U5 ( .A1(ref_1_maj_128_n24), .A2(ref_1_maj_128_n23), 
        .ZN(ref_1_maj_128_n25) );
  NAND2_X1 ref_1_maj_128_U4 ( .A1(ref_1_maj_128_n20), .A2(ref_1_maj_128_n19), 
        .ZN(ref_1_maj_128_n26) );
  NAND2_X1 ref_1_maj_128_U3 ( .A1(ref_1_maj_128_n26), .A2(ref_1_maj_128_n25), 
        .ZN(ref_1_maj_128_port_o) );
  XOR2_X1 ref_1_maj_128_U2 ( .A(ref_1_maj_128_n22), .B(ref_1_maj_128_n21), .Z(
        ref_1_maj_128_n23) );
  NAND2_X1 ref_1_maj_129_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_129_n18) );
  NAND2_X1 ref_1_maj_129_U14 ( .A1(ref_1_maj_129_n21), .A2(ref_1_maj_129_n22), 
        .ZN(ref_1_maj_129_n17) );
  NAND2_X1 ref_1_maj_129_U13 ( .A1(ref_1_maj_129_n18), .A2(ref_1_maj_129_n17), 
        .ZN(ref_1_maj_129_n19) );
  NAND2_X1 ref_1_maj_129_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_129_n16), .ZN(
        ref_1_maj_129_n14) );
  NAND2_X1 ref_1_maj_129_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_129_n15) );
  NAND2_X1 ref_1_maj_129_U10 ( .A1(ref_1_maj_129_n15), .A2(ref_1_maj_129_n14), 
        .ZN(ref_1_maj_129_n20) );
  XOR2_X1 ref_1_maj_129_U9 ( .A(ref_1_n35), .B(ref_1_maj_129_n16), .Z(
        ref_1_maj_129_n21) );
  XOR2_X1 ref_1_maj_129_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_129_n22) );
  XOR2_X1 ref_1_maj_129_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_129_n16) );
  OR2_X1 ref_1_maj_129_U6 ( .A1(ref_1_maj_129_n20), .A2(ref_1_maj_129_n19), 
        .ZN(ref_1_maj_129_n24) );
  NAND2_X1 ref_1_maj_129_U5 ( .A1(ref_1_maj_129_n24), .A2(ref_1_maj_129_n23), 
        .ZN(ref_1_maj_129_n25) );
  NAND2_X1 ref_1_maj_129_U4 ( .A1(ref_1_maj_129_n20), .A2(ref_1_maj_129_n19), 
        .ZN(ref_1_maj_129_n26) );
  NAND2_X1 ref_1_maj_129_U3 ( .A1(ref_1_maj_129_n26), .A2(ref_1_maj_129_n25), 
        .ZN(ref_1_maj_129_port_o) );
  XOR2_X1 ref_1_maj_129_U2 ( .A(ref_1_maj_129_n22), .B(ref_1_maj_129_n21), .Z(
        ref_1_maj_129_n23) );
  NAND2_X1 ref_1_maj_130_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_130_n18) );
  NAND2_X1 ref_1_maj_130_U14 ( .A1(ref_1_maj_130_n21), .A2(ref_1_maj_130_n22), 
        .ZN(ref_1_maj_130_n17) );
  NAND2_X1 ref_1_maj_130_U13 ( .A1(ref_1_maj_130_n18), .A2(ref_1_maj_130_n17), 
        .ZN(ref_1_maj_130_n19) );
  NAND2_X1 ref_1_maj_130_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_130_n16), .ZN(
        ref_1_maj_130_n14) );
  NAND2_X1 ref_1_maj_130_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_130_n15) );
  NAND2_X1 ref_1_maj_130_U10 ( .A1(ref_1_maj_130_n15), .A2(ref_1_maj_130_n14), 
        .ZN(ref_1_maj_130_n20) );
  XOR2_X1 ref_1_maj_130_U9 ( .A(ref_1_n35), .B(ref_1_maj_130_n16), .Z(
        ref_1_maj_130_n21) );
  XOR2_X1 ref_1_maj_130_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_130_n22) );
  XOR2_X1 ref_1_maj_130_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_130_n16) );
  OR2_X1 ref_1_maj_130_U6 ( .A1(ref_1_maj_130_n20), .A2(ref_1_maj_130_n19), 
        .ZN(ref_1_maj_130_n24) );
  NAND2_X1 ref_1_maj_130_U5 ( .A1(ref_1_maj_130_n24), .A2(ref_1_maj_130_n23), 
        .ZN(ref_1_maj_130_n25) );
  NAND2_X1 ref_1_maj_130_U4 ( .A1(ref_1_maj_130_n20), .A2(ref_1_maj_130_n19), 
        .ZN(ref_1_maj_130_n26) );
  NAND2_X1 ref_1_maj_130_U3 ( .A1(ref_1_maj_130_n26), .A2(ref_1_maj_130_n25), 
        .ZN(ref_1_maj_130_port_o) );
  XOR2_X1 ref_1_maj_130_U2 ( .A(ref_1_maj_130_n22), .B(ref_1_maj_130_n21), .Z(
        ref_1_maj_130_n23) );
  NAND2_X1 ref_1_maj_131_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_131_n18) );
  NAND2_X1 ref_1_maj_131_U14 ( .A1(ref_1_maj_131_n21), .A2(ref_1_maj_131_n22), 
        .ZN(ref_1_maj_131_n17) );
  NAND2_X1 ref_1_maj_131_U13 ( .A1(ref_1_maj_131_n18), .A2(ref_1_maj_131_n17), 
        .ZN(ref_1_maj_131_n19) );
  NAND2_X1 ref_1_maj_131_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_131_n16), .ZN(
        ref_1_maj_131_n14) );
  NAND2_X1 ref_1_maj_131_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_131_n15) );
  NAND2_X1 ref_1_maj_131_U10 ( .A1(ref_1_maj_131_n15), .A2(ref_1_maj_131_n14), 
        .ZN(ref_1_maj_131_n20) );
  XOR2_X1 ref_1_maj_131_U9 ( .A(ref_1_n35), .B(ref_1_maj_131_n16), .Z(
        ref_1_maj_131_n21) );
  XOR2_X1 ref_1_maj_131_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_131_n22) );
  XOR2_X1 ref_1_maj_131_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_131_n16) );
  OR2_X1 ref_1_maj_131_U6 ( .A1(ref_1_maj_131_n20), .A2(ref_1_maj_131_n19), 
        .ZN(ref_1_maj_131_n24) );
  NAND2_X1 ref_1_maj_131_U5 ( .A1(ref_1_maj_131_n24), .A2(ref_1_maj_131_n23), 
        .ZN(ref_1_maj_131_n25) );
  NAND2_X1 ref_1_maj_131_U4 ( .A1(ref_1_maj_131_n20), .A2(ref_1_maj_131_n19), 
        .ZN(ref_1_maj_131_n26) );
  NAND2_X1 ref_1_maj_131_U3 ( .A1(ref_1_maj_131_n26), .A2(ref_1_maj_131_n25), 
        .ZN(ref_1_maj_131_port_o) );
  XOR2_X1 ref_1_maj_131_U2 ( .A(ref_1_maj_131_n22), .B(ref_1_maj_131_n21), .Z(
        ref_1_maj_131_n23) );
  NAND2_X1 ref_1_maj_132_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_132_n18) );
  NAND2_X1 ref_1_maj_132_U14 ( .A1(ref_1_maj_132_n21), .A2(ref_1_maj_132_n22), 
        .ZN(ref_1_maj_132_n17) );
  NAND2_X1 ref_1_maj_132_U13 ( .A1(ref_1_maj_132_n18), .A2(ref_1_maj_132_n17), 
        .ZN(ref_1_maj_132_n19) );
  NAND2_X1 ref_1_maj_132_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_132_n16), .ZN(
        ref_1_maj_132_n14) );
  NAND2_X1 ref_1_maj_132_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_132_n15) );
  NAND2_X1 ref_1_maj_132_U10 ( .A1(ref_1_maj_132_n15), .A2(ref_1_maj_132_n14), 
        .ZN(ref_1_maj_132_n20) );
  XOR2_X1 ref_1_maj_132_U9 ( .A(ref_1_n25), .B(ref_1_maj_132_n16), .Z(
        ref_1_maj_132_n21) );
  XOR2_X1 ref_1_maj_132_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_132_n22) );
  XOR2_X1 ref_1_maj_132_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_132_n16) );
  OR2_X1 ref_1_maj_132_U6 ( .A1(ref_1_maj_132_n20), .A2(ref_1_maj_132_n19), 
        .ZN(ref_1_maj_132_n24) );
  NAND2_X1 ref_1_maj_132_U5 ( .A1(ref_1_maj_132_n24), .A2(ref_1_maj_132_n23), 
        .ZN(ref_1_maj_132_n25) );
  NAND2_X1 ref_1_maj_132_U4 ( .A1(ref_1_maj_132_n20), .A2(ref_1_maj_132_n19), 
        .ZN(ref_1_maj_132_n26) );
  NAND2_X1 ref_1_maj_132_U3 ( .A1(ref_1_maj_132_n26), .A2(ref_1_maj_132_n25), 
        .ZN(ref_1_maj_132_port_o) );
  XOR2_X1 ref_1_maj_132_U2 ( .A(ref_1_maj_132_n22), .B(ref_1_maj_132_n21), .Z(
        ref_1_maj_132_n23) );
  NAND2_X1 ref_1_maj_133_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_133_n18) );
  NAND2_X1 ref_1_maj_133_U14 ( .A1(ref_1_maj_133_n21), .A2(ref_1_maj_133_n22), 
        .ZN(ref_1_maj_133_n17) );
  NAND2_X1 ref_1_maj_133_U13 ( .A1(ref_1_maj_133_n18), .A2(ref_1_maj_133_n17), 
        .ZN(ref_1_maj_133_n19) );
  NAND2_X1 ref_1_maj_133_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_133_n16), .ZN(
        ref_1_maj_133_n14) );
  NAND2_X1 ref_1_maj_133_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_133_n15) );
  NAND2_X1 ref_1_maj_133_U10 ( .A1(ref_1_maj_133_n15), .A2(ref_1_maj_133_n14), 
        .ZN(ref_1_maj_133_n20) );
  XOR2_X1 ref_1_maj_133_U9 ( .A(ref_1_n25), .B(ref_1_maj_133_n16), .Z(
        ref_1_maj_133_n21) );
  XOR2_X1 ref_1_maj_133_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_133_n22) );
  XOR2_X1 ref_1_maj_133_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_133_n16) );
  OR2_X1 ref_1_maj_133_U6 ( .A1(ref_1_maj_133_n20), .A2(ref_1_maj_133_n19), 
        .ZN(ref_1_maj_133_n24) );
  NAND2_X1 ref_1_maj_133_U5 ( .A1(ref_1_maj_133_n24), .A2(ref_1_maj_133_n23), 
        .ZN(ref_1_maj_133_n25) );
  NAND2_X1 ref_1_maj_133_U4 ( .A1(ref_1_maj_133_n20), .A2(ref_1_maj_133_n19), 
        .ZN(ref_1_maj_133_n26) );
  NAND2_X1 ref_1_maj_133_U3 ( .A1(ref_1_maj_133_n26), .A2(ref_1_maj_133_n25), 
        .ZN(ref_1_maj_133_port_o) );
  XOR2_X1 ref_1_maj_133_U2 ( .A(ref_1_maj_133_n22), .B(ref_1_maj_133_n21), .Z(
        ref_1_maj_133_n23) );
  NAND2_X1 ref_1_maj_134_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_134_n18) );
  NAND2_X1 ref_1_maj_134_U14 ( .A1(ref_1_maj_134_n21), .A2(ref_1_maj_134_n22), 
        .ZN(ref_1_maj_134_n17) );
  NAND2_X1 ref_1_maj_134_U13 ( .A1(ref_1_maj_134_n18), .A2(ref_1_maj_134_n17), 
        .ZN(ref_1_maj_134_n19) );
  NAND2_X1 ref_1_maj_134_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_134_n16), .ZN(
        ref_1_maj_134_n14) );
  NAND2_X1 ref_1_maj_134_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_134_n15) );
  NAND2_X1 ref_1_maj_134_U10 ( .A1(ref_1_maj_134_n15), .A2(ref_1_maj_134_n14), 
        .ZN(ref_1_maj_134_n20) );
  XOR2_X1 ref_1_maj_134_U9 ( .A(ref_1_n25), .B(ref_1_maj_134_n16), .Z(
        ref_1_maj_134_n21) );
  XOR2_X1 ref_1_maj_134_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_134_n22) );
  XOR2_X1 ref_1_maj_134_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_134_n16) );
  OR2_X1 ref_1_maj_134_U6 ( .A1(ref_1_maj_134_n20), .A2(ref_1_maj_134_n19), 
        .ZN(ref_1_maj_134_n24) );
  NAND2_X1 ref_1_maj_134_U5 ( .A1(ref_1_maj_134_n24), .A2(ref_1_maj_134_n23), 
        .ZN(ref_1_maj_134_n25) );
  NAND2_X1 ref_1_maj_134_U4 ( .A1(ref_1_maj_134_n20), .A2(ref_1_maj_134_n19), 
        .ZN(ref_1_maj_134_n26) );
  NAND2_X1 ref_1_maj_134_U3 ( .A1(ref_1_maj_134_n26), .A2(ref_1_maj_134_n25), 
        .ZN(ref_1_maj_134_port_o) );
  XOR2_X1 ref_1_maj_134_U2 ( .A(ref_1_maj_134_n22), .B(ref_1_maj_134_n21), .Z(
        ref_1_maj_134_n23) );
  NAND2_X1 ref_1_maj_135_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_135_n18) );
  NAND2_X1 ref_1_maj_135_U14 ( .A1(ref_1_maj_135_n21), .A2(ref_1_maj_135_n22), 
        .ZN(ref_1_maj_135_n17) );
  NAND2_X1 ref_1_maj_135_U13 ( .A1(ref_1_maj_135_n18), .A2(ref_1_maj_135_n17), 
        .ZN(ref_1_maj_135_n19) );
  NAND2_X1 ref_1_maj_135_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_135_n16), .ZN(
        ref_1_maj_135_n14) );
  NAND2_X1 ref_1_maj_135_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_135_n15) );
  NAND2_X1 ref_1_maj_135_U10 ( .A1(ref_1_maj_135_n15), .A2(ref_1_maj_135_n14), 
        .ZN(ref_1_maj_135_n20) );
  XOR2_X1 ref_1_maj_135_U9 ( .A(ref_1_n25), .B(ref_1_maj_135_n16), .Z(
        ref_1_maj_135_n21) );
  XOR2_X1 ref_1_maj_135_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_135_n22) );
  XOR2_X1 ref_1_maj_135_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_135_n16) );
  OR2_X1 ref_1_maj_135_U6 ( .A1(ref_1_maj_135_n20), .A2(ref_1_maj_135_n19), 
        .ZN(ref_1_maj_135_n24) );
  NAND2_X1 ref_1_maj_135_U5 ( .A1(ref_1_maj_135_n24), .A2(ref_1_maj_135_n23), 
        .ZN(ref_1_maj_135_n25) );
  NAND2_X1 ref_1_maj_135_U4 ( .A1(ref_1_maj_135_n20), .A2(ref_1_maj_135_n19), 
        .ZN(ref_1_maj_135_n26) );
  NAND2_X1 ref_1_maj_135_U3 ( .A1(ref_1_maj_135_n26), .A2(ref_1_maj_135_n25), 
        .ZN(ref_1_maj_135_port_o) );
  XOR2_X1 ref_1_maj_135_U2 ( .A(ref_1_maj_135_n22), .B(ref_1_maj_135_n21), .Z(
        ref_1_maj_135_n23) );
  NAND2_X1 ref_1_maj_136_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_136_n18) );
  NAND2_X1 ref_1_maj_136_U14 ( .A1(ref_1_maj_136_n21), .A2(ref_1_maj_136_n22), 
        .ZN(ref_1_maj_136_n17) );
  NAND2_X1 ref_1_maj_136_U13 ( .A1(ref_1_maj_136_n18), .A2(ref_1_maj_136_n17), 
        .ZN(ref_1_maj_136_n19) );
  NAND2_X1 ref_1_maj_136_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_136_n16), .ZN(
        ref_1_maj_136_n14) );
  NAND2_X1 ref_1_maj_136_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_136_n15) );
  NAND2_X1 ref_1_maj_136_U10 ( .A1(ref_1_maj_136_n15), .A2(ref_1_maj_136_n14), 
        .ZN(ref_1_maj_136_n20) );
  XOR2_X1 ref_1_maj_136_U9 ( .A(ref_1_n15), .B(ref_1_maj_136_n16), .Z(
        ref_1_maj_136_n21) );
  XOR2_X1 ref_1_maj_136_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_136_n22) );
  XOR2_X1 ref_1_maj_136_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_136_n16) );
  OR2_X1 ref_1_maj_136_U6 ( .A1(ref_1_maj_136_n20), .A2(ref_1_maj_136_n19), 
        .ZN(ref_1_maj_136_n24) );
  NAND2_X1 ref_1_maj_136_U5 ( .A1(ref_1_maj_136_n24), .A2(ref_1_maj_136_n23), 
        .ZN(ref_1_maj_136_n25) );
  NAND2_X1 ref_1_maj_136_U4 ( .A1(ref_1_maj_136_n20), .A2(ref_1_maj_136_n19), 
        .ZN(ref_1_maj_136_n26) );
  NAND2_X1 ref_1_maj_136_U3 ( .A1(ref_1_maj_136_n26), .A2(ref_1_maj_136_n25), 
        .ZN(ref_1_maj_136_port_o) );
  XOR2_X1 ref_1_maj_136_U2 ( .A(ref_1_maj_136_n22), .B(ref_1_maj_136_n21), .Z(
        ref_1_maj_136_n23) );
  NAND2_X1 ref_1_maj_137_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_137_n18) );
  NAND2_X1 ref_1_maj_137_U14 ( .A1(ref_1_maj_137_n21), .A2(ref_1_maj_137_n22), 
        .ZN(ref_1_maj_137_n17) );
  NAND2_X1 ref_1_maj_137_U13 ( .A1(ref_1_maj_137_n18), .A2(ref_1_maj_137_n17), 
        .ZN(ref_1_maj_137_n19) );
  NAND2_X1 ref_1_maj_137_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_137_n16), .ZN(
        ref_1_maj_137_n14) );
  NAND2_X1 ref_1_maj_137_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_137_n15) );
  NAND2_X1 ref_1_maj_137_U10 ( .A1(ref_1_maj_137_n15), .A2(ref_1_maj_137_n14), 
        .ZN(ref_1_maj_137_n20) );
  XOR2_X1 ref_1_maj_137_U9 ( .A(ref_1_n15), .B(ref_1_maj_137_n16), .Z(
        ref_1_maj_137_n21) );
  XOR2_X1 ref_1_maj_137_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_137_n22) );
  XOR2_X1 ref_1_maj_137_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_137_n16) );
  OR2_X1 ref_1_maj_137_U6 ( .A1(ref_1_maj_137_n20), .A2(ref_1_maj_137_n19), 
        .ZN(ref_1_maj_137_n24) );
  NAND2_X1 ref_1_maj_137_U5 ( .A1(ref_1_maj_137_n24), .A2(ref_1_maj_137_n23), 
        .ZN(ref_1_maj_137_n25) );
  NAND2_X1 ref_1_maj_137_U4 ( .A1(ref_1_maj_137_n20), .A2(ref_1_maj_137_n19), 
        .ZN(ref_1_maj_137_n26) );
  NAND2_X1 ref_1_maj_137_U3 ( .A1(ref_1_maj_137_n26), .A2(ref_1_maj_137_n25), 
        .ZN(ref_1_maj_137_port_o) );
  XOR2_X1 ref_1_maj_137_U2 ( .A(ref_1_maj_137_n22), .B(ref_1_maj_137_n21), .Z(
        ref_1_maj_137_n23) );
  NAND2_X1 ref_1_maj_138_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_138_n18) );
  NAND2_X1 ref_1_maj_138_U14 ( .A1(ref_1_maj_138_n21), .A2(ref_1_maj_138_n22), 
        .ZN(ref_1_maj_138_n17) );
  NAND2_X1 ref_1_maj_138_U13 ( .A1(ref_1_maj_138_n18), .A2(ref_1_maj_138_n17), 
        .ZN(ref_1_maj_138_n19) );
  NAND2_X1 ref_1_maj_138_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_138_n16), .ZN(
        ref_1_maj_138_n14) );
  NAND2_X1 ref_1_maj_138_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_138_n15) );
  NAND2_X1 ref_1_maj_138_U10 ( .A1(ref_1_maj_138_n15), .A2(ref_1_maj_138_n14), 
        .ZN(ref_1_maj_138_n20) );
  XOR2_X1 ref_1_maj_138_U9 ( .A(ref_1_n15), .B(ref_1_maj_138_n16), .Z(
        ref_1_maj_138_n21) );
  XOR2_X1 ref_1_maj_138_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_138_n22) );
  XOR2_X1 ref_1_maj_138_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_138_n16) );
  OR2_X1 ref_1_maj_138_U6 ( .A1(ref_1_maj_138_n20), .A2(ref_1_maj_138_n19), 
        .ZN(ref_1_maj_138_n24) );
  NAND2_X1 ref_1_maj_138_U5 ( .A1(ref_1_maj_138_n24), .A2(ref_1_maj_138_n23), 
        .ZN(ref_1_maj_138_n25) );
  NAND2_X1 ref_1_maj_138_U4 ( .A1(ref_1_maj_138_n20), .A2(ref_1_maj_138_n19), 
        .ZN(ref_1_maj_138_n26) );
  NAND2_X1 ref_1_maj_138_U3 ( .A1(ref_1_maj_138_n26), .A2(ref_1_maj_138_n25), 
        .ZN(ref_1_maj_138_port_o) );
  XOR2_X1 ref_1_maj_138_U2 ( .A(ref_1_maj_138_n22), .B(ref_1_maj_138_n21), .Z(
        ref_1_maj_138_n23) );
  NAND2_X1 ref_1_maj_139_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_139_n18) );
  NAND2_X1 ref_1_maj_139_U14 ( .A1(ref_1_maj_139_n21), .A2(ref_1_maj_139_n22), 
        .ZN(ref_1_maj_139_n17) );
  NAND2_X1 ref_1_maj_139_U13 ( .A1(ref_1_maj_139_n18), .A2(ref_1_maj_139_n17), 
        .ZN(ref_1_maj_139_n19) );
  NAND2_X1 ref_1_maj_139_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_139_n16), .ZN(
        ref_1_maj_139_n14) );
  NAND2_X1 ref_1_maj_139_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_139_n15) );
  NAND2_X1 ref_1_maj_139_U10 ( .A1(ref_1_maj_139_n15), .A2(ref_1_maj_139_n14), 
        .ZN(ref_1_maj_139_n20) );
  XOR2_X1 ref_1_maj_139_U9 ( .A(ref_1_n15), .B(ref_1_maj_139_n16), .Z(
        ref_1_maj_139_n21) );
  XOR2_X1 ref_1_maj_139_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_139_n22) );
  XOR2_X1 ref_1_maj_139_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_139_n16) );
  OR2_X1 ref_1_maj_139_U6 ( .A1(ref_1_maj_139_n20), .A2(ref_1_maj_139_n19), 
        .ZN(ref_1_maj_139_n24) );
  NAND2_X1 ref_1_maj_139_U5 ( .A1(ref_1_maj_139_n24), .A2(ref_1_maj_139_n23), 
        .ZN(ref_1_maj_139_n25) );
  NAND2_X1 ref_1_maj_139_U4 ( .A1(ref_1_maj_139_n20), .A2(ref_1_maj_139_n19), 
        .ZN(ref_1_maj_139_n26) );
  NAND2_X1 ref_1_maj_139_U3 ( .A1(ref_1_maj_139_n26), .A2(ref_1_maj_139_n25), 
        .ZN(ref_1_maj_139_port_o) );
  XOR2_X1 ref_1_maj_139_U2 ( .A(ref_1_maj_139_n22), .B(ref_1_maj_139_n21), .Z(
        ref_1_maj_139_n23) );
  NAND2_X1 ref_1_maj_140_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_140_n18) );
  NAND2_X1 ref_1_maj_140_U14 ( .A1(ref_1_maj_140_n21), .A2(ref_1_maj_140_n22), 
        .ZN(ref_1_maj_140_n17) );
  NAND2_X1 ref_1_maj_140_U13 ( .A1(ref_1_maj_140_n18), .A2(ref_1_maj_140_n17), 
        .ZN(ref_1_maj_140_n19) );
  NAND2_X1 ref_1_maj_140_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_140_n16), .ZN(
        ref_1_maj_140_n14) );
  NAND2_X1 ref_1_maj_140_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_140_n15) );
  NAND2_X1 ref_1_maj_140_U10 ( .A1(ref_1_maj_140_n15), .A2(ref_1_maj_140_n14), 
        .ZN(ref_1_maj_140_n20) );
  XOR2_X1 ref_1_maj_140_U9 ( .A(ref_1_n5), .B(ref_1_maj_140_n16), .Z(
        ref_1_maj_140_n21) );
  XOR2_X1 ref_1_maj_140_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_140_n22)
         );
  XOR2_X1 ref_1_maj_140_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_140_n16)
         );
  OR2_X1 ref_1_maj_140_U6 ( .A1(ref_1_maj_140_n20), .A2(ref_1_maj_140_n19), 
        .ZN(ref_1_maj_140_n24) );
  NAND2_X1 ref_1_maj_140_U5 ( .A1(ref_1_maj_140_n24), .A2(ref_1_maj_140_n23), 
        .ZN(ref_1_maj_140_n25) );
  NAND2_X1 ref_1_maj_140_U4 ( .A1(ref_1_maj_140_n20), .A2(ref_1_maj_140_n19), 
        .ZN(ref_1_maj_140_n26) );
  NAND2_X1 ref_1_maj_140_U3 ( .A1(ref_1_maj_140_n26), .A2(ref_1_maj_140_n25), 
        .ZN(ref_1_maj_140_port_o) );
  XOR2_X1 ref_1_maj_140_U2 ( .A(ref_1_maj_140_n22), .B(ref_1_maj_140_n21), .Z(
        ref_1_maj_140_n23) );
  NAND2_X1 ref_1_maj_141_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_141_n18) );
  NAND2_X1 ref_1_maj_141_U14 ( .A1(ref_1_maj_141_n21), .A2(ref_1_maj_141_n22), 
        .ZN(ref_1_maj_141_n17) );
  NAND2_X1 ref_1_maj_141_U13 ( .A1(ref_1_maj_141_n18), .A2(ref_1_maj_141_n17), 
        .ZN(ref_1_maj_141_n19) );
  NAND2_X1 ref_1_maj_141_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_141_n16), .ZN(
        ref_1_maj_141_n14) );
  NAND2_X1 ref_1_maj_141_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_141_n15) );
  NAND2_X1 ref_1_maj_141_U10 ( .A1(ref_1_maj_141_n15), .A2(ref_1_maj_141_n14), 
        .ZN(ref_1_maj_141_n20) );
  XOR2_X1 ref_1_maj_141_U9 ( .A(ref_1_n5), .B(ref_1_maj_141_n16), .Z(
        ref_1_maj_141_n21) );
  XOR2_X1 ref_1_maj_141_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_141_n22)
         );
  XOR2_X1 ref_1_maj_141_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_141_n16)
         );
  OR2_X1 ref_1_maj_141_U6 ( .A1(ref_1_maj_141_n20), .A2(ref_1_maj_141_n19), 
        .ZN(ref_1_maj_141_n24) );
  NAND2_X1 ref_1_maj_141_U5 ( .A1(ref_1_maj_141_n24), .A2(ref_1_maj_141_n23), 
        .ZN(ref_1_maj_141_n25) );
  NAND2_X1 ref_1_maj_141_U4 ( .A1(ref_1_maj_141_n20), .A2(ref_1_maj_141_n19), 
        .ZN(ref_1_maj_141_n26) );
  NAND2_X1 ref_1_maj_141_U3 ( .A1(ref_1_maj_141_n26), .A2(ref_1_maj_141_n25), 
        .ZN(ref_1_maj_141_port_o) );
  XOR2_X1 ref_1_maj_141_U2 ( .A(ref_1_maj_141_n22), .B(ref_1_maj_141_n21), .Z(
        ref_1_maj_141_n23) );
  NAND2_X1 ref_1_maj_142_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_142_n18) );
  NAND2_X1 ref_1_maj_142_U14 ( .A1(ref_1_maj_142_n21), .A2(ref_1_maj_142_n22), 
        .ZN(ref_1_maj_142_n17) );
  NAND2_X1 ref_1_maj_142_U13 ( .A1(ref_1_maj_142_n18), .A2(ref_1_maj_142_n17), 
        .ZN(ref_1_maj_142_n19) );
  NAND2_X1 ref_1_maj_142_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_142_n16), .ZN(
        ref_1_maj_142_n14) );
  NAND2_X1 ref_1_maj_142_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_142_n15) );
  NAND2_X1 ref_1_maj_142_U10 ( .A1(ref_1_maj_142_n15), .A2(ref_1_maj_142_n14), 
        .ZN(ref_1_maj_142_n20) );
  XOR2_X1 ref_1_maj_142_U9 ( .A(ref_1_n5), .B(ref_1_maj_142_n16), .Z(
        ref_1_maj_142_n21) );
  XOR2_X1 ref_1_maj_142_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_142_n22)
         );
  XOR2_X1 ref_1_maj_142_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_142_n16)
         );
  OR2_X1 ref_1_maj_142_U6 ( .A1(ref_1_maj_142_n20), .A2(ref_1_maj_142_n19), 
        .ZN(ref_1_maj_142_n24) );
  NAND2_X1 ref_1_maj_142_U5 ( .A1(ref_1_maj_142_n24), .A2(ref_1_maj_142_n23), 
        .ZN(ref_1_maj_142_n25) );
  NAND2_X1 ref_1_maj_142_U4 ( .A1(ref_1_maj_142_n20), .A2(ref_1_maj_142_n19), 
        .ZN(ref_1_maj_142_n26) );
  NAND2_X1 ref_1_maj_142_U3 ( .A1(ref_1_maj_142_n26), .A2(ref_1_maj_142_n25), 
        .ZN(ref_1_maj_142_port_o) );
  XOR2_X1 ref_1_maj_142_U2 ( .A(ref_1_maj_142_n22), .B(ref_1_maj_142_n21), .Z(
        ref_1_maj_142_n23) );
  NAND2_X1 ref_1_maj_143_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_143_n18) );
  NAND2_X1 ref_1_maj_143_U14 ( .A1(ref_1_maj_143_n21), .A2(ref_1_maj_143_n22), 
        .ZN(ref_1_maj_143_n17) );
  NAND2_X1 ref_1_maj_143_U13 ( .A1(ref_1_maj_143_n18), .A2(ref_1_maj_143_n17), 
        .ZN(ref_1_maj_143_n19) );
  NAND2_X1 ref_1_maj_143_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_143_n16), .ZN(
        ref_1_maj_143_n14) );
  NAND2_X1 ref_1_maj_143_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_143_n15) );
  NAND2_X1 ref_1_maj_143_U10 ( .A1(ref_1_maj_143_n15), .A2(ref_1_maj_143_n14), 
        .ZN(ref_1_maj_143_n20) );
  XOR2_X1 ref_1_maj_143_U9 ( .A(ref_1_n5), .B(ref_1_maj_143_n16), .Z(
        ref_1_maj_143_n21) );
  XOR2_X1 ref_1_maj_143_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_143_n22)
         );
  XOR2_X1 ref_1_maj_143_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_143_n16)
         );
  OR2_X1 ref_1_maj_143_U6 ( .A1(ref_1_maj_143_n20), .A2(ref_1_maj_143_n19), 
        .ZN(ref_1_maj_143_n24) );
  NAND2_X1 ref_1_maj_143_U5 ( .A1(ref_1_maj_143_n24), .A2(ref_1_maj_143_n23), 
        .ZN(ref_1_maj_143_n25) );
  NAND2_X1 ref_1_maj_143_U4 ( .A1(ref_1_maj_143_n20), .A2(ref_1_maj_143_n19), 
        .ZN(ref_1_maj_143_n26) );
  NAND2_X1 ref_1_maj_143_U3 ( .A1(ref_1_maj_143_n26), .A2(ref_1_maj_143_n25), 
        .ZN(ref_1_maj_143_port_o) );
  XOR2_X1 ref_1_maj_143_U2 ( .A(ref_1_maj_143_n22), .B(ref_1_maj_143_n21), .Z(
        ref_1_maj_143_n23) );
  NAND2_X1 ref_1_maj_144_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_144_n18) );
  NAND2_X1 ref_1_maj_144_U14 ( .A1(ref_1_maj_144_n21), .A2(ref_1_maj_144_n22), 
        .ZN(ref_1_maj_144_n17) );
  NAND2_X1 ref_1_maj_144_U13 ( .A1(ref_1_maj_144_n18), .A2(ref_1_maj_144_n17), 
        .ZN(ref_1_maj_144_n19) );
  NAND2_X1 ref_1_maj_144_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_144_n16), .ZN(
        ref_1_maj_144_n14) );
  NAND2_X1 ref_1_maj_144_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_144_n15) );
  NAND2_X1 ref_1_maj_144_U10 ( .A1(ref_1_maj_144_n15), .A2(ref_1_maj_144_n14), 
        .ZN(ref_1_maj_144_n20) );
  XOR2_X1 ref_1_maj_144_U9 ( .A(ref_1_n35), .B(ref_1_maj_144_n16), .Z(
        ref_1_maj_144_n21) );
  XOR2_X1 ref_1_maj_144_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_144_n22) );
  XOR2_X1 ref_1_maj_144_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_144_n16) );
  OR2_X1 ref_1_maj_144_U6 ( .A1(ref_1_maj_144_n20), .A2(ref_1_maj_144_n19), 
        .ZN(ref_1_maj_144_n24) );
  NAND2_X1 ref_1_maj_144_U5 ( .A1(ref_1_maj_144_n24), .A2(ref_1_maj_144_n23), 
        .ZN(ref_1_maj_144_n25) );
  NAND2_X1 ref_1_maj_144_U4 ( .A1(ref_1_maj_144_n20), .A2(ref_1_maj_144_n19), 
        .ZN(ref_1_maj_144_n26) );
  NAND2_X1 ref_1_maj_144_U3 ( .A1(ref_1_maj_144_n26), .A2(ref_1_maj_144_n25), 
        .ZN(ref_1_maj_144_port_o) );
  XOR2_X1 ref_1_maj_144_U2 ( .A(ref_1_maj_144_n22), .B(ref_1_maj_144_n21), .Z(
        ref_1_maj_144_n23) );
  NAND2_X1 ref_1_maj_145_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_145_n18) );
  NAND2_X1 ref_1_maj_145_U14 ( .A1(ref_1_maj_145_n21), .A2(ref_1_maj_145_n22), 
        .ZN(ref_1_maj_145_n17) );
  NAND2_X1 ref_1_maj_145_U13 ( .A1(ref_1_maj_145_n18), .A2(ref_1_maj_145_n17), 
        .ZN(ref_1_maj_145_n19) );
  NAND2_X1 ref_1_maj_145_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_145_n16), .ZN(
        ref_1_maj_145_n14) );
  NAND2_X1 ref_1_maj_145_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_145_n15) );
  NAND2_X1 ref_1_maj_145_U10 ( .A1(ref_1_maj_145_n15), .A2(ref_1_maj_145_n14), 
        .ZN(ref_1_maj_145_n20) );
  XOR2_X1 ref_1_maj_145_U9 ( .A(ref_1_n36), .B(ref_1_maj_145_n16), .Z(
        ref_1_maj_145_n21) );
  XOR2_X1 ref_1_maj_145_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_145_n22) );
  XOR2_X1 ref_1_maj_145_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_145_n16) );
  OR2_X1 ref_1_maj_145_U6 ( .A1(ref_1_maj_145_n20), .A2(ref_1_maj_145_n19), 
        .ZN(ref_1_maj_145_n24) );
  NAND2_X1 ref_1_maj_145_U5 ( .A1(ref_1_maj_145_n24), .A2(ref_1_maj_145_n23), 
        .ZN(ref_1_maj_145_n25) );
  NAND2_X1 ref_1_maj_145_U4 ( .A1(ref_1_maj_145_n20), .A2(ref_1_maj_145_n19), 
        .ZN(ref_1_maj_145_n26) );
  NAND2_X1 ref_1_maj_145_U3 ( .A1(ref_1_maj_145_n26), .A2(ref_1_maj_145_n25), 
        .ZN(ref_1_maj_145_port_o) );
  XOR2_X1 ref_1_maj_145_U2 ( .A(ref_1_maj_145_n22), .B(ref_1_maj_145_n21), .Z(
        ref_1_maj_145_n23) );
  NAND2_X1 ref_1_maj_146_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_146_n18) );
  NAND2_X1 ref_1_maj_146_U14 ( .A1(ref_1_maj_146_n21), .A2(ref_1_maj_146_n22), 
        .ZN(ref_1_maj_146_n17) );
  NAND2_X1 ref_1_maj_146_U13 ( .A1(ref_1_maj_146_n18), .A2(ref_1_maj_146_n17), 
        .ZN(ref_1_maj_146_n19) );
  NAND2_X1 ref_1_maj_146_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_146_n16), .ZN(
        ref_1_maj_146_n14) );
  NAND2_X1 ref_1_maj_146_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_146_n15) );
  NAND2_X1 ref_1_maj_146_U10 ( .A1(ref_1_maj_146_n15), .A2(ref_1_maj_146_n14), 
        .ZN(ref_1_maj_146_n20) );
  XOR2_X1 ref_1_maj_146_U9 ( .A(ref_1_n36), .B(ref_1_maj_146_n16), .Z(
        ref_1_maj_146_n21) );
  XOR2_X1 ref_1_maj_146_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_146_n22) );
  XOR2_X1 ref_1_maj_146_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_146_n16) );
  OR2_X1 ref_1_maj_146_U6 ( .A1(ref_1_maj_146_n20), .A2(ref_1_maj_146_n19), 
        .ZN(ref_1_maj_146_n24) );
  NAND2_X1 ref_1_maj_146_U5 ( .A1(ref_1_maj_146_n24), .A2(ref_1_maj_146_n23), 
        .ZN(ref_1_maj_146_n25) );
  NAND2_X1 ref_1_maj_146_U4 ( .A1(ref_1_maj_146_n20), .A2(ref_1_maj_146_n19), 
        .ZN(ref_1_maj_146_n26) );
  NAND2_X1 ref_1_maj_146_U3 ( .A1(ref_1_maj_146_n26), .A2(ref_1_maj_146_n25), 
        .ZN(ref_1_maj_146_port_o) );
  XOR2_X1 ref_1_maj_146_U2 ( .A(ref_1_maj_146_n22), .B(ref_1_maj_146_n21), .Z(
        ref_1_maj_146_n23) );
  NAND2_X1 ref_1_maj_147_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_147_n18) );
  NAND2_X1 ref_1_maj_147_U14 ( .A1(ref_1_maj_147_n21), .A2(ref_1_maj_147_n22), 
        .ZN(ref_1_maj_147_n17) );
  NAND2_X1 ref_1_maj_147_U13 ( .A1(ref_1_maj_147_n18), .A2(ref_1_maj_147_n17), 
        .ZN(ref_1_maj_147_n19) );
  NAND2_X1 ref_1_maj_147_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_147_n16), .ZN(
        ref_1_maj_147_n14) );
  NAND2_X1 ref_1_maj_147_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_147_n15) );
  NAND2_X1 ref_1_maj_147_U10 ( .A1(ref_1_maj_147_n15), .A2(ref_1_maj_147_n14), 
        .ZN(ref_1_maj_147_n20) );
  XOR2_X1 ref_1_maj_147_U9 ( .A(ref_1_n36), .B(ref_1_maj_147_n16), .Z(
        ref_1_maj_147_n21) );
  XOR2_X1 ref_1_maj_147_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_147_n22) );
  XOR2_X1 ref_1_maj_147_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_147_n16) );
  OR2_X1 ref_1_maj_147_U6 ( .A1(ref_1_maj_147_n20), .A2(ref_1_maj_147_n19), 
        .ZN(ref_1_maj_147_n24) );
  NAND2_X1 ref_1_maj_147_U5 ( .A1(ref_1_maj_147_n24), .A2(ref_1_maj_147_n23), 
        .ZN(ref_1_maj_147_n25) );
  NAND2_X1 ref_1_maj_147_U4 ( .A1(ref_1_maj_147_n20), .A2(ref_1_maj_147_n19), 
        .ZN(ref_1_maj_147_n26) );
  NAND2_X1 ref_1_maj_147_U3 ( .A1(ref_1_maj_147_n26), .A2(ref_1_maj_147_n25), 
        .ZN(ref_1_maj_147_port_o) );
  XOR2_X1 ref_1_maj_147_U2 ( .A(ref_1_maj_147_n22), .B(ref_1_maj_147_n21), .Z(
        ref_1_maj_147_n23) );
  NAND2_X1 ref_1_maj_148_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_148_n18) );
  NAND2_X1 ref_1_maj_148_U14 ( .A1(ref_1_maj_148_n21), .A2(ref_1_maj_148_n22), 
        .ZN(ref_1_maj_148_n17) );
  NAND2_X1 ref_1_maj_148_U13 ( .A1(ref_1_maj_148_n18), .A2(ref_1_maj_148_n17), 
        .ZN(ref_1_maj_148_n19) );
  NAND2_X1 ref_1_maj_148_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_148_n16), .ZN(
        ref_1_maj_148_n14) );
  NAND2_X1 ref_1_maj_148_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_148_n15) );
  NAND2_X1 ref_1_maj_148_U10 ( .A1(ref_1_maj_148_n15), .A2(ref_1_maj_148_n14), 
        .ZN(ref_1_maj_148_n20) );
  XOR2_X1 ref_1_maj_148_U9 ( .A(ref_1_n26), .B(ref_1_maj_148_n16), .Z(
        ref_1_maj_148_n21) );
  XOR2_X1 ref_1_maj_148_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_148_n22) );
  XOR2_X1 ref_1_maj_148_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_148_n16) );
  OR2_X1 ref_1_maj_148_U6 ( .A1(ref_1_maj_148_n20), .A2(ref_1_maj_148_n19), 
        .ZN(ref_1_maj_148_n24) );
  NAND2_X1 ref_1_maj_148_U5 ( .A1(ref_1_maj_148_n24), .A2(ref_1_maj_148_n23), 
        .ZN(ref_1_maj_148_n25) );
  NAND2_X1 ref_1_maj_148_U4 ( .A1(ref_1_maj_148_n20), .A2(ref_1_maj_148_n19), 
        .ZN(ref_1_maj_148_n26) );
  NAND2_X1 ref_1_maj_148_U3 ( .A1(ref_1_maj_148_n26), .A2(ref_1_maj_148_n25), 
        .ZN(ref_1_maj_148_port_o) );
  XOR2_X1 ref_1_maj_148_U2 ( .A(ref_1_maj_148_n22), .B(ref_1_maj_148_n21), .Z(
        ref_1_maj_148_n23) );
  NAND2_X1 ref_1_maj_149_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_149_n18) );
  NAND2_X1 ref_1_maj_149_U14 ( .A1(ref_1_maj_149_n21), .A2(ref_1_maj_149_n22), 
        .ZN(ref_1_maj_149_n17) );
  NAND2_X1 ref_1_maj_149_U13 ( .A1(ref_1_maj_149_n18), .A2(ref_1_maj_149_n17), 
        .ZN(ref_1_maj_149_n19) );
  NAND2_X1 ref_1_maj_149_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_149_n16), .ZN(
        ref_1_maj_149_n14) );
  NAND2_X1 ref_1_maj_149_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_149_n15) );
  NAND2_X1 ref_1_maj_149_U10 ( .A1(ref_1_maj_149_n15), .A2(ref_1_maj_149_n14), 
        .ZN(ref_1_maj_149_n20) );
  XOR2_X1 ref_1_maj_149_U9 ( .A(ref_1_n26), .B(ref_1_maj_149_n16), .Z(
        ref_1_maj_149_n21) );
  XOR2_X1 ref_1_maj_149_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_149_n22) );
  XOR2_X1 ref_1_maj_149_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_149_n16) );
  OR2_X1 ref_1_maj_149_U6 ( .A1(ref_1_maj_149_n20), .A2(ref_1_maj_149_n19), 
        .ZN(ref_1_maj_149_n24) );
  NAND2_X1 ref_1_maj_149_U5 ( .A1(ref_1_maj_149_n24), .A2(ref_1_maj_149_n23), 
        .ZN(ref_1_maj_149_n25) );
  NAND2_X1 ref_1_maj_149_U4 ( .A1(ref_1_maj_149_n20), .A2(ref_1_maj_149_n19), 
        .ZN(ref_1_maj_149_n26) );
  NAND2_X1 ref_1_maj_149_U3 ( .A1(ref_1_maj_149_n26), .A2(ref_1_maj_149_n25), 
        .ZN(ref_1_maj_149_port_o) );
  XOR2_X1 ref_1_maj_149_U2 ( .A(ref_1_maj_149_n22), .B(ref_1_maj_149_n21), .Z(
        ref_1_maj_149_n23) );
  NAND2_X1 ref_1_maj_150_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_150_n18) );
  NAND2_X1 ref_1_maj_150_U14 ( .A1(ref_1_maj_150_n21), .A2(ref_1_maj_150_n22), 
        .ZN(ref_1_maj_150_n17) );
  NAND2_X1 ref_1_maj_150_U13 ( .A1(ref_1_maj_150_n18), .A2(ref_1_maj_150_n17), 
        .ZN(ref_1_maj_150_n19) );
  NAND2_X1 ref_1_maj_150_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_150_n16), .ZN(
        ref_1_maj_150_n14) );
  NAND2_X1 ref_1_maj_150_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_150_n15) );
  NAND2_X1 ref_1_maj_150_U10 ( .A1(ref_1_maj_150_n15), .A2(ref_1_maj_150_n14), 
        .ZN(ref_1_maj_150_n20) );
  XOR2_X1 ref_1_maj_150_U9 ( .A(ref_1_n26), .B(ref_1_maj_150_n16), .Z(
        ref_1_maj_150_n21) );
  XOR2_X1 ref_1_maj_150_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_150_n22) );
  XOR2_X1 ref_1_maj_150_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_150_n16) );
  OR2_X1 ref_1_maj_150_U6 ( .A1(ref_1_maj_150_n20), .A2(ref_1_maj_150_n19), 
        .ZN(ref_1_maj_150_n24) );
  NAND2_X1 ref_1_maj_150_U5 ( .A1(ref_1_maj_150_n24), .A2(ref_1_maj_150_n23), 
        .ZN(ref_1_maj_150_n25) );
  NAND2_X1 ref_1_maj_150_U4 ( .A1(ref_1_maj_150_n20), .A2(ref_1_maj_150_n19), 
        .ZN(ref_1_maj_150_n26) );
  NAND2_X1 ref_1_maj_150_U3 ( .A1(ref_1_maj_150_n26), .A2(ref_1_maj_150_n25), 
        .ZN(ref_1_maj_150_port_o) );
  XOR2_X1 ref_1_maj_150_U2 ( .A(ref_1_maj_150_n22), .B(ref_1_maj_150_n21), .Z(
        ref_1_maj_150_n23) );
  NAND2_X1 ref_1_maj_151_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_151_n18) );
  NAND2_X1 ref_1_maj_151_U14 ( .A1(ref_1_maj_151_n21), .A2(ref_1_maj_151_n22), 
        .ZN(ref_1_maj_151_n17) );
  NAND2_X1 ref_1_maj_151_U13 ( .A1(ref_1_maj_151_n18), .A2(ref_1_maj_151_n17), 
        .ZN(ref_1_maj_151_n19) );
  NAND2_X1 ref_1_maj_151_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_151_n16), .ZN(
        ref_1_maj_151_n14) );
  NAND2_X1 ref_1_maj_151_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_151_n15) );
  NAND2_X1 ref_1_maj_151_U10 ( .A1(ref_1_maj_151_n15), .A2(ref_1_maj_151_n14), 
        .ZN(ref_1_maj_151_n20) );
  XOR2_X1 ref_1_maj_151_U9 ( .A(ref_1_n26), .B(ref_1_maj_151_n16), .Z(
        ref_1_maj_151_n21) );
  XOR2_X1 ref_1_maj_151_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_151_n22) );
  XOR2_X1 ref_1_maj_151_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_151_n16) );
  OR2_X1 ref_1_maj_151_U6 ( .A1(ref_1_maj_151_n20), .A2(ref_1_maj_151_n19), 
        .ZN(ref_1_maj_151_n24) );
  NAND2_X1 ref_1_maj_151_U5 ( .A1(ref_1_maj_151_n24), .A2(ref_1_maj_151_n23), 
        .ZN(ref_1_maj_151_n25) );
  NAND2_X1 ref_1_maj_151_U4 ( .A1(ref_1_maj_151_n20), .A2(ref_1_maj_151_n19), 
        .ZN(ref_1_maj_151_n26) );
  NAND2_X1 ref_1_maj_151_U3 ( .A1(ref_1_maj_151_n26), .A2(ref_1_maj_151_n25), 
        .ZN(ref_1_maj_151_port_o) );
  XOR2_X1 ref_1_maj_151_U2 ( .A(ref_1_maj_151_n22), .B(ref_1_maj_151_n21), .Z(
        ref_1_maj_151_n23) );
  NAND2_X1 ref_1_maj_152_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_152_n18) );
  NAND2_X1 ref_1_maj_152_U14 ( .A1(ref_1_maj_152_n21), .A2(ref_1_maj_152_n22), 
        .ZN(ref_1_maj_152_n17) );
  NAND2_X1 ref_1_maj_152_U13 ( .A1(ref_1_maj_152_n18), .A2(ref_1_maj_152_n17), 
        .ZN(ref_1_maj_152_n19) );
  NAND2_X1 ref_1_maj_152_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_152_n16), .ZN(
        ref_1_maj_152_n14) );
  NAND2_X1 ref_1_maj_152_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_152_n15) );
  NAND2_X1 ref_1_maj_152_U10 ( .A1(ref_1_maj_152_n15), .A2(ref_1_maj_152_n14), 
        .ZN(ref_1_maj_152_n20) );
  XOR2_X1 ref_1_maj_152_U9 ( .A(ref_1_n16), .B(ref_1_maj_152_n16), .Z(
        ref_1_maj_152_n21) );
  XOR2_X1 ref_1_maj_152_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_152_n22) );
  XOR2_X1 ref_1_maj_152_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_152_n16) );
  OR2_X1 ref_1_maj_152_U6 ( .A1(ref_1_maj_152_n20), .A2(ref_1_maj_152_n19), 
        .ZN(ref_1_maj_152_n24) );
  NAND2_X1 ref_1_maj_152_U5 ( .A1(ref_1_maj_152_n24), .A2(ref_1_maj_152_n23), 
        .ZN(ref_1_maj_152_n25) );
  NAND2_X1 ref_1_maj_152_U4 ( .A1(ref_1_maj_152_n20), .A2(ref_1_maj_152_n19), 
        .ZN(ref_1_maj_152_n26) );
  NAND2_X1 ref_1_maj_152_U3 ( .A1(ref_1_maj_152_n26), .A2(ref_1_maj_152_n25), 
        .ZN(ref_1_maj_152_port_o) );
  XOR2_X1 ref_1_maj_152_U2 ( .A(ref_1_maj_152_n22), .B(ref_1_maj_152_n21), .Z(
        ref_1_maj_152_n23) );
  NAND2_X1 ref_1_maj_153_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_153_n18) );
  NAND2_X1 ref_1_maj_153_U14 ( .A1(ref_1_maj_153_n21), .A2(ref_1_maj_153_n22), 
        .ZN(ref_1_maj_153_n17) );
  NAND2_X1 ref_1_maj_153_U13 ( .A1(ref_1_maj_153_n18), .A2(ref_1_maj_153_n17), 
        .ZN(ref_1_maj_153_n19) );
  NAND2_X1 ref_1_maj_153_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_153_n16), .ZN(
        ref_1_maj_153_n14) );
  NAND2_X1 ref_1_maj_153_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_153_n15) );
  NAND2_X1 ref_1_maj_153_U10 ( .A1(ref_1_maj_153_n15), .A2(ref_1_maj_153_n14), 
        .ZN(ref_1_maj_153_n20) );
  XOR2_X1 ref_1_maj_153_U9 ( .A(ref_1_n16), .B(ref_1_maj_153_n16), .Z(
        ref_1_maj_153_n21) );
  XOR2_X1 ref_1_maj_153_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_153_n22) );
  XOR2_X1 ref_1_maj_153_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_153_n16) );
  OR2_X1 ref_1_maj_153_U6 ( .A1(ref_1_maj_153_n20), .A2(ref_1_maj_153_n19), 
        .ZN(ref_1_maj_153_n24) );
  NAND2_X1 ref_1_maj_153_U5 ( .A1(ref_1_maj_153_n24), .A2(ref_1_maj_153_n23), 
        .ZN(ref_1_maj_153_n25) );
  NAND2_X1 ref_1_maj_153_U4 ( .A1(ref_1_maj_153_n20), .A2(ref_1_maj_153_n19), 
        .ZN(ref_1_maj_153_n26) );
  NAND2_X1 ref_1_maj_153_U3 ( .A1(ref_1_maj_153_n26), .A2(ref_1_maj_153_n25), 
        .ZN(ref_1_maj_153_port_o) );
  XOR2_X1 ref_1_maj_153_U2 ( .A(ref_1_maj_153_n22), .B(ref_1_maj_153_n21), .Z(
        ref_1_maj_153_n23) );
  NAND2_X1 ref_1_maj_154_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_154_n18) );
  NAND2_X1 ref_1_maj_154_U14 ( .A1(ref_1_maj_154_n21), .A2(ref_1_maj_154_n22), 
        .ZN(ref_1_maj_154_n17) );
  NAND2_X1 ref_1_maj_154_U13 ( .A1(ref_1_maj_154_n18), .A2(ref_1_maj_154_n17), 
        .ZN(ref_1_maj_154_n19) );
  NAND2_X1 ref_1_maj_154_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_154_n16), .ZN(
        ref_1_maj_154_n14) );
  NAND2_X1 ref_1_maj_154_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_154_n15) );
  NAND2_X1 ref_1_maj_154_U10 ( .A1(ref_1_maj_154_n15), .A2(ref_1_maj_154_n14), 
        .ZN(ref_1_maj_154_n20) );
  XOR2_X1 ref_1_maj_154_U9 ( .A(ref_1_n16), .B(ref_1_maj_154_n16), .Z(
        ref_1_maj_154_n21) );
  XOR2_X1 ref_1_maj_154_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_154_n22) );
  XOR2_X1 ref_1_maj_154_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_154_n16) );
  OR2_X1 ref_1_maj_154_U6 ( .A1(ref_1_maj_154_n20), .A2(ref_1_maj_154_n19), 
        .ZN(ref_1_maj_154_n24) );
  NAND2_X1 ref_1_maj_154_U5 ( .A1(ref_1_maj_154_n24), .A2(ref_1_maj_154_n23), 
        .ZN(ref_1_maj_154_n25) );
  NAND2_X1 ref_1_maj_154_U4 ( .A1(ref_1_maj_154_n20), .A2(ref_1_maj_154_n19), 
        .ZN(ref_1_maj_154_n26) );
  NAND2_X1 ref_1_maj_154_U3 ( .A1(ref_1_maj_154_n26), .A2(ref_1_maj_154_n25), 
        .ZN(ref_1_maj_154_port_o) );
  XOR2_X1 ref_1_maj_154_U2 ( .A(ref_1_maj_154_n22), .B(ref_1_maj_154_n21), .Z(
        ref_1_maj_154_n23) );
  NAND2_X1 ref_1_maj_155_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_155_n18) );
  NAND2_X1 ref_1_maj_155_U14 ( .A1(ref_1_maj_155_n21), .A2(ref_1_maj_155_n22), 
        .ZN(ref_1_maj_155_n17) );
  NAND2_X1 ref_1_maj_155_U13 ( .A1(ref_1_maj_155_n18), .A2(ref_1_maj_155_n17), 
        .ZN(ref_1_maj_155_n19) );
  NAND2_X1 ref_1_maj_155_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_155_n16), .ZN(
        ref_1_maj_155_n14) );
  NAND2_X1 ref_1_maj_155_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_155_n15) );
  NAND2_X1 ref_1_maj_155_U10 ( .A1(ref_1_maj_155_n15), .A2(ref_1_maj_155_n14), 
        .ZN(ref_1_maj_155_n20) );
  XOR2_X1 ref_1_maj_155_U9 ( .A(ref_1_n16), .B(ref_1_maj_155_n16), .Z(
        ref_1_maj_155_n21) );
  XOR2_X1 ref_1_maj_155_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_155_n22) );
  XOR2_X1 ref_1_maj_155_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_155_n16) );
  OR2_X1 ref_1_maj_155_U6 ( .A1(ref_1_maj_155_n20), .A2(ref_1_maj_155_n19), 
        .ZN(ref_1_maj_155_n24) );
  NAND2_X1 ref_1_maj_155_U5 ( .A1(ref_1_maj_155_n24), .A2(ref_1_maj_155_n23), 
        .ZN(ref_1_maj_155_n25) );
  NAND2_X1 ref_1_maj_155_U4 ( .A1(ref_1_maj_155_n20), .A2(ref_1_maj_155_n19), 
        .ZN(ref_1_maj_155_n26) );
  NAND2_X1 ref_1_maj_155_U3 ( .A1(ref_1_maj_155_n26), .A2(ref_1_maj_155_n25), 
        .ZN(ref_1_maj_155_port_o) );
  XOR2_X1 ref_1_maj_155_U2 ( .A(ref_1_maj_155_n22), .B(ref_1_maj_155_n21), .Z(
        ref_1_maj_155_n23) );
  NAND2_X1 ref_1_maj_156_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_156_n18) );
  NAND2_X1 ref_1_maj_156_U14 ( .A1(ref_1_maj_156_n21), .A2(ref_1_maj_156_n22), 
        .ZN(ref_1_maj_156_n17) );
  NAND2_X1 ref_1_maj_156_U13 ( .A1(ref_1_maj_156_n18), .A2(ref_1_maj_156_n17), 
        .ZN(ref_1_maj_156_n19) );
  NAND2_X1 ref_1_maj_156_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_156_n16), .ZN(
        ref_1_maj_156_n14) );
  NAND2_X1 ref_1_maj_156_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_156_n15) );
  NAND2_X1 ref_1_maj_156_U10 ( .A1(ref_1_maj_156_n15), .A2(ref_1_maj_156_n14), 
        .ZN(ref_1_maj_156_n20) );
  XOR2_X1 ref_1_maj_156_U9 ( .A(ref_1_n6), .B(ref_1_maj_156_n16), .Z(
        ref_1_maj_156_n21) );
  XOR2_X1 ref_1_maj_156_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_156_n22) );
  XOR2_X1 ref_1_maj_156_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_156_n16)
         );
  OR2_X1 ref_1_maj_156_U6 ( .A1(ref_1_maj_156_n20), .A2(ref_1_maj_156_n19), 
        .ZN(ref_1_maj_156_n24) );
  NAND2_X1 ref_1_maj_156_U5 ( .A1(ref_1_maj_156_n24), .A2(ref_1_maj_156_n23), 
        .ZN(ref_1_maj_156_n25) );
  NAND2_X1 ref_1_maj_156_U4 ( .A1(ref_1_maj_156_n20), .A2(ref_1_maj_156_n19), 
        .ZN(ref_1_maj_156_n26) );
  NAND2_X1 ref_1_maj_156_U3 ( .A1(ref_1_maj_156_n26), .A2(ref_1_maj_156_n25), 
        .ZN(ref_1_maj_156_port_o) );
  XOR2_X1 ref_1_maj_156_U2 ( .A(ref_1_maj_156_n22), .B(ref_1_maj_156_n21), .Z(
        ref_1_maj_156_n23) );
  NAND2_X1 ref_1_maj_157_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_157_n18) );
  NAND2_X1 ref_1_maj_157_U14 ( .A1(ref_1_maj_157_n21), .A2(ref_1_maj_157_n22), 
        .ZN(ref_1_maj_157_n17) );
  NAND2_X1 ref_1_maj_157_U13 ( .A1(ref_1_maj_157_n18), .A2(ref_1_maj_157_n17), 
        .ZN(ref_1_maj_157_n19) );
  NAND2_X1 ref_1_maj_157_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_157_n16), .ZN(
        ref_1_maj_157_n14) );
  NAND2_X1 ref_1_maj_157_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_157_n15) );
  NAND2_X1 ref_1_maj_157_U10 ( .A1(ref_1_maj_157_n15), .A2(ref_1_maj_157_n14), 
        .ZN(ref_1_maj_157_n20) );
  XOR2_X1 ref_1_maj_157_U9 ( .A(ref_1_n6), .B(ref_1_maj_157_n16), .Z(
        ref_1_maj_157_n21) );
  XOR2_X1 ref_1_maj_157_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_157_n22) );
  XOR2_X1 ref_1_maj_157_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_157_n16)
         );
  OR2_X1 ref_1_maj_157_U6 ( .A1(ref_1_maj_157_n20), .A2(ref_1_maj_157_n19), 
        .ZN(ref_1_maj_157_n24) );
  NAND2_X1 ref_1_maj_157_U5 ( .A1(ref_1_maj_157_n24), .A2(ref_1_maj_157_n23), 
        .ZN(ref_1_maj_157_n25) );
  NAND2_X1 ref_1_maj_157_U4 ( .A1(ref_1_maj_157_n20), .A2(ref_1_maj_157_n19), 
        .ZN(ref_1_maj_157_n26) );
  NAND2_X1 ref_1_maj_157_U3 ( .A1(ref_1_maj_157_n26), .A2(ref_1_maj_157_n25), 
        .ZN(ref_1_maj_157_port_o) );
  XOR2_X1 ref_1_maj_157_U2 ( .A(ref_1_maj_157_n22), .B(ref_1_maj_157_n21), .Z(
        ref_1_maj_157_n23) );
  NAND2_X1 ref_1_maj_158_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_158_n18) );
  NAND2_X1 ref_1_maj_158_U14 ( .A1(ref_1_maj_158_n21), .A2(ref_1_maj_158_n22), 
        .ZN(ref_1_maj_158_n17) );
  NAND2_X1 ref_1_maj_158_U13 ( .A1(ref_1_maj_158_n18), .A2(ref_1_maj_158_n17), 
        .ZN(ref_1_maj_158_n19) );
  NAND2_X1 ref_1_maj_158_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_158_n16), .ZN(
        ref_1_maj_158_n14) );
  NAND2_X1 ref_1_maj_158_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_158_n15) );
  NAND2_X1 ref_1_maj_158_U10 ( .A1(ref_1_maj_158_n15), .A2(ref_1_maj_158_n14), 
        .ZN(ref_1_maj_158_n20) );
  XOR2_X1 ref_1_maj_158_U9 ( .A(ref_1_n6), .B(ref_1_maj_158_n16), .Z(
        ref_1_maj_158_n21) );
  XOR2_X1 ref_1_maj_158_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_158_n22) );
  XOR2_X1 ref_1_maj_158_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_158_n16)
         );
  OR2_X1 ref_1_maj_158_U6 ( .A1(ref_1_maj_158_n20), .A2(ref_1_maj_158_n19), 
        .ZN(ref_1_maj_158_n24) );
  NAND2_X1 ref_1_maj_158_U5 ( .A1(ref_1_maj_158_n24), .A2(ref_1_maj_158_n23), 
        .ZN(ref_1_maj_158_n25) );
  NAND2_X1 ref_1_maj_158_U4 ( .A1(ref_1_maj_158_n20), .A2(ref_1_maj_158_n19), 
        .ZN(ref_1_maj_158_n26) );
  NAND2_X1 ref_1_maj_158_U3 ( .A1(ref_1_maj_158_n26), .A2(ref_1_maj_158_n25), 
        .ZN(ref_1_maj_158_port_o) );
  XOR2_X1 ref_1_maj_158_U2 ( .A(ref_1_maj_158_n22), .B(ref_1_maj_158_n21), .Z(
        ref_1_maj_158_n23) );
  NAND2_X1 ref_1_maj_159_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_159_n18) );
  NAND2_X1 ref_1_maj_159_U14 ( .A1(ref_1_maj_159_n21), .A2(ref_1_maj_159_n22), 
        .ZN(ref_1_maj_159_n17) );
  NAND2_X1 ref_1_maj_159_U13 ( .A1(ref_1_maj_159_n18), .A2(ref_1_maj_159_n17), 
        .ZN(ref_1_maj_159_n19) );
  NAND2_X1 ref_1_maj_159_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_159_n16), .ZN(
        ref_1_maj_159_n14) );
  NAND2_X1 ref_1_maj_159_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_159_n15) );
  NAND2_X1 ref_1_maj_159_U10 ( .A1(ref_1_maj_159_n15), .A2(ref_1_maj_159_n14), 
        .ZN(ref_1_maj_159_n20) );
  XOR2_X1 ref_1_maj_159_U9 ( .A(ref_1_n6), .B(ref_1_maj_159_n16), .Z(
        ref_1_maj_159_n21) );
  XOR2_X1 ref_1_maj_159_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_159_n22) );
  XOR2_X1 ref_1_maj_159_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_159_n16)
         );
  OR2_X1 ref_1_maj_159_U6 ( .A1(ref_1_maj_159_n20), .A2(ref_1_maj_159_n19), 
        .ZN(ref_1_maj_159_n24) );
  NAND2_X1 ref_1_maj_159_U5 ( .A1(ref_1_maj_159_n24), .A2(ref_1_maj_159_n23), 
        .ZN(ref_1_maj_159_n25) );
  NAND2_X1 ref_1_maj_159_U4 ( .A1(ref_1_maj_159_n20), .A2(ref_1_maj_159_n19), 
        .ZN(ref_1_maj_159_n26) );
  NAND2_X1 ref_1_maj_159_U3 ( .A1(ref_1_maj_159_n26), .A2(ref_1_maj_159_n25), 
        .ZN(ref_1_maj_159_port_o) );
  XOR2_X1 ref_1_maj_159_U2 ( .A(ref_1_maj_159_n22), .B(ref_1_maj_159_n21), .Z(
        ref_1_maj_159_n23) );
endmodule

