
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i0_s5, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, 
        io_i1_s5, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, 
        p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, 
        p_rand_12, p_rand_13, p_rand_14, io_o0_s0, io_o0_s1, io_o0_s2, 
        io_o0_s3, io_o0_s4, io_o0_s5 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i0_s5, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, io_i1_s5,
         p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6,
         p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12,
         p_rand_13, p_rand_14;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5;
  wire   n_dom_0_n78, n_dom_0_n77, n_dom_0_n76, n_dom_0_n75, n_dom_0_n74,
         n_dom_0_n73, n_dom_0_n72, n_dom_0_n71, n_dom_0_n70, n_dom_0_n69,
         n_dom_0_n68, n_dom_0_n67, n_dom_0_n66, n_dom_0_n65, n_dom_0_n64,
         n_dom_0_n63, n_dom_0_n62, n_dom_0_n61, n_dom_0_n60, n_dom_0_n59,
         n_dom_0_n58, n_dom_0_n57, n_dom_0_n56, n_dom_0_n55, n_dom_0_n54,
         n_dom_0_n53, n_dom_0_n52, n_dom_0_n51, n_dom_0_n50, n_dom_0_n49,
         n_dom_0_n48, n_dom_0_n47, n_dom_0_n46, n_dom_0_n45, n_dom_0_n44,
         n_dom_0_n43, n_dom_0_n42, n_dom_0_n41, n_dom_0_n40, n_dom_0_n39,
         n_dom_0_n38, n_dom_0_n37, n_dom_0_n36, n_dom_0_n35, n_dom_0_n34,
         n_dom_0_n33, n_dom_0_n32, n_dom_0_n31, n_dom_0_n30, n_dom_0_n29,
         n_dom_0_n28, n_dom_0_n27, n_dom_0_n26, n_dom_0_n25, n_dom_0_n24,
         n_dom_0_n23, n_dom_0_n22, n_dom_0_n21, n_dom_0_n20, n_dom_0_n19,
         n_dom_0_n18, n_dom_0_n17, n_dom_0_n16, n_dom_0_n15, n_dom_0_n14,
         n_dom_0_n13, n_dom_0_n12, n_dom_0_n11, n_dom_0_n10, n_dom_0_n9,
         n_dom_0_n8, n_dom_0_n7, n_dom_0_n6, n_dom_0_n5, n_dom_0_n4,
         n_dom_0_n3, n_dom_0_n2, n_dom_0_n1, n_dom_0_N41, n_dom_0_N40,
         n_dom_0_N39, n_dom_0_N38, n_dom_0_N37, n_dom_0_N36, n_dom_0_N35,
         n_dom_0__dom_inter5_2, n_dom_0_reg_pipeline, n_dom_0_N34,
         n_dom_0__dom_inter4_7, n_dom_0_reg_pipeline_4, n_dom_0_N33,
         n_dom_0__dom_inter3_12, n_dom_0_reg_pipeline_9, n_dom_0_N32,
         n_dom_0__dom_inter2_17, n_dom_0_reg_pipeline_14, n_dom_0_N31,
         n_dom_0__dom_inter1_22, n_dom_0_reg_pipeline_19, n_dom_0_N30,
         n_dom_0__dom_inter0_27, n_dom_0_reg_pipeline_24, n_dom_0_N29,
         n_dom_0_N28, n_dom_0_N27, n_dom_0_N26, n_dom_0_N25, n_dom_0_N24,
         n_dom_0_N23, n_dom_0_N22, n_dom_0_N21, n_dom_0_N20, n_dom_0_N19,
         n_dom_0_N18, n_dom_0_N17, n_dom_0_N16, n_dom_0_N15, n_dom_0_N14,
         n_dom_0_N13, n_dom_0_N12, n_dom_0_N11, n_dom_0_N10, n_dom_0_N9,
         n_dom_0_N8, n_dom_0_N7, n_dom_0_N6, n_dom_0_N5, n_dom_0_N4,
         n_dom_0_N3, n_dom_0_N2, n_dom_0_N1, n_dom_0_N0;

  NAND2_X1 u_dom_0_U98 ( .A1(io_i0_s0), .A2(io_i1_s5), .ZN(n_dom_0_n54) );
  XNOR2_X1 u_dom_0_U97 ( .A(p_rand_4), .B(n_dom_0_n54), .ZN(n_dom_0_N0) );
  NAND2_X1 u_dom_0_U96 ( .A1(io_i0_s0), .A2(io_i1_s4), .ZN(n_dom_0_n53) );
  XNOR2_X1 u_dom_0_U95 ( .A(p_rand_3), .B(n_dom_0_n53), .ZN(n_dom_0_N1) );
  NAND2_X1 u_dom_0_U94 ( .A1(io_i0_s2), .A2(io_i1_s5), .ZN(n_dom_0_n52) );
  XNOR2_X1 u_dom_0_U93 ( .A(p_rand_11), .B(n_dom_0_n52), .ZN(n_dom_0_N10) );
  NAND2_X1 u_dom_0_U92 ( .A1(io_i0_s2), .A2(io_i1_s4), .ZN(n_dom_0_n51) );
  XNOR2_X1 u_dom_0_U91 ( .A(p_rand_10), .B(n_dom_0_n51), .ZN(n_dom_0_N11) );
  NAND2_X1 u_dom_0_U90 ( .A1(io_i0_s2), .A2(io_i1_s3), .ZN(n_dom_0_n50) );
  XNOR2_X1 u_dom_0_U89 ( .A(p_rand_9), .B(n_dom_0_n50), .ZN(n_dom_0_N12) );
  NAND2_X1 u_dom_0_U88 ( .A1(io_i0_s2), .A2(io_i1_s1), .ZN(n_dom_0_n49) );
  XNOR2_X1 u_dom_0_U87 ( .A(p_rand_5), .B(n_dom_0_n49), .ZN(n_dom_0_N13) );
  NAND2_X1 u_dom_0_U86 ( .A1(io_i0_s2), .A2(io_i1_s0), .ZN(n_dom_0_n48) );
  XNOR2_X1 u_dom_0_U85 ( .A(p_rand_1), .B(n_dom_0_n48), .ZN(n_dom_0_N14) );
  NAND2_X1 u_dom_0_U84 ( .A1(io_i0_s3), .A2(io_i1_s5), .ZN(n_dom_0_n47) );
  XNOR2_X1 u_dom_0_U83 ( .A(p_rand_13), .B(n_dom_0_n47), .ZN(n_dom_0_N15) );
  NAND2_X1 u_dom_0_U82 ( .A1(io_i0_s3), .A2(io_i1_s4), .ZN(n_dom_0_n46) );
  XNOR2_X1 u_dom_0_U81 ( .A(p_rand_12), .B(n_dom_0_n46), .ZN(n_dom_0_N16) );
  NAND2_X1 u_dom_0_U80 ( .A1(io_i0_s3), .A2(io_i1_s2), .ZN(n_dom_0_n45) );
  XNOR2_X1 u_dom_0_U79 ( .A(p_rand_9), .B(n_dom_0_n45), .ZN(n_dom_0_N17) );
  NAND2_X1 u_dom_0_U78 ( .A1(io_i1_s1), .A2(io_i0_s3), .ZN(n_dom_0_n44) );
  XNOR2_X1 u_dom_0_U77 ( .A(p_rand_6), .B(n_dom_0_n44), .ZN(n_dom_0_N18) );
  NAND2_X1 u_dom_0_U76 ( .A1(io_i0_s3), .A2(io_i1_s0), .ZN(n_dom_0_n43) );
  XNOR2_X1 u_dom_0_U75 ( .A(p_rand_2), .B(n_dom_0_n43), .ZN(n_dom_0_N19) );
  NAND2_X1 u_dom_0_U74 ( .A1(io_i0_s0), .A2(io_i1_s3), .ZN(n_dom_0_n42) );
  XNOR2_X1 u_dom_0_U73 ( .A(p_rand_2), .B(n_dom_0_n42), .ZN(n_dom_0_N2) );
  NAND2_X1 u_dom_0_U72 ( .A1(io_i0_s4), .A2(io_i1_s5), .ZN(n_dom_0_n41) );
  XNOR2_X1 u_dom_0_U71 ( .A(p_rand_14), .B(n_dom_0_n41), .ZN(n_dom_0_N20) );
  NAND2_X1 u_dom_0_U70 ( .A1(io_i0_s4), .A2(io_i1_s3), .ZN(n_dom_0_n40) );
  XNOR2_X1 u_dom_0_U69 ( .A(p_rand_12), .B(n_dom_0_n40), .ZN(n_dom_0_N21) );
  NAND2_X1 u_dom_0_U68 ( .A1(io_i0_s4), .A2(io_i1_s2), .ZN(n_dom_0_n39) );
  XNOR2_X1 u_dom_0_U67 ( .A(p_rand_10), .B(n_dom_0_n39), .ZN(n_dom_0_N22) );
  NAND2_X1 u_dom_0_U66 ( .A1(io_i1_s1), .A2(io_i0_s4), .ZN(n_dom_0_n38) );
  XNOR2_X1 u_dom_0_U65 ( .A(p_rand_7), .B(n_dom_0_n38), .ZN(n_dom_0_N23) );
  NAND2_X1 u_dom_0_U64 ( .A1(io_i0_s4), .A2(io_i1_s0), .ZN(n_dom_0_n37) );
  XNOR2_X1 u_dom_0_U63 ( .A(p_rand_3), .B(n_dom_0_n37), .ZN(n_dom_0_N24) );
  NAND2_X1 u_dom_0_U62 ( .A1(io_i0_s5), .A2(io_i1_s4), .ZN(n_dom_0_n36) );
  XNOR2_X1 u_dom_0_U61 ( .A(p_rand_14), .B(n_dom_0_n36), .ZN(n_dom_0_N25) );
  NAND2_X1 u_dom_0_U60 ( .A1(io_i0_s5), .A2(io_i1_s3), .ZN(n_dom_0_n35) );
  XNOR2_X1 u_dom_0_U59 ( .A(p_rand_13), .B(n_dom_0_n35), .ZN(n_dom_0_N26) );
  NAND2_X1 u_dom_0_U58 ( .A1(io_i0_s5), .A2(io_i1_s2), .ZN(n_dom_0_n34) );
  XNOR2_X1 u_dom_0_U57 ( .A(p_rand_11), .B(n_dom_0_n34), .ZN(n_dom_0_N27) );
  NAND2_X1 u_dom_0_U56 ( .A1(io_i0_s5), .A2(io_i1_s1), .ZN(n_dom_0_n33) );
  XNOR2_X1 u_dom_0_U55 ( .A(p_rand_8), .B(n_dom_0_n33), .ZN(n_dom_0_N28) );
  NAND2_X1 u_dom_0_U54 ( .A1(io_i0_s5), .A2(io_i1_s0), .ZN(n_dom_0_n32) );
  XNOR2_X1 u_dom_0_U53 ( .A(p_rand_4), .B(n_dom_0_n32), .ZN(n_dom_0_N29) );
  NAND2_X1 u_dom_0_U52 ( .A1(io_i0_s0), .A2(io_i1_s2), .ZN(n_dom_0_n31) );
  XNOR2_X1 u_dom_0_U51 ( .A(p_rand_1), .B(n_dom_0_n31), .ZN(n_dom_0_N3) );
  XOR2_X1 u_dom_0_U50 ( .A(n_dom_0__dom_inter0_27), .B(n_dom_0_n77), .Z(
        n_dom_0_n30) );
  XOR2_X1 u_dom_0_U49 ( .A(n_dom_0_n30), .B(n_dom_0_n78), .Z(n_dom_0_n27) );
  XOR2_X1 u_dom_0_U48 ( .A(n_dom_0_reg_pipeline_24), .B(n_dom_0_n75), .Z(
        n_dom_0_n29) );
  XOR2_X1 u_dom_0_U47 ( .A(n_dom_0_n76), .B(n_dom_0_n29), .Z(n_dom_0_n28) );
  XOR2_X1 u_dom_0_U46 ( .A(n_dom_0_n27), .B(n_dom_0_n28), .Z(n_dom_0_N30) );
  XOR2_X1 u_dom_0_U45 ( .A(n_dom_0__dom_inter1_22), .B(n_dom_0_n73), .Z(
        n_dom_0_n26) );
  XOR2_X1 u_dom_0_U44 ( .A(n_dom_0_n26), .B(n_dom_0_n74), .Z(n_dom_0_n23) );
  XOR2_X1 u_dom_0_U43 ( .A(n_dom_0_reg_pipeline_19), .B(n_dom_0_n71), .Z(
        n_dom_0_n25) );
  XOR2_X1 u_dom_0_U42 ( .A(n_dom_0_n72), .B(n_dom_0_n25), .Z(n_dom_0_n24) );
  XOR2_X1 u_dom_0_U41 ( .A(n_dom_0_n23), .B(n_dom_0_n24), .Z(n_dom_0_N31) );
  XOR2_X1 u_dom_0_U40 ( .A(n_dom_0__dom_inter2_17), .B(n_dom_0_n69), .Z(
        n_dom_0_n22) );
  XOR2_X1 u_dom_0_U39 ( .A(n_dom_0_n22), .B(n_dom_0_n70), .Z(n_dom_0_n19) );
  XOR2_X1 u_dom_0_U38 ( .A(n_dom_0_reg_pipeline_14), .B(n_dom_0_n67), .Z(
        n_dom_0_n21) );
  XOR2_X1 u_dom_0_U37 ( .A(n_dom_0_n68), .B(n_dom_0_n21), .Z(n_dom_0_n20) );
  XOR2_X1 u_dom_0_U36 ( .A(n_dom_0_n19), .B(n_dom_0_n20), .Z(n_dom_0_N32) );
  XOR2_X1 u_dom_0_U35 ( .A(n_dom_0__dom_inter3_12), .B(n_dom_0_n65), .Z(
        n_dom_0_n18) );
  XOR2_X1 u_dom_0_U34 ( .A(n_dom_0_n18), .B(n_dom_0_n66), .Z(n_dom_0_n15) );
  XOR2_X1 u_dom_0_U33 ( .A(n_dom_0_reg_pipeline_9), .B(n_dom_0_n63), .Z(
        n_dom_0_n17) );
  XOR2_X1 u_dom_0_U32 ( .A(n_dom_0_n64), .B(n_dom_0_n17), .Z(n_dom_0_n16) );
  XOR2_X1 u_dom_0_U31 ( .A(n_dom_0_n15), .B(n_dom_0_n16), .Z(n_dom_0_N33) );
  XOR2_X1 u_dom_0_U30 ( .A(n_dom_0__dom_inter4_7), .B(n_dom_0_n61), .Z(
        n_dom_0_n14) );
  XOR2_X1 u_dom_0_U29 ( .A(n_dom_0_n14), .B(n_dom_0_n62), .Z(n_dom_0_n11) );
  XOR2_X1 u_dom_0_U28 ( .A(n_dom_0_reg_pipeline_4), .B(n_dom_0_n59), .Z(
        n_dom_0_n13) );
  XOR2_X1 u_dom_0_U27 ( .A(n_dom_0_n60), .B(n_dom_0_n13), .Z(n_dom_0_n12) );
  XOR2_X1 u_dom_0_U26 ( .A(n_dom_0_n11), .B(n_dom_0_n12), .Z(n_dom_0_N34) );
  XOR2_X1 u_dom_0_U25 ( .A(n_dom_0__dom_inter5_2), .B(n_dom_0_n57), .Z(
        n_dom_0_n10) );
  XOR2_X1 u_dom_0_U24 ( .A(n_dom_0_n10), .B(n_dom_0_n58), .Z(n_dom_0_n7) );
  XOR2_X1 u_dom_0_U23 ( .A(n_dom_0_reg_pipeline), .B(n_dom_0_n55), .Z(
        n_dom_0_n9) );
  XOR2_X1 u_dom_0_U22 ( .A(n_dom_0_n56), .B(n_dom_0_n9), .Z(n_dom_0_n8) );
  XOR2_X1 u_dom_0_U21 ( .A(n_dom_0_n7), .B(n_dom_0_n8), .Z(n_dom_0_N35) );
  AND2_X1 u_dom_0_U20 ( .A1(io_i1_s5), .A2(io_i0_s5), .ZN(n_dom_0_N36) );
  AND2_X1 u_dom_0_U19 ( .A1(io_i1_s2), .A2(io_i0_s2), .ZN(n_dom_0_N37) );
  AND2_X1 u_dom_0_U18 ( .A1(io_i0_s1), .A2(io_i1_s1), .ZN(n_dom_0_N38) );
  AND2_X1 u_dom_0_U17 ( .A1(io_i1_s0), .A2(io_i0_s0), .ZN(n_dom_0_N39) );
  NAND2_X1 u_dom_0_U16 ( .A1(io_i1_s1), .A2(io_i0_s0), .ZN(n_dom_0_n6) );
  XNOR2_X1 u_dom_0_U15 ( .A(p_rand_0), .B(n_dom_0_n6), .ZN(n_dom_0_N4) );
  AND2_X1 u_dom_0_U14 ( .A1(io_i1_s4), .A2(io_i0_s4), .ZN(n_dom_0_N40) );
  AND2_X1 u_dom_0_U13 ( .A1(io_i1_s3), .A2(io_i0_s3), .ZN(n_dom_0_N41) );
  NAND2_X1 u_dom_0_U12 ( .A1(io_i1_s5), .A2(io_i0_s1), .ZN(n_dom_0_n5) );
  XNOR2_X1 u_dom_0_U11 ( .A(p_rand_8), .B(n_dom_0_n5), .ZN(n_dom_0_N5) );
  NAND2_X1 u_dom_0_U10 ( .A1(io_i1_s4), .A2(io_i0_s1), .ZN(n_dom_0_n4) );
  XNOR2_X1 u_dom_0_U9 ( .A(p_rand_7), .B(n_dom_0_n4), .ZN(n_dom_0_N6) );
  NAND2_X1 u_dom_0_U8 ( .A1(io_i1_s3), .A2(io_i0_s1), .ZN(n_dom_0_n3) );
  XNOR2_X1 u_dom_0_U7 ( .A(p_rand_6), .B(n_dom_0_n3), .ZN(n_dom_0_N7) );
  NAND2_X1 u_dom_0_U6 ( .A1(io_i1_s2), .A2(io_i0_s1), .ZN(n_dom_0_n2) );
  XNOR2_X1 u_dom_0_U5 ( .A(p_rand_5), .B(n_dom_0_n2), .ZN(n_dom_0_N8) );
  NAND2_X1 u_dom_0_U4 ( .A1(io_i1_s0), .A2(io_i0_s1), .ZN(n_dom_0_n1) );
  XNOR2_X1 u_dom_0_U3 ( .A(p_rand_0), .B(n_dom_0_n1), .ZN(n_dom_0_N9) );
  DFF_X1 u_dom_0_dom_out4_reg ( .D(n_dom_0_N34), .CK(clock_0), .Q(io_o0_s4), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter4_8_reg ( .D(n_dom_0_N24), .CK(clock_0), .Q(), .QN(
        n_dom_0_n62) );
  DFF_X1 u_dom_0_dom_out5_reg ( .D(n_dom_0_N35), .CK(clock_0), .Q(io_o0_s5), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter5_reg ( .D(n_dom_0_N25), .CK(clock_0), .Q(), .QN(
        n_dom_0_n55) );
  DFF_X1 u_dom_0_dom_out3_reg ( .D(n_dom_0_N33), .CK(clock_0), .Q(io_o0_s3), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter3_11_reg ( .D(n_dom_0_N17), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n65) );
  DFF_X1 u_dom_0__dom_inter5_0_reg ( .D(n_dom_0_N26), .CK(clock_0), .Q(), .QN(
        n_dom_0_n56) );
  DFF_X1 u_dom_0__dom_inter4_5_reg ( .D(n_dom_0_N21), .CK(clock_0), .Q(), .QN(
        n_dom_0_n60) );
  DFF_X1 u_dom_0_dom_out2_reg ( .D(n_dom_0_N32), .CK(clock_0), .Q(io_o0_s2), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter2_reg ( .D(n_dom_0_N10), .CK(clock_0), .Q(), .QN(
        n_dom_0_n67) );
  DFF_X1 u_dom_0__dom_inter5_1_reg ( .D(n_dom_0_N27), .CK(clock_0), .Q(), .QN(
        n_dom_0_n57) );
  DFF_X1 u_dom_0__dom_inter5_2_reg ( .D(n_dom_0_N28), .CK(clock_0), .Q(
        n_dom_0__dom_inter5_2), .QN() );
  DFF_X1 u_dom_0__dom_inter5_3_reg ( .D(n_dom_0_N29), .CK(clock_0), .Q(), .QN(
        n_dom_0_n58) );
  DFF_X1 u_dom_0__dom_inter3_reg ( .D(n_dom_0_N15), .CK(clock_0), .Q(), .QN(
        n_dom_0_n63) );
  DFF_X1 u_dom_0_reg_pipeline_9_reg ( .D(n_dom_0_N41), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_9), .QN() );
  DFF_X1 u_dom_0__dom_inter3_12_reg ( .D(n_dom_0_N18), .CK(clock_0), .Q(
        n_dom_0__dom_inter3_12), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_4_reg ( .D(n_dom_0_N40), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_4), .QN() );
  DFF_X1 u_dom_0_dom_out1_reg ( .D(n_dom_0_N31), .CK(clock_0), .Q(io_o0_s1), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter1_22_reg ( .D(n_dom_0_N8), .CK(clock_0), .Q(
        n_dom_0__dom_inter1_22), .QN() );
  DFF_X1 u_dom_0_dom_out0_reg ( .D(n_dom_0_N30), .CK(clock_0), .Q(io_o0_s0), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter0_26_reg ( .D(n_dom_0_N2), .CK(clock_0), .Q(), .QN(
        n_dom_0_n77) );
  DFF_X1 u_dom_0_reg_pipeline_24_reg ( .D(n_dom_0_N39), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_24), .QN() );
  DFF_X1 u_dom_0__dom_inter1_20_reg ( .D(n_dom_0_N6), .CK(clock_0), .Q(), .QN(
        n_dom_0_n72) );
  DFF_X1 u_dom_0_reg_pipeline_19_reg ( .D(n_dom_0_N38), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_19), .QN() );
  DFF_X1 u_dom_0__dom_inter2_17_reg ( .D(n_dom_0_N13), .CK(clock_0), .Q(
        n_dom_0__dom_inter2_17), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_14_reg ( .D(n_dom_0_N37), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_14), .QN() );
  DFF_X1 u_dom_0__dom_inter3_10_reg ( .D(n_dom_0_N16), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n64) );
  DFF_X1 u_dom_0_reg_pipeline_reg ( .D(n_dom_0_N36), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline), .QN() );
  DFF_X1 u_dom_0__dom_inter3_13_reg ( .D(n_dom_0_N19), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n66) );
  DFF_X1 u_dom_0__dom_inter4_6_reg ( .D(n_dom_0_N22), .CK(clock_0), .Q(), .QN(
        n_dom_0_n61) );
  DFF_X1 u_dom_0__dom_inter0_28_reg ( .D(n_dom_0_N4), .CK(clock_0), .Q(), .QN(
        n_dom_0_n78) );
  DFF_X1 u_dom_0__dom_inter2_16_reg ( .D(n_dom_0_N12), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n69) );
  DFF_X1 u_dom_0__dom_inter1_reg ( .D(n_dom_0_N5), .CK(clock_0), .Q(), .QN(
        n_dom_0_n71) );
  DFF_X1 u_dom_0__dom_inter2_18_reg ( .D(n_dom_0_N14), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n70) );
  DFF_X1 u_dom_0__dom_inter0_27_reg ( .D(n_dom_0_N3), .CK(clock_0), .Q(
        n_dom_0__dom_inter0_27), .QN() );
  DFF_X1 u_dom_0__dom_inter0_reg ( .D(n_dom_0_N0), .CK(clock_0), .Q(), .QN(
        n_dom_0_n75) );
  DFF_X1 u_dom_0__dom_inter2_15_reg ( .D(n_dom_0_N11), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n68) );
  DFF_X1 u_dom_0__dom_inter4_reg ( .D(n_dom_0_N20), .CK(clock_0), .Q(), .QN(
        n_dom_0_n59) );
  DFF_X1 u_dom_0__dom_inter1_23_reg ( .D(n_dom_0_N9), .CK(clock_0), .Q(), .QN(
        n_dom_0_n74) );
  DFF_X1 u_dom_0__dom_inter4_7_reg ( .D(n_dom_0_N23), .CK(clock_0), .Q(
        n_dom_0__dom_inter4_7), .QN() );
  DFF_X1 u_dom_0__dom_inter0_25_reg ( .D(n_dom_0_N1), .CK(clock_0), .Q(), .QN(
        n_dom_0_n76) );
  DFF_X1 u_dom_0__dom_inter1_21_reg ( .D(n_dom_0_N7), .CK(clock_0), .Q(), .QN(
        n_dom_0_n73) );
endmodule

