module PresentSbox_keyAdd ( clock, reset, io_state, io_key, io_out );
  input [3:0] io_state;
  input [3:0] io_key;
  output [3:0] io_out;
  input clock, reset;
  wire   sbox_io_o0, sbox_io_o1, sbox_io_o2, sbox_io_o3, sbox_n18, sbox_n17,
         sbox_n16, sbox_n15, sbox_n14, sbox_n13, sbox_n12, sbox_n11, sbox_n10,
         sbox_n9, sbox_n8, sbox_n7, sbox_n6, sbox_n5, sbox_n4, sbox_n3,
         sbox_n2, sbox_n1;

  XOR2_X1 U5 ( .A(sbox_io_o3), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 U6 ( .A(sbox_io_o2), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 U7 ( .A(sbox_io_o1), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 U8 ( .A(sbox_io_o0), .B(io_key[0]), .Z(io_out[0]) );
  INV_X1 sbox_U22 ( .A(io_state[1]), .ZN(sbox_n18) );
  NOR2_X1 sbox_U21 ( .A1(sbox_n18), .A2(io_state[2]), .ZN(sbox_n1) );
  AND2_X1 sbox_U20 ( .A1(io_state[2]), .A2(sbox_n18), .ZN(sbox_n17) );
  OR2_X1 sbox_U19 ( .A1(sbox_n1), .A2(sbox_n17), .ZN(sbox_n13) );
  INV_X1 sbox_U18 ( .A(io_state[3]), .ZN(sbox_n12) );
  XNOR2_X1 sbox_U17 ( .A(sbox_n13), .B(sbox_n12), .ZN(sbox_n15) );
  NOR2_X1 sbox_U16 ( .A1(sbox_n13), .A2(io_state[0]), .ZN(sbox_n11) );
  OR2_X1 sbox_U15 ( .A1(sbox_n11), .A2(sbox_n1), .ZN(sbox_n14) );
  XNOR2_X1 sbox_U14 ( .A(io_state[0]), .B(io_state[2]), .ZN(sbox_n4) );
  XOR2_X1 sbox_U13 ( .A(sbox_n14), .B(sbox_n4), .Z(sbox_n16) );
  NAND2_X1 sbox_U12 ( .A1(sbox_n15), .A2(sbox_n16), .ZN(sbox_n3) );
  XNOR2_X1 sbox_U11 ( .A(sbox_n14), .B(io_state[3]), .ZN(sbox_n6) );
  XOR2_X1 sbox_U10 ( .A(sbox_n3), .B(sbox_n6), .Z(sbox_io_o0) );
  XNOR2_X1 sbox_U9 ( .A(io_state[0]), .B(sbox_n12), .ZN(sbox_n2) );
  XOR2_X1 sbox_U8 ( .A(sbox_n13), .B(sbox_n2), .Z(sbox_n8) );
  NOR2_X1 sbox_U7 ( .A1(sbox_n11), .A2(sbox_n12), .ZN(sbox_n10) );
  XOR2_X1 sbox_U6 ( .A(sbox_n4), .B(sbox_n10), .Z(sbox_n9) );
  NAND2_X1 sbox_U5 ( .A1(sbox_n8), .A2(sbox_n9), .ZN(sbox_n7) );
  XOR2_X1 sbox_U4 ( .A(sbox_n7), .B(io_state[2]), .Z(sbox_n5) );
  XOR2_X1 sbox_U3 ( .A(sbox_n5), .B(sbox_n6), .Z(sbox_io_o1) );
  XOR2_X1 sbox_U2 ( .A(sbox_n3), .B(sbox_n4), .Z(sbox_io_o2) );
  XOR2_X1 sbox_U1 ( .A(sbox_n1), .B(sbox_n2), .Z(sbox_io_o3) );
endmodule