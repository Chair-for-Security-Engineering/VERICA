
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i1_s0, 
        io_i1_s1, io_i1_s2, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, 
        p_rand_5, io_o0_s0, io_o0_s1, io_o0_s2 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i1_s0, io_i1_s1,
         io_i1_s2, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5;
  output io_o0_s0, io_o0_s1, io_o0_s2;
  wire   n_hpc2_0_n21, n_hpc2_0_n20, n_hpc2_0_n19, n_hpc2_0_n18, n_hpc2_0_n17,
         n_hpc2_0_n16, n_hpc2_0_n15, n_hpc2_0_n14, n_hpc2_0_n13, n_hpc2_0_n12,
         n_hpc2_0_n11, n_hpc2_0_n10, n_hpc2_0_n9, n_hpc2_0_n8, n_hpc2_0_n7,
         n_hpc2_0_n6, n_hpc2_0_n5, n_hpc2_0_n4, n_hpc2_0_n3, n_hpc2_0_n2,
         n_hpc2_0_n1, n_hpc2_0_N11, n_hpc2_0_N10, n_hpc2_0_N9, n_hpc2_0_N8,
         n_hpc2_0_N7, n_hpc2_0_N6, n_hpc2_0_N5, n_hpc2_0_N4, n_hpc2_0_N3,
         n_hpc2_0_reg_pipeline_4, n_hpc2_0_reg_pipeline_3,
         n_hpc2_0_reg_pipeline_2, n_hpc2_0_reg_pipeline_1,
         n_hpc2_0_reg_pipeline_0, n_hpc2_0_reg_pipeline, n_hpc2_0_N2,
         n_hpc2_0_N1, n_hpc2_0_N0, n_hpc2_0__hpc1_z21, n_hpc2_0__hpc1_z11,
         n_hpc2_0__hpc1_z01;

  XOR2_X1 u_hpc2_0_U29 ( .A(io_i1_s0), .B(p_rand_1), .Z(n_hpc2_0_n15) );
  XOR2_X1 u_hpc2_0_U28 ( .A(p_rand_0), .B(n_hpc2_0_n15), .Z(n_hpc2_0_N0) );
  XOR2_X1 u_hpc2_0_U27 ( .A(io_i1_s1), .B(p_rand_2), .Z(n_hpc2_0_n14) );
  XOR2_X1 u_hpc2_0_U26 ( .A(p_rand_0), .B(n_hpc2_0_n14), .Z(n_hpc2_0_N1) );
  NAND2_X1 u_hpc2_0_U25 ( .A1(n_hpc2_0_reg_pipeline_4), .A2(n_hpc2_0_n3), .ZN(
        n_hpc2_0_n13) );
  XNOR2_X1 u_hpc2_0_U24 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N10) );
  AND2_X1 u_hpc2_0_U23 ( .A1(n_hpc2_0_n2), .A2(n_hpc2_0_reg_pipeline_4), .ZN(
        n_hpc2_0_N11) );
  XOR2_X1 u_hpc2_0_U22 ( .A(io_i1_s2), .B(p_rand_2), .Z(n_hpc2_0_n12) );
  XOR2_X1 u_hpc2_0_U21 ( .A(p_rand_1), .B(n_hpc2_0_n12), .Z(n_hpc2_0_N2) );
  AND2_X1 u_hpc2_0_U20 ( .A1(n_hpc2_0_n1), .A2(n_hpc2_0_reg_pipeline), .ZN(
        n_hpc2_0_N3) );
  NAND2_X1 u_hpc2_0_U19 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n3), .ZN(
        n_hpc2_0_n11) );
  XNOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N4) );
  NAND2_X1 u_hpc2_0_U17 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n10) );
  XNOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N5) );
  NAND2_X1 u_hpc2_0_U15 ( .A1(n_hpc2_0_reg_pipeline_2), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n9) );
  XNOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N6) );
  AND2_X1 u_hpc2_0_U13 ( .A1(n_hpc2_0_n3), .A2(n_hpc2_0_reg_pipeline_2), .ZN(
        n_hpc2_0_N7) );
  NAND2_X1 u_hpc2_0_U12 ( .A1(n_hpc2_0_reg_pipeline_2), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n8) );
  XNOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N8) );
  NAND2_X1 u_hpc2_0_U10 ( .A1(n_hpc2_0_reg_pipeline_4), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n7) );
  XNOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N9) );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0__hpc1_z01), .B(n_hpc2_0_n20), .Z(
        n_hpc2_0_n6) );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0_n6), .B(n_hpc2_0_n21), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0__hpc1_z11), .B(n_hpc2_0_n18), .Z(
        n_hpc2_0_n5) );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0_n5), .B(n_hpc2_0_n19), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0__hpc1_z21), .B(n_hpc2_0_n16), .Z(
        n_hpc2_0_n4) );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n4), .B(n_hpc2_0_n17), .Z(io_o0_s2) );
  DFF_X1 u_hpc2_0__hpc1_z12_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n19) );
  DFF_X1 u_hpc2_0__hpc1_z11_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z11), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z10_reg ( .D(n_hpc2_0_N6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n18) );
  DFF_X1 u_hpc2_0__hpc1_z02_reg ( .D(n_hpc2_0_N5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n21) );
  DFF_X1 u_hpc2_0__hpc1_z01_reg ( .D(n_hpc2_0_N4), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z01), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z00_reg ( .D(n_hpc2_0_N3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n20) );
  DFF_X1 u_hpc2_0__hpc1_z21_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z21), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z22_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n17) );
  DFF_X1 u_hpc2_0__hpc1_z20_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n16) );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(io_i0_s2), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_4), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(io_i0_s0), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v1_reg ( .D(n_hpc2_0_N1), .CK(clock_0), .Q(
        n_hpc2_0_n3), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(p_rand_4), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_1), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(p_rand_5), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_3), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v0_reg ( .D(n_hpc2_0_N0), .CK(clock_0), .Q(
        n_hpc2_0_n1), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(io_i0_s1), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_2), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v2_reg ( .D(n_hpc2_0_N2), .CK(clock_0), .Q(
        n_hpc2_0_n2), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(p_rand_3), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_0), .QN() );
endmodule

