
module ICINI4 ( port_a_0, port_a_1, port_a_2, port_a_3, port_b_0, port_b_1, 
        port_b_2, port_b_3, port_c_0, port_c_1, port_c_2, port_c_3, 
        port_rand_ref, port_rand_mul_0, port_rand_mul_1, port_rand_mul_2, 
        port_rand_mul_3, port_rand_mul_4, port_rand_mul_5, clk, reset );
  input [4:0] port_a_0;
  input [4:0] port_a_1;
  input [4:0] port_a_2;
  input [4:0] port_a_3;
  input [4:0] port_b_0;
  input [4:0] port_b_1;
  input [4:0] port_b_2;
  input [4:0] port_b_3;
  output [4:0] port_c_0;
  output [4:0] port_c_1;
  output [4:0] port_c_2;
  output [4:0] port_c_3;
  input [11:0] port_rand_ref;
  input [1:0] port_rand_mul_0;
  input [1:0] port_rand_mul_1;
  input [1:0] port_rand_mul_2;
  input [1:0] port_rand_mul_3;
  input [1:0] port_rand_mul_4;
  input [1:0] port_rand_mul_5;
  input clk, reset;
  wire   simpleXor_240_port_a0, simpleXor_240_port_z, simpleXor_241_port_z,
         simpleXor_242_port_a0, simpleXor_242_port_z, simpleXor_243_port_z,
         simpleXor_244_port_a0, simpleXor_244_port_z, simpleXor_245_port_z,
         simpleXor_246_port_a0, simpleXor_246_port_z, simpleXor_247_port_z,
         simpleXor_248_port_a0, simpleXor_248_port_z, simpleXor_249_port_z,
         simpleXor_250_port_a0, simpleXor_250_port_z, simpleXor_251_port_z,
         simpleXor_252_port_a0, simpleXor_252_port_z, simpleXor_253_port_z,
         simpleXor_254_port_a0, simpleXor_254_port_z, simpleXor_255_port_z,
         simpleXor_256_port_a0, simpleXor_256_port_z, simpleXor_257_port_z,
         simpleXor_258_port_a0, simpleXor_258_port_z, simpleXor_259_port_z,
         simpleXor_260_port_a0, simpleXor_260_port_z, simpleXor_261_port_z,
         simpleXor_262_port_a0, simpleXor_262_port_z, simpleXor_263_port_z,
         simpleXor_264_port_a0, simpleXor_264_port_z, simpleXor_265_port_z,
         simpleXor_266_port_a0, simpleXor_266_port_z, simpleXor_267_port_z,
         simpleXor_268_port_a0, simpleXor_268_port_z, simpleXor_269_port_z,
         simpleXor_270_port_a0, simpleXor_270_port_z, simpleXor_271_port_z,
         simpleXor_272_port_a0, simpleXor_272_port_z, simpleXor_273_port_z,
         simpleXor_274_port_a0, simpleXor_274_port_z, simpleXor_275_port_z,
         simpleXor_276_port_a0, simpleXor_276_port_z, simpleXor_277_port_z,
         simpleXor_278_port_a0, simpleXor_278_port_z, simpleXor_279_port_z,
         simpleXor_280_port_a0, simpleXor_280_port_z, simpleXor_281_port_z,
         simpleXor_282_port_a0, simpleXor_282_port_z, simpleXor_283_port_z,
         simpleXor_284_port_a0, simpleXor_284_port_z, simpleXor_285_port_z,
         simpleXor_286_port_a0, simpleXor_286_port_z, simpleXor_287_port_z,
         simpleXor_288_port_a0, simpleXor_288_port_z, simpleXor_289_port_z,
         simpleXor_290_port_a0, simpleXor_290_port_z, simpleXor_291_port_z,
         simpleXor_292_port_a0, simpleXor_292_port_z, simpleXor_293_port_z,
         simpleXor_294_port_a0, simpleXor_294_port_z, simpleXor_295_port_z,
         simpleXor_296_port_a0, simpleXor_296_port_z, simpleXor_297_port_z,
         simpleXor_298_port_a0, simpleXor_298_port_z, simpleXor_299_port_z,
         simpleXor_300_port_a0, simpleXor_300_port_z, simpleXor_301_port_z,
         simpleXor_302_port_a0, simpleXor_302_port_z, simpleXor_303_port_z,
         simpleXor_304_port_a0, simpleXor_304_port_z, simpleXor_305_port_z,
         simpleXor_306_port_a0, simpleXor_306_port_z, simpleXor_307_port_z,
         simpleXor_308_port_a0, simpleXor_308_port_z, simpleXor_309_port_z,
         simpleXor_310_port_a0, simpleXor_310_port_z, simpleXor_311_port_z,
         simpleXor_312_port_a0, simpleXor_312_port_z, simpleXor_313_port_z,
         simpleXor_314_port_a0, simpleXor_314_port_z, simpleXor_315_port_z,
         simpleXor_316_port_a0, simpleXor_316_port_z, simpleXor_317_port_z,
         simpleXor_318_port_a0, simpleXor_318_port_z, simpleXor_319_port_z,
         simpleXor_320_port_a0, simpleXor_320_port_z, simpleXor_321_port_z,
         simpleXor_322_port_a0, simpleXor_322_port_z, simpleXor_323_port_z,
         simpleXor_324_port_a0, simpleXor_324_port_z, simpleXor_325_port_z,
         simpleXor_326_port_a0, simpleXor_326_port_z, simpleXor_327_port_z,
         simpleXor_328_port_a0, simpleXor_328_port_z, simpleXor_329_port_z,
         simpleXor_330_port_a0, simpleXor_330_port_z, simpleXor_331_port_z,
         simpleXor_332_port_a0, simpleXor_332_port_z, simpleXor_333_port_z,
         simpleXor_334_port_a0, simpleXor_334_port_z, simpleXor_335_port_z,
         simpleXor_336_port_a0, simpleXor_336_port_z, simpleXor_337_port_z,
         simpleXor_338_port_a0, simpleXor_338_port_z, simpleXor_339_port_z,
         simpleXor_340_port_a0, simpleXor_340_port_z, simpleXor_341_port_z,
         simpleXor_342_port_a0, simpleXor_342_port_z, simpleXor_343_port_z,
         simpleXor_344_port_a0, simpleXor_344_port_z, simpleXor_345_port_z,
         simpleXor_346_port_a0, simpleXor_346_port_z, simpleXor_347_port_z,
         simpleXor_348_port_a0, simpleXor_348_port_z, simpleXor_349_port_z,
         simpleXor_350_port_a0, simpleXor_350_port_z, simpleXor_351_port_z,
         simpleXor_352_port_a0, simpleXor_352_port_z, simpleXor_353_port_z,
         simpleXor_354_port_a0, simpleXor_354_port_z, simpleXor_355_port_z,
         simpleXor_356_port_a0, simpleXor_356_port_z, simpleXor_357_port_z,
         simpleXor_358_port_a0, simpleXor_358_port_z, simpleXor_359_port_z, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         ref_1_n40, ref_1_n39, ref_1_n38, ref_1_n37, ref_1_n36, ref_1_n35,
         ref_1_n34, ref_1_n33, ref_1_n32, ref_1_n31, ref_1_n30, ref_1_n29,
         ref_1_n28, ref_1_n27, ref_1_n26, ref_1_n25, ref_1_n24, ref_1_n23,
         ref_1_n22, ref_1_n21, ref_1_n20, ref_1_n19, ref_1_n18, ref_1_n17,
         ref_1_n16, ref_1_n15, ref_1_n14, ref_1_n13, ref_1_n12, ref_1_n11,
         ref_1_n10, ref_1_n9, ref_1_n8, ref_1_n7, ref_1_n6, ref_1_n5, ref_1_n4,
         ref_1_n3, ref_1_n2, ref_1_n1, ref_1_maj_159_port_o,
         ref_1_maj_158_port_o, ref_1_maj_157_port_o, ref_1_maj_156_port_o,
         ref_1_maj_155_port_o, ref_1_maj_154_port_o, ref_1_maj_153_port_o,
         ref_1_maj_152_port_o, ref_1_maj_151_port_o, ref_1_maj_150_port_o,
         ref_1_maj_149_port_o, ref_1_maj_148_port_o, ref_1_maj_147_port_o,
         ref_1_maj_146_port_o, ref_1_maj_145_port_o, ref_1_maj_144_port_o,
         ref_1_maj_143_port_o, ref_1_maj_142_port_o, ref_1_maj_141_port_o,
         ref_1_maj_140_port_o, ref_1_maj_139_port_o, ref_1_maj_138_port_o,
         ref_1_maj_137_port_o, ref_1_maj_136_port_o, ref_1_maj_135_port_o,
         ref_1_maj_134_port_o, ref_1_maj_133_port_o, ref_1_maj_132_port_o,
         ref_1_maj_131_port_o, ref_1_maj_130_port_o, ref_1_maj_129_port_o,
         ref_1_maj_128_port_o, ref_1_maj_127_port_o, ref_1_maj_126_port_o,
         ref_1_maj_125_port_o, ref_1_maj_124_port_o, ref_1_maj_123_port_o,
         ref_1_maj_122_port_o, ref_1_maj_121_port_o, ref_1_maj_120_port_o,
         ref_1_maj_119_port_o, ref_1_maj_118_port_o, ref_1_maj_117_port_o,
         ref_1_maj_116_port_o, ref_1_maj_115_port_o, ref_1_maj_114_port_o,
         ref_1_maj_113_port_o, ref_1_maj_112_port_o, ref_1_maj_111_port_o,
         ref_1_maj_110_port_o, ref_1_maj_109_port_o, ref_1_maj_108_port_o,
         ref_1_maj_107_port_o, ref_1_maj_106_port_o, ref_1_maj_105_port_o,
         ref_1_maj_104_port_o, ref_1_maj_103_port_o, ref_1_maj_102_port_o,
         ref_1_maj_101_port_o, ref_1_maj_100_port_o, ref_1_maj_99_port_o,
         ref_1_maj_98_port_o, ref_1_maj_97_port_o, ref_1_maj_96_port_o,
         ref_1_maj_95_port_o, ref_1_maj_94_port_o, ref_1_maj_93_port_o,
         ref_1_maj_92_port_o, ref_1_refreshed_3_0_, ref_1_refreshed_3_1_,
         ref_1_refreshed_3_2_, ref_1_refreshed_3_3_, ref_1_refreshed_3_4_,
         ref_1_maj_91_port_o, ref_1_maj_90_port_o, ref_1_maj_89_port_o,
         ref_1_maj_88_port_o, ref_1_refreshed_2_0_, ref_1_refreshed_2_1_,
         ref_1_refreshed_2_2_, ref_1_refreshed_2_3_, ref_1_refreshed_2_4_,
         ref_1_maj_87_port_o, ref_1_maj_86_port_o, ref_1_maj_85_port_o,
         ref_1_maj_84_port_o, ref_1_refreshed_1_0_, ref_1_refreshed_1_1_,
         ref_1_refreshed_1_2_, ref_1_refreshed_1_3_, ref_1_refreshed_1_4_,
         ref_1_maj_83_port_o, ref_1_maj_82_port_o, ref_1_maj_81_port_o,
         ref_1_maj_80_port_o, ref_1_refreshed_0_0_, ref_1_refreshed_0_1_,
         ref_1_refreshed_0_2_, ref_1_refreshed_0_3_, ref_1_refreshed_0_4_,
         ref_1_simpleXor_358_port_z, ref_1_simpleXor_357_port_z,
         ref_1_simpleXor_356_port_z, ref_1_simpleXor_355_port_z,
         ref_1_simpleXor_354_port_z, ref_1_simpleXor_352_port_z,
         ref_1_simpleXor_351_port_z, ref_1_simpleXor_350_port_z,
         ref_1_simpleXor_349_port_z, ref_1_simpleXor_348_port_z,
         ref_1_simpleXor_346_port_z, ref_1_simpleXor_345_port_z,
         ref_1_simpleXor_344_port_z, ref_1_simpleXor_343_port_z,
         ref_1_simpleXor_342_port_z, ref_1_simpleXor_340_port_z,
         ref_1_simpleXor_339_port_z, ref_1_simpleXor_338_port_z,
         ref_1_simpleXor_337_port_z, ref_1_simpleXor_336_port_z,
         ref_1_simpleXor_334_port_z, ref_1_simpleXor_333_port_z,
         ref_1_simpleXor_332_port_z, ref_1_simpleXor_331_port_z,
         ref_1_simpleXor_330_port_z, ref_1_simpleXor_328_port_z,
         ref_1_simpleXor_327_port_z, ref_1_simpleXor_326_port_z,
         ref_1_simpleXor_325_port_z, ref_1_simpleXor_324_port_z,
         ref_1_simpleXor_322_port_z, ref_1_simpleXor_321_port_z,
         ref_1_simpleXor_320_port_z, ref_1_simpleXor_319_port_z,
         ref_1_simpleXor_318_port_z, ref_1_simpleXor_316_port_z,
         ref_1_simpleXor_315_port_z, ref_1_simpleXor_314_port_z,
         ref_1_simpleXor_313_port_z, ref_1_simpleXor_312_port_z,
         ref_1_simpleXor_310_port_z, ref_1_simpleXor_309_port_z,
         ref_1_simpleXor_308_port_z, ref_1_simpleXor_307_port_z,
         ref_1_simpleXor_306_port_z, ref_1_simpleXor_304_port_z,
         ref_1_simpleXor_303_port_z, ref_1_simpleXor_302_port_z,
         ref_1_simpleXor_301_port_z, ref_1_simpleXor_300_port_z,
         ref_1_simpleXor_298_port_z, ref_1_simpleXor_297_port_z,
         ref_1_simpleXor_296_port_z, ref_1_simpleXor_295_port_z,
         ref_1_simpleXor_294_port_z, ref_1_simpleXor_292_port_z,
         ref_1_simpleXor_291_port_z, ref_1_simpleXor_290_port_z,
         ref_1_simpleXor_289_port_z, ref_1_simpleXor_288_port_z,
         ref_1_simpleXor_286_port_z, ref_1_simpleXor_285_port_z,
         ref_1_simpleXor_284_port_z, ref_1_simpleXor_283_port_z,
         ref_1_simpleXor_282_port_z, ref_1_simpleXor_280_port_z,
         ref_1_simpleXor_279_port_z, ref_1_simpleXor_278_port_z,
         ref_1_simpleXor_277_port_z, ref_1_simpleXor_276_port_z,
         ref_1_simpleXor_274_port_z, ref_1_simpleXor_273_port_z,
         ref_1_simpleXor_272_port_z, ref_1_simpleXor_271_port_z,
         ref_1_simpleXor_270_port_z, ref_1_simpleXor_268_port_z,
         ref_1_simpleXor_267_port_z, ref_1_simpleXor_266_port_z,
         ref_1_simpleXor_265_port_z, ref_1_simpleXor_264_port_z,
         ref_1_simpleXor_262_port_z, ref_1_simpleXor_261_port_z,
         ref_1_simpleXor_260_port_z, ref_1_simpleXor_259_port_z,
         ref_1_simpleXor_258_port_z, ref_1_simpleXor_256_port_z,
         ref_1_simpleXor_255_port_z, ref_1_simpleXor_254_port_z,
         ref_1_simpleXor_253_port_z, ref_1_simpleXor_252_port_z,
         ref_1_simpleXor_250_port_z, ref_1_simpleXor_249_port_z,
         ref_1_simpleXor_248_port_z, ref_1_simpleXor_247_port_z,
         ref_1_simpleXor_246_port_z, ref_1_simpleXor_244_port_z,
         ref_1_simpleXor_243_port_z, ref_1_simpleXor_242_port_z,
         ref_1_simpleXor_241_port_z, ref_1_simpleXor_240_port_z,
         ref_1_maj_80_n13, ref_1_maj_80_n12, ref_1_maj_80_n11,
         ref_1_maj_80_n10, ref_1_maj_80_n9, ref_1_maj_80_n8, ref_1_maj_80_n7,
         ref_1_maj_80_n6, ref_1_maj_80_n5, ref_1_maj_80_n4, ref_1_maj_80_n3,
         ref_1_maj_80_n2, ref_1_maj_80_n1, ref_1_maj_81_n26, ref_1_maj_81_n25,
         ref_1_maj_81_n24, ref_1_maj_81_n23, ref_1_maj_81_n22,
         ref_1_maj_81_n21, ref_1_maj_81_n20, ref_1_maj_81_n19,
         ref_1_maj_81_n18, ref_1_maj_81_n17, ref_1_maj_81_n16,
         ref_1_maj_81_n15, ref_1_maj_81_n14, ref_1_maj_82_n26,
         ref_1_maj_82_n25, ref_1_maj_82_n24, ref_1_maj_82_n23,
         ref_1_maj_82_n22, ref_1_maj_82_n21, ref_1_maj_82_n20,
         ref_1_maj_82_n19, ref_1_maj_82_n18, ref_1_maj_82_n17,
         ref_1_maj_82_n16, ref_1_maj_82_n15, ref_1_maj_82_n14,
         ref_1_maj_83_n26, ref_1_maj_83_n25, ref_1_maj_83_n24,
         ref_1_maj_83_n23, ref_1_maj_83_n22, ref_1_maj_83_n21,
         ref_1_maj_83_n20, ref_1_maj_83_n19, ref_1_maj_83_n18,
         ref_1_maj_83_n17, ref_1_maj_83_n16, ref_1_maj_83_n15,
         ref_1_maj_83_n14, ref_1_maj_84_n26, ref_1_maj_84_n25,
         ref_1_maj_84_n24, ref_1_maj_84_n23, ref_1_maj_84_n22,
         ref_1_maj_84_n21, ref_1_maj_84_n20, ref_1_maj_84_n19,
         ref_1_maj_84_n18, ref_1_maj_84_n17, ref_1_maj_84_n16,
         ref_1_maj_84_n15, ref_1_maj_84_n14, ref_1_maj_85_n26,
         ref_1_maj_85_n25, ref_1_maj_85_n24, ref_1_maj_85_n23,
         ref_1_maj_85_n22, ref_1_maj_85_n21, ref_1_maj_85_n20,
         ref_1_maj_85_n19, ref_1_maj_85_n18, ref_1_maj_85_n17,
         ref_1_maj_85_n16, ref_1_maj_85_n15, ref_1_maj_85_n14,
         ref_1_maj_86_n26, ref_1_maj_86_n25, ref_1_maj_86_n24,
         ref_1_maj_86_n23, ref_1_maj_86_n22, ref_1_maj_86_n21,
         ref_1_maj_86_n20, ref_1_maj_86_n19, ref_1_maj_86_n18,
         ref_1_maj_86_n17, ref_1_maj_86_n16, ref_1_maj_86_n15,
         ref_1_maj_86_n14, ref_1_maj_87_n26, ref_1_maj_87_n25,
         ref_1_maj_87_n24, ref_1_maj_87_n23, ref_1_maj_87_n22,
         ref_1_maj_87_n21, ref_1_maj_87_n20, ref_1_maj_87_n19,
         ref_1_maj_87_n18, ref_1_maj_87_n17, ref_1_maj_87_n16,
         ref_1_maj_87_n15, ref_1_maj_87_n14, ref_1_maj_88_n26,
         ref_1_maj_88_n25, ref_1_maj_88_n24, ref_1_maj_88_n23,
         ref_1_maj_88_n22, ref_1_maj_88_n21, ref_1_maj_88_n20,
         ref_1_maj_88_n19, ref_1_maj_88_n18, ref_1_maj_88_n17,
         ref_1_maj_88_n16, ref_1_maj_88_n15, ref_1_maj_88_n14,
         ref_1_maj_89_n26, ref_1_maj_89_n25, ref_1_maj_89_n24,
         ref_1_maj_89_n23, ref_1_maj_89_n22, ref_1_maj_89_n21,
         ref_1_maj_89_n20, ref_1_maj_89_n19, ref_1_maj_89_n18,
         ref_1_maj_89_n17, ref_1_maj_89_n16, ref_1_maj_89_n15,
         ref_1_maj_89_n14, ref_1_maj_90_n26, ref_1_maj_90_n25,
         ref_1_maj_90_n24, ref_1_maj_90_n23, ref_1_maj_90_n22,
         ref_1_maj_90_n21, ref_1_maj_90_n20, ref_1_maj_90_n19,
         ref_1_maj_90_n18, ref_1_maj_90_n17, ref_1_maj_90_n16,
         ref_1_maj_90_n15, ref_1_maj_90_n14, ref_1_maj_91_n26,
         ref_1_maj_91_n25, ref_1_maj_91_n24, ref_1_maj_91_n23,
         ref_1_maj_91_n22, ref_1_maj_91_n21, ref_1_maj_91_n20,
         ref_1_maj_91_n19, ref_1_maj_91_n18, ref_1_maj_91_n17,
         ref_1_maj_91_n16, ref_1_maj_91_n15, ref_1_maj_91_n14,
         ref_1_maj_92_n26, ref_1_maj_92_n25, ref_1_maj_92_n24,
         ref_1_maj_92_n23, ref_1_maj_92_n22, ref_1_maj_92_n21,
         ref_1_maj_92_n20, ref_1_maj_92_n19, ref_1_maj_92_n18,
         ref_1_maj_92_n17, ref_1_maj_92_n16, ref_1_maj_92_n15,
         ref_1_maj_92_n14, ref_1_maj_93_n26, ref_1_maj_93_n25,
         ref_1_maj_93_n24, ref_1_maj_93_n23, ref_1_maj_93_n22,
         ref_1_maj_93_n21, ref_1_maj_93_n20, ref_1_maj_93_n19,
         ref_1_maj_93_n18, ref_1_maj_93_n17, ref_1_maj_93_n16,
         ref_1_maj_93_n15, ref_1_maj_93_n14, ref_1_maj_94_n26,
         ref_1_maj_94_n25, ref_1_maj_94_n24, ref_1_maj_94_n23,
         ref_1_maj_94_n22, ref_1_maj_94_n21, ref_1_maj_94_n20,
         ref_1_maj_94_n19, ref_1_maj_94_n18, ref_1_maj_94_n17,
         ref_1_maj_94_n16, ref_1_maj_94_n15, ref_1_maj_94_n14,
         ref_1_maj_95_n26, ref_1_maj_95_n25, ref_1_maj_95_n24,
         ref_1_maj_95_n23, ref_1_maj_95_n22, ref_1_maj_95_n21,
         ref_1_maj_95_n20, ref_1_maj_95_n19, ref_1_maj_95_n18,
         ref_1_maj_95_n17, ref_1_maj_95_n16, ref_1_maj_95_n15,
         ref_1_maj_95_n14, ref_1_maj_96_n26, ref_1_maj_96_n25,
         ref_1_maj_96_n24, ref_1_maj_96_n23, ref_1_maj_96_n22,
         ref_1_maj_96_n21, ref_1_maj_96_n20, ref_1_maj_96_n19,
         ref_1_maj_96_n18, ref_1_maj_96_n17, ref_1_maj_96_n16,
         ref_1_maj_96_n15, ref_1_maj_96_n14, ref_1_maj_97_n26,
         ref_1_maj_97_n25, ref_1_maj_97_n24, ref_1_maj_97_n23,
         ref_1_maj_97_n22, ref_1_maj_97_n21, ref_1_maj_97_n20,
         ref_1_maj_97_n19, ref_1_maj_97_n18, ref_1_maj_97_n17,
         ref_1_maj_97_n16, ref_1_maj_97_n15, ref_1_maj_97_n14,
         ref_1_maj_98_n26, ref_1_maj_98_n25, ref_1_maj_98_n24,
         ref_1_maj_98_n23, ref_1_maj_98_n22, ref_1_maj_98_n21,
         ref_1_maj_98_n20, ref_1_maj_98_n19, ref_1_maj_98_n18,
         ref_1_maj_98_n17, ref_1_maj_98_n16, ref_1_maj_98_n15,
         ref_1_maj_98_n14, ref_1_maj_99_n26, ref_1_maj_99_n25,
         ref_1_maj_99_n24, ref_1_maj_99_n23, ref_1_maj_99_n22,
         ref_1_maj_99_n21, ref_1_maj_99_n20, ref_1_maj_99_n19,
         ref_1_maj_99_n18, ref_1_maj_99_n17, ref_1_maj_99_n16,
         ref_1_maj_99_n15, ref_1_maj_99_n14, ref_1_maj_100_n26,
         ref_1_maj_100_n25, ref_1_maj_100_n24, ref_1_maj_100_n23,
         ref_1_maj_100_n22, ref_1_maj_100_n21, ref_1_maj_100_n20,
         ref_1_maj_100_n19, ref_1_maj_100_n18, ref_1_maj_100_n17,
         ref_1_maj_100_n16, ref_1_maj_100_n15, ref_1_maj_100_n14,
         ref_1_maj_101_n26, ref_1_maj_101_n25, ref_1_maj_101_n24,
         ref_1_maj_101_n23, ref_1_maj_101_n22, ref_1_maj_101_n21,
         ref_1_maj_101_n20, ref_1_maj_101_n19, ref_1_maj_101_n18,
         ref_1_maj_101_n17, ref_1_maj_101_n16, ref_1_maj_101_n15,
         ref_1_maj_101_n14, ref_1_maj_102_n26, ref_1_maj_102_n25,
         ref_1_maj_102_n24, ref_1_maj_102_n23, ref_1_maj_102_n22,
         ref_1_maj_102_n21, ref_1_maj_102_n20, ref_1_maj_102_n19,
         ref_1_maj_102_n18, ref_1_maj_102_n17, ref_1_maj_102_n16,
         ref_1_maj_102_n15, ref_1_maj_102_n14, ref_1_maj_103_n26,
         ref_1_maj_103_n25, ref_1_maj_103_n24, ref_1_maj_103_n23,
         ref_1_maj_103_n22, ref_1_maj_103_n21, ref_1_maj_103_n20,
         ref_1_maj_103_n19, ref_1_maj_103_n18, ref_1_maj_103_n17,
         ref_1_maj_103_n16, ref_1_maj_103_n15, ref_1_maj_103_n14,
         ref_1_maj_104_n26, ref_1_maj_104_n25, ref_1_maj_104_n24,
         ref_1_maj_104_n23, ref_1_maj_104_n22, ref_1_maj_104_n21,
         ref_1_maj_104_n20, ref_1_maj_104_n19, ref_1_maj_104_n18,
         ref_1_maj_104_n17, ref_1_maj_104_n16, ref_1_maj_104_n15,
         ref_1_maj_104_n14, ref_1_maj_105_n26, ref_1_maj_105_n25,
         ref_1_maj_105_n24, ref_1_maj_105_n23, ref_1_maj_105_n22,
         ref_1_maj_105_n21, ref_1_maj_105_n20, ref_1_maj_105_n19,
         ref_1_maj_105_n18, ref_1_maj_105_n17, ref_1_maj_105_n16,
         ref_1_maj_105_n15, ref_1_maj_105_n14, ref_1_maj_106_n26,
         ref_1_maj_106_n25, ref_1_maj_106_n24, ref_1_maj_106_n23,
         ref_1_maj_106_n22, ref_1_maj_106_n21, ref_1_maj_106_n20,
         ref_1_maj_106_n19, ref_1_maj_106_n18, ref_1_maj_106_n17,
         ref_1_maj_106_n16, ref_1_maj_106_n15, ref_1_maj_106_n14,
         ref_1_maj_107_n26, ref_1_maj_107_n25, ref_1_maj_107_n24,
         ref_1_maj_107_n23, ref_1_maj_107_n22, ref_1_maj_107_n21,
         ref_1_maj_107_n20, ref_1_maj_107_n19, ref_1_maj_107_n18,
         ref_1_maj_107_n17, ref_1_maj_107_n16, ref_1_maj_107_n15,
         ref_1_maj_107_n14, ref_1_maj_108_n26, ref_1_maj_108_n25,
         ref_1_maj_108_n24, ref_1_maj_108_n23, ref_1_maj_108_n22,
         ref_1_maj_108_n21, ref_1_maj_108_n20, ref_1_maj_108_n19,
         ref_1_maj_108_n18, ref_1_maj_108_n17, ref_1_maj_108_n16,
         ref_1_maj_108_n15, ref_1_maj_108_n14, ref_1_maj_109_n26,
         ref_1_maj_109_n25, ref_1_maj_109_n24, ref_1_maj_109_n23,
         ref_1_maj_109_n22, ref_1_maj_109_n21, ref_1_maj_109_n20,
         ref_1_maj_109_n19, ref_1_maj_109_n18, ref_1_maj_109_n17,
         ref_1_maj_109_n16, ref_1_maj_109_n15, ref_1_maj_109_n14,
         ref_1_maj_110_n26, ref_1_maj_110_n25, ref_1_maj_110_n24,
         ref_1_maj_110_n23, ref_1_maj_110_n22, ref_1_maj_110_n21,
         ref_1_maj_110_n20, ref_1_maj_110_n19, ref_1_maj_110_n18,
         ref_1_maj_110_n17, ref_1_maj_110_n16, ref_1_maj_110_n15,
         ref_1_maj_110_n14, ref_1_maj_111_n26, ref_1_maj_111_n25,
         ref_1_maj_111_n24, ref_1_maj_111_n23, ref_1_maj_111_n22,
         ref_1_maj_111_n21, ref_1_maj_111_n20, ref_1_maj_111_n19,
         ref_1_maj_111_n18, ref_1_maj_111_n17, ref_1_maj_111_n16,
         ref_1_maj_111_n15, ref_1_maj_111_n14, ref_1_maj_112_n26,
         ref_1_maj_112_n25, ref_1_maj_112_n24, ref_1_maj_112_n23,
         ref_1_maj_112_n22, ref_1_maj_112_n21, ref_1_maj_112_n20,
         ref_1_maj_112_n19, ref_1_maj_112_n18, ref_1_maj_112_n17,
         ref_1_maj_112_n16, ref_1_maj_112_n15, ref_1_maj_112_n14,
         ref_1_maj_113_n26, ref_1_maj_113_n25, ref_1_maj_113_n24,
         ref_1_maj_113_n23, ref_1_maj_113_n22, ref_1_maj_113_n21,
         ref_1_maj_113_n20, ref_1_maj_113_n19, ref_1_maj_113_n18,
         ref_1_maj_113_n17, ref_1_maj_113_n16, ref_1_maj_113_n15,
         ref_1_maj_113_n14, ref_1_maj_114_n26, ref_1_maj_114_n25,
         ref_1_maj_114_n24, ref_1_maj_114_n23, ref_1_maj_114_n22,
         ref_1_maj_114_n21, ref_1_maj_114_n20, ref_1_maj_114_n19,
         ref_1_maj_114_n18, ref_1_maj_114_n17, ref_1_maj_114_n16,
         ref_1_maj_114_n15, ref_1_maj_114_n14, ref_1_maj_115_n26,
         ref_1_maj_115_n25, ref_1_maj_115_n24, ref_1_maj_115_n23,
         ref_1_maj_115_n22, ref_1_maj_115_n21, ref_1_maj_115_n20,
         ref_1_maj_115_n19, ref_1_maj_115_n18, ref_1_maj_115_n17,
         ref_1_maj_115_n16, ref_1_maj_115_n15, ref_1_maj_115_n14,
         ref_1_maj_116_n26, ref_1_maj_116_n25, ref_1_maj_116_n24,
         ref_1_maj_116_n23, ref_1_maj_116_n22, ref_1_maj_116_n21,
         ref_1_maj_116_n20, ref_1_maj_116_n19, ref_1_maj_116_n18,
         ref_1_maj_116_n17, ref_1_maj_116_n16, ref_1_maj_116_n15,
         ref_1_maj_116_n14, ref_1_maj_117_n26, ref_1_maj_117_n25,
         ref_1_maj_117_n24, ref_1_maj_117_n23, ref_1_maj_117_n22,
         ref_1_maj_117_n21, ref_1_maj_117_n20, ref_1_maj_117_n19,
         ref_1_maj_117_n18, ref_1_maj_117_n17, ref_1_maj_117_n16,
         ref_1_maj_117_n15, ref_1_maj_117_n14, ref_1_maj_118_n26,
         ref_1_maj_118_n25, ref_1_maj_118_n24, ref_1_maj_118_n23,
         ref_1_maj_118_n22, ref_1_maj_118_n21, ref_1_maj_118_n20,
         ref_1_maj_118_n19, ref_1_maj_118_n18, ref_1_maj_118_n17,
         ref_1_maj_118_n16, ref_1_maj_118_n15, ref_1_maj_118_n14,
         ref_1_maj_119_n26, ref_1_maj_119_n25, ref_1_maj_119_n24,
         ref_1_maj_119_n23, ref_1_maj_119_n22, ref_1_maj_119_n21,
         ref_1_maj_119_n20, ref_1_maj_119_n19, ref_1_maj_119_n18,
         ref_1_maj_119_n17, ref_1_maj_119_n16, ref_1_maj_119_n15,
         ref_1_maj_119_n14, ref_1_maj_120_n26, ref_1_maj_120_n25,
         ref_1_maj_120_n24, ref_1_maj_120_n23, ref_1_maj_120_n22,
         ref_1_maj_120_n21, ref_1_maj_120_n20, ref_1_maj_120_n19,
         ref_1_maj_120_n18, ref_1_maj_120_n17, ref_1_maj_120_n16,
         ref_1_maj_120_n15, ref_1_maj_120_n14, ref_1_maj_121_n26,
         ref_1_maj_121_n25, ref_1_maj_121_n24, ref_1_maj_121_n23,
         ref_1_maj_121_n22, ref_1_maj_121_n21, ref_1_maj_121_n20,
         ref_1_maj_121_n19, ref_1_maj_121_n18, ref_1_maj_121_n17,
         ref_1_maj_121_n16, ref_1_maj_121_n15, ref_1_maj_121_n14,
         ref_1_maj_122_n26, ref_1_maj_122_n25, ref_1_maj_122_n24,
         ref_1_maj_122_n23, ref_1_maj_122_n22, ref_1_maj_122_n21,
         ref_1_maj_122_n20, ref_1_maj_122_n19, ref_1_maj_122_n18,
         ref_1_maj_122_n17, ref_1_maj_122_n16, ref_1_maj_122_n15,
         ref_1_maj_122_n14, ref_1_maj_123_n26, ref_1_maj_123_n25,
         ref_1_maj_123_n24, ref_1_maj_123_n23, ref_1_maj_123_n22,
         ref_1_maj_123_n21, ref_1_maj_123_n20, ref_1_maj_123_n19,
         ref_1_maj_123_n18, ref_1_maj_123_n17, ref_1_maj_123_n16,
         ref_1_maj_123_n15, ref_1_maj_123_n14, ref_1_maj_124_n26,
         ref_1_maj_124_n25, ref_1_maj_124_n24, ref_1_maj_124_n23,
         ref_1_maj_124_n22, ref_1_maj_124_n21, ref_1_maj_124_n20,
         ref_1_maj_124_n19, ref_1_maj_124_n18, ref_1_maj_124_n17,
         ref_1_maj_124_n16, ref_1_maj_124_n15, ref_1_maj_124_n14,
         ref_1_maj_125_n26, ref_1_maj_125_n25, ref_1_maj_125_n24,
         ref_1_maj_125_n23, ref_1_maj_125_n22, ref_1_maj_125_n21,
         ref_1_maj_125_n20, ref_1_maj_125_n19, ref_1_maj_125_n18,
         ref_1_maj_125_n17, ref_1_maj_125_n16, ref_1_maj_125_n15,
         ref_1_maj_125_n14, ref_1_maj_126_n26, ref_1_maj_126_n25,
         ref_1_maj_126_n24, ref_1_maj_126_n23, ref_1_maj_126_n22,
         ref_1_maj_126_n21, ref_1_maj_126_n20, ref_1_maj_126_n19,
         ref_1_maj_126_n18, ref_1_maj_126_n17, ref_1_maj_126_n16,
         ref_1_maj_126_n15, ref_1_maj_126_n14, ref_1_maj_127_n26,
         ref_1_maj_127_n25, ref_1_maj_127_n24, ref_1_maj_127_n23,
         ref_1_maj_127_n22, ref_1_maj_127_n21, ref_1_maj_127_n20,
         ref_1_maj_127_n19, ref_1_maj_127_n18, ref_1_maj_127_n17,
         ref_1_maj_127_n16, ref_1_maj_127_n15, ref_1_maj_127_n14,
         ref_1_maj_128_n26, ref_1_maj_128_n25, ref_1_maj_128_n24,
         ref_1_maj_128_n23, ref_1_maj_128_n22, ref_1_maj_128_n21,
         ref_1_maj_128_n20, ref_1_maj_128_n19, ref_1_maj_128_n18,
         ref_1_maj_128_n17, ref_1_maj_128_n16, ref_1_maj_128_n15,
         ref_1_maj_128_n14, ref_1_maj_129_n26, ref_1_maj_129_n25,
         ref_1_maj_129_n24, ref_1_maj_129_n23, ref_1_maj_129_n22,
         ref_1_maj_129_n21, ref_1_maj_129_n20, ref_1_maj_129_n19,
         ref_1_maj_129_n18, ref_1_maj_129_n17, ref_1_maj_129_n16,
         ref_1_maj_129_n15, ref_1_maj_129_n14, ref_1_maj_130_n26,
         ref_1_maj_130_n25, ref_1_maj_130_n24, ref_1_maj_130_n23,
         ref_1_maj_130_n22, ref_1_maj_130_n21, ref_1_maj_130_n20,
         ref_1_maj_130_n19, ref_1_maj_130_n18, ref_1_maj_130_n17,
         ref_1_maj_130_n16, ref_1_maj_130_n15, ref_1_maj_130_n14,
         ref_1_maj_131_n26, ref_1_maj_131_n25, ref_1_maj_131_n24,
         ref_1_maj_131_n23, ref_1_maj_131_n22, ref_1_maj_131_n21,
         ref_1_maj_131_n20, ref_1_maj_131_n19, ref_1_maj_131_n18,
         ref_1_maj_131_n17, ref_1_maj_131_n16, ref_1_maj_131_n15,
         ref_1_maj_131_n14, ref_1_maj_132_n26, ref_1_maj_132_n25,
         ref_1_maj_132_n24, ref_1_maj_132_n23, ref_1_maj_132_n22,
         ref_1_maj_132_n21, ref_1_maj_132_n20, ref_1_maj_132_n19,
         ref_1_maj_132_n18, ref_1_maj_132_n17, ref_1_maj_132_n16,
         ref_1_maj_132_n15, ref_1_maj_132_n14, ref_1_maj_133_n26,
         ref_1_maj_133_n25, ref_1_maj_133_n24, ref_1_maj_133_n23,
         ref_1_maj_133_n22, ref_1_maj_133_n21, ref_1_maj_133_n20,
         ref_1_maj_133_n19, ref_1_maj_133_n18, ref_1_maj_133_n17,
         ref_1_maj_133_n16, ref_1_maj_133_n15, ref_1_maj_133_n14,
         ref_1_maj_134_n26, ref_1_maj_134_n25, ref_1_maj_134_n24,
         ref_1_maj_134_n23, ref_1_maj_134_n22, ref_1_maj_134_n21,
         ref_1_maj_134_n20, ref_1_maj_134_n19, ref_1_maj_134_n18,
         ref_1_maj_134_n17, ref_1_maj_134_n16, ref_1_maj_134_n15,
         ref_1_maj_134_n14, ref_1_maj_135_n26, ref_1_maj_135_n25,
         ref_1_maj_135_n24, ref_1_maj_135_n23, ref_1_maj_135_n22,
         ref_1_maj_135_n21, ref_1_maj_135_n20, ref_1_maj_135_n19,
         ref_1_maj_135_n18, ref_1_maj_135_n17, ref_1_maj_135_n16,
         ref_1_maj_135_n15, ref_1_maj_135_n14, ref_1_maj_136_n26,
         ref_1_maj_136_n25, ref_1_maj_136_n24, ref_1_maj_136_n23,
         ref_1_maj_136_n22, ref_1_maj_136_n21, ref_1_maj_136_n20,
         ref_1_maj_136_n19, ref_1_maj_136_n18, ref_1_maj_136_n17,
         ref_1_maj_136_n16, ref_1_maj_136_n15, ref_1_maj_136_n14,
         ref_1_maj_137_n26, ref_1_maj_137_n25, ref_1_maj_137_n24,
         ref_1_maj_137_n23, ref_1_maj_137_n22, ref_1_maj_137_n21,
         ref_1_maj_137_n20, ref_1_maj_137_n19, ref_1_maj_137_n18,
         ref_1_maj_137_n17, ref_1_maj_137_n16, ref_1_maj_137_n15,
         ref_1_maj_137_n14, ref_1_maj_138_n26, ref_1_maj_138_n25,
         ref_1_maj_138_n24, ref_1_maj_138_n23, ref_1_maj_138_n22,
         ref_1_maj_138_n21, ref_1_maj_138_n20, ref_1_maj_138_n19,
         ref_1_maj_138_n18, ref_1_maj_138_n17, ref_1_maj_138_n16,
         ref_1_maj_138_n15, ref_1_maj_138_n14, ref_1_maj_139_n26,
         ref_1_maj_139_n25, ref_1_maj_139_n24, ref_1_maj_139_n23,
         ref_1_maj_139_n22, ref_1_maj_139_n21, ref_1_maj_139_n20,
         ref_1_maj_139_n19, ref_1_maj_139_n18, ref_1_maj_139_n17,
         ref_1_maj_139_n16, ref_1_maj_139_n15, ref_1_maj_139_n14,
         ref_1_maj_140_n26, ref_1_maj_140_n25, ref_1_maj_140_n24,
         ref_1_maj_140_n23, ref_1_maj_140_n22, ref_1_maj_140_n21,
         ref_1_maj_140_n20, ref_1_maj_140_n19, ref_1_maj_140_n18,
         ref_1_maj_140_n17, ref_1_maj_140_n16, ref_1_maj_140_n15,
         ref_1_maj_140_n14, ref_1_maj_141_n26, ref_1_maj_141_n25,
         ref_1_maj_141_n24, ref_1_maj_141_n23, ref_1_maj_141_n22,
         ref_1_maj_141_n21, ref_1_maj_141_n20, ref_1_maj_141_n19,
         ref_1_maj_141_n18, ref_1_maj_141_n17, ref_1_maj_141_n16,
         ref_1_maj_141_n15, ref_1_maj_141_n14, ref_1_maj_142_n26,
         ref_1_maj_142_n25, ref_1_maj_142_n24, ref_1_maj_142_n23,
         ref_1_maj_142_n22, ref_1_maj_142_n21, ref_1_maj_142_n20,
         ref_1_maj_142_n19, ref_1_maj_142_n18, ref_1_maj_142_n17,
         ref_1_maj_142_n16, ref_1_maj_142_n15, ref_1_maj_142_n14,
         ref_1_maj_143_n26, ref_1_maj_143_n25, ref_1_maj_143_n24,
         ref_1_maj_143_n23, ref_1_maj_143_n22, ref_1_maj_143_n21,
         ref_1_maj_143_n20, ref_1_maj_143_n19, ref_1_maj_143_n18,
         ref_1_maj_143_n17, ref_1_maj_143_n16, ref_1_maj_143_n15,
         ref_1_maj_143_n14, ref_1_maj_144_n26, ref_1_maj_144_n25,
         ref_1_maj_144_n24, ref_1_maj_144_n23, ref_1_maj_144_n22,
         ref_1_maj_144_n21, ref_1_maj_144_n20, ref_1_maj_144_n19,
         ref_1_maj_144_n18, ref_1_maj_144_n17, ref_1_maj_144_n16,
         ref_1_maj_144_n15, ref_1_maj_144_n14, ref_1_maj_145_n26,
         ref_1_maj_145_n25, ref_1_maj_145_n24, ref_1_maj_145_n23,
         ref_1_maj_145_n22, ref_1_maj_145_n21, ref_1_maj_145_n20,
         ref_1_maj_145_n19, ref_1_maj_145_n18, ref_1_maj_145_n17,
         ref_1_maj_145_n16, ref_1_maj_145_n15, ref_1_maj_145_n14,
         ref_1_maj_146_n26, ref_1_maj_146_n25, ref_1_maj_146_n24,
         ref_1_maj_146_n23, ref_1_maj_146_n22, ref_1_maj_146_n21,
         ref_1_maj_146_n20, ref_1_maj_146_n19, ref_1_maj_146_n18,
         ref_1_maj_146_n17, ref_1_maj_146_n16, ref_1_maj_146_n15,
         ref_1_maj_146_n14, ref_1_maj_147_n26, ref_1_maj_147_n25,
         ref_1_maj_147_n24, ref_1_maj_147_n23, ref_1_maj_147_n22,
         ref_1_maj_147_n21, ref_1_maj_147_n20, ref_1_maj_147_n19,
         ref_1_maj_147_n18, ref_1_maj_147_n17, ref_1_maj_147_n16,
         ref_1_maj_147_n15, ref_1_maj_147_n14, ref_1_maj_148_n26,
         ref_1_maj_148_n25, ref_1_maj_148_n24, ref_1_maj_148_n23,
         ref_1_maj_148_n22, ref_1_maj_148_n21, ref_1_maj_148_n20,
         ref_1_maj_148_n19, ref_1_maj_148_n18, ref_1_maj_148_n17,
         ref_1_maj_148_n16, ref_1_maj_148_n15, ref_1_maj_148_n14,
         ref_1_maj_149_n26, ref_1_maj_149_n25, ref_1_maj_149_n24,
         ref_1_maj_149_n23, ref_1_maj_149_n22, ref_1_maj_149_n21,
         ref_1_maj_149_n20, ref_1_maj_149_n19, ref_1_maj_149_n18,
         ref_1_maj_149_n17, ref_1_maj_149_n16, ref_1_maj_149_n15,
         ref_1_maj_149_n14, ref_1_maj_150_n26, ref_1_maj_150_n25,
         ref_1_maj_150_n24, ref_1_maj_150_n23, ref_1_maj_150_n22,
         ref_1_maj_150_n21, ref_1_maj_150_n20, ref_1_maj_150_n19,
         ref_1_maj_150_n18, ref_1_maj_150_n17, ref_1_maj_150_n16,
         ref_1_maj_150_n15, ref_1_maj_150_n14, ref_1_maj_151_n26,
         ref_1_maj_151_n25, ref_1_maj_151_n24, ref_1_maj_151_n23,
         ref_1_maj_151_n22, ref_1_maj_151_n21, ref_1_maj_151_n20,
         ref_1_maj_151_n19, ref_1_maj_151_n18, ref_1_maj_151_n17,
         ref_1_maj_151_n16, ref_1_maj_151_n15, ref_1_maj_151_n14,
         ref_1_maj_152_n26, ref_1_maj_152_n25, ref_1_maj_152_n24,
         ref_1_maj_152_n23, ref_1_maj_152_n22, ref_1_maj_152_n21,
         ref_1_maj_152_n20, ref_1_maj_152_n19, ref_1_maj_152_n18,
         ref_1_maj_152_n17, ref_1_maj_152_n16, ref_1_maj_152_n15,
         ref_1_maj_152_n14, ref_1_maj_153_n26, ref_1_maj_153_n25,
         ref_1_maj_153_n24, ref_1_maj_153_n23, ref_1_maj_153_n22,
         ref_1_maj_153_n21, ref_1_maj_153_n20, ref_1_maj_153_n19,
         ref_1_maj_153_n18, ref_1_maj_153_n17, ref_1_maj_153_n16,
         ref_1_maj_153_n15, ref_1_maj_153_n14, ref_1_maj_154_n26,
         ref_1_maj_154_n25, ref_1_maj_154_n24, ref_1_maj_154_n23,
         ref_1_maj_154_n22, ref_1_maj_154_n21, ref_1_maj_154_n20,
         ref_1_maj_154_n19, ref_1_maj_154_n18, ref_1_maj_154_n17,
         ref_1_maj_154_n16, ref_1_maj_154_n15, ref_1_maj_154_n14,
         ref_1_maj_155_n26, ref_1_maj_155_n25, ref_1_maj_155_n24,
         ref_1_maj_155_n23, ref_1_maj_155_n22, ref_1_maj_155_n21,
         ref_1_maj_155_n20, ref_1_maj_155_n19, ref_1_maj_155_n18,
         ref_1_maj_155_n17, ref_1_maj_155_n16, ref_1_maj_155_n15,
         ref_1_maj_155_n14, ref_1_maj_156_n26, ref_1_maj_156_n25,
         ref_1_maj_156_n24, ref_1_maj_156_n23, ref_1_maj_156_n22,
         ref_1_maj_156_n21, ref_1_maj_156_n20, ref_1_maj_156_n19,
         ref_1_maj_156_n18, ref_1_maj_156_n17, ref_1_maj_156_n16,
         ref_1_maj_156_n15, ref_1_maj_156_n14, ref_1_maj_157_n26,
         ref_1_maj_157_n25, ref_1_maj_157_n24, ref_1_maj_157_n23,
         ref_1_maj_157_n22, ref_1_maj_157_n21, ref_1_maj_157_n20,
         ref_1_maj_157_n19, ref_1_maj_157_n18, ref_1_maj_157_n17,
         ref_1_maj_157_n16, ref_1_maj_157_n15, ref_1_maj_157_n14,
         ref_1_maj_158_n26, ref_1_maj_158_n25, ref_1_maj_158_n24,
         ref_1_maj_158_n23, ref_1_maj_158_n22, ref_1_maj_158_n21,
         ref_1_maj_158_n20, ref_1_maj_158_n19, ref_1_maj_158_n18,
         ref_1_maj_158_n17, ref_1_maj_158_n16, ref_1_maj_158_n15,
         ref_1_maj_158_n14, ref_1_maj_159_n26, ref_1_maj_159_n25,
         ref_1_maj_159_n24, ref_1_maj_159_n23, ref_1_maj_159_n22,
         ref_1_maj_159_n21, ref_1_maj_159_n20, ref_1_maj_159_n19,
         ref_1_maj_159_n18, ref_1_maj_159_n17, ref_1_maj_159_n16,
         ref_1_maj_159_n15, ref_1_maj_159_n14;
  wire   [4:0] ref_1_port_o_0_0;
  wire   [4:0] ref_1_port_o_0_1;
  wire   [4:0] ref_1_port_o_0_2;
  wire   [4:0] ref_1_port_o_0_3;
  wire   [4:0] ref_1_port_o_1_0;
  wire   [4:0] ref_1_port_o_1_1;
  wire   [4:0] ref_1_port_o_1_2;
  wire   [4:0] ref_1_port_o_1_3;
  wire   [4:0] ref_1_port_o_2_0;
  wire   [4:0] ref_1_port_o_2_1;
  wire   [4:0] ref_1_port_o_2_2;
  wire   [4:0] ref_1_port_o_2_3;
  wire   [4:0] ref_1_port_o_3_0;
  wire   [4:0] ref_1_port_o_3_1;
  wire   [4:0] ref_1_port_o_3_2;
  wire   [4:0] ref_1_port_o_3_3;
  wire   [4:0] temp_0_0;
  wire   [4:0] mult_ab_0_1;
  wire   [4:0] mult_ab_0_2;
  wire   [4:0] mult_ab_0_3;
  wire   [4:0] temp_0_1;
  wire   [4:0] mult_ab_1_0;
  wire   [4:0] mult_ab_1_2;
  wire   [4:0] mult_ab_1_3;
  wire   [4:0] temp_0_2;
  wire   [4:0] mult_ab_2_0;
  wire   [4:0] mult_ab_2_1;
  wire   [4:0] mult_ab_2_3;
  wire   [4:0] temp_0_3;
  wire   [4:0] mult_ab_3_0;
  wire   [4:0] mult_ab_3_1;
  wire   [4:0] mult_ab_3_2;

  DFF_X1 mult_ab_3_2_reg_4_ ( .D(simpleXor_359_port_z), .CK(clk), .Q(
        mult_ab_3_2[4]), .QN() );
  DFF_X1 mult_ab_3_2_reg_3_ ( .D(simpleXor_335_port_z), .CK(clk), .Q(
        mult_ab_3_2[3]), .QN() );
  DFF_X1 mult_ab_3_2_reg_2_ ( .D(simpleXor_311_port_z), .CK(clk), .Q(
        mult_ab_3_2[2]), .QN() );
  DFF_X1 mult_ab_3_2_reg_1_ ( .D(simpleXor_287_port_z), .CK(clk), .Q(
        mult_ab_3_2[1]), .QN() );
  DFF_X1 mult_ab_3_2_reg_0_ ( .D(simpleXor_263_port_z), .CK(clk), .Q(
        mult_ab_3_2[0]), .QN() );
  DFF_X1 mult_ab_3_3_reg_4_ ( .D(N19), .CK(clk), .Q(temp_0_3[4]), .QN() );
  DFF_X1 mult_ab_3_3_reg_3_ ( .D(N15), .CK(clk), .Q(temp_0_3[3]), .QN() );
  DFF_X1 mult_ab_3_3_reg_2_ ( .D(N11), .CK(clk), .Q(temp_0_3[2]), .QN() );
  DFF_X1 mult_ab_3_3_reg_1_ ( .D(N7), .CK(clk), .Q(temp_0_3[1]), .QN() );
  DFF_X1 mult_ab_3_3_reg_0_ ( .D(N3), .CK(clk), .Q(temp_0_3[0]), .QN() );
  DFF_X1 mult_ab_3_0_reg_4_ ( .D(simpleXor_355_port_z), .CK(clk), .Q(
        mult_ab_3_0[4]), .QN() );
  DFF_X1 mult_ab_3_0_reg_3_ ( .D(simpleXor_331_port_z), .CK(clk), .Q(
        mult_ab_3_0[3]), .QN() );
  DFF_X1 mult_ab_3_0_reg_2_ ( .D(simpleXor_307_port_z), .CK(clk), .Q(
        mult_ab_3_0[2]), .QN() );
  DFF_X1 mult_ab_3_0_reg_1_ ( .D(simpleXor_283_port_z), .CK(clk), .Q(
        mult_ab_3_0[1]), .QN() );
  DFF_X1 mult_ab_3_0_reg_0_ ( .D(simpleXor_259_port_z), .CK(clk), .Q(
        mult_ab_3_0[0]), .QN() );
  DFF_X1 mult_ab_3_1_reg_4_ ( .D(simpleXor_357_port_z), .CK(clk), .Q(
        mult_ab_3_1[4]), .QN() );
  DFF_X1 mult_ab_3_1_reg_3_ ( .D(simpleXor_333_port_z), .CK(clk), .Q(
        mult_ab_3_1[3]), .QN() );
  DFF_X1 mult_ab_3_1_reg_2_ ( .D(simpleXor_309_port_z), .CK(clk), .Q(
        mult_ab_3_1[2]), .QN() );
  DFF_X1 mult_ab_3_1_reg_1_ ( .D(simpleXor_285_port_z), .CK(clk), .Q(
        mult_ab_3_1[1]), .QN() );
  DFF_X1 mult_ab_3_1_reg_0_ ( .D(simpleXor_261_port_z), .CK(clk), .Q(
        mult_ab_3_1[0]), .QN() );
  DFF_X1 mult_ab_2_2_reg_4_ ( .D(N18), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 mult_ab_2_2_reg_3_ ( .D(N14), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 mult_ab_2_2_reg_2_ ( .D(N10), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 mult_ab_2_2_reg_1_ ( .D(N6), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 mult_ab_2_2_reg_0_ ( .D(N2), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 mult_ab_2_3_reg_4_ ( .D(simpleXor_353_port_z), .CK(clk), .Q(
        mult_ab_2_3[4]), .QN() );
  DFF_X1 mult_ab_2_3_reg_3_ ( .D(simpleXor_329_port_z), .CK(clk), .Q(
        mult_ab_2_3[3]), .QN() );
  DFF_X1 mult_ab_2_3_reg_2_ ( .D(simpleXor_305_port_z), .CK(clk), .Q(
        mult_ab_2_3[2]), .QN() );
  DFF_X1 mult_ab_2_3_reg_1_ ( .D(simpleXor_281_port_z), .CK(clk), .Q(
        mult_ab_2_3[1]), .QN() );
  DFF_X1 mult_ab_2_3_reg_0_ ( .D(simpleXor_257_port_z), .CK(clk), .Q(
        mult_ab_2_3[0]), .QN() );
  DFF_X1 mult_ab_2_0_reg_4_ ( .D(simpleXor_349_port_z), .CK(clk), .Q(
        mult_ab_2_0[4]), .QN() );
  DFF_X1 mult_ab_2_0_reg_3_ ( .D(simpleXor_325_port_z), .CK(clk), .Q(
        mult_ab_2_0[3]), .QN() );
  DFF_X1 mult_ab_2_0_reg_2_ ( .D(simpleXor_301_port_z), .CK(clk), .Q(
        mult_ab_2_0[2]), .QN() );
  DFF_X1 mult_ab_2_0_reg_1_ ( .D(simpleXor_277_port_z), .CK(clk), .Q(
        mult_ab_2_0[1]), .QN() );
  DFF_X1 mult_ab_2_0_reg_0_ ( .D(simpleXor_253_port_z), .CK(clk), .Q(
        mult_ab_2_0[0]), .QN() );
  DFF_X1 mult_ab_2_1_reg_4_ ( .D(simpleXor_351_port_z), .CK(clk), .Q(
        mult_ab_2_1[4]), .QN() );
  DFF_X1 mult_ab_2_1_reg_3_ ( .D(simpleXor_327_port_z), .CK(clk), .Q(
        mult_ab_2_1[3]), .QN() );
  DFF_X1 mult_ab_2_1_reg_2_ ( .D(simpleXor_303_port_z), .CK(clk), .Q(
        mult_ab_2_1[2]), .QN() );
  DFF_X1 mult_ab_2_1_reg_1_ ( .D(simpleXor_279_port_z), .CK(clk), .Q(
        mult_ab_2_1[1]), .QN() );
  DFF_X1 mult_ab_2_1_reg_0_ ( .D(simpleXor_255_port_z), .CK(clk), .Q(
        mult_ab_2_1[0]), .QN() );
  DFF_X1 mult_ab_0_0_reg_4_ ( .D(N16), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 mult_ab_0_0_reg_3_ ( .D(N12), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 mult_ab_0_0_reg_2_ ( .D(N8), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 mult_ab_0_0_reg_1_ ( .D(N4), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 mult_ab_0_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 mult_ab_0_1_reg_4_ ( .D(simpleXor_337_port_z), .CK(clk), .Q(
        mult_ab_0_1[4]), .QN() );
  DFF_X1 mult_ab_0_1_reg_3_ ( .D(simpleXor_313_port_z), .CK(clk), .Q(
        mult_ab_0_1[3]), .QN() );
  DFF_X1 mult_ab_0_1_reg_2_ ( .D(simpleXor_289_port_z), .CK(clk), .Q(
        mult_ab_0_1[2]), .QN() );
  DFF_X1 mult_ab_0_1_reg_1_ ( .D(simpleXor_265_port_z), .CK(clk), .Q(
        mult_ab_0_1[1]), .QN() );
  DFF_X1 mult_ab_0_1_reg_0_ ( .D(simpleXor_241_port_z), .CK(clk), .Q(
        mult_ab_0_1[0]), .QN() );
  DFF_X1 mult_ab_0_2_reg_4_ ( .D(simpleXor_339_port_z), .CK(clk), .Q(
        mult_ab_0_2[4]), .QN() );
  DFF_X1 mult_ab_0_2_reg_3_ ( .D(simpleXor_315_port_z), .CK(clk), .Q(
        mult_ab_0_2[3]), .QN() );
  DFF_X1 mult_ab_0_2_reg_2_ ( .D(simpleXor_291_port_z), .CK(clk), .Q(
        mult_ab_0_2[2]), .QN() );
  DFF_X1 mult_ab_0_2_reg_1_ ( .D(simpleXor_267_port_z), .CK(clk), .Q(
        mult_ab_0_2[1]), .QN() );
  DFF_X1 mult_ab_0_2_reg_0_ ( .D(simpleXor_243_port_z), .CK(clk), .Q(
        mult_ab_0_2[0]), .QN() );
  DFF_X1 mult_ab_0_3_reg_4_ ( .D(simpleXor_341_port_z), .CK(clk), .Q(
        mult_ab_0_3[4]), .QN() );
  DFF_X1 mult_ab_0_3_reg_3_ ( .D(simpleXor_317_port_z), .CK(clk), .Q(
        mult_ab_0_3[3]), .QN() );
  DFF_X1 mult_ab_0_3_reg_2_ ( .D(simpleXor_293_port_z), .CK(clk), .Q(
        mult_ab_0_3[2]), .QN() );
  DFF_X1 mult_ab_0_3_reg_1_ ( .D(simpleXor_269_port_z), .CK(clk), .Q(
        mult_ab_0_3[1]), .QN() );
  DFF_X1 mult_ab_0_3_reg_0_ ( .D(simpleXor_245_port_z), .CK(clk), .Q(
        mult_ab_0_3[0]), .QN() );
  DFF_X1 mult_ab_1_0_reg_4_ ( .D(simpleXor_343_port_z), .CK(clk), .Q(
        mult_ab_1_0[4]), .QN() );
  DFF_X1 mult_ab_1_0_reg_3_ ( .D(simpleXor_319_port_z), .CK(clk), .Q(
        mult_ab_1_0[3]), .QN() );
  DFF_X1 mult_ab_1_0_reg_2_ ( .D(simpleXor_295_port_z), .CK(clk), .Q(
        mult_ab_1_0[2]), .QN() );
  DFF_X1 mult_ab_1_0_reg_1_ ( .D(simpleXor_271_port_z), .CK(clk), .Q(
        mult_ab_1_0[1]), .QN() );
  DFF_X1 mult_ab_1_0_reg_0_ ( .D(simpleXor_247_port_z), .CK(clk), .Q(
        mult_ab_1_0[0]), .QN() );
  DFF_X1 mult_ab_1_1_reg_4_ ( .D(N17), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 mult_ab_1_1_reg_3_ ( .D(N13), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 mult_ab_1_1_reg_2_ ( .D(N9), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 mult_ab_1_1_reg_1_ ( .D(N5), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 mult_ab_1_1_reg_0_ ( .D(N1), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 mult_ab_1_2_reg_4_ ( .D(simpleXor_345_port_z), .CK(clk), .Q(
        mult_ab_1_2[4]), .QN() );
  DFF_X1 mult_ab_1_2_reg_3_ ( .D(simpleXor_321_port_z), .CK(clk), .Q(
        mult_ab_1_2[3]), .QN() );
  DFF_X1 mult_ab_1_2_reg_2_ ( .D(simpleXor_297_port_z), .CK(clk), .Q(
        mult_ab_1_2[2]), .QN() );
  DFF_X1 mult_ab_1_2_reg_1_ ( .D(simpleXor_273_port_z), .CK(clk), .Q(
        mult_ab_1_2[1]), .QN() );
  DFF_X1 mult_ab_1_2_reg_0_ ( .D(simpleXor_249_port_z), .CK(clk), .Q(
        mult_ab_1_2[0]), .QN() );
  DFF_X1 mult_ab_1_3_reg_4_ ( .D(simpleXor_347_port_z), .CK(clk), .Q(
        mult_ab_1_3[4]), .QN() );
  DFF_X1 mult_ab_1_3_reg_3_ ( .D(simpleXor_323_port_z), .CK(clk), .Q(
        mult_ab_1_3[3]), .QN() );
  DFF_X1 mult_ab_1_3_reg_2_ ( .D(simpleXor_299_port_z), .CK(clk), .Q(
        mult_ab_1_3[2]), .QN() );
  DFF_X1 mult_ab_1_3_reg_1_ ( .D(simpleXor_275_port_z), .CK(clk), .Q(
        mult_ab_1_3[1]), .QN() );
  DFF_X1 mult_ab_1_3_reg_0_ ( .D(simpleXor_251_port_z), .CK(clk), .Q(
        mult_ab_1_3[0]), .QN() );
  AND2_X1 U143 ( .A1(ref_1_port_o_1_3[0]), .A2(port_a_1[0]), .ZN(
        simpleXor_250_port_a0) );
  AND2_X1 U144 ( .A1(ref_1_port_o_1_3[1]), .A2(port_a_1[1]), .ZN(
        simpleXor_274_port_a0) );
  AND2_X1 U145 ( .A1(ref_1_port_o_1_3[2]), .A2(port_a_1[2]), .ZN(
        simpleXor_298_port_a0) );
  AND2_X1 U146 ( .A1(ref_1_port_o_1_3[3]), .A2(port_a_1[3]), .ZN(
        simpleXor_322_port_a0) );
  AND2_X1 U147 ( .A1(ref_1_port_o_1_3[4]), .A2(port_a_1[4]), .ZN(
        simpleXor_346_port_a0) );
  AND2_X1 U148 ( .A1(ref_1_port_o_1_2[0]), .A2(port_a_1[0]), .ZN(
        simpleXor_248_port_a0) );
  AND2_X1 U149 ( .A1(ref_1_port_o_1_2[1]), .A2(port_a_1[1]), .ZN(
        simpleXor_272_port_a0) );
  AND2_X1 U150 ( .A1(ref_1_port_o_1_2[2]), .A2(port_a_1[2]), .ZN(
        simpleXor_296_port_a0) );
  AND2_X1 U151 ( .A1(ref_1_port_o_1_2[3]), .A2(port_a_1[3]), .ZN(
        simpleXor_320_port_a0) );
  AND2_X1 U152 ( .A1(ref_1_port_o_1_2[4]), .A2(port_a_1[4]), .ZN(
        simpleXor_344_port_a0) );
  AND2_X1 U153 ( .A1(ref_1_port_o_1_0[0]), .A2(port_a_1[0]), .ZN(
        simpleXor_246_port_a0) );
  AND2_X1 U154 ( .A1(ref_1_port_o_1_0[1]), .A2(port_a_1[1]), .ZN(
        simpleXor_270_port_a0) );
  AND2_X1 U155 ( .A1(ref_1_port_o_1_0[2]), .A2(port_a_1[2]), .ZN(
        simpleXor_294_port_a0) );
  AND2_X1 U156 ( .A1(ref_1_port_o_1_0[3]), .A2(port_a_1[3]), .ZN(
        simpleXor_318_port_a0) );
  AND2_X1 U157 ( .A1(ref_1_port_o_1_0[4]), .A2(port_a_1[4]), .ZN(
        simpleXor_342_port_a0) );
  AND2_X1 U158 ( .A1(ref_1_port_o_0_3[0]), .A2(port_a_0[0]), .ZN(
        simpleXor_244_port_a0) );
  AND2_X1 U159 ( .A1(ref_1_port_o_0_3[1]), .A2(port_a_0[1]), .ZN(
        simpleXor_268_port_a0) );
  AND2_X1 U160 ( .A1(ref_1_port_o_0_3[2]), .A2(port_a_0[2]), .ZN(
        simpleXor_292_port_a0) );
  AND2_X1 U161 ( .A1(ref_1_port_o_0_3[3]), .A2(port_a_0[3]), .ZN(
        simpleXor_316_port_a0) );
  AND2_X1 U162 ( .A1(ref_1_port_o_0_3[4]), .A2(port_a_0[4]), .ZN(
        simpleXor_340_port_a0) );
  AND2_X1 U163 ( .A1(ref_1_port_o_0_2[0]), .A2(port_a_0[0]), .ZN(
        simpleXor_242_port_a0) );
  AND2_X1 U164 ( .A1(ref_1_port_o_0_2[1]), .A2(port_a_0[1]), .ZN(
        simpleXor_266_port_a0) );
  AND2_X1 U165 ( .A1(ref_1_port_o_0_2[2]), .A2(port_a_0[2]), .ZN(
        simpleXor_290_port_a0) );
  AND2_X1 U166 ( .A1(ref_1_port_o_0_2[3]), .A2(port_a_0[3]), .ZN(
        simpleXor_314_port_a0) );
  AND2_X1 U167 ( .A1(ref_1_port_o_0_2[4]), .A2(port_a_0[4]), .ZN(
        simpleXor_338_port_a0) );
  AND2_X1 U168 ( .A1(ref_1_port_o_0_1[0]), .A2(port_a_0[0]), .ZN(
        simpleXor_240_port_a0) );
  AND2_X1 U169 ( .A1(ref_1_port_o_0_1[1]), .A2(port_a_0[1]), .ZN(
        simpleXor_264_port_a0) );
  AND2_X1 U170 ( .A1(ref_1_port_o_0_1[2]), .A2(port_a_0[2]), .ZN(
        simpleXor_288_port_a0) );
  AND2_X1 U171 ( .A1(ref_1_port_o_0_1[3]), .A2(port_a_0[3]), .ZN(
        simpleXor_312_port_a0) );
  AND2_X1 U172 ( .A1(ref_1_port_o_0_1[4]), .A2(port_a_0[4]), .ZN(
        simpleXor_336_port_a0) );
  AND2_X1 U173 ( .A1(ref_1_port_o_2_1[0]), .A2(port_a_2[0]), .ZN(
        simpleXor_254_port_a0) );
  AND2_X1 U174 ( .A1(ref_1_port_o_2_1[1]), .A2(port_a_2[1]), .ZN(
        simpleXor_278_port_a0) );
  AND2_X1 U175 ( .A1(ref_1_port_o_2_1[2]), .A2(port_a_2[2]), .ZN(
        simpleXor_302_port_a0) );
  AND2_X1 U176 ( .A1(ref_1_port_o_2_1[3]), .A2(port_a_2[3]), .ZN(
        simpleXor_326_port_a0) );
  AND2_X1 U177 ( .A1(ref_1_port_o_2_1[4]), .A2(port_a_2[4]), .ZN(
        simpleXor_350_port_a0) );
  AND2_X1 U178 ( .A1(ref_1_port_o_2_0[0]), .A2(port_a_2[0]), .ZN(
        simpleXor_252_port_a0) );
  AND2_X1 U179 ( .A1(ref_1_port_o_2_0[1]), .A2(port_a_2[1]), .ZN(
        simpleXor_276_port_a0) );
  AND2_X1 U180 ( .A1(ref_1_port_o_2_0[2]), .A2(port_a_2[2]), .ZN(
        simpleXor_300_port_a0) );
  AND2_X1 U181 ( .A1(ref_1_port_o_2_0[3]), .A2(port_a_2[3]), .ZN(
        simpleXor_324_port_a0) );
  AND2_X1 U182 ( .A1(ref_1_port_o_2_0[4]), .A2(port_a_2[4]), .ZN(
        simpleXor_348_port_a0) );
  AND2_X1 U183 ( .A1(ref_1_port_o_2_3[0]), .A2(port_a_2[0]), .ZN(
        simpleXor_256_port_a0) );
  AND2_X1 U184 ( .A1(ref_1_port_o_2_3[1]), .A2(port_a_2[1]), .ZN(
        simpleXor_280_port_a0) );
  AND2_X1 U185 ( .A1(ref_1_port_o_2_3[2]), .A2(port_a_2[2]), .ZN(
        simpleXor_304_port_a0) );
  AND2_X1 U186 ( .A1(ref_1_port_o_2_3[3]), .A2(port_a_2[3]), .ZN(
        simpleXor_328_port_a0) );
  AND2_X1 U187 ( .A1(ref_1_port_o_2_3[4]), .A2(port_a_2[4]), .ZN(
        simpleXor_352_port_a0) );
  AND2_X1 U188 ( .A1(ref_1_port_o_3_1[0]), .A2(port_a_3[0]), .ZN(
        simpleXor_260_port_a0) );
  AND2_X1 U189 ( .A1(ref_1_port_o_3_1[1]), .A2(port_a_3[1]), .ZN(
        simpleXor_284_port_a0) );
  AND2_X1 U190 ( .A1(ref_1_port_o_3_1[2]), .A2(port_a_3[2]), .ZN(
        simpleXor_308_port_a0) );
  AND2_X1 U191 ( .A1(ref_1_port_o_3_1[3]), .A2(port_a_3[3]), .ZN(
        simpleXor_332_port_a0) );
  AND2_X1 U192 ( .A1(ref_1_port_o_3_1[4]), .A2(port_a_3[4]), .ZN(
        simpleXor_356_port_a0) );
  AND2_X1 U193 ( .A1(ref_1_port_o_3_0[0]), .A2(port_a_3[0]), .ZN(
        simpleXor_258_port_a0) );
  AND2_X1 U194 ( .A1(ref_1_port_o_3_0[1]), .A2(port_a_3[1]), .ZN(
        simpleXor_282_port_a0) );
  AND2_X1 U195 ( .A1(ref_1_port_o_3_0[2]), .A2(port_a_3[2]), .ZN(
        simpleXor_306_port_a0) );
  AND2_X1 U196 ( .A1(ref_1_port_o_3_0[3]), .A2(port_a_3[3]), .ZN(
        simpleXor_330_port_a0) );
  AND2_X1 U197 ( .A1(ref_1_port_o_3_0[4]), .A2(port_a_3[4]), .ZN(
        simpleXor_354_port_a0) );
  AND2_X1 U198 ( .A1(ref_1_port_o_3_2[0]), .A2(port_a_3[0]), .ZN(
        simpleXor_262_port_a0) );
  AND2_X1 U199 ( .A1(ref_1_port_o_3_2[1]), .A2(port_a_3[1]), .ZN(
        simpleXor_286_port_a0) );
  AND2_X1 U200 ( .A1(ref_1_port_o_3_2[2]), .A2(port_a_3[2]), .ZN(
        simpleXor_310_port_a0) );
  AND2_X1 U201 ( .A1(ref_1_port_o_3_2[3]), .A2(port_a_3[3]), .ZN(
        simpleXor_334_port_a0) );
  AND2_X1 U202 ( .A1(ref_1_port_o_3_2[4]), .A2(port_a_3[4]), .ZN(
        simpleXor_358_port_a0) );
  AND2_X1 U203 ( .A1(ref_1_port_o_1_1[0]), .A2(port_a_1[0]), .ZN(N1) );
  AND2_X1 U204 ( .A1(ref_1_port_o_1_1[1]), .A2(port_a_1[1]), .ZN(N5) );
  AND2_X1 U205 ( .A1(ref_1_port_o_1_1[2]), .A2(port_a_1[2]), .ZN(N9) );
  AND2_X1 U206 ( .A1(ref_1_port_o_1_1[3]), .A2(port_a_1[3]), .ZN(N13) );
  AND2_X1 U207 ( .A1(ref_1_port_o_1_1[4]), .A2(port_a_1[4]), .ZN(N17) );
  AND2_X1 U208 ( .A1(ref_1_port_o_0_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U209 ( .A1(ref_1_port_o_0_0[1]), .A2(port_a_0[1]), .ZN(N4) );
  AND2_X1 U210 ( .A1(ref_1_port_o_0_0[2]), .A2(port_a_0[2]), .ZN(N8) );
  AND2_X1 U211 ( .A1(ref_1_port_o_0_0[3]), .A2(port_a_0[3]), .ZN(N12) );
  AND2_X1 U212 ( .A1(ref_1_port_o_0_0[4]), .A2(port_a_0[4]), .ZN(N16) );
  AND2_X1 U213 ( .A1(ref_1_port_o_2_2[0]), .A2(port_a_2[0]), .ZN(N2) );
  AND2_X1 U214 ( .A1(ref_1_port_o_2_2[1]), .A2(port_a_2[1]), .ZN(N6) );
  AND2_X1 U215 ( .A1(ref_1_port_o_2_2[2]), .A2(port_a_2[2]), .ZN(N10) );
  AND2_X1 U216 ( .A1(ref_1_port_o_2_2[3]), .A2(port_a_2[3]), .ZN(N14) );
  AND2_X1 U217 ( .A1(ref_1_port_o_2_2[4]), .A2(port_a_2[4]), .ZN(N18) );
  AND2_X1 U218 ( .A1(ref_1_port_o_3_3[0]), .A2(port_a_3[0]), .ZN(N3) );
  AND2_X1 U219 ( .A1(ref_1_port_o_3_3[1]), .A2(port_a_3[1]), .ZN(N7) );
  AND2_X1 U220 ( .A1(ref_1_port_o_3_3[2]), .A2(port_a_3[2]), .ZN(N11) );
  AND2_X1 U221 ( .A1(ref_1_port_o_3_3[3]), .A2(port_a_3[3]), .ZN(N15) );
  AND2_X1 U222 ( .A1(ref_1_port_o_3_3[4]), .A2(port_a_3[4]), .ZN(N19) );
  XOR2_X1 U223 ( .A(n9), .B(n10), .Z(port_c_3[0]) );
  XNOR2_X1 U224 ( .A(temp_0_3[0]), .B(mult_ab_3_2[0]), .ZN(n9) );
  XNOR2_X1 U225 ( .A(mult_ab_3_1[0]), .B(mult_ab_3_0[0]), .ZN(n10) );
  XOR2_X1 U226 ( .A(n7), .B(n8), .Z(port_c_3[1]) );
  XNOR2_X1 U227 ( .A(temp_0_3[1]), .B(mult_ab_3_2[1]), .ZN(n7) );
  XNOR2_X1 U228 ( .A(mult_ab_3_1[1]), .B(mult_ab_3_0[1]), .ZN(n8) );
  XOR2_X1 U229 ( .A(n5), .B(n6), .Z(port_c_3[2]) );
  XNOR2_X1 U230 ( .A(temp_0_3[2]), .B(mult_ab_3_2[2]), .ZN(n5) );
  XNOR2_X1 U231 ( .A(mult_ab_3_1[2]), .B(mult_ab_3_0[2]), .ZN(n6) );
  XOR2_X1 U232 ( .A(n3), .B(n4), .Z(port_c_3[3]) );
  XNOR2_X1 U233 ( .A(temp_0_3[3]), .B(mult_ab_3_2[3]), .ZN(n3) );
  XNOR2_X1 U234 ( .A(mult_ab_3_1[3]), .B(mult_ab_3_0[3]), .ZN(n4) );
  XOR2_X1 U235 ( .A(n1), .B(n2), .Z(port_c_3[4]) );
  XNOR2_X1 U236 ( .A(temp_0_3[4]), .B(mult_ab_3_2[4]), .ZN(n1) );
  XNOR2_X1 U237 ( .A(mult_ab_3_1[4]), .B(mult_ab_3_0[4]), .ZN(n2) );
  XOR2_X1 U238 ( .A(n19), .B(n20), .Z(port_c_2[0]) );
  XNOR2_X1 U239 ( .A(temp_0_2[0]), .B(mult_ab_2_3[0]), .ZN(n19) );
  XNOR2_X1 U240 ( .A(mult_ab_2_1[0]), .B(mult_ab_2_0[0]), .ZN(n20) );
  XOR2_X1 U241 ( .A(n17), .B(n18), .Z(port_c_2[1]) );
  XNOR2_X1 U242 ( .A(temp_0_2[1]), .B(mult_ab_2_3[1]), .ZN(n17) );
  XNOR2_X1 U243 ( .A(mult_ab_2_1[1]), .B(mult_ab_2_0[1]), .ZN(n18) );
  XOR2_X1 U244 ( .A(n15), .B(n16), .Z(port_c_2[2]) );
  XNOR2_X1 U245 ( .A(temp_0_2[2]), .B(mult_ab_2_3[2]), .ZN(n15) );
  XNOR2_X1 U246 ( .A(mult_ab_2_1[2]), .B(mult_ab_2_0[2]), .ZN(n16) );
  XOR2_X1 U247 ( .A(n13), .B(n14), .Z(port_c_2[3]) );
  XNOR2_X1 U248 ( .A(temp_0_2[3]), .B(mult_ab_2_3[3]), .ZN(n13) );
  XNOR2_X1 U249 ( .A(mult_ab_2_1[3]), .B(mult_ab_2_0[3]), .ZN(n14) );
  XOR2_X1 U250 ( .A(n11), .B(n12), .Z(port_c_2[4]) );
  XNOR2_X1 U251 ( .A(temp_0_2[4]), .B(mult_ab_2_3[4]), .ZN(n11) );
  XNOR2_X1 U252 ( .A(mult_ab_2_1[4]), .B(mult_ab_2_0[4]), .ZN(n12) );
  XOR2_X1 U253 ( .A(n29), .B(n30), .Z(port_c_1[0]) );
  XNOR2_X1 U254 ( .A(temp_0_1[0]), .B(mult_ab_1_3[0]), .ZN(n29) );
  XNOR2_X1 U255 ( .A(mult_ab_1_2[0]), .B(mult_ab_1_0[0]), .ZN(n30) );
  XOR2_X1 U256 ( .A(n27), .B(n28), .Z(port_c_1[1]) );
  XNOR2_X1 U257 ( .A(temp_0_1[1]), .B(mult_ab_1_3[1]), .ZN(n27) );
  XNOR2_X1 U258 ( .A(mult_ab_1_2[1]), .B(mult_ab_1_0[1]), .ZN(n28) );
  XOR2_X1 U259 ( .A(n25), .B(n26), .Z(port_c_1[2]) );
  XNOR2_X1 U260 ( .A(temp_0_1[2]), .B(mult_ab_1_3[2]), .ZN(n25) );
  XNOR2_X1 U261 ( .A(mult_ab_1_2[2]), .B(mult_ab_1_0[2]), .ZN(n26) );
  XOR2_X1 U262 ( .A(n23), .B(n24), .Z(port_c_1[3]) );
  XNOR2_X1 U263 ( .A(temp_0_1[3]), .B(mult_ab_1_3[3]), .ZN(n23) );
  XNOR2_X1 U264 ( .A(mult_ab_1_2[3]), .B(mult_ab_1_0[3]), .ZN(n24) );
  XOR2_X1 U265 ( .A(n21), .B(n22), .Z(port_c_1[4]) );
  XNOR2_X1 U266 ( .A(temp_0_1[4]), .B(mult_ab_1_3[4]), .ZN(n21) );
  XNOR2_X1 U267 ( .A(mult_ab_1_2[4]), .B(mult_ab_1_0[4]), .ZN(n22) );
  XOR2_X1 U268 ( .A(n39), .B(n40), .Z(port_c_0[0]) );
  XNOR2_X1 U269 ( .A(temp_0_0[0]), .B(mult_ab_0_3[0]), .ZN(n39) );
  XNOR2_X1 U270 ( .A(mult_ab_0_2[0]), .B(mult_ab_0_1[0]), .ZN(n40) );
  XOR2_X1 U271 ( .A(n37), .B(n38), .Z(port_c_0[1]) );
  XNOR2_X1 U272 ( .A(temp_0_0[1]), .B(mult_ab_0_3[1]), .ZN(n37) );
  XNOR2_X1 U273 ( .A(mult_ab_0_2[1]), .B(mult_ab_0_1[1]), .ZN(n38) );
  XOR2_X1 U274 ( .A(n35), .B(n36), .Z(port_c_0[2]) );
  XNOR2_X1 U275 ( .A(temp_0_0[2]), .B(mult_ab_0_3[2]), .ZN(n35) );
  XNOR2_X1 U276 ( .A(mult_ab_0_2[2]), .B(mult_ab_0_1[2]), .ZN(n36) );
  XOR2_X1 U277 ( .A(n33), .B(n34), .Z(port_c_0[3]) );
  XNOR2_X1 U278 ( .A(temp_0_0[3]), .B(mult_ab_0_3[3]), .ZN(n33) );
  XNOR2_X1 U279 ( .A(mult_ab_0_2[3]), .B(mult_ab_0_1[3]), .ZN(n34) );
  XOR2_X1 U280 ( .A(n31), .B(n32), .Z(port_c_0[4]) );
  XNOR2_X1 U281 ( .A(temp_0_0[4]), .B(mult_ab_0_3[4]), .ZN(n31) );
  XNOR2_X1 U282 ( .A(mult_ab_0_2[4]), .B(mult_ab_0_1[4]), .ZN(n32) );
  BUF_X1 ref_1_U42 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n40) );
  BUF_X1 ref_1_U41 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n39) );
  BUF_X1 ref_1_U40 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n38) );
  BUF_X1 ref_1_U39 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n37) );
  BUF_X1 ref_1_U38 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n36) );
  BUF_X1 ref_1_U37 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n35) );
  BUF_X1 ref_1_U36 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n34) );
  BUF_X1 ref_1_U35 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n33) );
  BUF_X1 ref_1_U34 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n32) );
  BUF_X1 ref_1_U33 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n31) );
  BUF_X1 ref_1_U32 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n30) );
  BUF_X1 ref_1_U31 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n29) );
  BUF_X1 ref_1_U30 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n28) );
  BUF_X1 ref_1_U29 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n27) );
  BUF_X1 ref_1_U28 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n26) );
  BUF_X1 ref_1_U27 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n25) );
  BUF_X1 ref_1_U26 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n24) );
  BUF_X1 ref_1_U25 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n23) );
  BUF_X1 ref_1_U24 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n22) );
  BUF_X1 ref_1_U23 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n21) );
  BUF_X1 ref_1_U22 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n20) );
  BUF_X1 ref_1_U21 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n19) );
  BUF_X1 ref_1_U20 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n18) );
  BUF_X1 ref_1_U19 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n17) );
  BUF_X1 ref_1_U18 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n16) );
  BUF_X1 ref_1_U17 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n15) );
  BUF_X1 ref_1_U16 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n14) );
  BUF_X1 ref_1_U15 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n13) );
  BUF_X1 ref_1_U14 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n12) );
  BUF_X1 ref_1_U13 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n11) );
  BUF_X1 ref_1_U12 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n10) );
  BUF_X1 ref_1_U11 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n9) );
  BUF_X1 ref_1_U10 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n8) );
  BUF_X1 ref_1_U9 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n7) );
  BUF_X1 ref_1_U8 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n6) );
  BUF_X1 ref_1_U7 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n5) );
  BUF_X1 ref_1_U6 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n4) );
  BUF_X1 ref_1_U5 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n3) );
  BUF_X1 ref_1_U4 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n2) );
  BUF_X1 ref_1_U3 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n1) );
  DFF_X1 ref_1_reg_out_3_3_reg_0_ ( .D(ref_1_maj_95_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_1_ ( .D(ref_1_maj_111_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_2_ ( .D(ref_1_maj_127_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_3_ ( .D(ref_1_maj_143_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_4_ ( .D(ref_1_maj_159_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_0_ ( .D(ref_1_maj_94_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_1_ ( .D(ref_1_maj_110_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_2_ ( .D(ref_1_maj_126_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_3_ ( .D(ref_1_maj_142_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_4_ ( .D(ref_1_maj_158_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_0_ ( .D(ref_1_maj_93_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_1_ ( .D(ref_1_maj_109_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_2_ ( .D(ref_1_maj_125_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_3_ ( .D(ref_1_maj_141_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_4_ ( .D(ref_1_maj_157_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_0_ ( .D(ref_1_maj_92_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_1_ ( .D(ref_1_maj_108_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_2_ ( .D(ref_1_maj_124_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_3_ ( .D(ref_1_maj_140_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_4_ ( .D(ref_1_maj_156_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_0_ ( .D(ref_1_maj_91_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_1_ ( .D(ref_1_maj_107_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_2_ ( .D(ref_1_maj_123_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_3_ ( .D(ref_1_maj_139_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_4_ ( .D(ref_1_maj_155_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_0_ ( .D(ref_1_maj_90_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_1_ ( .D(ref_1_maj_106_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_2_ ( .D(ref_1_maj_122_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_3_ ( .D(ref_1_maj_138_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_4_ ( .D(ref_1_maj_154_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_0_ ( .D(ref_1_maj_89_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_1_ ( .D(ref_1_maj_105_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_2_ ( .D(ref_1_maj_121_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_3_ ( .D(ref_1_maj_137_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_4_ ( .D(ref_1_maj_153_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_0_ ( .D(ref_1_maj_88_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_1_ ( .D(ref_1_maj_104_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_2_ ( .D(ref_1_maj_120_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_3_ ( .D(ref_1_maj_136_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_4_ ( .D(ref_1_maj_152_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_0_ ( .D(ref_1_maj_87_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_1_ ( .D(ref_1_maj_103_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_2_ ( .D(ref_1_maj_119_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_3_ ( .D(ref_1_maj_135_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_4_ ( .D(ref_1_maj_151_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_0_ ( .D(ref_1_maj_86_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_1_ ( .D(ref_1_maj_102_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_2_ ( .D(ref_1_maj_118_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_3_ ( .D(ref_1_maj_134_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_4_ ( .D(ref_1_maj_150_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_0_ ( .D(ref_1_maj_85_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_1_ ( .D(ref_1_maj_101_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_2_ ( .D(ref_1_maj_117_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_3_ ( .D(ref_1_maj_133_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_4_ ( .D(ref_1_maj_149_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_0_ ( .D(ref_1_maj_84_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_1_ ( .D(ref_1_maj_100_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_2_ ( .D(ref_1_maj_116_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_3_ ( .D(ref_1_maj_132_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_4_ ( .D(ref_1_maj_148_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_0_ ( .D(ref_1_maj_83_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_1_ ( .D(ref_1_maj_99_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_2_ ( .D(ref_1_maj_115_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_3_ ( .D(ref_1_maj_131_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_4_ ( .D(ref_1_maj_147_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_0_ ( .D(ref_1_maj_82_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_1_ ( .D(ref_1_maj_98_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_2_ ( .D(ref_1_maj_114_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_3_ ( .D(ref_1_maj_130_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_4_ ( .D(ref_1_maj_146_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_0_ ( .D(ref_1_maj_81_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_1_ ( .D(ref_1_maj_97_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_2_ ( .D(ref_1_maj_113_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_3_ ( .D(ref_1_maj_129_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_4_ ( .D(ref_1_maj_145_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_0_ ( .D(ref_1_maj_80_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_1_ ( .D(ref_1_maj_96_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_2_ ( .D(ref_1_maj_112_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_3_ ( .D(ref_1_maj_128_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_4_ ( .D(ref_1_maj_144_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[4]), .QN() );
  XOR2_X1 ref_1_simpleXor_240_U1 ( .A(port_rand_ref[0]), .B(port_b_0[0]), .Z(
        ref_1_simpleXor_240_port_z) );
  XOR2_X1 ref_1_simpleXor_241_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_240_port_z), .Z(ref_1_simpleXor_241_port_z) );
  XOR2_X1 ref_1_simpleXor_242_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_241_port_z), .Z(ref_1_simpleXor_242_port_z) );
  XOR2_X1 ref_1_simpleXor_243_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_242_port_z), .Z(ref_1_simpleXor_243_port_z) );
  XOR2_X1 ref_1_simpleXor_244_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_243_port_z), .Z(ref_1_simpleXor_244_port_z) );
  XOR2_X1 ref_1_simpleXor_245_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_244_port_z), .Z(ref_1_refreshed_0_0_) );
  XOR2_X1 ref_1_simpleXor_246_U1 ( .A(port_rand_ref[0]), .B(port_b_1[0]), .Z(
        ref_1_simpleXor_246_port_z) );
  XOR2_X1 ref_1_simpleXor_247_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_246_port_z), .Z(ref_1_simpleXor_247_port_z) );
  XOR2_X1 ref_1_simpleXor_248_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_247_port_z), .Z(ref_1_simpleXor_248_port_z) );
  XOR2_X1 ref_1_simpleXor_249_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_248_port_z), .Z(ref_1_simpleXor_249_port_z) );
  XOR2_X1 ref_1_simpleXor_250_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_249_port_z), .Z(ref_1_simpleXor_250_port_z) );
  XOR2_X1 ref_1_simpleXor_251_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_250_port_z), .Z(ref_1_refreshed_1_0_) );
  XOR2_X1 ref_1_simpleXor_252_U1 ( .A(port_rand_ref[2]), .B(port_b_2[0]), .Z(
        ref_1_simpleXor_252_port_z) );
  XOR2_X1 ref_1_simpleXor_253_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_252_port_z), .Z(ref_1_simpleXor_253_port_z) );
  XOR2_X1 ref_1_simpleXor_254_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_253_port_z), .Z(ref_1_simpleXor_254_port_z) );
  XOR2_X1 ref_1_simpleXor_255_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_254_port_z), .Z(ref_1_simpleXor_255_port_z) );
  XOR2_X1 ref_1_simpleXor_256_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_255_port_z), .Z(ref_1_simpleXor_256_port_z) );
  XOR2_X1 ref_1_simpleXor_257_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_256_port_z), .Z(ref_1_refreshed_2_0_) );
  XOR2_X1 ref_1_simpleXor_258_U1 ( .A(port_rand_ref[4]), .B(port_b_3[0]), .Z(
        ref_1_simpleXor_258_port_z) );
  XOR2_X1 ref_1_simpleXor_259_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_258_port_z), .Z(ref_1_simpleXor_259_port_z) );
  XOR2_X1 ref_1_simpleXor_260_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_259_port_z), .Z(ref_1_simpleXor_260_port_z) );
  XOR2_X1 ref_1_simpleXor_261_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_260_port_z), .Z(ref_1_simpleXor_261_port_z) );
  XOR2_X1 ref_1_simpleXor_262_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_261_port_z), .Z(ref_1_simpleXor_262_port_z) );
  XOR2_X1 ref_1_simpleXor_263_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_262_port_z), .Z(ref_1_refreshed_3_0_) );
  XOR2_X1 ref_1_simpleXor_264_U1 ( .A(port_rand_ref[0]), .B(port_b_0[1]), .Z(
        ref_1_simpleXor_264_port_z) );
  XOR2_X1 ref_1_simpleXor_265_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_264_port_z), .Z(ref_1_simpleXor_265_port_z) );
  XOR2_X1 ref_1_simpleXor_266_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_265_port_z), .Z(ref_1_simpleXor_266_port_z) );
  XOR2_X1 ref_1_simpleXor_267_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_266_port_z), .Z(ref_1_simpleXor_267_port_z) );
  XOR2_X1 ref_1_simpleXor_268_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_267_port_z), .Z(ref_1_simpleXor_268_port_z) );
  XOR2_X1 ref_1_simpleXor_269_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_268_port_z), .Z(ref_1_refreshed_0_1_) );
  XOR2_X1 ref_1_simpleXor_270_U1 ( .A(port_rand_ref[0]), .B(port_b_1[1]), .Z(
        ref_1_simpleXor_270_port_z) );
  XOR2_X1 ref_1_simpleXor_271_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_270_port_z), .Z(ref_1_simpleXor_271_port_z) );
  XOR2_X1 ref_1_simpleXor_272_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_271_port_z), .Z(ref_1_simpleXor_272_port_z) );
  XOR2_X1 ref_1_simpleXor_273_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_272_port_z), .Z(ref_1_simpleXor_273_port_z) );
  XOR2_X1 ref_1_simpleXor_274_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_273_port_z), .Z(ref_1_simpleXor_274_port_z) );
  XOR2_X1 ref_1_simpleXor_275_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_274_port_z), .Z(ref_1_refreshed_1_1_) );
  XOR2_X1 ref_1_simpleXor_276_U1 ( .A(port_rand_ref[2]), .B(port_b_2[1]), .Z(
        ref_1_simpleXor_276_port_z) );
  XOR2_X1 ref_1_simpleXor_277_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_276_port_z), .Z(ref_1_simpleXor_277_port_z) );
  XOR2_X1 ref_1_simpleXor_278_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_277_port_z), .Z(ref_1_simpleXor_278_port_z) );
  XOR2_X1 ref_1_simpleXor_279_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_278_port_z), .Z(ref_1_simpleXor_279_port_z) );
  XOR2_X1 ref_1_simpleXor_280_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_279_port_z), .Z(ref_1_simpleXor_280_port_z) );
  XOR2_X1 ref_1_simpleXor_281_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_280_port_z), .Z(ref_1_refreshed_2_1_) );
  XOR2_X1 ref_1_simpleXor_282_U1 ( .A(port_rand_ref[4]), .B(port_b_3[1]), .Z(
        ref_1_simpleXor_282_port_z) );
  XOR2_X1 ref_1_simpleXor_283_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_282_port_z), .Z(ref_1_simpleXor_283_port_z) );
  XOR2_X1 ref_1_simpleXor_284_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_283_port_z), .Z(ref_1_simpleXor_284_port_z) );
  XOR2_X1 ref_1_simpleXor_285_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_284_port_z), .Z(ref_1_simpleXor_285_port_z) );
  XOR2_X1 ref_1_simpleXor_286_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_285_port_z), .Z(ref_1_simpleXor_286_port_z) );
  XOR2_X1 ref_1_simpleXor_287_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_286_port_z), .Z(ref_1_refreshed_3_1_) );
  XOR2_X1 ref_1_simpleXor_288_U1 ( .A(port_rand_ref[0]), .B(port_b_0[2]), .Z(
        ref_1_simpleXor_288_port_z) );
  XOR2_X1 ref_1_simpleXor_289_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_288_port_z), .Z(ref_1_simpleXor_289_port_z) );
  XOR2_X1 ref_1_simpleXor_290_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_289_port_z), .Z(ref_1_simpleXor_290_port_z) );
  XOR2_X1 ref_1_simpleXor_291_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_290_port_z), .Z(ref_1_simpleXor_291_port_z) );
  XOR2_X1 ref_1_simpleXor_292_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_291_port_z), .Z(ref_1_simpleXor_292_port_z) );
  XOR2_X1 ref_1_simpleXor_293_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_292_port_z), .Z(ref_1_refreshed_0_2_) );
  XOR2_X1 ref_1_simpleXor_294_U1 ( .A(port_rand_ref[0]), .B(port_b_1[2]), .Z(
        ref_1_simpleXor_294_port_z) );
  XOR2_X1 ref_1_simpleXor_295_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_294_port_z), .Z(ref_1_simpleXor_295_port_z) );
  XOR2_X1 ref_1_simpleXor_296_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_295_port_z), .Z(ref_1_simpleXor_296_port_z) );
  XOR2_X1 ref_1_simpleXor_297_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_296_port_z), .Z(ref_1_simpleXor_297_port_z) );
  XOR2_X1 ref_1_simpleXor_298_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_297_port_z), .Z(ref_1_simpleXor_298_port_z) );
  XOR2_X1 ref_1_simpleXor_299_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_298_port_z), .Z(ref_1_refreshed_1_2_) );
  XOR2_X1 ref_1_simpleXor_300_U1 ( .A(port_rand_ref[2]), .B(port_b_2[2]), .Z(
        ref_1_simpleXor_300_port_z) );
  XOR2_X1 ref_1_simpleXor_301_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_300_port_z), .Z(ref_1_simpleXor_301_port_z) );
  XOR2_X1 ref_1_simpleXor_302_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_301_port_z), .Z(ref_1_simpleXor_302_port_z) );
  XOR2_X1 ref_1_simpleXor_303_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_302_port_z), .Z(ref_1_simpleXor_303_port_z) );
  XOR2_X1 ref_1_simpleXor_304_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_303_port_z), .Z(ref_1_simpleXor_304_port_z) );
  XOR2_X1 ref_1_simpleXor_305_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_304_port_z), .Z(ref_1_refreshed_2_2_) );
  XOR2_X1 ref_1_simpleXor_306_U1 ( .A(port_rand_ref[4]), .B(port_b_3[2]), .Z(
        ref_1_simpleXor_306_port_z) );
  XOR2_X1 ref_1_simpleXor_307_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_306_port_z), .Z(ref_1_simpleXor_307_port_z) );
  XOR2_X1 ref_1_simpleXor_308_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_307_port_z), .Z(ref_1_simpleXor_308_port_z) );
  XOR2_X1 ref_1_simpleXor_309_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_308_port_z), .Z(ref_1_simpleXor_309_port_z) );
  XOR2_X1 ref_1_simpleXor_310_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_309_port_z), .Z(ref_1_simpleXor_310_port_z) );
  XOR2_X1 ref_1_simpleXor_311_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_310_port_z), .Z(ref_1_refreshed_3_2_) );
  XOR2_X1 ref_1_simpleXor_312_U1 ( .A(port_rand_ref[0]), .B(port_b_0[3]), .Z(
        ref_1_simpleXor_312_port_z) );
  XOR2_X1 ref_1_simpleXor_313_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_312_port_z), .Z(ref_1_simpleXor_313_port_z) );
  XOR2_X1 ref_1_simpleXor_314_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_313_port_z), .Z(ref_1_simpleXor_314_port_z) );
  XOR2_X1 ref_1_simpleXor_315_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_314_port_z), .Z(ref_1_simpleXor_315_port_z) );
  XOR2_X1 ref_1_simpleXor_316_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_315_port_z), .Z(ref_1_simpleXor_316_port_z) );
  XOR2_X1 ref_1_simpleXor_317_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_316_port_z), .Z(ref_1_refreshed_0_3_) );
  XOR2_X1 ref_1_simpleXor_318_U1 ( .A(port_rand_ref[0]), .B(port_b_1[3]), .Z(
        ref_1_simpleXor_318_port_z) );
  XOR2_X1 ref_1_simpleXor_319_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_318_port_z), .Z(ref_1_simpleXor_319_port_z) );
  XOR2_X1 ref_1_simpleXor_320_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_319_port_z), .Z(ref_1_simpleXor_320_port_z) );
  XOR2_X1 ref_1_simpleXor_321_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_320_port_z), .Z(ref_1_simpleXor_321_port_z) );
  XOR2_X1 ref_1_simpleXor_322_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_321_port_z), .Z(ref_1_simpleXor_322_port_z) );
  XOR2_X1 ref_1_simpleXor_323_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_322_port_z), .Z(ref_1_refreshed_1_3_) );
  XOR2_X1 ref_1_simpleXor_324_U1 ( .A(port_rand_ref[2]), .B(port_b_2[3]), .Z(
        ref_1_simpleXor_324_port_z) );
  XOR2_X1 ref_1_simpleXor_325_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_324_port_z), .Z(ref_1_simpleXor_325_port_z) );
  XOR2_X1 ref_1_simpleXor_326_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_325_port_z), .Z(ref_1_simpleXor_326_port_z) );
  XOR2_X1 ref_1_simpleXor_327_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_326_port_z), .Z(ref_1_simpleXor_327_port_z) );
  XOR2_X1 ref_1_simpleXor_328_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_327_port_z), .Z(ref_1_simpleXor_328_port_z) );
  XOR2_X1 ref_1_simpleXor_329_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_328_port_z), .Z(ref_1_refreshed_2_3_) );
  XOR2_X1 ref_1_simpleXor_330_U1 ( .A(port_rand_ref[4]), .B(port_b_3[3]), .Z(
        ref_1_simpleXor_330_port_z) );
  XOR2_X1 ref_1_simpleXor_331_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_330_port_z), .Z(ref_1_simpleXor_331_port_z) );
  XOR2_X1 ref_1_simpleXor_332_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_331_port_z), .Z(ref_1_simpleXor_332_port_z) );
  XOR2_X1 ref_1_simpleXor_333_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_332_port_z), .Z(ref_1_simpleXor_333_port_z) );
  XOR2_X1 ref_1_simpleXor_334_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_333_port_z), .Z(ref_1_simpleXor_334_port_z) );
  XOR2_X1 ref_1_simpleXor_335_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_334_port_z), .Z(ref_1_refreshed_3_3_) );
  XOR2_X1 ref_1_simpleXor_336_U1 ( .A(port_rand_ref[0]), .B(port_b_0[4]), .Z(
        ref_1_simpleXor_336_port_z) );
  XOR2_X1 ref_1_simpleXor_337_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_336_port_z), .Z(ref_1_simpleXor_337_port_z) );
  XOR2_X1 ref_1_simpleXor_338_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_337_port_z), .Z(ref_1_simpleXor_338_port_z) );
  XOR2_X1 ref_1_simpleXor_339_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_338_port_z), .Z(ref_1_simpleXor_339_port_z) );
  XOR2_X1 ref_1_simpleXor_340_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_339_port_z), .Z(ref_1_simpleXor_340_port_z) );
  XOR2_X1 ref_1_simpleXor_341_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_340_port_z), .Z(ref_1_refreshed_0_4_) );
  XOR2_X1 ref_1_simpleXor_342_U1 ( .A(port_rand_ref[0]), .B(port_b_1[4]), .Z(
        ref_1_simpleXor_342_port_z) );
  XOR2_X1 ref_1_simpleXor_343_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_342_port_z), .Z(ref_1_simpleXor_343_port_z) );
  XOR2_X1 ref_1_simpleXor_344_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_343_port_z), .Z(ref_1_simpleXor_344_port_z) );
  XOR2_X1 ref_1_simpleXor_345_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_344_port_z), .Z(ref_1_simpleXor_345_port_z) );
  XOR2_X1 ref_1_simpleXor_346_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_345_port_z), .Z(ref_1_simpleXor_346_port_z) );
  XOR2_X1 ref_1_simpleXor_347_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_346_port_z), .Z(ref_1_refreshed_1_4_) );
  XOR2_X1 ref_1_simpleXor_348_U1 ( .A(port_rand_ref[2]), .B(port_b_2[4]), .Z(
        ref_1_simpleXor_348_port_z) );
  XOR2_X1 ref_1_simpleXor_349_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_348_port_z), .Z(ref_1_simpleXor_349_port_z) );
  XOR2_X1 ref_1_simpleXor_350_U1 ( .A(port_rand_ref[6]), .B(
        ref_1_simpleXor_349_port_z), .Z(ref_1_simpleXor_350_port_z) );
  XOR2_X1 ref_1_simpleXor_351_U1 ( .A(port_rand_ref[7]), .B(
        ref_1_simpleXor_350_port_z), .Z(ref_1_simpleXor_351_port_z) );
  XOR2_X1 ref_1_simpleXor_352_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_351_port_z), .Z(ref_1_simpleXor_352_port_z) );
  XOR2_X1 ref_1_simpleXor_353_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_352_port_z), .Z(ref_1_refreshed_2_4_) );
  XOR2_X1 ref_1_simpleXor_354_U1 ( .A(port_rand_ref[4]), .B(port_b_3[4]), .Z(
        ref_1_simpleXor_354_port_z) );
  XOR2_X1 ref_1_simpleXor_355_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_354_port_z), .Z(ref_1_simpleXor_355_port_z) );
  XOR2_X1 ref_1_simpleXor_356_U1 ( .A(port_rand_ref[8]), .B(
        ref_1_simpleXor_355_port_z), .Z(ref_1_simpleXor_356_port_z) );
  XOR2_X1 ref_1_simpleXor_357_U1 ( .A(port_rand_ref[9]), .B(
        ref_1_simpleXor_356_port_z), .Z(ref_1_simpleXor_357_port_z) );
  XOR2_X1 ref_1_simpleXor_358_U1 ( .A(port_rand_ref[10]), .B(
        ref_1_simpleXor_357_port_z), .Z(ref_1_simpleXor_358_port_z) );
  XOR2_X1 ref_1_simpleXor_359_U1 ( .A(port_rand_ref[11]), .B(
        ref_1_simpleXor_358_port_z), .Z(ref_1_refreshed_3_4_) );
  NAND2_X1 ref_1_maj_80_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_80_n9) );
  NAND2_X1 ref_1_maj_80_U14 ( .A1(ref_1_maj_80_n6), .A2(ref_1_maj_80_n5), .ZN(
        ref_1_maj_80_n10) );
  NAND2_X1 ref_1_maj_80_U13 ( .A1(ref_1_maj_80_n9), .A2(ref_1_maj_80_n10), 
        .ZN(ref_1_maj_80_n8) );
  NAND2_X1 ref_1_maj_80_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_80_n11), .ZN(
        ref_1_maj_80_n13) );
  NAND2_X1 ref_1_maj_80_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_80_n12) );
  NAND2_X1 ref_1_maj_80_U10 ( .A1(ref_1_maj_80_n12), .A2(ref_1_maj_80_n13), 
        .ZN(ref_1_maj_80_n7) );
  XOR2_X1 ref_1_maj_80_U9 ( .A(ref_1_n36), .B(ref_1_maj_80_n11), .Z(
        ref_1_maj_80_n6) );
  XOR2_X1 ref_1_maj_80_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_80_n5)
         );
  XOR2_X1 ref_1_maj_80_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_80_n11)
         );
  OR2_X1 ref_1_maj_80_U6 ( .A1(ref_1_maj_80_n7), .A2(ref_1_maj_80_n8), .ZN(
        ref_1_maj_80_n3) );
  NAND2_X1 ref_1_maj_80_U5 ( .A1(ref_1_maj_80_n3), .A2(ref_1_maj_80_n4), .ZN(
        ref_1_maj_80_n2) );
  NAND2_X1 ref_1_maj_80_U4 ( .A1(ref_1_maj_80_n7), .A2(ref_1_maj_80_n8), .ZN(
        ref_1_maj_80_n1) );
  NAND2_X1 ref_1_maj_80_U3 ( .A1(ref_1_maj_80_n1), .A2(ref_1_maj_80_n2), .ZN(
        ref_1_maj_80_port_o) );
  XOR2_X1 ref_1_maj_80_U2 ( .A(ref_1_maj_80_n5), .B(ref_1_maj_80_n6), .Z(
        ref_1_maj_80_n4) );
  NAND2_X1 ref_1_maj_81_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_81_n18) );
  NAND2_X1 ref_1_maj_81_U14 ( .A1(ref_1_maj_81_n21), .A2(ref_1_maj_81_n22), 
        .ZN(ref_1_maj_81_n17) );
  NAND2_X1 ref_1_maj_81_U13 ( .A1(ref_1_maj_81_n18), .A2(ref_1_maj_81_n17), 
        .ZN(ref_1_maj_81_n19) );
  NAND2_X1 ref_1_maj_81_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_81_n16), .ZN(
        ref_1_maj_81_n14) );
  NAND2_X1 ref_1_maj_81_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_81_n15) );
  NAND2_X1 ref_1_maj_81_U10 ( .A1(ref_1_maj_81_n15), .A2(ref_1_maj_81_n14), 
        .ZN(ref_1_maj_81_n20) );
  XOR2_X1 ref_1_maj_81_U9 ( .A(ref_1_n36), .B(ref_1_maj_81_n16), .Z(
        ref_1_maj_81_n21) );
  XOR2_X1 ref_1_maj_81_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_81_n22)
         );
  XOR2_X1 ref_1_maj_81_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_81_n16)
         );
  OR2_X1 ref_1_maj_81_U6 ( .A1(ref_1_maj_81_n20), .A2(ref_1_maj_81_n19), .ZN(
        ref_1_maj_81_n24) );
  NAND2_X1 ref_1_maj_81_U5 ( .A1(ref_1_maj_81_n24), .A2(ref_1_maj_81_n23), 
        .ZN(ref_1_maj_81_n25) );
  NAND2_X1 ref_1_maj_81_U4 ( .A1(ref_1_maj_81_n20), .A2(ref_1_maj_81_n19), 
        .ZN(ref_1_maj_81_n26) );
  NAND2_X1 ref_1_maj_81_U3 ( .A1(ref_1_maj_81_n26), .A2(ref_1_maj_81_n25), 
        .ZN(ref_1_maj_81_port_o) );
  XOR2_X1 ref_1_maj_81_U2 ( .A(ref_1_maj_81_n22), .B(ref_1_maj_81_n21), .Z(
        ref_1_maj_81_n23) );
  NAND2_X1 ref_1_maj_82_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_82_n18) );
  NAND2_X1 ref_1_maj_82_U14 ( .A1(ref_1_maj_82_n21), .A2(ref_1_maj_82_n22), 
        .ZN(ref_1_maj_82_n17) );
  NAND2_X1 ref_1_maj_82_U13 ( .A1(ref_1_maj_82_n18), .A2(ref_1_maj_82_n17), 
        .ZN(ref_1_maj_82_n19) );
  NAND2_X1 ref_1_maj_82_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_82_n16), 
        .ZN(ref_1_maj_82_n14) );
  NAND2_X1 ref_1_maj_82_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_82_n15) );
  NAND2_X1 ref_1_maj_82_U10 ( .A1(ref_1_maj_82_n15), .A2(ref_1_maj_82_n14), 
        .ZN(ref_1_maj_82_n20) );
  XOR2_X1 ref_1_maj_82_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_82_n16), 
        .Z(ref_1_maj_82_n21) );
  XOR2_X1 ref_1_maj_82_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_82_n22) );
  XOR2_X1 ref_1_maj_82_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), 
        .Z(ref_1_maj_82_n16) );
  OR2_X1 ref_1_maj_82_U6 ( .A1(ref_1_maj_82_n20), .A2(ref_1_maj_82_n19), .ZN(
        ref_1_maj_82_n24) );
  NAND2_X1 ref_1_maj_82_U5 ( .A1(ref_1_maj_82_n24), .A2(ref_1_maj_82_n23), 
        .ZN(ref_1_maj_82_n25) );
  NAND2_X1 ref_1_maj_82_U4 ( .A1(ref_1_maj_82_n20), .A2(ref_1_maj_82_n19), 
        .ZN(ref_1_maj_82_n26) );
  NAND2_X1 ref_1_maj_82_U3 ( .A1(ref_1_maj_82_n26), .A2(ref_1_maj_82_n25), 
        .ZN(ref_1_maj_82_port_o) );
  XOR2_X1 ref_1_maj_82_U2 ( .A(ref_1_maj_82_n22), .B(ref_1_maj_82_n21), .Z(
        ref_1_maj_82_n23) );
  NAND2_X1 ref_1_maj_83_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_83_n18) );
  NAND2_X1 ref_1_maj_83_U14 ( .A1(ref_1_maj_83_n21), .A2(ref_1_maj_83_n22), 
        .ZN(ref_1_maj_83_n17) );
  NAND2_X1 ref_1_maj_83_U13 ( .A1(ref_1_maj_83_n18), .A2(ref_1_maj_83_n17), 
        .ZN(ref_1_maj_83_n19) );
  NAND2_X1 ref_1_maj_83_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_83_n16), 
        .ZN(ref_1_maj_83_n14) );
  NAND2_X1 ref_1_maj_83_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_83_n15) );
  NAND2_X1 ref_1_maj_83_U10 ( .A1(ref_1_maj_83_n15), .A2(ref_1_maj_83_n14), 
        .ZN(ref_1_maj_83_n20) );
  XOR2_X1 ref_1_maj_83_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_83_n16), 
        .Z(ref_1_maj_83_n21) );
  XOR2_X1 ref_1_maj_83_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_83_n22) );
  XOR2_X1 ref_1_maj_83_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), 
        .Z(ref_1_maj_83_n16) );
  OR2_X1 ref_1_maj_83_U6 ( .A1(ref_1_maj_83_n20), .A2(ref_1_maj_83_n19), .ZN(
        ref_1_maj_83_n24) );
  NAND2_X1 ref_1_maj_83_U5 ( .A1(ref_1_maj_83_n24), .A2(ref_1_maj_83_n23), 
        .ZN(ref_1_maj_83_n25) );
  NAND2_X1 ref_1_maj_83_U4 ( .A1(ref_1_maj_83_n20), .A2(ref_1_maj_83_n19), 
        .ZN(ref_1_maj_83_n26) );
  NAND2_X1 ref_1_maj_83_U3 ( .A1(ref_1_maj_83_n26), .A2(ref_1_maj_83_n25), 
        .ZN(ref_1_maj_83_port_o) );
  XOR2_X1 ref_1_maj_83_U2 ( .A(ref_1_maj_83_n22), .B(ref_1_maj_83_n21), .Z(
        ref_1_maj_83_n23) );
  NAND2_X1 ref_1_maj_84_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_84_n18) );
  NAND2_X1 ref_1_maj_84_U14 ( .A1(ref_1_maj_84_n21), .A2(ref_1_maj_84_n22), 
        .ZN(ref_1_maj_84_n17) );
  NAND2_X1 ref_1_maj_84_U13 ( .A1(ref_1_maj_84_n18), .A2(ref_1_maj_84_n17), 
        .ZN(ref_1_maj_84_n19) );
  NAND2_X1 ref_1_maj_84_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_84_n16), .ZN(
        ref_1_maj_84_n14) );
  NAND2_X1 ref_1_maj_84_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_84_n15) );
  NAND2_X1 ref_1_maj_84_U10 ( .A1(ref_1_maj_84_n15), .A2(ref_1_maj_84_n14), 
        .ZN(ref_1_maj_84_n20) );
  XOR2_X1 ref_1_maj_84_U9 ( .A(ref_1_n26), .B(ref_1_maj_84_n16), .Z(
        ref_1_maj_84_n21) );
  XOR2_X1 ref_1_maj_84_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_84_n22)
         );
  XOR2_X1 ref_1_maj_84_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(ref_1_maj_84_n16)
         );
  OR2_X1 ref_1_maj_84_U6 ( .A1(ref_1_maj_84_n20), .A2(ref_1_maj_84_n19), .ZN(
        ref_1_maj_84_n24) );
  NAND2_X1 ref_1_maj_84_U5 ( .A1(ref_1_maj_84_n24), .A2(ref_1_maj_84_n23), 
        .ZN(ref_1_maj_84_n25) );
  NAND2_X1 ref_1_maj_84_U4 ( .A1(ref_1_maj_84_n20), .A2(ref_1_maj_84_n19), 
        .ZN(ref_1_maj_84_n26) );
  NAND2_X1 ref_1_maj_84_U3 ( .A1(ref_1_maj_84_n26), .A2(ref_1_maj_84_n25), 
        .ZN(ref_1_maj_84_port_o) );
  XOR2_X1 ref_1_maj_84_U2 ( .A(ref_1_maj_84_n22), .B(ref_1_maj_84_n21), .Z(
        ref_1_maj_84_n23) );
  NAND2_X1 ref_1_maj_85_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_85_n18) );
  NAND2_X1 ref_1_maj_85_U14 ( .A1(ref_1_maj_85_n21), .A2(ref_1_maj_85_n22), 
        .ZN(ref_1_maj_85_n17) );
  NAND2_X1 ref_1_maj_85_U13 ( .A1(ref_1_maj_85_n18), .A2(ref_1_maj_85_n17), 
        .ZN(ref_1_maj_85_n19) );
  NAND2_X1 ref_1_maj_85_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_85_n16), 
        .ZN(ref_1_maj_85_n14) );
  NAND2_X1 ref_1_maj_85_U11 ( .A1(ref_1_refreshed_1_0_), .A2(
        ref_1_refreshed_1_1_), .ZN(ref_1_maj_85_n15) );
  NAND2_X1 ref_1_maj_85_U10 ( .A1(ref_1_maj_85_n15), .A2(ref_1_maj_85_n14), 
        .ZN(ref_1_maj_85_n20) );
  XOR2_X1 ref_1_maj_85_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_85_n16), 
        .Z(ref_1_maj_85_n21) );
  XOR2_X1 ref_1_maj_85_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_85_n22) );
  XOR2_X1 ref_1_maj_85_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_refreshed_1_1_), 
        .Z(ref_1_maj_85_n16) );
  OR2_X1 ref_1_maj_85_U6 ( .A1(ref_1_maj_85_n20), .A2(ref_1_maj_85_n19), .ZN(
        ref_1_maj_85_n24) );
  NAND2_X1 ref_1_maj_85_U5 ( .A1(ref_1_maj_85_n24), .A2(ref_1_maj_85_n23), 
        .ZN(ref_1_maj_85_n25) );
  NAND2_X1 ref_1_maj_85_U4 ( .A1(ref_1_maj_85_n20), .A2(ref_1_maj_85_n19), 
        .ZN(ref_1_maj_85_n26) );
  NAND2_X1 ref_1_maj_85_U3 ( .A1(ref_1_maj_85_n26), .A2(ref_1_maj_85_n25), 
        .ZN(ref_1_maj_85_port_o) );
  XOR2_X1 ref_1_maj_85_U2 ( .A(ref_1_maj_85_n22), .B(ref_1_maj_85_n21), .Z(
        ref_1_maj_85_n23) );
  NAND2_X1 ref_1_maj_86_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_86_n18) );
  NAND2_X1 ref_1_maj_86_U14 ( .A1(ref_1_maj_86_n21), .A2(ref_1_maj_86_n22), 
        .ZN(ref_1_maj_86_n17) );
  NAND2_X1 ref_1_maj_86_U13 ( .A1(ref_1_maj_86_n18), .A2(ref_1_maj_86_n17), 
        .ZN(ref_1_maj_86_n19) );
  NAND2_X1 ref_1_maj_86_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_86_n16), 
        .ZN(ref_1_maj_86_n14) );
  NAND2_X1 ref_1_maj_86_U11 ( .A1(ref_1_refreshed_1_0_), .A2(
        ref_1_refreshed_1_1_), .ZN(ref_1_maj_86_n15) );
  NAND2_X1 ref_1_maj_86_U10 ( .A1(ref_1_maj_86_n15), .A2(ref_1_maj_86_n14), 
        .ZN(ref_1_maj_86_n20) );
  XOR2_X1 ref_1_maj_86_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_86_n16), 
        .Z(ref_1_maj_86_n21) );
  XOR2_X1 ref_1_maj_86_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_86_n22) );
  XOR2_X1 ref_1_maj_86_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_refreshed_1_1_), 
        .Z(ref_1_maj_86_n16) );
  OR2_X1 ref_1_maj_86_U6 ( .A1(ref_1_maj_86_n20), .A2(ref_1_maj_86_n19), .ZN(
        ref_1_maj_86_n24) );
  NAND2_X1 ref_1_maj_86_U5 ( .A1(ref_1_maj_86_n24), .A2(ref_1_maj_86_n23), 
        .ZN(ref_1_maj_86_n25) );
  NAND2_X1 ref_1_maj_86_U4 ( .A1(ref_1_maj_86_n20), .A2(ref_1_maj_86_n19), 
        .ZN(ref_1_maj_86_n26) );
  NAND2_X1 ref_1_maj_86_U3 ( .A1(ref_1_maj_86_n26), .A2(ref_1_maj_86_n25), 
        .ZN(ref_1_maj_86_port_o) );
  XOR2_X1 ref_1_maj_86_U2 ( .A(ref_1_maj_86_n22), .B(ref_1_maj_86_n21), .Z(
        ref_1_maj_86_n23) );
  NAND2_X1 ref_1_maj_87_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_87_n18) );
  NAND2_X1 ref_1_maj_87_U14 ( .A1(ref_1_maj_87_n21), .A2(ref_1_maj_87_n22), 
        .ZN(ref_1_maj_87_n17) );
  NAND2_X1 ref_1_maj_87_U13 ( .A1(ref_1_maj_87_n18), .A2(ref_1_maj_87_n17), 
        .ZN(ref_1_maj_87_n19) );
  NAND2_X1 ref_1_maj_87_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_87_n16), 
        .ZN(ref_1_maj_87_n14) );
  NAND2_X1 ref_1_maj_87_U11 ( .A1(ref_1_refreshed_1_0_), .A2(
        ref_1_refreshed_1_1_), .ZN(ref_1_maj_87_n15) );
  NAND2_X1 ref_1_maj_87_U10 ( .A1(ref_1_maj_87_n15), .A2(ref_1_maj_87_n14), 
        .ZN(ref_1_maj_87_n20) );
  XOR2_X1 ref_1_maj_87_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_87_n16), 
        .Z(ref_1_maj_87_n21) );
  XOR2_X1 ref_1_maj_87_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_87_n22) );
  XOR2_X1 ref_1_maj_87_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_refreshed_1_1_), 
        .Z(ref_1_maj_87_n16) );
  OR2_X1 ref_1_maj_87_U6 ( .A1(ref_1_maj_87_n20), .A2(ref_1_maj_87_n19), .ZN(
        ref_1_maj_87_n24) );
  NAND2_X1 ref_1_maj_87_U5 ( .A1(ref_1_maj_87_n24), .A2(ref_1_maj_87_n23), 
        .ZN(ref_1_maj_87_n25) );
  NAND2_X1 ref_1_maj_87_U4 ( .A1(ref_1_maj_87_n20), .A2(ref_1_maj_87_n19), 
        .ZN(ref_1_maj_87_n26) );
  NAND2_X1 ref_1_maj_87_U3 ( .A1(ref_1_maj_87_n26), .A2(ref_1_maj_87_n25), 
        .ZN(ref_1_maj_87_port_o) );
  XOR2_X1 ref_1_maj_87_U2 ( .A(ref_1_maj_87_n22), .B(ref_1_maj_87_n21), .Z(
        ref_1_maj_87_n23) );
  NAND2_X1 ref_1_maj_88_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_88_n18) );
  NAND2_X1 ref_1_maj_88_U14 ( .A1(ref_1_maj_88_n21), .A2(ref_1_maj_88_n22), 
        .ZN(ref_1_maj_88_n17) );
  NAND2_X1 ref_1_maj_88_U13 ( .A1(ref_1_maj_88_n18), .A2(ref_1_maj_88_n17), 
        .ZN(ref_1_maj_88_n19) );
  NAND2_X1 ref_1_maj_88_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_88_n16), .ZN(
        ref_1_maj_88_n14) );
  NAND2_X1 ref_1_maj_88_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_88_n15) );
  NAND2_X1 ref_1_maj_88_U10 ( .A1(ref_1_maj_88_n15), .A2(ref_1_maj_88_n14), 
        .ZN(ref_1_maj_88_n20) );
  XOR2_X1 ref_1_maj_88_U9 ( .A(ref_1_n16), .B(ref_1_maj_88_n16), .Z(
        ref_1_maj_88_n21) );
  XOR2_X1 ref_1_maj_88_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_88_n22)
         );
  XOR2_X1 ref_1_maj_88_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(ref_1_maj_88_n16)
         );
  OR2_X1 ref_1_maj_88_U6 ( .A1(ref_1_maj_88_n20), .A2(ref_1_maj_88_n19), .ZN(
        ref_1_maj_88_n24) );
  NAND2_X1 ref_1_maj_88_U5 ( .A1(ref_1_maj_88_n24), .A2(ref_1_maj_88_n23), 
        .ZN(ref_1_maj_88_n25) );
  NAND2_X1 ref_1_maj_88_U4 ( .A1(ref_1_maj_88_n20), .A2(ref_1_maj_88_n19), 
        .ZN(ref_1_maj_88_n26) );
  NAND2_X1 ref_1_maj_88_U3 ( .A1(ref_1_maj_88_n26), .A2(ref_1_maj_88_n25), 
        .ZN(ref_1_maj_88_port_o) );
  XOR2_X1 ref_1_maj_88_U2 ( .A(ref_1_maj_88_n22), .B(ref_1_maj_88_n21), .Z(
        ref_1_maj_88_n23) );
  NAND2_X1 ref_1_maj_89_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_89_n18) );
  NAND2_X1 ref_1_maj_89_U14 ( .A1(ref_1_maj_89_n21), .A2(ref_1_maj_89_n22), 
        .ZN(ref_1_maj_89_n17) );
  NAND2_X1 ref_1_maj_89_U13 ( .A1(ref_1_maj_89_n18), .A2(ref_1_maj_89_n17), 
        .ZN(ref_1_maj_89_n19) );
  NAND2_X1 ref_1_maj_89_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_89_n16), 
        .ZN(ref_1_maj_89_n14) );
  NAND2_X1 ref_1_maj_89_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_89_n15) );
  NAND2_X1 ref_1_maj_89_U10 ( .A1(ref_1_maj_89_n15), .A2(ref_1_maj_89_n14), 
        .ZN(ref_1_maj_89_n20) );
  XOR2_X1 ref_1_maj_89_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_89_n16), 
        .Z(ref_1_maj_89_n21) );
  XOR2_X1 ref_1_maj_89_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_89_n22) );
  XOR2_X1 ref_1_maj_89_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), 
        .Z(ref_1_maj_89_n16) );
  OR2_X1 ref_1_maj_89_U6 ( .A1(ref_1_maj_89_n20), .A2(ref_1_maj_89_n19), .ZN(
        ref_1_maj_89_n24) );
  NAND2_X1 ref_1_maj_89_U5 ( .A1(ref_1_maj_89_n24), .A2(ref_1_maj_89_n23), 
        .ZN(ref_1_maj_89_n25) );
  NAND2_X1 ref_1_maj_89_U4 ( .A1(ref_1_maj_89_n20), .A2(ref_1_maj_89_n19), 
        .ZN(ref_1_maj_89_n26) );
  NAND2_X1 ref_1_maj_89_U3 ( .A1(ref_1_maj_89_n26), .A2(ref_1_maj_89_n25), 
        .ZN(ref_1_maj_89_port_o) );
  XOR2_X1 ref_1_maj_89_U2 ( .A(ref_1_maj_89_n22), .B(ref_1_maj_89_n21), .Z(
        ref_1_maj_89_n23) );
  NAND2_X1 ref_1_maj_90_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_90_n18) );
  NAND2_X1 ref_1_maj_90_U14 ( .A1(ref_1_maj_90_n21), .A2(ref_1_maj_90_n22), 
        .ZN(ref_1_maj_90_n17) );
  NAND2_X1 ref_1_maj_90_U13 ( .A1(ref_1_maj_90_n18), .A2(ref_1_maj_90_n17), 
        .ZN(ref_1_maj_90_n19) );
  NAND2_X1 ref_1_maj_90_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_90_n16), 
        .ZN(ref_1_maj_90_n14) );
  NAND2_X1 ref_1_maj_90_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_90_n15) );
  NAND2_X1 ref_1_maj_90_U10 ( .A1(ref_1_maj_90_n15), .A2(ref_1_maj_90_n14), 
        .ZN(ref_1_maj_90_n20) );
  XOR2_X1 ref_1_maj_90_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_90_n16), 
        .Z(ref_1_maj_90_n21) );
  XOR2_X1 ref_1_maj_90_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_90_n22) );
  XOR2_X1 ref_1_maj_90_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), 
        .Z(ref_1_maj_90_n16) );
  OR2_X1 ref_1_maj_90_U6 ( .A1(ref_1_maj_90_n20), .A2(ref_1_maj_90_n19), .ZN(
        ref_1_maj_90_n24) );
  NAND2_X1 ref_1_maj_90_U5 ( .A1(ref_1_maj_90_n24), .A2(ref_1_maj_90_n23), 
        .ZN(ref_1_maj_90_n25) );
  NAND2_X1 ref_1_maj_90_U4 ( .A1(ref_1_maj_90_n20), .A2(ref_1_maj_90_n19), 
        .ZN(ref_1_maj_90_n26) );
  NAND2_X1 ref_1_maj_90_U3 ( .A1(ref_1_maj_90_n26), .A2(ref_1_maj_90_n25), 
        .ZN(ref_1_maj_90_port_o) );
  XOR2_X1 ref_1_maj_90_U2 ( .A(ref_1_maj_90_n22), .B(ref_1_maj_90_n21), .Z(
        ref_1_maj_90_n23) );
  NAND2_X1 ref_1_maj_91_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_91_n18) );
  NAND2_X1 ref_1_maj_91_U14 ( .A1(ref_1_maj_91_n21), .A2(ref_1_maj_91_n22), 
        .ZN(ref_1_maj_91_n17) );
  NAND2_X1 ref_1_maj_91_U13 ( .A1(ref_1_maj_91_n18), .A2(ref_1_maj_91_n17), 
        .ZN(ref_1_maj_91_n19) );
  NAND2_X1 ref_1_maj_91_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_91_n16), 
        .ZN(ref_1_maj_91_n14) );
  NAND2_X1 ref_1_maj_91_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_91_n15) );
  NAND2_X1 ref_1_maj_91_U10 ( .A1(ref_1_maj_91_n15), .A2(ref_1_maj_91_n14), 
        .ZN(ref_1_maj_91_n20) );
  XOR2_X1 ref_1_maj_91_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_91_n16), 
        .Z(ref_1_maj_91_n21) );
  XOR2_X1 ref_1_maj_91_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_91_n22) );
  XOR2_X1 ref_1_maj_91_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), 
        .Z(ref_1_maj_91_n16) );
  OR2_X1 ref_1_maj_91_U6 ( .A1(ref_1_maj_91_n20), .A2(ref_1_maj_91_n19), .ZN(
        ref_1_maj_91_n24) );
  NAND2_X1 ref_1_maj_91_U5 ( .A1(ref_1_maj_91_n24), .A2(ref_1_maj_91_n23), 
        .ZN(ref_1_maj_91_n25) );
  NAND2_X1 ref_1_maj_91_U4 ( .A1(ref_1_maj_91_n20), .A2(ref_1_maj_91_n19), 
        .ZN(ref_1_maj_91_n26) );
  NAND2_X1 ref_1_maj_91_U3 ( .A1(ref_1_maj_91_n26), .A2(ref_1_maj_91_n25), 
        .ZN(ref_1_maj_91_port_o) );
  XOR2_X1 ref_1_maj_91_U2 ( .A(ref_1_maj_91_n22), .B(ref_1_maj_91_n21), .Z(
        ref_1_maj_91_n23) );
  NAND2_X1 ref_1_maj_92_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_92_n18) );
  NAND2_X1 ref_1_maj_92_U14 ( .A1(ref_1_maj_92_n21), .A2(ref_1_maj_92_n22), 
        .ZN(ref_1_maj_92_n17) );
  NAND2_X1 ref_1_maj_92_U13 ( .A1(ref_1_maj_92_n18), .A2(ref_1_maj_92_n17), 
        .ZN(ref_1_maj_92_n19) );
  NAND2_X1 ref_1_maj_92_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_92_n16), .ZN(
        ref_1_maj_92_n14) );
  NAND2_X1 ref_1_maj_92_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_92_n15) );
  NAND2_X1 ref_1_maj_92_U10 ( .A1(ref_1_maj_92_n15), .A2(ref_1_maj_92_n14), 
        .ZN(ref_1_maj_92_n20) );
  XOR2_X1 ref_1_maj_92_U9 ( .A(ref_1_n6), .B(ref_1_maj_92_n16), .Z(
        ref_1_maj_92_n21) );
  XOR2_X1 ref_1_maj_92_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_92_n22)
         );
  XOR2_X1 ref_1_maj_92_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_92_n16)
         );
  OR2_X1 ref_1_maj_92_U6 ( .A1(ref_1_maj_92_n20), .A2(ref_1_maj_92_n19), .ZN(
        ref_1_maj_92_n24) );
  NAND2_X1 ref_1_maj_92_U5 ( .A1(ref_1_maj_92_n24), .A2(ref_1_maj_92_n23), 
        .ZN(ref_1_maj_92_n25) );
  NAND2_X1 ref_1_maj_92_U4 ( .A1(ref_1_maj_92_n20), .A2(ref_1_maj_92_n19), 
        .ZN(ref_1_maj_92_n26) );
  NAND2_X1 ref_1_maj_92_U3 ( .A1(ref_1_maj_92_n26), .A2(ref_1_maj_92_n25), 
        .ZN(ref_1_maj_92_port_o) );
  XOR2_X1 ref_1_maj_92_U2 ( .A(ref_1_maj_92_n22), .B(ref_1_maj_92_n21), .Z(
        ref_1_maj_92_n23) );
  NAND2_X1 ref_1_maj_93_U15 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_93_n18) );
  NAND2_X1 ref_1_maj_93_U14 ( .A1(ref_1_maj_93_n21), .A2(ref_1_maj_93_n22), 
        .ZN(ref_1_maj_93_n17) );
  NAND2_X1 ref_1_maj_93_U13 ( .A1(ref_1_maj_93_n18), .A2(ref_1_maj_93_n17), 
        .ZN(ref_1_maj_93_n19) );
  NAND2_X1 ref_1_maj_93_U12 ( .A1(ref_1_refreshed_3_2_), .A2(ref_1_maj_93_n16), 
        .ZN(ref_1_maj_93_n14) );
  NAND2_X1 ref_1_maj_93_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_93_n15) );
  NAND2_X1 ref_1_maj_93_U10 ( .A1(ref_1_maj_93_n15), .A2(ref_1_maj_93_n14), 
        .ZN(ref_1_maj_93_n20) );
  XOR2_X1 ref_1_maj_93_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_93_n16), 
        .Z(ref_1_maj_93_n21) );
  XOR2_X1 ref_1_maj_93_U8 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), 
        .Z(ref_1_maj_93_n22) );
  XOR2_X1 ref_1_maj_93_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), 
        .Z(ref_1_maj_93_n16) );
  OR2_X1 ref_1_maj_93_U6 ( .A1(ref_1_maj_93_n20), .A2(ref_1_maj_93_n19), .ZN(
        ref_1_maj_93_n24) );
  NAND2_X1 ref_1_maj_93_U5 ( .A1(ref_1_maj_93_n24), .A2(ref_1_maj_93_n23), 
        .ZN(ref_1_maj_93_n25) );
  NAND2_X1 ref_1_maj_93_U4 ( .A1(ref_1_maj_93_n20), .A2(ref_1_maj_93_n19), 
        .ZN(ref_1_maj_93_n26) );
  NAND2_X1 ref_1_maj_93_U3 ( .A1(ref_1_maj_93_n26), .A2(ref_1_maj_93_n25), 
        .ZN(ref_1_maj_93_port_o) );
  XOR2_X1 ref_1_maj_93_U2 ( .A(ref_1_maj_93_n22), .B(ref_1_maj_93_n21), .Z(
        ref_1_maj_93_n23) );
  NAND2_X1 ref_1_maj_94_U15 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_94_n18) );
  NAND2_X1 ref_1_maj_94_U14 ( .A1(ref_1_maj_94_n21), .A2(ref_1_maj_94_n22), 
        .ZN(ref_1_maj_94_n17) );
  NAND2_X1 ref_1_maj_94_U13 ( .A1(ref_1_maj_94_n18), .A2(ref_1_maj_94_n17), 
        .ZN(ref_1_maj_94_n19) );
  NAND2_X1 ref_1_maj_94_U12 ( .A1(ref_1_refreshed_3_2_), .A2(ref_1_maj_94_n16), 
        .ZN(ref_1_maj_94_n14) );
  NAND2_X1 ref_1_maj_94_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_94_n15) );
  NAND2_X1 ref_1_maj_94_U10 ( .A1(ref_1_maj_94_n15), .A2(ref_1_maj_94_n14), 
        .ZN(ref_1_maj_94_n20) );
  XOR2_X1 ref_1_maj_94_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_94_n16), 
        .Z(ref_1_maj_94_n21) );
  XOR2_X1 ref_1_maj_94_U8 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), 
        .Z(ref_1_maj_94_n22) );
  XOR2_X1 ref_1_maj_94_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), 
        .Z(ref_1_maj_94_n16) );
  OR2_X1 ref_1_maj_94_U6 ( .A1(ref_1_maj_94_n20), .A2(ref_1_maj_94_n19), .ZN(
        ref_1_maj_94_n24) );
  NAND2_X1 ref_1_maj_94_U5 ( .A1(ref_1_maj_94_n24), .A2(ref_1_maj_94_n23), 
        .ZN(ref_1_maj_94_n25) );
  NAND2_X1 ref_1_maj_94_U4 ( .A1(ref_1_maj_94_n20), .A2(ref_1_maj_94_n19), 
        .ZN(ref_1_maj_94_n26) );
  NAND2_X1 ref_1_maj_94_U3 ( .A1(ref_1_maj_94_n26), .A2(ref_1_maj_94_n25), 
        .ZN(ref_1_maj_94_port_o) );
  XOR2_X1 ref_1_maj_94_U2 ( .A(ref_1_maj_94_n22), .B(ref_1_maj_94_n21), .Z(
        ref_1_maj_94_n23) );
  NAND2_X1 ref_1_maj_95_U15 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_95_n18) );
  NAND2_X1 ref_1_maj_95_U14 ( .A1(ref_1_maj_95_n21), .A2(ref_1_maj_95_n22), 
        .ZN(ref_1_maj_95_n17) );
  NAND2_X1 ref_1_maj_95_U13 ( .A1(ref_1_maj_95_n18), .A2(ref_1_maj_95_n17), 
        .ZN(ref_1_maj_95_n19) );
  NAND2_X1 ref_1_maj_95_U12 ( .A1(ref_1_refreshed_3_2_), .A2(ref_1_maj_95_n16), 
        .ZN(ref_1_maj_95_n14) );
  NAND2_X1 ref_1_maj_95_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_95_n15) );
  NAND2_X1 ref_1_maj_95_U10 ( .A1(ref_1_maj_95_n15), .A2(ref_1_maj_95_n14), 
        .ZN(ref_1_maj_95_n20) );
  XOR2_X1 ref_1_maj_95_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_95_n16), 
        .Z(ref_1_maj_95_n21) );
  XOR2_X1 ref_1_maj_95_U8 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), 
        .Z(ref_1_maj_95_n22) );
  XOR2_X1 ref_1_maj_95_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), 
        .Z(ref_1_maj_95_n16) );
  OR2_X1 ref_1_maj_95_U6 ( .A1(ref_1_maj_95_n20), .A2(ref_1_maj_95_n19), .ZN(
        ref_1_maj_95_n24) );
  NAND2_X1 ref_1_maj_95_U5 ( .A1(ref_1_maj_95_n24), .A2(ref_1_maj_95_n23), 
        .ZN(ref_1_maj_95_n25) );
  NAND2_X1 ref_1_maj_95_U4 ( .A1(ref_1_maj_95_n20), .A2(ref_1_maj_95_n19), 
        .ZN(ref_1_maj_95_n26) );
  NAND2_X1 ref_1_maj_95_U3 ( .A1(ref_1_maj_95_n26), .A2(ref_1_maj_95_n25), 
        .ZN(ref_1_maj_95_port_o) );
  XOR2_X1 ref_1_maj_95_U2 ( .A(ref_1_maj_95_n22), .B(ref_1_maj_95_n21), .Z(
        ref_1_maj_95_n23) );
  NAND2_X1 ref_1_maj_96_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_96_n18) );
  NAND2_X1 ref_1_maj_96_U14 ( .A1(ref_1_maj_96_n21), .A2(ref_1_maj_96_n22), 
        .ZN(ref_1_maj_96_n17) );
  NAND2_X1 ref_1_maj_96_U13 ( .A1(ref_1_maj_96_n18), .A2(ref_1_maj_96_n17), 
        .ZN(ref_1_maj_96_n19) );
  NAND2_X1 ref_1_maj_96_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_96_n16), 
        .ZN(ref_1_maj_96_n14) );
  NAND2_X1 ref_1_maj_96_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_96_n15) );
  NAND2_X1 ref_1_maj_96_U10 ( .A1(ref_1_maj_96_n15), .A2(ref_1_maj_96_n14), 
        .ZN(ref_1_maj_96_n20) );
  XOR2_X1 ref_1_maj_96_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_96_n16), 
        .Z(ref_1_maj_96_n21) );
  XOR2_X1 ref_1_maj_96_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_96_n22) );
  XOR2_X1 ref_1_maj_96_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), 
        .Z(ref_1_maj_96_n16) );
  OR2_X1 ref_1_maj_96_U6 ( .A1(ref_1_maj_96_n20), .A2(ref_1_maj_96_n19), .ZN(
        ref_1_maj_96_n24) );
  NAND2_X1 ref_1_maj_96_U5 ( .A1(ref_1_maj_96_n24), .A2(ref_1_maj_96_n23), 
        .ZN(ref_1_maj_96_n25) );
  NAND2_X1 ref_1_maj_96_U4 ( .A1(ref_1_maj_96_n20), .A2(ref_1_maj_96_n19), 
        .ZN(ref_1_maj_96_n26) );
  NAND2_X1 ref_1_maj_96_U3 ( .A1(ref_1_maj_96_n26), .A2(ref_1_maj_96_n25), 
        .ZN(ref_1_maj_96_port_o) );
  XOR2_X1 ref_1_maj_96_U2 ( .A(ref_1_maj_96_n22), .B(ref_1_maj_96_n21), .Z(
        ref_1_maj_96_n23) );
  NAND2_X1 ref_1_maj_97_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_97_n18) );
  NAND2_X1 ref_1_maj_97_U14 ( .A1(ref_1_maj_97_n21), .A2(ref_1_maj_97_n22), 
        .ZN(ref_1_maj_97_n17) );
  NAND2_X1 ref_1_maj_97_U13 ( .A1(ref_1_maj_97_n18), .A2(ref_1_maj_97_n17), 
        .ZN(ref_1_maj_97_n19) );
  NAND2_X1 ref_1_maj_97_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_97_n16), .ZN(
        ref_1_maj_97_n14) );
  NAND2_X1 ref_1_maj_97_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_97_n15) );
  NAND2_X1 ref_1_maj_97_U10 ( .A1(ref_1_maj_97_n15), .A2(ref_1_maj_97_n14), 
        .ZN(ref_1_maj_97_n20) );
  XOR2_X1 ref_1_maj_97_U9 ( .A(ref_1_n35), .B(ref_1_maj_97_n16), .Z(
        ref_1_maj_97_n21) );
  XOR2_X1 ref_1_maj_97_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(ref_1_maj_97_n22)
         );
  XOR2_X1 ref_1_maj_97_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(ref_1_maj_97_n16)
         );
  OR2_X1 ref_1_maj_97_U6 ( .A1(ref_1_maj_97_n20), .A2(ref_1_maj_97_n19), .ZN(
        ref_1_maj_97_n24) );
  NAND2_X1 ref_1_maj_97_U5 ( .A1(ref_1_maj_97_n24), .A2(ref_1_maj_97_n23), 
        .ZN(ref_1_maj_97_n25) );
  NAND2_X1 ref_1_maj_97_U4 ( .A1(ref_1_maj_97_n20), .A2(ref_1_maj_97_n19), 
        .ZN(ref_1_maj_97_n26) );
  NAND2_X1 ref_1_maj_97_U3 ( .A1(ref_1_maj_97_n26), .A2(ref_1_maj_97_n25), 
        .ZN(ref_1_maj_97_port_o) );
  XOR2_X1 ref_1_maj_97_U2 ( .A(ref_1_maj_97_n22), .B(ref_1_maj_97_n21), .Z(
        ref_1_maj_97_n23) );
  NAND2_X1 ref_1_maj_98_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_98_n18) );
  NAND2_X1 ref_1_maj_98_U14 ( .A1(ref_1_maj_98_n21), .A2(ref_1_maj_98_n22), 
        .ZN(ref_1_maj_98_n17) );
  NAND2_X1 ref_1_maj_98_U13 ( .A1(ref_1_maj_98_n18), .A2(ref_1_maj_98_n17), 
        .ZN(ref_1_maj_98_n19) );
  NAND2_X1 ref_1_maj_98_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_98_n16), .ZN(
        ref_1_maj_98_n14) );
  NAND2_X1 ref_1_maj_98_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_98_n15) );
  NAND2_X1 ref_1_maj_98_U10 ( .A1(ref_1_maj_98_n15), .A2(ref_1_maj_98_n14), 
        .ZN(ref_1_maj_98_n20) );
  XOR2_X1 ref_1_maj_98_U9 ( .A(ref_1_n36), .B(ref_1_maj_98_n16), .Z(
        ref_1_maj_98_n21) );
  XOR2_X1 ref_1_maj_98_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_98_n22)
         );
  XOR2_X1 ref_1_maj_98_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_98_n16)
         );
  OR2_X1 ref_1_maj_98_U6 ( .A1(ref_1_maj_98_n20), .A2(ref_1_maj_98_n19), .ZN(
        ref_1_maj_98_n24) );
  NAND2_X1 ref_1_maj_98_U5 ( .A1(ref_1_maj_98_n24), .A2(ref_1_maj_98_n23), 
        .ZN(ref_1_maj_98_n25) );
  NAND2_X1 ref_1_maj_98_U4 ( .A1(ref_1_maj_98_n20), .A2(ref_1_maj_98_n19), 
        .ZN(ref_1_maj_98_n26) );
  NAND2_X1 ref_1_maj_98_U3 ( .A1(ref_1_maj_98_n26), .A2(ref_1_maj_98_n25), 
        .ZN(ref_1_maj_98_port_o) );
  XOR2_X1 ref_1_maj_98_U2 ( .A(ref_1_maj_98_n22), .B(ref_1_maj_98_n21), .Z(
        ref_1_maj_98_n23) );
  NAND2_X1 ref_1_maj_99_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_99_n18) );
  NAND2_X1 ref_1_maj_99_U14 ( .A1(ref_1_maj_99_n21), .A2(ref_1_maj_99_n22), 
        .ZN(ref_1_maj_99_n17) );
  NAND2_X1 ref_1_maj_99_U13 ( .A1(ref_1_maj_99_n18), .A2(ref_1_maj_99_n17), 
        .ZN(ref_1_maj_99_n19) );
  NAND2_X1 ref_1_maj_99_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_99_n16), .ZN(
        ref_1_maj_99_n14) );
  NAND2_X1 ref_1_maj_99_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_99_n15) );
  NAND2_X1 ref_1_maj_99_U10 ( .A1(ref_1_maj_99_n15), .A2(ref_1_maj_99_n14), 
        .ZN(ref_1_maj_99_n20) );
  XOR2_X1 ref_1_maj_99_U9 ( .A(ref_1_n36), .B(ref_1_maj_99_n16), .Z(
        ref_1_maj_99_n21) );
  XOR2_X1 ref_1_maj_99_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(ref_1_maj_99_n22)
         );
  XOR2_X1 ref_1_maj_99_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(ref_1_maj_99_n16)
         );
  OR2_X1 ref_1_maj_99_U6 ( .A1(ref_1_maj_99_n20), .A2(ref_1_maj_99_n19), .ZN(
        ref_1_maj_99_n24) );
  NAND2_X1 ref_1_maj_99_U5 ( .A1(ref_1_maj_99_n24), .A2(ref_1_maj_99_n23), 
        .ZN(ref_1_maj_99_n25) );
  NAND2_X1 ref_1_maj_99_U4 ( .A1(ref_1_maj_99_n20), .A2(ref_1_maj_99_n19), 
        .ZN(ref_1_maj_99_n26) );
  NAND2_X1 ref_1_maj_99_U3 ( .A1(ref_1_maj_99_n26), .A2(ref_1_maj_99_n25), 
        .ZN(ref_1_maj_99_port_o) );
  XOR2_X1 ref_1_maj_99_U2 ( .A(ref_1_maj_99_n22), .B(ref_1_maj_99_n21), .Z(
        ref_1_maj_99_n23) );
  NAND2_X1 ref_1_maj_100_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_100_n18) );
  NAND2_X1 ref_1_maj_100_U14 ( .A1(ref_1_maj_100_n21), .A2(ref_1_maj_100_n22), 
        .ZN(ref_1_maj_100_n17) );
  NAND2_X1 ref_1_maj_100_U13 ( .A1(ref_1_maj_100_n18), .A2(ref_1_maj_100_n17), 
        .ZN(ref_1_maj_100_n19) );
  NAND2_X1 ref_1_maj_100_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_100_n16), .ZN(
        ref_1_maj_100_n14) );
  NAND2_X1 ref_1_maj_100_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_100_n15) );
  NAND2_X1 ref_1_maj_100_U10 ( .A1(ref_1_maj_100_n15), .A2(ref_1_maj_100_n14), 
        .ZN(ref_1_maj_100_n20) );
  XOR2_X1 ref_1_maj_100_U9 ( .A(ref_1_n25), .B(ref_1_maj_100_n16), .Z(
        ref_1_maj_100_n21) );
  XOR2_X1 ref_1_maj_100_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_100_n22) );
  XOR2_X1 ref_1_maj_100_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_100_n16) );
  OR2_X1 ref_1_maj_100_U6 ( .A1(ref_1_maj_100_n20), .A2(ref_1_maj_100_n19), 
        .ZN(ref_1_maj_100_n24) );
  NAND2_X1 ref_1_maj_100_U5 ( .A1(ref_1_maj_100_n24), .A2(ref_1_maj_100_n23), 
        .ZN(ref_1_maj_100_n25) );
  NAND2_X1 ref_1_maj_100_U4 ( .A1(ref_1_maj_100_n20), .A2(ref_1_maj_100_n19), 
        .ZN(ref_1_maj_100_n26) );
  NAND2_X1 ref_1_maj_100_U3 ( .A1(ref_1_maj_100_n26), .A2(ref_1_maj_100_n25), 
        .ZN(ref_1_maj_100_port_o) );
  XOR2_X1 ref_1_maj_100_U2 ( .A(ref_1_maj_100_n22), .B(ref_1_maj_100_n21), .Z(
        ref_1_maj_100_n23) );
  NAND2_X1 ref_1_maj_101_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_101_n18) );
  NAND2_X1 ref_1_maj_101_U14 ( .A1(ref_1_maj_101_n21), .A2(ref_1_maj_101_n22), 
        .ZN(ref_1_maj_101_n17) );
  NAND2_X1 ref_1_maj_101_U13 ( .A1(ref_1_maj_101_n18), .A2(ref_1_maj_101_n17), 
        .ZN(ref_1_maj_101_n19) );
  NAND2_X1 ref_1_maj_101_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_101_n16), .ZN(
        ref_1_maj_101_n14) );
  NAND2_X1 ref_1_maj_101_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_101_n15) );
  NAND2_X1 ref_1_maj_101_U10 ( .A1(ref_1_maj_101_n15), .A2(ref_1_maj_101_n14), 
        .ZN(ref_1_maj_101_n20) );
  XOR2_X1 ref_1_maj_101_U9 ( .A(ref_1_n26), .B(ref_1_maj_101_n16), .Z(
        ref_1_maj_101_n21) );
  XOR2_X1 ref_1_maj_101_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_101_n22) );
  XOR2_X1 ref_1_maj_101_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_101_n16) );
  OR2_X1 ref_1_maj_101_U6 ( .A1(ref_1_maj_101_n20), .A2(ref_1_maj_101_n19), 
        .ZN(ref_1_maj_101_n24) );
  NAND2_X1 ref_1_maj_101_U5 ( .A1(ref_1_maj_101_n24), .A2(ref_1_maj_101_n23), 
        .ZN(ref_1_maj_101_n25) );
  NAND2_X1 ref_1_maj_101_U4 ( .A1(ref_1_maj_101_n20), .A2(ref_1_maj_101_n19), 
        .ZN(ref_1_maj_101_n26) );
  NAND2_X1 ref_1_maj_101_U3 ( .A1(ref_1_maj_101_n26), .A2(ref_1_maj_101_n25), 
        .ZN(ref_1_maj_101_port_o) );
  XOR2_X1 ref_1_maj_101_U2 ( .A(ref_1_maj_101_n22), .B(ref_1_maj_101_n21), .Z(
        ref_1_maj_101_n23) );
  NAND2_X1 ref_1_maj_102_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_102_n18) );
  NAND2_X1 ref_1_maj_102_U14 ( .A1(ref_1_maj_102_n21), .A2(ref_1_maj_102_n22), 
        .ZN(ref_1_maj_102_n17) );
  NAND2_X1 ref_1_maj_102_U13 ( .A1(ref_1_maj_102_n18), .A2(ref_1_maj_102_n17), 
        .ZN(ref_1_maj_102_n19) );
  NAND2_X1 ref_1_maj_102_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_102_n16), .ZN(
        ref_1_maj_102_n14) );
  NAND2_X1 ref_1_maj_102_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_102_n15) );
  NAND2_X1 ref_1_maj_102_U10 ( .A1(ref_1_maj_102_n15), .A2(ref_1_maj_102_n14), 
        .ZN(ref_1_maj_102_n20) );
  XOR2_X1 ref_1_maj_102_U9 ( .A(ref_1_n26), .B(ref_1_maj_102_n16), .Z(
        ref_1_maj_102_n21) );
  XOR2_X1 ref_1_maj_102_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_102_n22) );
  XOR2_X1 ref_1_maj_102_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_102_n16) );
  OR2_X1 ref_1_maj_102_U6 ( .A1(ref_1_maj_102_n20), .A2(ref_1_maj_102_n19), 
        .ZN(ref_1_maj_102_n24) );
  NAND2_X1 ref_1_maj_102_U5 ( .A1(ref_1_maj_102_n24), .A2(ref_1_maj_102_n23), 
        .ZN(ref_1_maj_102_n25) );
  NAND2_X1 ref_1_maj_102_U4 ( .A1(ref_1_maj_102_n20), .A2(ref_1_maj_102_n19), 
        .ZN(ref_1_maj_102_n26) );
  NAND2_X1 ref_1_maj_102_U3 ( .A1(ref_1_maj_102_n26), .A2(ref_1_maj_102_n25), 
        .ZN(ref_1_maj_102_port_o) );
  XOR2_X1 ref_1_maj_102_U2 ( .A(ref_1_maj_102_n22), .B(ref_1_maj_102_n21), .Z(
        ref_1_maj_102_n23) );
  NAND2_X1 ref_1_maj_103_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_103_n18) );
  NAND2_X1 ref_1_maj_103_U14 ( .A1(ref_1_maj_103_n21), .A2(ref_1_maj_103_n22), 
        .ZN(ref_1_maj_103_n17) );
  NAND2_X1 ref_1_maj_103_U13 ( .A1(ref_1_maj_103_n18), .A2(ref_1_maj_103_n17), 
        .ZN(ref_1_maj_103_n19) );
  NAND2_X1 ref_1_maj_103_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_103_n16), .ZN(
        ref_1_maj_103_n14) );
  NAND2_X1 ref_1_maj_103_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_103_n15) );
  NAND2_X1 ref_1_maj_103_U10 ( .A1(ref_1_maj_103_n15), .A2(ref_1_maj_103_n14), 
        .ZN(ref_1_maj_103_n20) );
  XOR2_X1 ref_1_maj_103_U9 ( .A(ref_1_n25), .B(ref_1_maj_103_n16), .Z(
        ref_1_maj_103_n21) );
  XOR2_X1 ref_1_maj_103_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_103_n22) );
  XOR2_X1 ref_1_maj_103_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_103_n16) );
  OR2_X1 ref_1_maj_103_U6 ( .A1(ref_1_maj_103_n20), .A2(ref_1_maj_103_n19), 
        .ZN(ref_1_maj_103_n24) );
  NAND2_X1 ref_1_maj_103_U5 ( .A1(ref_1_maj_103_n24), .A2(ref_1_maj_103_n23), 
        .ZN(ref_1_maj_103_n25) );
  NAND2_X1 ref_1_maj_103_U4 ( .A1(ref_1_maj_103_n20), .A2(ref_1_maj_103_n19), 
        .ZN(ref_1_maj_103_n26) );
  NAND2_X1 ref_1_maj_103_U3 ( .A1(ref_1_maj_103_n26), .A2(ref_1_maj_103_n25), 
        .ZN(ref_1_maj_103_port_o) );
  XOR2_X1 ref_1_maj_103_U2 ( .A(ref_1_maj_103_n22), .B(ref_1_maj_103_n21), .Z(
        ref_1_maj_103_n23) );
  NAND2_X1 ref_1_maj_104_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_104_n18) );
  NAND2_X1 ref_1_maj_104_U14 ( .A1(ref_1_maj_104_n21), .A2(ref_1_maj_104_n22), 
        .ZN(ref_1_maj_104_n17) );
  NAND2_X1 ref_1_maj_104_U13 ( .A1(ref_1_maj_104_n18), .A2(ref_1_maj_104_n17), 
        .ZN(ref_1_maj_104_n19) );
  NAND2_X1 ref_1_maj_104_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_104_n16), .ZN(
        ref_1_maj_104_n14) );
  NAND2_X1 ref_1_maj_104_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_104_n15) );
  NAND2_X1 ref_1_maj_104_U10 ( .A1(ref_1_maj_104_n15), .A2(ref_1_maj_104_n14), 
        .ZN(ref_1_maj_104_n20) );
  XOR2_X1 ref_1_maj_104_U9 ( .A(ref_1_n15), .B(ref_1_maj_104_n16), .Z(
        ref_1_maj_104_n21) );
  XOR2_X1 ref_1_maj_104_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_104_n22) );
  XOR2_X1 ref_1_maj_104_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_104_n16) );
  OR2_X1 ref_1_maj_104_U6 ( .A1(ref_1_maj_104_n20), .A2(ref_1_maj_104_n19), 
        .ZN(ref_1_maj_104_n24) );
  NAND2_X1 ref_1_maj_104_U5 ( .A1(ref_1_maj_104_n24), .A2(ref_1_maj_104_n23), 
        .ZN(ref_1_maj_104_n25) );
  NAND2_X1 ref_1_maj_104_U4 ( .A1(ref_1_maj_104_n20), .A2(ref_1_maj_104_n19), 
        .ZN(ref_1_maj_104_n26) );
  NAND2_X1 ref_1_maj_104_U3 ( .A1(ref_1_maj_104_n26), .A2(ref_1_maj_104_n25), 
        .ZN(ref_1_maj_104_port_o) );
  XOR2_X1 ref_1_maj_104_U2 ( .A(ref_1_maj_104_n22), .B(ref_1_maj_104_n21), .Z(
        ref_1_maj_104_n23) );
  NAND2_X1 ref_1_maj_105_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_105_n18) );
  NAND2_X1 ref_1_maj_105_U14 ( .A1(ref_1_maj_105_n21), .A2(ref_1_maj_105_n22), 
        .ZN(ref_1_maj_105_n17) );
  NAND2_X1 ref_1_maj_105_U13 ( .A1(ref_1_maj_105_n18), .A2(ref_1_maj_105_n17), 
        .ZN(ref_1_maj_105_n19) );
  NAND2_X1 ref_1_maj_105_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_105_n16), .ZN(
        ref_1_maj_105_n14) );
  NAND2_X1 ref_1_maj_105_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_105_n15) );
  NAND2_X1 ref_1_maj_105_U10 ( .A1(ref_1_maj_105_n15), .A2(ref_1_maj_105_n14), 
        .ZN(ref_1_maj_105_n20) );
  XOR2_X1 ref_1_maj_105_U9 ( .A(ref_1_n16), .B(ref_1_maj_105_n16), .Z(
        ref_1_maj_105_n21) );
  XOR2_X1 ref_1_maj_105_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_105_n22) );
  XOR2_X1 ref_1_maj_105_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_105_n16) );
  OR2_X1 ref_1_maj_105_U6 ( .A1(ref_1_maj_105_n20), .A2(ref_1_maj_105_n19), 
        .ZN(ref_1_maj_105_n24) );
  NAND2_X1 ref_1_maj_105_U5 ( .A1(ref_1_maj_105_n24), .A2(ref_1_maj_105_n23), 
        .ZN(ref_1_maj_105_n25) );
  NAND2_X1 ref_1_maj_105_U4 ( .A1(ref_1_maj_105_n20), .A2(ref_1_maj_105_n19), 
        .ZN(ref_1_maj_105_n26) );
  NAND2_X1 ref_1_maj_105_U3 ( .A1(ref_1_maj_105_n26), .A2(ref_1_maj_105_n25), 
        .ZN(ref_1_maj_105_port_o) );
  XOR2_X1 ref_1_maj_105_U2 ( .A(ref_1_maj_105_n22), .B(ref_1_maj_105_n21), .Z(
        ref_1_maj_105_n23) );
  NAND2_X1 ref_1_maj_106_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_106_n18) );
  NAND2_X1 ref_1_maj_106_U14 ( .A1(ref_1_maj_106_n21), .A2(ref_1_maj_106_n22), 
        .ZN(ref_1_maj_106_n17) );
  NAND2_X1 ref_1_maj_106_U13 ( .A1(ref_1_maj_106_n18), .A2(ref_1_maj_106_n17), 
        .ZN(ref_1_maj_106_n19) );
  NAND2_X1 ref_1_maj_106_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_106_n16), .ZN(
        ref_1_maj_106_n14) );
  NAND2_X1 ref_1_maj_106_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_106_n15) );
  NAND2_X1 ref_1_maj_106_U10 ( .A1(ref_1_maj_106_n15), .A2(ref_1_maj_106_n14), 
        .ZN(ref_1_maj_106_n20) );
  XOR2_X1 ref_1_maj_106_U9 ( .A(ref_1_n16), .B(ref_1_maj_106_n16), .Z(
        ref_1_maj_106_n21) );
  XOR2_X1 ref_1_maj_106_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_106_n22) );
  XOR2_X1 ref_1_maj_106_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_106_n16) );
  OR2_X1 ref_1_maj_106_U6 ( .A1(ref_1_maj_106_n20), .A2(ref_1_maj_106_n19), 
        .ZN(ref_1_maj_106_n24) );
  NAND2_X1 ref_1_maj_106_U5 ( .A1(ref_1_maj_106_n24), .A2(ref_1_maj_106_n23), 
        .ZN(ref_1_maj_106_n25) );
  NAND2_X1 ref_1_maj_106_U4 ( .A1(ref_1_maj_106_n20), .A2(ref_1_maj_106_n19), 
        .ZN(ref_1_maj_106_n26) );
  NAND2_X1 ref_1_maj_106_U3 ( .A1(ref_1_maj_106_n26), .A2(ref_1_maj_106_n25), 
        .ZN(ref_1_maj_106_port_o) );
  XOR2_X1 ref_1_maj_106_U2 ( .A(ref_1_maj_106_n22), .B(ref_1_maj_106_n21), .Z(
        ref_1_maj_106_n23) );
  NAND2_X1 ref_1_maj_107_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_107_n18) );
  NAND2_X1 ref_1_maj_107_U14 ( .A1(ref_1_maj_107_n21), .A2(ref_1_maj_107_n22), 
        .ZN(ref_1_maj_107_n17) );
  NAND2_X1 ref_1_maj_107_U13 ( .A1(ref_1_maj_107_n18), .A2(ref_1_maj_107_n17), 
        .ZN(ref_1_maj_107_n19) );
  NAND2_X1 ref_1_maj_107_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_107_n16), .ZN(
        ref_1_maj_107_n14) );
  NAND2_X1 ref_1_maj_107_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_107_n15) );
  NAND2_X1 ref_1_maj_107_U10 ( .A1(ref_1_maj_107_n15), .A2(ref_1_maj_107_n14), 
        .ZN(ref_1_maj_107_n20) );
  XOR2_X1 ref_1_maj_107_U9 ( .A(ref_1_n15), .B(ref_1_maj_107_n16), .Z(
        ref_1_maj_107_n21) );
  XOR2_X1 ref_1_maj_107_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_107_n22) );
  XOR2_X1 ref_1_maj_107_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_107_n16) );
  OR2_X1 ref_1_maj_107_U6 ( .A1(ref_1_maj_107_n20), .A2(ref_1_maj_107_n19), 
        .ZN(ref_1_maj_107_n24) );
  NAND2_X1 ref_1_maj_107_U5 ( .A1(ref_1_maj_107_n24), .A2(ref_1_maj_107_n23), 
        .ZN(ref_1_maj_107_n25) );
  NAND2_X1 ref_1_maj_107_U4 ( .A1(ref_1_maj_107_n20), .A2(ref_1_maj_107_n19), 
        .ZN(ref_1_maj_107_n26) );
  NAND2_X1 ref_1_maj_107_U3 ( .A1(ref_1_maj_107_n26), .A2(ref_1_maj_107_n25), 
        .ZN(ref_1_maj_107_port_o) );
  XOR2_X1 ref_1_maj_107_U2 ( .A(ref_1_maj_107_n22), .B(ref_1_maj_107_n21), .Z(
        ref_1_maj_107_n23) );
  NAND2_X1 ref_1_maj_108_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_108_n18) );
  NAND2_X1 ref_1_maj_108_U14 ( .A1(ref_1_maj_108_n21), .A2(ref_1_maj_108_n22), 
        .ZN(ref_1_maj_108_n17) );
  NAND2_X1 ref_1_maj_108_U13 ( .A1(ref_1_maj_108_n18), .A2(ref_1_maj_108_n17), 
        .ZN(ref_1_maj_108_n19) );
  NAND2_X1 ref_1_maj_108_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_108_n16), .ZN(
        ref_1_maj_108_n14) );
  NAND2_X1 ref_1_maj_108_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_108_n15) );
  NAND2_X1 ref_1_maj_108_U10 ( .A1(ref_1_maj_108_n15), .A2(ref_1_maj_108_n14), 
        .ZN(ref_1_maj_108_n20) );
  XOR2_X1 ref_1_maj_108_U9 ( .A(ref_1_n5), .B(ref_1_maj_108_n16), .Z(
        ref_1_maj_108_n21) );
  XOR2_X1 ref_1_maj_108_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_108_n22)
         );
  XOR2_X1 ref_1_maj_108_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_108_n16)
         );
  OR2_X1 ref_1_maj_108_U6 ( .A1(ref_1_maj_108_n20), .A2(ref_1_maj_108_n19), 
        .ZN(ref_1_maj_108_n24) );
  NAND2_X1 ref_1_maj_108_U5 ( .A1(ref_1_maj_108_n24), .A2(ref_1_maj_108_n23), 
        .ZN(ref_1_maj_108_n25) );
  NAND2_X1 ref_1_maj_108_U4 ( .A1(ref_1_maj_108_n20), .A2(ref_1_maj_108_n19), 
        .ZN(ref_1_maj_108_n26) );
  NAND2_X1 ref_1_maj_108_U3 ( .A1(ref_1_maj_108_n26), .A2(ref_1_maj_108_n25), 
        .ZN(ref_1_maj_108_port_o) );
  XOR2_X1 ref_1_maj_108_U2 ( .A(ref_1_maj_108_n22), .B(ref_1_maj_108_n21), .Z(
        ref_1_maj_108_n23) );
  NAND2_X1 ref_1_maj_109_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_109_n18) );
  NAND2_X1 ref_1_maj_109_U14 ( .A1(ref_1_maj_109_n21), .A2(ref_1_maj_109_n22), 
        .ZN(ref_1_maj_109_n17) );
  NAND2_X1 ref_1_maj_109_U13 ( .A1(ref_1_maj_109_n18), .A2(ref_1_maj_109_n17), 
        .ZN(ref_1_maj_109_n19) );
  NAND2_X1 ref_1_maj_109_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_109_n16), .ZN(
        ref_1_maj_109_n14) );
  NAND2_X1 ref_1_maj_109_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_109_n15) );
  NAND2_X1 ref_1_maj_109_U10 ( .A1(ref_1_maj_109_n15), .A2(ref_1_maj_109_n14), 
        .ZN(ref_1_maj_109_n20) );
  XOR2_X1 ref_1_maj_109_U9 ( .A(ref_1_n6), .B(ref_1_maj_109_n16), .Z(
        ref_1_maj_109_n21) );
  XOR2_X1 ref_1_maj_109_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_109_n22) );
  XOR2_X1 ref_1_maj_109_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_109_n16)
         );
  OR2_X1 ref_1_maj_109_U6 ( .A1(ref_1_maj_109_n20), .A2(ref_1_maj_109_n19), 
        .ZN(ref_1_maj_109_n24) );
  NAND2_X1 ref_1_maj_109_U5 ( .A1(ref_1_maj_109_n24), .A2(ref_1_maj_109_n23), 
        .ZN(ref_1_maj_109_n25) );
  NAND2_X1 ref_1_maj_109_U4 ( .A1(ref_1_maj_109_n20), .A2(ref_1_maj_109_n19), 
        .ZN(ref_1_maj_109_n26) );
  NAND2_X1 ref_1_maj_109_U3 ( .A1(ref_1_maj_109_n26), .A2(ref_1_maj_109_n25), 
        .ZN(ref_1_maj_109_port_o) );
  XOR2_X1 ref_1_maj_109_U2 ( .A(ref_1_maj_109_n22), .B(ref_1_maj_109_n21), .Z(
        ref_1_maj_109_n23) );
  NAND2_X1 ref_1_maj_110_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_110_n18) );
  NAND2_X1 ref_1_maj_110_U14 ( .A1(ref_1_maj_110_n21), .A2(ref_1_maj_110_n22), 
        .ZN(ref_1_maj_110_n17) );
  NAND2_X1 ref_1_maj_110_U13 ( .A1(ref_1_maj_110_n18), .A2(ref_1_maj_110_n17), 
        .ZN(ref_1_maj_110_n19) );
  NAND2_X1 ref_1_maj_110_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_110_n16), .ZN(
        ref_1_maj_110_n14) );
  NAND2_X1 ref_1_maj_110_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_110_n15) );
  NAND2_X1 ref_1_maj_110_U10 ( .A1(ref_1_maj_110_n15), .A2(ref_1_maj_110_n14), 
        .ZN(ref_1_maj_110_n20) );
  XOR2_X1 ref_1_maj_110_U9 ( .A(ref_1_n6), .B(ref_1_maj_110_n16), .Z(
        ref_1_maj_110_n21) );
  XOR2_X1 ref_1_maj_110_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_110_n22) );
  XOR2_X1 ref_1_maj_110_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_110_n16)
         );
  OR2_X1 ref_1_maj_110_U6 ( .A1(ref_1_maj_110_n20), .A2(ref_1_maj_110_n19), 
        .ZN(ref_1_maj_110_n24) );
  NAND2_X1 ref_1_maj_110_U5 ( .A1(ref_1_maj_110_n24), .A2(ref_1_maj_110_n23), 
        .ZN(ref_1_maj_110_n25) );
  NAND2_X1 ref_1_maj_110_U4 ( .A1(ref_1_maj_110_n20), .A2(ref_1_maj_110_n19), 
        .ZN(ref_1_maj_110_n26) );
  NAND2_X1 ref_1_maj_110_U3 ( .A1(ref_1_maj_110_n26), .A2(ref_1_maj_110_n25), 
        .ZN(ref_1_maj_110_port_o) );
  XOR2_X1 ref_1_maj_110_U2 ( .A(ref_1_maj_110_n22), .B(ref_1_maj_110_n21), .Z(
        ref_1_maj_110_n23) );
  NAND2_X1 ref_1_maj_111_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_111_n18) );
  NAND2_X1 ref_1_maj_111_U14 ( .A1(ref_1_maj_111_n21), .A2(ref_1_maj_111_n22), 
        .ZN(ref_1_maj_111_n17) );
  NAND2_X1 ref_1_maj_111_U13 ( .A1(ref_1_maj_111_n18), .A2(ref_1_maj_111_n17), 
        .ZN(ref_1_maj_111_n19) );
  NAND2_X1 ref_1_maj_111_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_111_n16), .ZN(
        ref_1_maj_111_n14) );
  NAND2_X1 ref_1_maj_111_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_111_n15) );
  NAND2_X1 ref_1_maj_111_U10 ( .A1(ref_1_maj_111_n15), .A2(ref_1_maj_111_n14), 
        .ZN(ref_1_maj_111_n20) );
  XOR2_X1 ref_1_maj_111_U9 ( .A(ref_1_n5), .B(ref_1_maj_111_n16), .Z(
        ref_1_maj_111_n21) );
  XOR2_X1 ref_1_maj_111_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_111_n22)
         );
  XOR2_X1 ref_1_maj_111_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_111_n16)
         );
  OR2_X1 ref_1_maj_111_U6 ( .A1(ref_1_maj_111_n20), .A2(ref_1_maj_111_n19), 
        .ZN(ref_1_maj_111_n24) );
  NAND2_X1 ref_1_maj_111_U5 ( .A1(ref_1_maj_111_n24), .A2(ref_1_maj_111_n23), 
        .ZN(ref_1_maj_111_n25) );
  NAND2_X1 ref_1_maj_111_U4 ( .A1(ref_1_maj_111_n20), .A2(ref_1_maj_111_n19), 
        .ZN(ref_1_maj_111_n26) );
  NAND2_X1 ref_1_maj_111_U3 ( .A1(ref_1_maj_111_n26), .A2(ref_1_maj_111_n25), 
        .ZN(ref_1_maj_111_port_o) );
  XOR2_X1 ref_1_maj_111_U2 ( .A(ref_1_maj_111_n22), .B(ref_1_maj_111_n21), .Z(
        ref_1_maj_111_n23) );
  NAND2_X1 ref_1_maj_112_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_112_n18) );
  NAND2_X1 ref_1_maj_112_U14 ( .A1(ref_1_maj_112_n21), .A2(ref_1_maj_112_n22), 
        .ZN(ref_1_maj_112_n17) );
  NAND2_X1 ref_1_maj_112_U13 ( .A1(ref_1_maj_112_n18), .A2(ref_1_maj_112_n17), 
        .ZN(ref_1_maj_112_n19) );
  NAND2_X1 ref_1_maj_112_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_112_n16), .ZN(
        ref_1_maj_112_n14) );
  NAND2_X1 ref_1_maj_112_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_112_n15) );
  NAND2_X1 ref_1_maj_112_U10 ( .A1(ref_1_maj_112_n15), .A2(ref_1_maj_112_n14), 
        .ZN(ref_1_maj_112_n20) );
  XOR2_X1 ref_1_maj_112_U9 ( .A(ref_1_n35), .B(ref_1_maj_112_n16), .Z(
        ref_1_maj_112_n21) );
  XOR2_X1 ref_1_maj_112_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_112_n22) );
  XOR2_X1 ref_1_maj_112_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_112_n16) );
  OR2_X1 ref_1_maj_112_U6 ( .A1(ref_1_maj_112_n20), .A2(ref_1_maj_112_n19), 
        .ZN(ref_1_maj_112_n24) );
  NAND2_X1 ref_1_maj_112_U5 ( .A1(ref_1_maj_112_n24), .A2(ref_1_maj_112_n23), 
        .ZN(ref_1_maj_112_n25) );
  NAND2_X1 ref_1_maj_112_U4 ( .A1(ref_1_maj_112_n20), .A2(ref_1_maj_112_n19), 
        .ZN(ref_1_maj_112_n26) );
  NAND2_X1 ref_1_maj_112_U3 ( .A1(ref_1_maj_112_n26), .A2(ref_1_maj_112_n25), 
        .ZN(ref_1_maj_112_port_o) );
  XOR2_X1 ref_1_maj_112_U2 ( .A(ref_1_maj_112_n22), .B(ref_1_maj_112_n21), .Z(
        ref_1_maj_112_n23) );
  NAND2_X1 ref_1_maj_113_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_113_n18) );
  NAND2_X1 ref_1_maj_113_U14 ( .A1(ref_1_maj_113_n21), .A2(ref_1_maj_113_n22), 
        .ZN(ref_1_maj_113_n17) );
  NAND2_X1 ref_1_maj_113_U13 ( .A1(ref_1_maj_113_n18), .A2(ref_1_maj_113_n17), 
        .ZN(ref_1_maj_113_n19) );
  NAND2_X1 ref_1_maj_113_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_113_n16), .ZN(
        ref_1_maj_113_n14) );
  NAND2_X1 ref_1_maj_113_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_113_n15) );
  NAND2_X1 ref_1_maj_113_U10 ( .A1(ref_1_maj_113_n15), .A2(ref_1_maj_113_n14), 
        .ZN(ref_1_maj_113_n20) );
  XOR2_X1 ref_1_maj_113_U9 ( .A(ref_1_n36), .B(ref_1_maj_113_n16), .Z(
        ref_1_maj_113_n21) );
  XOR2_X1 ref_1_maj_113_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_113_n22) );
  XOR2_X1 ref_1_maj_113_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_113_n16) );
  OR2_X1 ref_1_maj_113_U6 ( .A1(ref_1_maj_113_n20), .A2(ref_1_maj_113_n19), 
        .ZN(ref_1_maj_113_n24) );
  NAND2_X1 ref_1_maj_113_U5 ( .A1(ref_1_maj_113_n24), .A2(ref_1_maj_113_n23), 
        .ZN(ref_1_maj_113_n25) );
  NAND2_X1 ref_1_maj_113_U4 ( .A1(ref_1_maj_113_n20), .A2(ref_1_maj_113_n19), 
        .ZN(ref_1_maj_113_n26) );
  NAND2_X1 ref_1_maj_113_U3 ( .A1(ref_1_maj_113_n26), .A2(ref_1_maj_113_n25), 
        .ZN(ref_1_maj_113_port_o) );
  XOR2_X1 ref_1_maj_113_U2 ( .A(ref_1_maj_113_n22), .B(ref_1_maj_113_n21), .Z(
        ref_1_maj_113_n23) );
  NAND2_X1 ref_1_maj_114_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_114_n18) );
  NAND2_X1 ref_1_maj_114_U14 ( .A1(ref_1_maj_114_n21), .A2(ref_1_maj_114_n22), 
        .ZN(ref_1_maj_114_n17) );
  NAND2_X1 ref_1_maj_114_U13 ( .A1(ref_1_maj_114_n18), .A2(ref_1_maj_114_n17), 
        .ZN(ref_1_maj_114_n19) );
  NAND2_X1 ref_1_maj_114_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_114_n16), .ZN(
        ref_1_maj_114_n14) );
  NAND2_X1 ref_1_maj_114_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_114_n15) );
  NAND2_X1 ref_1_maj_114_U10 ( .A1(ref_1_maj_114_n15), .A2(ref_1_maj_114_n14), 
        .ZN(ref_1_maj_114_n20) );
  XOR2_X1 ref_1_maj_114_U9 ( .A(ref_1_n35), .B(ref_1_maj_114_n16), .Z(
        ref_1_maj_114_n21) );
  XOR2_X1 ref_1_maj_114_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_114_n22) );
  XOR2_X1 ref_1_maj_114_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_114_n16) );
  OR2_X1 ref_1_maj_114_U6 ( .A1(ref_1_maj_114_n20), .A2(ref_1_maj_114_n19), 
        .ZN(ref_1_maj_114_n24) );
  NAND2_X1 ref_1_maj_114_U5 ( .A1(ref_1_maj_114_n24), .A2(ref_1_maj_114_n23), 
        .ZN(ref_1_maj_114_n25) );
  NAND2_X1 ref_1_maj_114_U4 ( .A1(ref_1_maj_114_n20), .A2(ref_1_maj_114_n19), 
        .ZN(ref_1_maj_114_n26) );
  NAND2_X1 ref_1_maj_114_U3 ( .A1(ref_1_maj_114_n26), .A2(ref_1_maj_114_n25), 
        .ZN(ref_1_maj_114_port_o) );
  XOR2_X1 ref_1_maj_114_U2 ( .A(ref_1_maj_114_n22), .B(ref_1_maj_114_n21), .Z(
        ref_1_maj_114_n23) );
  NAND2_X1 ref_1_maj_115_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_115_n18) );
  NAND2_X1 ref_1_maj_115_U14 ( .A1(ref_1_maj_115_n21), .A2(ref_1_maj_115_n22), 
        .ZN(ref_1_maj_115_n17) );
  NAND2_X1 ref_1_maj_115_U13 ( .A1(ref_1_maj_115_n18), .A2(ref_1_maj_115_n17), 
        .ZN(ref_1_maj_115_n19) );
  NAND2_X1 ref_1_maj_115_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_115_n16), .ZN(
        ref_1_maj_115_n14) );
  NAND2_X1 ref_1_maj_115_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_115_n15) );
  NAND2_X1 ref_1_maj_115_U10 ( .A1(ref_1_maj_115_n15), .A2(ref_1_maj_115_n14), 
        .ZN(ref_1_maj_115_n20) );
  XOR2_X1 ref_1_maj_115_U9 ( .A(ref_1_n36), .B(ref_1_maj_115_n16), .Z(
        ref_1_maj_115_n21) );
  XOR2_X1 ref_1_maj_115_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_115_n22) );
  XOR2_X1 ref_1_maj_115_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_115_n16) );
  OR2_X1 ref_1_maj_115_U6 ( .A1(ref_1_maj_115_n20), .A2(ref_1_maj_115_n19), 
        .ZN(ref_1_maj_115_n24) );
  NAND2_X1 ref_1_maj_115_U5 ( .A1(ref_1_maj_115_n24), .A2(ref_1_maj_115_n23), 
        .ZN(ref_1_maj_115_n25) );
  NAND2_X1 ref_1_maj_115_U4 ( .A1(ref_1_maj_115_n20), .A2(ref_1_maj_115_n19), 
        .ZN(ref_1_maj_115_n26) );
  NAND2_X1 ref_1_maj_115_U3 ( .A1(ref_1_maj_115_n26), .A2(ref_1_maj_115_n25), 
        .ZN(ref_1_maj_115_port_o) );
  XOR2_X1 ref_1_maj_115_U2 ( .A(ref_1_maj_115_n22), .B(ref_1_maj_115_n21), .Z(
        ref_1_maj_115_n23) );
  NAND2_X1 ref_1_maj_116_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_116_n18) );
  NAND2_X1 ref_1_maj_116_U14 ( .A1(ref_1_maj_116_n21), .A2(ref_1_maj_116_n22), 
        .ZN(ref_1_maj_116_n17) );
  NAND2_X1 ref_1_maj_116_U13 ( .A1(ref_1_maj_116_n18), .A2(ref_1_maj_116_n17), 
        .ZN(ref_1_maj_116_n19) );
  NAND2_X1 ref_1_maj_116_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_116_n16), .ZN(
        ref_1_maj_116_n14) );
  NAND2_X1 ref_1_maj_116_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_116_n15) );
  NAND2_X1 ref_1_maj_116_U10 ( .A1(ref_1_maj_116_n15), .A2(ref_1_maj_116_n14), 
        .ZN(ref_1_maj_116_n20) );
  XOR2_X1 ref_1_maj_116_U9 ( .A(ref_1_n26), .B(ref_1_maj_116_n16), .Z(
        ref_1_maj_116_n21) );
  XOR2_X1 ref_1_maj_116_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_116_n22) );
  XOR2_X1 ref_1_maj_116_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_116_n16) );
  OR2_X1 ref_1_maj_116_U6 ( .A1(ref_1_maj_116_n20), .A2(ref_1_maj_116_n19), 
        .ZN(ref_1_maj_116_n24) );
  NAND2_X1 ref_1_maj_116_U5 ( .A1(ref_1_maj_116_n24), .A2(ref_1_maj_116_n23), 
        .ZN(ref_1_maj_116_n25) );
  NAND2_X1 ref_1_maj_116_U4 ( .A1(ref_1_maj_116_n20), .A2(ref_1_maj_116_n19), 
        .ZN(ref_1_maj_116_n26) );
  NAND2_X1 ref_1_maj_116_U3 ( .A1(ref_1_maj_116_n26), .A2(ref_1_maj_116_n25), 
        .ZN(ref_1_maj_116_port_o) );
  XOR2_X1 ref_1_maj_116_U2 ( .A(ref_1_maj_116_n22), .B(ref_1_maj_116_n21), .Z(
        ref_1_maj_116_n23) );
  NAND2_X1 ref_1_maj_117_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_117_n18) );
  NAND2_X1 ref_1_maj_117_U14 ( .A1(ref_1_maj_117_n21), .A2(ref_1_maj_117_n22), 
        .ZN(ref_1_maj_117_n17) );
  NAND2_X1 ref_1_maj_117_U13 ( .A1(ref_1_maj_117_n18), .A2(ref_1_maj_117_n17), 
        .ZN(ref_1_maj_117_n19) );
  NAND2_X1 ref_1_maj_117_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_117_n16), .ZN(
        ref_1_maj_117_n14) );
  NAND2_X1 ref_1_maj_117_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_117_n15) );
  NAND2_X1 ref_1_maj_117_U10 ( .A1(ref_1_maj_117_n15), .A2(ref_1_maj_117_n14), 
        .ZN(ref_1_maj_117_n20) );
  XOR2_X1 ref_1_maj_117_U9 ( .A(ref_1_n25), .B(ref_1_maj_117_n16), .Z(
        ref_1_maj_117_n21) );
  XOR2_X1 ref_1_maj_117_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_117_n22) );
  XOR2_X1 ref_1_maj_117_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_117_n16) );
  OR2_X1 ref_1_maj_117_U6 ( .A1(ref_1_maj_117_n20), .A2(ref_1_maj_117_n19), 
        .ZN(ref_1_maj_117_n24) );
  NAND2_X1 ref_1_maj_117_U5 ( .A1(ref_1_maj_117_n24), .A2(ref_1_maj_117_n23), 
        .ZN(ref_1_maj_117_n25) );
  NAND2_X1 ref_1_maj_117_U4 ( .A1(ref_1_maj_117_n20), .A2(ref_1_maj_117_n19), 
        .ZN(ref_1_maj_117_n26) );
  NAND2_X1 ref_1_maj_117_U3 ( .A1(ref_1_maj_117_n26), .A2(ref_1_maj_117_n25), 
        .ZN(ref_1_maj_117_port_o) );
  XOR2_X1 ref_1_maj_117_U2 ( .A(ref_1_maj_117_n22), .B(ref_1_maj_117_n21), .Z(
        ref_1_maj_117_n23) );
  NAND2_X1 ref_1_maj_118_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_118_n18) );
  NAND2_X1 ref_1_maj_118_U14 ( .A1(ref_1_maj_118_n21), .A2(ref_1_maj_118_n22), 
        .ZN(ref_1_maj_118_n17) );
  NAND2_X1 ref_1_maj_118_U13 ( .A1(ref_1_maj_118_n18), .A2(ref_1_maj_118_n17), 
        .ZN(ref_1_maj_118_n19) );
  NAND2_X1 ref_1_maj_118_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_118_n16), .ZN(
        ref_1_maj_118_n14) );
  NAND2_X1 ref_1_maj_118_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_118_n15) );
  NAND2_X1 ref_1_maj_118_U10 ( .A1(ref_1_maj_118_n15), .A2(ref_1_maj_118_n14), 
        .ZN(ref_1_maj_118_n20) );
  XOR2_X1 ref_1_maj_118_U9 ( .A(ref_1_n26), .B(ref_1_maj_118_n16), .Z(
        ref_1_maj_118_n21) );
  XOR2_X1 ref_1_maj_118_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_118_n22) );
  XOR2_X1 ref_1_maj_118_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_118_n16) );
  OR2_X1 ref_1_maj_118_U6 ( .A1(ref_1_maj_118_n20), .A2(ref_1_maj_118_n19), 
        .ZN(ref_1_maj_118_n24) );
  NAND2_X1 ref_1_maj_118_U5 ( .A1(ref_1_maj_118_n24), .A2(ref_1_maj_118_n23), 
        .ZN(ref_1_maj_118_n25) );
  NAND2_X1 ref_1_maj_118_U4 ( .A1(ref_1_maj_118_n20), .A2(ref_1_maj_118_n19), 
        .ZN(ref_1_maj_118_n26) );
  NAND2_X1 ref_1_maj_118_U3 ( .A1(ref_1_maj_118_n26), .A2(ref_1_maj_118_n25), 
        .ZN(ref_1_maj_118_port_o) );
  XOR2_X1 ref_1_maj_118_U2 ( .A(ref_1_maj_118_n22), .B(ref_1_maj_118_n21), .Z(
        ref_1_maj_118_n23) );
  NAND2_X1 ref_1_maj_119_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_119_n18) );
  NAND2_X1 ref_1_maj_119_U14 ( .A1(ref_1_maj_119_n21), .A2(ref_1_maj_119_n22), 
        .ZN(ref_1_maj_119_n17) );
  NAND2_X1 ref_1_maj_119_U13 ( .A1(ref_1_maj_119_n18), .A2(ref_1_maj_119_n17), 
        .ZN(ref_1_maj_119_n19) );
  NAND2_X1 ref_1_maj_119_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_119_n16), .ZN(
        ref_1_maj_119_n14) );
  NAND2_X1 ref_1_maj_119_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_119_n15) );
  NAND2_X1 ref_1_maj_119_U10 ( .A1(ref_1_maj_119_n15), .A2(ref_1_maj_119_n14), 
        .ZN(ref_1_maj_119_n20) );
  XOR2_X1 ref_1_maj_119_U9 ( .A(ref_1_n25), .B(ref_1_maj_119_n16), .Z(
        ref_1_maj_119_n21) );
  XOR2_X1 ref_1_maj_119_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_119_n22) );
  XOR2_X1 ref_1_maj_119_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_119_n16) );
  OR2_X1 ref_1_maj_119_U6 ( .A1(ref_1_maj_119_n20), .A2(ref_1_maj_119_n19), 
        .ZN(ref_1_maj_119_n24) );
  NAND2_X1 ref_1_maj_119_U5 ( .A1(ref_1_maj_119_n24), .A2(ref_1_maj_119_n23), 
        .ZN(ref_1_maj_119_n25) );
  NAND2_X1 ref_1_maj_119_U4 ( .A1(ref_1_maj_119_n20), .A2(ref_1_maj_119_n19), 
        .ZN(ref_1_maj_119_n26) );
  NAND2_X1 ref_1_maj_119_U3 ( .A1(ref_1_maj_119_n26), .A2(ref_1_maj_119_n25), 
        .ZN(ref_1_maj_119_port_o) );
  XOR2_X1 ref_1_maj_119_U2 ( .A(ref_1_maj_119_n22), .B(ref_1_maj_119_n21), .Z(
        ref_1_maj_119_n23) );
  NAND2_X1 ref_1_maj_120_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_120_n18) );
  NAND2_X1 ref_1_maj_120_U14 ( .A1(ref_1_maj_120_n21), .A2(ref_1_maj_120_n22), 
        .ZN(ref_1_maj_120_n17) );
  NAND2_X1 ref_1_maj_120_U13 ( .A1(ref_1_maj_120_n18), .A2(ref_1_maj_120_n17), 
        .ZN(ref_1_maj_120_n19) );
  NAND2_X1 ref_1_maj_120_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_120_n16), .ZN(
        ref_1_maj_120_n14) );
  NAND2_X1 ref_1_maj_120_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_120_n15) );
  NAND2_X1 ref_1_maj_120_U10 ( .A1(ref_1_maj_120_n15), .A2(ref_1_maj_120_n14), 
        .ZN(ref_1_maj_120_n20) );
  XOR2_X1 ref_1_maj_120_U9 ( .A(ref_1_n16), .B(ref_1_maj_120_n16), .Z(
        ref_1_maj_120_n21) );
  XOR2_X1 ref_1_maj_120_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_120_n22) );
  XOR2_X1 ref_1_maj_120_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_120_n16) );
  OR2_X1 ref_1_maj_120_U6 ( .A1(ref_1_maj_120_n20), .A2(ref_1_maj_120_n19), 
        .ZN(ref_1_maj_120_n24) );
  NAND2_X1 ref_1_maj_120_U5 ( .A1(ref_1_maj_120_n24), .A2(ref_1_maj_120_n23), 
        .ZN(ref_1_maj_120_n25) );
  NAND2_X1 ref_1_maj_120_U4 ( .A1(ref_1_maj_120_n20), .A2(ref_1_maj_120_n19), 
        .ZN(ref_1_maj_120_n26) );
  NAND2_X1 ref_1_maj_120_U3 ( .A1(ref_1_maj_120_n26), .A2(ref_1_maj_120_n25), 
        .ZN(ref_1_maj_120_port_o) );
  XOR2_X1 ref_1_maj_120_U2 ( .A(ref_1_maj_120_n22), .B(ref_1_maj_120_n21), .Z(
        ref_1_maj_120_n23) );
  NAND2_X1 ref_1_maj_121_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_121_n18) );
  NAND2_X1 ref_1_maj_121_U14 ( .A1(ref_1_maj_121_n21), .A2(ref_1_maj_121_n22), 
        .ZN(ref_1_maj_121_n17) );
  NAND2_X1 ref_1_maj_121_U13 ( .A1(ref_1_maj_121_n18), .A2(ref_1_maj_121_n17), 
        .ZN(ref_1_maj_121_n19) );
  NAND2_X1 ref_1_maj_121_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_121_n16), .ZN(
        ref_1_maj_121_n14) );
  NAND2_X1 ref_1_maj_121_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_121_n15) );
  NAND2_X1 ref_1_maj_121_U10 ( .A1(ref_1_maj_121_n15), .A2(ref_1_maj_121_n14), 
        .ZN(ref_1_maj_121_n20) );
  XOR2_X1 ref_1_maj_121_U9 ( .A(ref_1_n15), .B(ref_1_maj_121_n16), .Z(
        ref_1_maj_121_n21) );
  XOR2_X1 ref_1_maj_121_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_121_n22) );
  XOR2_X1 ref_1_maj_121_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_121_n16) );
  OR2_X1 ref_1_maj_121_U6 ( .A1(ref_1_maj_121_n20), .A2(ref_1_maj_121_n19), 
        .ZN(ref_1_maj_121_n24) );
  NAND2_X1 ref_1_maj_121_U5 ( .A1(ref_1_maj_121_n24), .A2(ref_1_maj_121_n23), 
        .ZN(ref_1_maj_121_n25) );
  NAND2_X1 ref_1_maj_121_U4 ( .A1(ref_1_maj_121_n20), .A2(ref_1_maj_121_n19), 
        .ZN(ref_1_maj_121_n26) );
  NAND2_X1 ref_1_maj_121_U3 ( .A1(ref_1_maj_121_n26), .A2(ref_1_maj_121_n25), 
        .ZN(ref_1_maj_121_port_o) );
  XOR2_X1 ref_1_maj_121_U2 ( .A(ref_1_maj_121_n22), .B(ref_1_maj_121_n21), .Z(
        ref_1_maj_121_n23) );
  NAND2_X1 ref_1_maj_122_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_122_n18) );
  NAND2_X1 ref_1_maj_122_U14 ( .A1(ref_1_maj_122_n21), .A2(ref_1_maj_122_n22), 
        .ZN(ref_1_maj_122_n17) );
  NAND2_X1 ref_1_maj_122_U13 ( .A1(ref_1_maj_122_n18), .A2(ref_1_maj_122_n17), 
        .ZN(ref_1_maj_122_n19) );
  NAND2_X1 ref_1_maj_122_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_122_n16), .ZN(
        ref_1_maj_122_n14) );
  NAND2_X1 ref_1_maj_122_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_122_n15) );
  NAND2_X1 ref_1_maj_122_U10 ( .A1(ref_1_maj_122_n15), .A2(ref_1_maj_122_n14), 
        .ZN(ref_1_maj_122_n20) );
  XOR2_X1 ref_1_maj_122_U9 ( .A(ref_1_n16), .B(ref_1_maj_122_n16), .Z(
        ref_1_maj_122_n21) );
  XOR2_X1 ref_1_maj_122_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_122_n22) );
  XOR2_X1 ref_1_maj_122_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_122_n16) );
  OR2_X1 ref_1_maj_122_U6 ( .A1(ref_1_maj_122_n20), .A2(ref_1_maj_122_n19), 
        .ZN(ref_1_maj_122_n24) );
  NAND2_X1 ref_1_maj_122_U5 ( .A1(ref_1_maj_122_n24), .A2(ref_1_maj_122_n23), 
        .ZN(ref_1_maj_122_n25) );
  NAND2_X1 ref_1_maj_122_U4 ( .A1(ref_1_maj_122_n20), .A2(ref_1_maj_122_n19), 
        .ZN(ref_1_maj_122_n26) );
  NAND2_X1 ref_1_maj_122_U3 ( .A1(ref_1_maj_122_n26), .A2(ref_1_maj_122_n25), 
        .ZN(ref_1_maj_122_port_o) );
  XOR2_X1 ref_1_maj_122_U2 ( .A(ref_1_maj_122_n22), .B(ref_1_maj_122_n21), .Z(
        ref_1_maj_122_n23) );
  NAND2_X1 ref_1_maj_123_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_123_n18) );
  NAND2_X1 ref_1_maj_123_U14 ( .A1(ref_1_maj_123_n21), .A2(ref_1_maj_123_n22), 
        .ZN(ref_1_maj_123_n17) );
  NAND2_X1 ref_1_maj_123_U13 ( .A1(ref_1_maj_123_n18), .A2(ref_1_maj_123_n17), 
        .ZN(ref_1_maj_123_n19) );
  NAND2_X1 ref_1_maj_123_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_123_n16), .ZN(
        ref_1_maj_123_n14) );
  NAND2_X1 ref_1_maj_123_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_123_n15) );
  NAND2_X1 ref_1_maj_123_U10 ( .A1(ref_1_maj_123_n15), .A2(ref_1_maj_123_n14), 
        .ZN(ref_1_maj_123_n20) );
  XOR2_X1 ref_1_maj_123_U9 ( .A(ref_1_n15), .B(ref_1_maj_123_n16), .Z(
        ref_1_maj_123_n21) );
  XOR2_X1 ref_1_maj_123_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_123_n22) );
  XOR2_X1 ref_1_maj_123_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_123_n16) );
  OR2_X1 ref_1_maj_123_U6 ( .A1(ref_1_maj_123_n20), .A2(ref_1_maj_123_n19), 
        .ZN(ref_1_maj_123_n24) );
  NAND2_X1 ref_1_maj_123_U5 ( .A1(ref_1_maj_123_n24), .A2(ref_1_maj_123_n23), 
        .ZN(ref_1_maj_123_n25) );
  NAND2_X1 ref_1_maj_123_U4 ( .A1(ref_1_maj_123_n20), .A2(ref_1_maj_123_n19), 
        .ZN(ref_1_maj_123_n26) );
  NAND2_X1 ref_1_maj_123_U3 ( .A1(ref_1_maj_123_n26), .A2(ref_1_maj_123_n25), 
        .ZN(ref_1_maj_123_port_o) );
  XOR2_X1 ref_1_maj_123_U2 ( .A(ref_1_maj_123_n22), .B(ref_1_maj_123_n21), .Z(
        ref_1_maj_123_n23) );
  NAND2_X1 ref_1_maj_124_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_124_n18) );
  NAND2_X1 ref_1_maj_124_U14 ( .A1(ref_1_maj_124_n21), .A2(ref_1_maj_124_n22), 
        .ZN(ref_1_maj_124_n17) );
  NAND2_X1 ref_1_maj_124_U13 ( .A1(ref_1_maj_124_n18), .A2(ref_1_maj_124_n17), 
        .ZN(ref_1_maj_124_n19) );
  NAND2_X1 ref_1_maj_124_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_124_n16), .ZN(
        ref_1_maj_124_n14) );
  NAND2_X1 ref_1_maj_124_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_124_n15) );
  NAND2_X1 ref_1_maj_124_U10 ( .A1(ref_1_maj_124_n15), .A2(ref_1_maj_124_n14), 
        .ZN(ref_1_maj_124_n20) );
  XOR2_X1 ref_1_maj_124_U9 ( .A(ref_1_n6), .B(ref_1_maj_124_n16), .Z(
        ref_1_maj_124_n21) );
  XOR2_X1 ref_1_maj_124_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_124_n22) );
  XOR2_X1 ref_1_maj_124_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_124_n16)
         );
  OR2_X1 ref_1_maj_124_U6 ( .A1(ref_1_maj_124_n20), .A2(ref_1_maj_124_n19), 
        .ZN(ref_1_maj_124_n24) );
  NAND2_X1 ref_1_maj_124_U5 ( .A1(ref_1_maj_124_n24), .A2(ref_1_maj_124_n23), 
        .ZN(ref_1_maj_124_n25) );
  NAND2_X1 ref_1_maj_124_U4 ( .A1(ref_1_maj_124_n20), .A2(ref_1_maj_124_n19), 
        .ZN(ref_1_maj_124_n26) );
  NAND2_X1 ref_1_maj_124_U3 ( .A1(ref_1_maj_124_n26), .A2(ref_1_maj_124_n25), 
        .ZN(ref_1_maj_124_port_o) );
  XOR2_X1 ref_1_maj_124_U2 ( .A(ref_1_maj_124_n22), .B(ref_1_maj_124_n21), .Z(
        ref_1_maj_124_n23) );
  NAND2_X1 ref_1_maj_125_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_125_n18) );
  NAND2_X1 ref_1_maj_125_U14 ( .A1(ref_1_maj_125_n21), .A2(ref_1_maj_125_n22), 
        .ZN(ref_1_maj_125_n17) );
  NAND2_X1 ref_1_maj_125_U13 ( .A1(ref_1_maj_125_n18), .A2(ref_1_maj_125_n17), 
        .ZN(ref_1_maj_125_n19) );
  NAND2_X1 ref_1_maj_125_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_125_n16), .ZN(
        ref_1_maj_125_n14) );
  NAND2_X1 ref_1_maj_125_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_125_n15) );
  NAND2_X1 ref_1_maj_125_U10 ( .A1(ref_1_maj_125_n15), .A2(ref_1_maj_125_n14), 
        .ZN(ref_1_maj_125_n20) );
  XOR2_X1 ref_1_maj_125_U9 ( .A(ref_1_n5), .B(ref_1_maj_125_n16), .Z(
        ref_1_maj_125_n21) );
  XOR2_X1 ref_1_maj_125_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_125_n22)
         );
  XOR2_X1 ref_1_maj_125_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_125_n16)
         );
  OR2_X1 ref_1_maj_125_U6 ( .A1(ref_1_maj_125_n20), .A2(ref_1_maj_125_n19), 
        .ZN(ref_1_maj_125_n24) );
  NAND2_X1 ref_1_maj_125_U5 ( .A1(ref_1_maj_125_n24), .A2(ref_1_maj_125_n23), 
        .ZN(ref_1_maj_125_n25) );
  NAND2_X1 ref_1_maj_125_U4 ( .A1(ref_1_maj_125_n20), .A2(ref_1_maj_125_n19), 
        .ZN(ref_1_maj_125_n26) );
  NAND2_X1 ref_1_maj_125_U3 ( .A1(ref_1_maj_125_n26), .A2(ref_1_maj_125_n25), 
        .ZN(ref_1_maj_125_port_o) );
  XOR2_X1 ref_1_maj_125_U2 ( .A(ref_1_maj_125_n22), .B(ref_1_maj_125_n21), .Z(
        ref_1_maj_125_n23) );
  NAND2_X1 ref_1_maj_126_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_126_n18) );
  NAND2_X1 ref_1_maj_126_U14 ( .A1(ref_1_maj_126_n21), .A2(ref_1_maj_126_n22), 
        .ZN(ref_1_maj_126_n17) );
  NAND2_X1 ref_1_maj_126_U13 ( .A1(ref_1_maj_126_n18), .A2(ref_1_maj_126_n17), 
        .ZN(ref_1_maj_126_n19) );
  NAND2_X1 ref_1_maj_126_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_126_n16), .ZN(
        ref_1_maj_126_n14) );
  NAND2_X1 ref_1_maj_126_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_126_n15) );
  NAND2_X1 ref_1_maj_126_U10 ( .A1(ref_1_maj_126_n15), .A2(ref_1_maj_126_n14), 
        .ZN(ref_1_maj_126_n20) );
  XOR2_X1 ref_1_maj_126_U9 ( .A(ref_1_n6), .B(ref_1_maj_126_n16), .Z(
        ref_1_maj_126_n21) );
  XOR2_X1 ref_1_maj_126_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_126_n22) );
  XOR2_X1 ref_1_maj_126_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_126_n16)
         );
  OR2_X1 ref_1_maj_126_U6 ( .A1(ref_1_maj_126_n20), .A2(ref_1_maj_126_n19), 
        .ZN(ref_1_maj_126_n24) );
  NAND2_X1 ref_1_maj_126_U5 ( .A1(ref_1_maj_126_n24), .A2(ref_1_maj_126_n23), 
        .ZN(ref_1_maj_126_n25) );
  NAND2_X1 ref_1_maj_126_U4 ( .A1(ref_1_maj_126_n20), .A2(ref_1_maj_126_n19), 
        .ZN(ref_1_maj_126_n26) );
  NAND2_X1 ref_1_maj_126_U3 ( .A1(ref_1_maj_126_n26), .A2(ref_1_maj_126_n25), 
        .ZN(ref_1_maj_126_port_o) );
  XOR2_X1 ref_1_maj_126_U2 ( .A(ref_1_maj_126_n22), .B(ref_1_maj_126_n21), .Z(
        ref_1_maj_126_n23) );
  NAND2_X1 ref_1_maj_127_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_127_n18) );
  NAND2_X1 ref_1_maj_127_U14 ( .A1(ref_1_maj_127_n21), .A2(ref_1_maj_127_n22), 
        .ZN(ref_1_maj_127_n17) );
  NAND2_X1 ref_1_maj_127_U13 ( .A1(ref_1_maj_127_n18), .A2(ref_1_maj_127_n17), 
        .ZN(ref_1_maj_127_n19) );
  NAND2_X1 ref_1_maj_127_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_127_n16), .ZN(
        ref_1_maj_127_n14) );
  NAND2_X1 ref_1_maj_127_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_127_n15) );
  NAND2_X1 ref_1_maj_127_U10 ( .A1(ref_1_maj_127_n15), .A2(ref_1_maj_127_n14), 
        .ZN(ref_1_maj_127_n20) );
  XOR2_X1 ref_1_maj_127_U9 ( .A(ref_1_n5), .B(ref_1_maj_127_n16), .Z(
        ref_1_maj_127_n21) );
  XOR2_X1 ref_1_maj_127_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_127_n22)
         );
  XOR2_X1 ref_1_maj_127_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_127_n16)
         );
  OR2_X1 ref_1_maj_127_U6 ( .A1(ref_1_maj_127_n20), .A2(ref_1_maj_127_n19), 
        .ZN(ref_1_maj_127_n24) );
  NAND2_X1 ref_1_maj_127_U5 ( .A1(ref_1_maj_127_n24), .A2(ref_1_maj_127_n23), 
        .ZN(ref_1_maj_127_n25) );
  NAND2_X1 ref_1_maj_127_U4 ( .A1(ref_1_maj_127_n20), .A2(ref_1_maj_127_n19), 
        .ZN(ref_1_maj_127_n26) );
  NAND2_X1 ref_1_maj_127_U3 ( .A1(ref_1_maj_127_n26), .A2(ref_1_maj_127_n25), 
        .ZN(ref_1_maj_127_port_o) );
  XOR2_X1 ref_1_maj_127_U2 ( .A(ref_1_maj_127_n22), .B(ref_1_maj_127_n21), .Z(
        ref_1_maj_127_n23) );
  NAND2_X1 ref_1_maj_128_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_128_n18) );
  NAND2_X1 ref_1_maj_128_U14 ( .A1(ref_1_maj_128_n21), .A2(ref_1_maj_128_n22), 
        .ZN(ref_1_maj_128_n17) );
  NAND2_X1 ref_1_maj_128_U13 ( .A1(ref_1_maj_128_n18), .A2(ref_1_maj_128_n17), 
        .ZN(ref_1_maj_128_n19) );
  NAND2_X1 ref_1_maj_128_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_128_n16), .ZN(
        ref_1_maj_128_n14) );
  NAND2_X1 ref_1_maj_128_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_128_n15) );
  NAND2_X1 ref_1_maj_128_U10 ( .A1(ref_1_maj_128_n15), .A2(ref_1_maj_128_n14), 
        .ZN(ref_1_maj_128_n20) );
  XOR2_X1 ref_1_maj_128_U9 ( .A(ref_1_n35), .B(ref_1_maj_128_n16), .Z(
        ref_1_maj_128_n21) );
  XOR2_X1 ref_1_maj_128_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_128_n22) );
  XOR2_X1 ref_1_maj_128_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_128_n16) );
  OR2_X1 ref_1_maj_128_U6 ( .A1(ref_1_maj_128_n20), .A2(ref_1_maj_128_n19), 
        .ZN(ref_1_maj_128_n24) );
  NAND2_X1 ref_1_maj_128_U5 ( .A1(ref_1_maj_128_n24), .A2(ref_1_maj_128_n23), 
        .ZN(ref_1_maj_128_n25) );
  NAND2_X1 ref_1_maj_128_U4 ( .A1(ref_1_maj_128_n20), .A2(ref_1_maj_128_n19), 
        .ZN(ref_1_maj_128_n26) );
  NAND2_X1 ref_1_maj_128_U3 ( .A1(ref_1_maj_128_n26), .A2(ref_1_maj_128_n25), 
        .ZN(ref_1_maj_128_port_o) );
  XOR2_X1 ref_1_maj_128_U2 ( .A(ref_1_maj_128_n22), .B(ref_1_maj_128_n21), .Z(
        ref_1_maj_128_n23) );
  NAND2_X1 ref_1_maj_129_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_129_n18) );
  NAND2_X1 ref_1_maj_129_U14 ( .A1(ref_1_maj_129_n21), .A2(ref_1_maj_129_n22), 
        .ZN(ref_1_maj_129_n17) );
  NAND2_X1 ref_1_maj_129_U13 ( .A1(ref_1_maj_129_n18), .A2(ref_1_maj_129_n17), 
        .ZN(ref_1_maj_129_n19) );
  NAND2_X1 ref_1_maj_129_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_129_n16), .ZN(
        ref_1_maj_129_n14) );
  NAND2_X1 ref_1_maj_129_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_129_n15) );
  NAND2_X1 ref_1_maj_129_U10 ( .A1(ref_1_maj_129_n15), .A2(ref_1_maj_129_n14), 
        .ZN(ref_1_maj_129_n20) );
  XOR2_X1 ref_1_maj_129_U9 ( .A(ref_1_n35), .B(ref_1_maj_129_n16), .Z(
        ref_1_maj_129_n21) );
  XOR2_X1 ref_1_maj_129_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_129_n22) );
  XOR2_X1 ref_1_maj_129_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_129_n16) );
  OR2_X1 ref_1_maj_129_U6 ( .A1(ref_1_maj_129_n20), .A2(ref_1_maj_129_n19), 
        .ZN(ref_1_maj_129_n24) );
  NAND2_X1 ref_1_maj_129_U5 ( .A1(ref_1_maj_129_n24), .A2(ref_1_maj_129_n23), 
        .ZN(ref_1_maj_129_n25) );
  NAND2_X1 ref_1_maj_129_U4 ( .A1(ref_1_maj_129_n20), .A2(ref_1_maj_129_n19), 
        .ZN(ref_1_maj_129_n26) );
  NAND2_X1 ref_1_maj_129_U3 ( .A1(ref_1_maj_129_n26), .A2(ref_1_maj_129_n25), 
        .ZN(ref_1_maj_129_port_o) );
  XOR2_X1 ref_1_maj_129_U2 ( .A(ref_1_maj_129_n22), .B(ref_1_maj_129_n21), .Z(
        ref_1_maj_129_n23) );
  NAND2_X1 ref_1_maj_130_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_130_n18) );
  NAND2_X1 ref_1_maj_130_U14 ( .A1(ref_1_maj_130_n21), .A2(ref_1_maj_130_n22), 
        .ZN(ref_1_maj_130_n17) );
  NAND2_X1 ref_1_maj_130_U13 ( .A1(ref_1_maj_130_n18), .A2(ref_1_maj_130_n17), 
        .ZN(ref_1_maj_130_n19) );
  NAND2_X1 ref_1_maj_130_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_130_n16), .ZN(
        ref_1_maj_130_n14) );
  NAND2_X1 ref_1_maj_130_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_130_n15) );
  NAND2_X1 ref_1_maj_130_U10 ( .A1(ref_1_maj_130_n15), .A2(ref_1_maj_130_n14), 
        .ZN(ref_1_maj_130_n20) );
  XOR2_X1 ref_1_maj_130_U9 ( .A(ref_1_n35), .B(ref_1_maj_130_n16), .Z(
        ref_1_maj_130_n21) );
  XOR2_X1 ref_1_maj_130_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_130_n22) );
  XOR2_X1 ref_1_maj_130_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_130_n16) );
  OR2_X1 ref_1_maj_130_U6 ( .A1(ref_1_maj_130_n20), .A2(ref_1_maj_130_n19), 
        .ZN(ref_1_maj_130_n24) );
  NAND2_X1 ref_1_maj_130_U5 ( .A1(ref_1_maj_130_n24), .A2(ref_1_maj_130_n23), 
        .ZN(ref_1_maj_130_n25) );
  NAND2_X1 ref_1_maj_130_U4 ( .A1(ref_1_maj_130_n20), .A2(ref_1_maj_130_n19), 
        .ZN(ref_1_maj_130_n26) );
  NAND2_X1 ref_1_maj_130_U3 ( .A1(ref_1_maj_130_n26), .A2(ref_1_maj_130_n25), 
        .ZN(ref_1_maj_130_port_o) );
  XOR2_X1 ref_1_maj_130_U2 ( .A(ref_1_maj_130_n22), .B(ref_1_maj_130_n21), .Z(
        ref_1_maj_130_n23) );
  NAND2_X1 ref_1_maj_131_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_131_n18) );
  NAND2_X1 ref_1_maj_131_U14 ( .A1(ref_1_maj_131_n21), .A2(ref_1_maj_131_n22), 
        .ZN(ref_1_maj_131_n17) );
  NAND2_X1 ref_1_maj_131_U13 ( .A1(ref_1_maj_131_n18), .A2(ref_1_maj_131_n17), 
        .ZN(ref_1_maj_131_n19) );
  NAND2_X1 ref_1_maj_131_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_131_n16), .ZN(
        ref_1_maj_131_n14) );
  NAND2_X1 ref_1_maj_131_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_131_n15) );
  NAND2_X1 ref_1_maj_131_U10 ( .A1(ref_1_maj_131_n15), .A2(ref_1_maj_131_n14), 
        .ZN(ref_1_maj_131_n20) );
  XOR2_X1 ref_1_maj_131_U9 ( .A(ref_1_n35), .B(ref_1_maj_131_n16), .Z(
        ref_1_maj_131_n21) );
  XOR2_X1 ref_1_maj_131_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_131_n22) );
  XOR2_X1 ref_1_maj_131_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_131_n16) );
  OR2_X1 ref_1_maj_131_U6 ( .A1(ref_1_maj_131_n20), .A2(ref_1_maj_131_n19), 
        .ZN(ref_1_maj_131_n24) );
  NAND2_X1 ref_1_maj_131_U5 ( .A1(ref_1_maj_131_n24), .A2(ref_1_maj_131_n23), 
        .ZN(ref_1_maj_131_n25) );
  NAND2_X1 ref_1_maj_131_U4 ( .A1(ref_1_maj_131_n20), .A2(ref_1_maj_131_n19), 
        .ZN(ref_1_maj_131_n26) );
  NAND2_X1 ref_1_maj_131_U3 ( .A1(ref_1_maj_131_n26), .A2(ref_1_maj_131_n25), 
        .ZN(ref_1_maj_131_port_o) );
  XOR2_X1 ref_1_maj_131_U2 ( .A(ref_1_maj_131_n22), .B(ref_1_maj_131_n21), .Z(
        ref_1_maj_131_n23) );
  NAND2_X1 ref_1_maj_132_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_132_n18) );
  NAND2_X1 ref_1_maj_132_U14 ( .A1(ref_1_maj_132_n21), .A2(ref_1_maj_132_n22), 
        .ZN(ref_1_maj_132_n17) );
  NAND2_X1 ref_1_maj_132_U13 ( .A1(ref_1_maj_132_n18), .A2(ref_1_maj_132_n17), 
        .ZN(ref_1_maj_132_n19) );
  NAND2_X1 ref_1_maj_132_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_132_n16), .ZN(
        ref_1_maj_132_n14) );
  NAND2_X1 ref_1_maj_132_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_132_n15) );
  NAND2_X1 ref_1_maj_132_U10 ( .A1(ref_1_maj_132_n15), .A2(ref_1_maj_132_n14), 
        .ZN(ref_1_maj_132_n20) );
  XOR2_X1 ref_1_maj_132_U9 ( .A(ref_1_n25), .B(ref_1_maj_132_n16), .Z(
        ref_1_maj_132_n21) );
  XOR2_X1 ref_1_maj_132_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_132_n22) );
  XOR2_X1 ref_1_maj_132_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_132_n16) );
  OR2_X1 ref_1_maj_132_U6 ( .A1(ref_1_maj_132_n20), .A2(ref_1_maj_132_n19), 
        .ZN(ref_1_maj_132_n24) );
  NAND2_X1 ref_1_maj_132_U5 ( .A1(ref_1_maj_132_n24), .A2(ref_1_maj_132_n23), 
        .ZN(ref_1_maj_132_n25) );
  NAND2_X1 ref_1_maj_132_U4 ( .A1(ref_1_maj_132_n20), .A2(ref_1_maj_132_n19), 
        .ZN(ref_1_maj_132_n26) );
  NAND2_X1 ref_1_maj_132_U3 ( .A1(ref_1_maj_132_n26), .A2(ref_1_maj_132_n25), 
        .ZN(ref_1_maj_132_port_o) );
  XOR2_X1 ref_1_maj_132_U2 ( .A(ref_1_maj_132_n22), .B(ref_1_maj_132_n21), .Z(
        ref_1_maj_132_n23) );
  NAND2_X1 ref_1_maj_133_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_133_n18) );
  NAND2_X1 ref_1_maj_133_U14 ( .A1(ref_1_maj_133_n21), .A2(ref_1_maj_133_n22), 
        .ZN(ref_1_maj_133_n17) );
  NAND2_X1 ref_1_maj_133_U13 ( .A1(ref_1_maj_133_n18), .A2(ref_1_maj_133_n17), 
        .ZN(ref_1_maj_133_n19) );
  NAND2_X1 ref_1_maj_133_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_133_n16), .ZN(
        ref_1_maj_133_n14) );
  NAND2_X1 ref_1_maj_133_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_133_n15) );
  NAND2_X1 ref_1_maj_133_U10 ( .A1(ref_1_maj_133_n15), .A2(ref_1_maj_133_n14), 
        .ZN(ref_1_maj_133_n20) );
  XOR2_X1 ref_1_maj_133_U9 ( .A(ref_1_n25), .B(ref_1_maj_133_n16), .Z(
        ref_1_maj_133_n21) );
  XOR2_X1 ref_1_maj_133_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_133_n22) );
  XOR2_X1 ref_1_maj_133_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_133_n16) );
  OR2_X1 ref_1_maj_133_U6 ( .A1(ref_1_maj_133_n20), .A2(ref_1_maj_133_n19), 
        .ZN(ref_1_maj_133_n24) );
  NAND2_X1 ref_1_maj_133_U5 ( .A1(ref_1_maj_133_n24), .A2(ref_1_maj_133_n23), 
        .ZN(ref_1_maj_133_n25) );
  NAND2_X1 ref_1_maj_133_U4 ( .A1(ref_1_maj_133_n20), .A2(ref_1_maj_133_n19), 
        .ZN(ref_1_maj_133_n26) );
  NAND2_X1 ref_1_maj_133_U3 ( .A1(ref_1_maj_133_n26), .A2(ref_1_maj_133_n25), 
        .ZN(ref_1_maj_133_port_o) );
  XOR2_X1 ref_1_maj_133_U2 ( .A(ref_1_maj_133_n22), .B(ref_1_maj_133_n21), .Z(
        ref_1_maj_133_n23) );
  NAND2_X1 ref_1_maj_134_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_134_n18) );
  NAND2_X1 ref_1_maj_134_U14 ( .A1(ref_1_maj_134_n21), .A2(ref_1_maj_134_n22), 
        .ZN(ref_1_maj_134_n17) );
  NAND2_X1 ref_1_maj_134_U13 ( .A1(ref_1_maj_134_n18), .A2(ref_1_maj_134_n17), 
        .ZN(ref_1_maj_134_n19) );
  NAND2_X1 ref_1_maj_134_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_134_n16), .ZN(
        ref_1_maj_134_n14) );
  NAND2_X1 ref_1_maj_134_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_134_n15) );
  NAND2_X1 ref_1_maj_134_U10 ( .A1(ref_1_maj_134_n15), .A2(ref_1_maj_134_n14), 
        .ZN(ref_1_maj_134_n20) );
  XOR2_X1 ref_1_maj_134_U9 ( .A(ref_1_n25), .B(ref_1_maj_134_n16), .Z(
        ref_1_maj_134_n21) );
  XOR2_X1 ref_1_maj_134_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_134_n22) );
  XOR2_X1 ref_1_maj_134_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_134_n16) );
  OR2_X1 ref_1_maj_134_U6 ( .A1(ref_1_maj_134_n20), .A2(ref_1_maj_134_n19), 
        .ZN(ref_1_maj_134_n24) );
  NAND2_X1 ref_1_maj_134_U5 ( .A1(ref_1_maj_134_n24), .A2(ref_1_maj_134_n23), 
        .ZN(ref_1_maj_134_n25) );
  NAND2_X1 ref_1_maj_134_U4 ( .A1(ref_1_maj_134_n20), .A2(ref_1_maj_134_n19), 
        .ZN(ref_1_maj_134_n26) );
  NAND2_X1 ref_1_maj_134_U3 ( .A1(ref_1_maj_134_n26), .A2(ref_1_maj_134_n25), 
        .ZN(ref_1_maj_134_port_o) );
  XOR2_X1 ref_1_maj_134_U2 ( .A(ref_1_maj_134_n22), .B(ref_1_maj_134_n21), .Z(
        ref_1_maj_134_n23) );
  NAND2_X1 ref_1_maj_135_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_135_n18) );
  NAND2_X1 ref_1_maj_135_U14 ( .A1(ref_1_maj_135_n21), .A2(ref_1_maj_135_n22), 
        .ZN(ref_1_maj_135_n17) );
  NAND2_X1 ref_1_maj_135_U13 ( .A1(ref_1_maj_135_n18), .A2(ref_1_maj_135_n17), 
        .ZN(ref_1_maj_135_n19) );
  NAND2_X1 ref_1_maj_135_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_135_n16), .ZN(
        ref_1_maj_135_n14) );
  NAND2_X1 ref_1_maj_135_U11 ( .A1(ref_1_n21), .A2(ref_1_n23), .ZN(
        ref_1_maj_135_n15) );
  NAND2_X1 ref_1_maj_135_U10 ( .A1(ref_1_maj_135_n15), .A2(ref_1_maj_135_n14), 
        .ZN(ref_1_maj_135_n20) );
  XOR2_X1 ref_1_maj_135_U9 ( .A(ref_1_n25), .B(ref_1_maj_135_n16), .Z(
        ref_1_maj_135_n21) );
  XOR2_X1 ref_1_maj_135_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(
        ref_1_maj_135_n22) );
  XOR2_X1 ref_1_maj_135_U7 ( .A(ref_1_n21), .B(ref_1_n23), .Z(
        ref_1_maj_135_n16) );
  OR2_X1 ref_1_maj_135_U6 ( .A1(ref_1_maj_135_n20), .A2(ref_1_maj_135_n19), 
        .ZN(ref_1_maj_135_n24) );
  NAND2_X1 ref_1_maj_135_U5 ( .A1(ref_1_maj_135_n24), .A2(ref_1_maj_135_n23), 
        .ZN(ref_1_maj_135_n25) );
  NAND2_X1 ref_1_maj_135_U4 ( .A1(ref_1_maj_135_n20), .A2(ref_1_maj_135_n19), 
        .ZN(ref_1_maj_135_n26) );
  NAND2_X1 ref_1_maj_135_U3 ( .A1(ref_1_maj_135_n26), .A2(ref_1_maj_135_n25), 
        .ZN(ref_1_maj_135_port_o) );
  XOR2_X1 ref_1_maj_135_U2 ( .A(ref_1_maj_135_n22), .B(ref_1_maj_135_n21), .Z(
        ref_1_maj_135_n23) );
  NAND2_X1 ref_1_maj_136_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_136_n18) );
  NAND2_X1 ref_1_maj_136_U14 ( .A1(ref_1_maj_136_n21), .A2(ref_1_maj_136_n22), 
        .ZN(ref_1_maj_136_n17) );
  NAND2_X1 ref_1_maj_136_U13 ( .A1(ref_1_maj_136_n18), .A2(ref_1_maj_136_n17), 
        .ZN(ref_1_maj_136_n19) );
  NAND2_X1 ref_1_maj_136_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_136_n16), .ZN(
        ref_1_maj_136_n14) );
  NAND2_X1 ref_1_maj_136_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_136_n15) );
  NAND2_X1 ref_1_maj_136_U10 ( .A1(ref_1_maj_136_n15), .A2(ref_1_maj_136_n14), 
        .ZN(ref_1_maj_136_n20) );
  XOR2_X1 ref_1_maj_136_U9 ( .A(ref_1_n15), .B(ref_1_maj_136_n16), .Z(
        ref_1_maj_136_n21) );
  XOR2_X1 ref_1_maj_136_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_136_n22) );
  XOR2_X1 ref_1_maj_136_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_136_n16) );
  OR2_X1 ref_1_maj_136_U6 ( .A1(ref_1_maj_136_n20), .A2(ref_1_maj_136_n19), 
        .ZN(ref_1_maj_136_n24) );
  NAND2_X1 ref_1_maj_136_U5 ( .A1(ref_1_maj_136_n24), .A2(ref_1_maj_136_n23), 
        .ZN(ref_1_maj_136_n25) );
  NAND2_X1 ref_1_maj_136_U4 ( .A1(ref_1_maj_136_n20), .A2(ref_1_maj_136_n19), 
        .ZN(ref_1_maj_136_n26) );
  NAND2_X1 ref_1_maj_136_U3 ( .A1(ref_1_maj_136_n26), .A2(ref_1_maj_136_n25), 
        .ZN(ref_1_maj_136_port_o) );
  XOR2_X1 ref_1_maj_136_U2 ( .A(ref_1_maj_136_n22), .B(ref_1_maj_136_n21), .Z(
        ref_1_maj_136_n23) );
  NAND2_X1 ref_1_maj_137_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_137_n18) );
  NAND2_X1 ref_1_maj_137_U14 ( .A1(ref_1_maj_137_n21), .A2(ref_1_maj_137_n22), 
        .ZN(ref_1_maj_137_n17) );
  NAND2_X1 ref_1_maj_137_U13 ( .A1(ref_1_maj_137_n18), .A2(ref_1_maj_137_n17), 
        .ZN(ref_1_maj_137_n19) );
  NAND2_X1 ref_1_maj_137_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_137_n16), .ZN(
        ref_1_maj_137_n14) );
  NAND2_X1 ref_1_maj_137_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_137_n15) );
  NAND2_X1 ref_1_maj_137_U10 ( .A1(ref_1_maj_137_n15), .A2(ref_1_maj_137_n14), 
        .ZN(ref_1_maj_137_n20) );
  XOR2_X1 ref_1_maj_137_U9 ( .A(ref_1_n15), .B(ref_1_maj_137_n16), .Z(
        ref_1_maj_137_n21) );
  XOR2_X1 ref_1_maj_137_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_137_n22) );
  XOR2_X1 ref_1_maj_137_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_137_n16) );
  OR2_X1 ref_1_maj_137_U6 ( .A1(ref_1_maj_137_n20), .A2(ref_1_maj_137_n19), 
        .ZN(ref_1_maj_137_n24) );
  NAND2_X1 ref_1_maj_137_U5 ( .A1(ref_1_maj_137_n24), .A2(ref_1_maj_137_n23), 
        .ZN(ref_1_maj_137_n25) );
  NAND2_X1 ref_1_maj_137_U4 ( .A1(ref_1_maj_137_n20), .A2(ref_1_maj_137_n19), 
        .ZN(ref_1_maj_137_n26) );
  NAND2_X1 ref_1_maj_137_U3 ( .A1(ref_1_maj_137_n26), .A2(ref_1_maj_137_n25), 
        .ZN(ref_1_maj_137_port_o) );
  XOR2_X1 ref_1_maj_137_U2 ( .A(ref_1_maj_137_n22), .B(ref_1_maj_137_n21), .Z(
        ref_1_maj_137_n23) );
  NAND2_X1 ref_1_maj_138_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_138_n18) );
  NAND2_X1 ref_1_maj_138_U14 ( .A1(ref_1_maj_138_n21), .A2(ref_1_maj_138_n22), 
        .ZN(ref_1_maj_138_n17) );
  NAND2_X1 ref_1_maj_138_U13 ( .A1(ref_1_maj_138_n18), .A2(ref_1_maj_138_n17), 
        .ZN(ref_1_maj_138_n19) );
  NAND2_X1 ref_1_maj_138_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_138_n16), .ZN(
        ref_1_maj_138_n14) );
  NAND2_X1 ref_1_maj_138_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_138_n15) );
  NAND2_X1 ref_1_maj_138_U10 ( .A1(ref_1_maj_138_n15), .A2(ref_1_maj_138_n14), 
        .ZN(ref_1_maj_138_n20) );
  XOR2_X1 ref_1_maj_138_U9 ( .A(ref_1_n15), .B(ref_1_maj_138_n16), .Z(
        ref_1_maj_138_n21) );
  XOR2_X1 ref_1_maj_138_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_138_n22) );
  XOR2_X1 ref_1_maj_138_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_138_n16) );
  OR2_X1 ref_1_maj_138_U6 ( .A1(ref_1_maj_138_n20), .A2(ref_1_maj_138_n19), 
        .ZN(ref_1_maj_138_n24) );
  NAND2_X1 ref_1_maj_138_U5 ( .A1(ref_1_maj_138_n24), .A2(ref_1_maj_138_n23), 
        .ZN(ref_1_maj_138_n25) );
  NAND2_X1 ref_1_maj_138_U4 ( .A1(ref_1_maj_138_n20), .A2(ref_1_maj_138_n19), 
        .ZN(ref_1_maj_138_n26) );
  NAND2_X1 ref_1_maj_138_U3 ( .A1(ref_1_maj_138_n26), .A2(ref_1_maj_138_n25), 
        .ZN(ref_1_maj_138_port_o) );
  XOR2_X1 ref_1_maj_138_U2 ( .A(ref_1_maj_138_n22), .B(ref_1_maj_138_n21), .Z(
        ref_1_maj_138_n23) );
  NAND2_X1 ref_1_maj_139_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_139_n18) );
  NAND2_X1 ref_1_maj_139_U14 ( .A1(ref_1_maj_139_n21), .A2(ref_1_maj_139_n22), 
        .ZN(ref_1_maj_139_n17) );
  NAND2_X1 ref_1_maj_139_U13 ( .A1(ref_1_maj_139_n18), .A2(ref_1_maj_139_n17), 
        .ZN(ref_1_maj_139_n19) );
  NAND2_X1 ref_1_maj_139_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_139_n16), .ZN(
        ref_1_maj_139_n14) );
  NAND2_X1 ref_1_maj_139_U11 ( .A1(ref_1_n11), .A2(ref_1_n13), .ZN(
        ref_1_maj_139_n15) );
  NAND2_X1 ref_1_maj_139_U10 ( .A1(ref_1_maj_139_n15), .A2(ref_1_maj_139_n14), 
        .ZN(ref_1_maj_139_n20) );
  XOR2_X1 ref_1_maj_139_U9 ( .A(ref_1_n15), .B(ref_1_maj_139_n16), .Z(
        ref_1_maj_139_n21) );
  XOR2_X1 ref_1_maj_139_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(
        ref_1_maj_139_n22) );
  XOR2_X1 ref_1_maj_139_U7 ( .A(ref_1_n11), .B(ref_1_n13), .Z(
        ref_1_maj_139_n16) );
  OR2_X1 ref_1_maj_139_U6 ( .A1(ref_1_maj_139_n20), .A2(ref_1_maj_139_n19), 
        .ZN(ref_1_maj_139_n24) );
  NAND2_X1 ref_1_maj_139_U5 ( .A1(ref_1_maj_139_n24), .A2(ref_1_maj_139_n23), 
        .ZN(ref_1_maj_139_n25) );
  NAND2_X1 ref_1_maj_139_U4 ( .A1(ref_1_maj_139_n20), .A2(ref_1_maj_139_n19), 
        .ZN(ref_1_maj_139_n26) );
  NAND2_X1 ref_1_maj_139_U3 ( .A1(ref_1_maj_139_n26), .A2(ref_1_maj_139_n25), 
        .ZN(ref_1_maj_139_port_o) );
  XOR2_X1 ref_1_maj_139_U2 ( .A(ref_1_maj_139_n22), .B(ref_1_maj_139_n21), .Z(
        ref_1_maj_139_n23) );
  NAND2_X1 ref_1_maj_140_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_140_n18) );
  NAND2_X1 ref_1_maj_140_U14 ( .A1(ref_1_maj_140_n21), .A2(ref_1_maj_140_n22), 
        .ZN(ref_1_maj_140_n17) );
  NAND2_X1 ref_1_maj_140_U13 ( .A1(ref_1_maj_140_n18), .A2(ref_1_maj_140_n17), 
        .ZN(ref_1_maj_140_n19) );
  NAND2_X1 ref_1_maj_140_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_140_n16), .ZN(
        ref_1_maj_140_n14) );
  NAND2_X1 ref_1_maj_140_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_140_n15) );
  NAND2_X1 ref_1_maj_140_U10 ( .A1(ref_1_maj_140_n15), .A2(ref_1_maj_140_n14), 
        .ZN(ref_1_maj_140_n20) );
  XOR2_X1 ref_1_maj_140_U9 ( .A(ref_1_n5), .B(ref_1_maj_140_n16), .Z(
        ref_1_maj_140_n21) );
  XOR2_X1 ref_1_maj_140_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_140_n22)
         );
  XOR2_X1 ref_1_maj_140_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_140_n16)
         );
  OR2_X1 ref_1_maj_140_U6 ( .A1(ref_1_maj_140_n20), .A2(ref_1_maj_140_n19), 
        .ZN(ref_1_maj_140_n24) );
  NAND2_X1 ref_1_maj_140_U5 ( .A1(ref_1_maj_140_n24), .A2(ref_1_maj_140_n23), 
        .ZN(ref_1_maj_140_n25) );
  NAND2_X1 ref_1_maj_140_U4 ( .A1(ref_1_maj_140_n20), .A2(ref_1_maj_140_n19), 
        .ZN(ref_1_maj_140_n26) );
  NAND2_X1 ref_1_maj_140_U3 ( .A1(ref_1_maj_140_n26), .A2(ref_1_maj_140_n25), 
        .ZN(ref_1_maj_140_port_o) );
  XOR2_X1 ref_1_maj_140_U2 ( .A(ref_1_maj_140_n22), .B(ref_1_maj_140_n21), .Z(
        ref_1_maj_140_n23) );
  NAND2_X1 ref_1_maj_141_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_141_n18) );
  NAND2_X1 ref_1_maj_141_U14 ( .A1(ref_1_maj_141_n21), .A2(ref_1_maj_141_n22), 
        .ZN(ref_1_maj_141_n17) );
  NAND2_X1 ref_1_maj_141_U13 ( .A1(ref_1_maj_141_n18), .A2(ref_1_maj_141_n17), 
        .ZN(ref_1_maj_141_n19) );
  NAND2_X1 ref_1_maj_141_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_141_n16), .ZN(
        ref_1_maj_141_n14) );
  NAND2_X1 ref_1_maj_141_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_141_n15) );
  NAND2_X1 ref_1_maj_141_U10 ( .A1(ref_1_maj_141_n15), .A2(ref_1_maj_141_n14), 
        .ZN(ref_1_maj_141_n20) );
  XOR2_X1 ref_1_maj_141_U9 ( .A(ref_1_n5), .B(ref_1_maj_141_n16), .Z(
        ref_1_maj_141_n21) );
  XOR2_X1 ref_1_maj_141_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_141_n22)
         );
  XOR2_X1 ref_1_maj_141_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_141_n16)
         );
  OR2_X1 ref_1_maj_141_U6 ( .A1(ref_1_maj_141_n20), .A2(ref_1_maj_141_n19), 
        .ZN(ref_1_maj_141_n24) );
  NAND2_X1 ref_1_maj_141_U5 ( .A1(ref_1_maj_141_n24), .A2(ref_1_maj_141_n23), 
        .ZN(ref_1_maj_141_n25) );
  NAND2_X1 ref_1_maj_141_U4 ( .A1(ref_1_maj_141_n20), .A2(ref_1_maj_141_n19), 
        .ZN(ref_1_maj_141_n26) );
  NAND2_X1 ref_1_maj_141_U3 ( .A1(ref_1_maj_141_n26), .A2(ref_1_maj_141_n25), 
        .ZN(ref_1_maj_141_port_o) );
  XOR2_X1 ref_1_maj_141_U2 ( .A(ref_1_maj_141_n22), .B(ref_1_maj_141_n21), .Z(
        ref_1_maj_141_n23) );
  NAND2_X1 ref_1_maj_142_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_142_n18) );
  NAND2_X1 ref_1_maj_142_U14 ( .A1(ref_1_maj_142_n21), .A2(ref_1_maj_142_n22), 
        .ZN(ref_1_maj_142_n17) );
  NAND2_X1 ref_1_maj_142_U13 ( .A1(ref_1_maj_142_n18), .A2(ref_1_maj_142_n17), 
        .ZN(ref_1_maj_142_n19) );
  NAND2_X1 ref_1_maj_142_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_142_n16), .ZN(
        ref_1_maj_142_n14) );
  NAND2_X1 ref_1_maj_142_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_142_n15) );
  NAND2_X1 ref_1_maj_142_U10 ( .A1(ref_1_maj_142_n15), .A2(ref_1_maj_142_n14), 
        .ZN(ref_1_maj_142_n20) );
  XOR2_X1 ref_1_maj_142_U9 ( .A(ref_1_n5), .B(ref_1_maj_142_n16), .Z(
        ref_1_maj_142_n21) );
  XOR2_X1 ref_1_maj_142_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_142_n22)
         );
  XOR2_X1 ref_1_maj_142_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_142_n16)
         );
  OR2_X1 ref_1_maj_142_U6 ( .A1(ref_1_maj_142_n20), .A2(ref_1_maj_142_n19), 
        .ZN(ref_1_maj_142_n24) );
  NAND2_X1 ref_1_maj_142_U5 ( .A1(ref_1_maj_142_n24), .A2(ref_1_maj_142_n23), 
        .ZN(ref_1_maj_142_n25) );
  NAND2_X1 ref_1_maj_142_U4 ( .A1(ref_1_maj_142_n20), .A2(ref_1_maj_142_n19), 
        .ZN(ref_1_maj_142_n26) );
  NAND2_X1 ref_1_maj_142_U3 ( .A1(ref_1_maj_142_n26), .A2(ref_1_maj_142_n25), 
        .ZN(ref_1_maj_142_port_o) );
  XOR2_X1 ref_1_maj_142_U2 ( .A(ref_1_maj_142_n22), .B(ref_1_maj_142_n21), .Z(
        ref_1_maj_142_n23) );
  NAND2_X1 ref_1_maj_143_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_143_n18) );
  NAND2_X1 ref_1_maj_143_U14 ( .A1(ref_1_maj_143_n21), .A2(ref_1_maj_143_n22), 
        .ZN(ref_1_maj_143_n17) );
  NAND2_X1 ref_1_maj_143_U13 ( .A1(ref_1_maj_143_n18), .A2(ref_1_maj_143_n17), 
        .ZN(ref_1_maj_143_n19) );
  NAND2_X1 ref_1_maj_143_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_143_n16), .ZN(
        ref_1_maj_143_n14) );
  NAND2_X1 ref_1_maj_143_U11 ( .A1(ref_1_n1), .A2(ref_1_n3), .ZN(
        ref_1_maj_143_n15) );
  NAND2_X1 ref_1_maj_143_U10 ( .A1(ref_1_maj_143_n15), .A2(ref_1_maj_143_n14), 
        .ZN(ref_1_maj_143_n20) );
  XOR2_X1 ref_1_maj_143_U9 ( .A(ref_1_n5), .B(ref_1_maj_143_n16), .Z(
        ref_1_maj_143_n21) );
  XOR2_X1 ref_1_maj_143_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_143_n22)
         );
  XOR2_X1 ref_1_maj_143_U7 ( .A(ref_1_n1), .B(ref_1_n3), .Z(ref_1_maj_143_n16)
         );
  OR2_X1 ref_1_maj_143_U6 ( .A1(ref_1_maj_143_n20), .A2(ref_1_maj_143_n19), 
        .ZN(ref_1_maj_143_n24) );
  NAND2_X1 ref_1_maj_143_U5 ( .A1(ref_1_maj_143_n24), .A2(ref_1_maj_143_n23), 
        .ZN(ref_1_maj_143_n25) );
  NAND2_X1 ref_1_maj_143_U4 ( .A1(ref_1_maj_143_n20), .A2(ref_1_maj_143_n19), 
        .ZN(ref_1_maj_143_n26) );
  NAND2_X1 ref_1_maj_143_U3 ( .A1(ref_1_maj_143_n26), .A2(ref_1_maj_143_n25), 
        .ZN(ref_1_maj_143_port_o) );
  XOR2_X1 ref_1_maj_143_U2 ( .A(ref_1_maj_143_n22), .B(ref_1_maj_143_n21), .Z(
        ref_1_maj_143_n23) );
  NAND2_X1 ref_1_maj_144_U15 ( .A1(ref_1_n37), .A2(ref_1_n39), .ZN(
        ref_1_maj_144_n18) );
  NAND2_X1 ref_1_maj_144_U14 ( .A1(ref_1_maj_144_n21), .A2(ref_1_maj_144_n22), 
        .ZN(ref_1_maj_144_n17) );
  NAND2_X1 ref_1_maj_144_U13 ( .A1(ref_1_maj_144_n18), .A2(ref_1_maj_144_n17), 
        .ZN(ref_1_maj_144_n19) );
  NAND2_X1 ref_1_maj_144_U12 ( .A1(ref_1_n35), .A2(ref_1_maj_144_n16), .ZN(
        ref_1_maj_144_n14) );
  NAND2_X1 ref_1_maj_144_U11 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_144_n15) );
  NAND2_X1 ref_1_maj_144_U10 ( .A1(ref_1_maj_144_n15), .A2(ref_1_maj_144_n14), 
        .ZN(ref_1_maj_144_n20) );
  XOR2_X1 ref_1_maj_144_U9 ( .A(ref_1_n35), .B(ref_1_maj_144_n16), .Z(
        ref_1_maj_144_n21) );
  XOR2_X1 ref_1_maj_144_U8 ( .A(ref_1_n37), .B(ref_1_n39), .Z(
        ref_1_maj_144_n22) );
  XOR2_X1 ref_1_maj_144_U7 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_144_n16) );
  OR2_X1 ref_1_maj_144_U6 ( .A1(ref_1_maj_144_n20), .A2(ref_1_maj_144_n19), 
        .ZN(ref_1_maj_144_n24) );
  NAND2_X1 ref_1_maj_144_U5 ( .A1(ref_1_maj_144_n24), .A2(ref_1_maj_144_n23), 
        .ZN(ref_1_maj_144_n25) );
  NAND2_X1 ref_1_maj_144_U4 ( .A1(ref_1_maj_144_n20), .A2(ref_1_maj_144_n19), 
        .ZN(ref_1_maj_144_n26) );
  NAND2_X1 ref_1_maj_144_U3 ( .A1(ref_1_maj_144_n26), .A2(ref_1_maj_144_n25), 
        .ZN(ref_1_maj_144_port_o) );
  XOR2_X1 ref_1_maj_144_U2 ( .A(ref_1_maj_144_n22), .B(ref_1_maj_144_n21), .Z(
        ref_1_maj_144_n23) );
  NAND2_X1 ref_1_maj_145_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_145_n18) );
  NAND2_X1 ref_1_maj_145_U14 ( .A1(ref_1_maj_145_n21), .A2(ref_1_maj_145_n22), 
        .ZN(ref_1_maj_145_n17) );
  NAND2_X1 ref_1_maj_145_U13 ( .A1(ref_1_maj_145_n18), .A2(ref_1_maj_145_n17), 
        .ZN(ref_1_maj_145_n19) );
  NAND2_X1 ref_1_maj_145_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_145_n16), .ZN(
        ref_1_maj_145_n14) );
  NAND2_X1 ref_1_maj_145_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_145_n15) );
  NAND2_X1 ref_1_maj_145_U10 ( .A1(ref_1_maj_145_n15), .A2(ref_1_maj_145_n14), 
        .ZN(ref_1_maj_145_n20) );
  XOR2_X1 ref_1_maj_145_U9 ( .A(ref_1_n36), .B(ref_1_maj_145_n16), .Z(
        ref_1_maj_145_n21) );
  XOR2_X1 ref_1_maj_145_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_145_n22) );
  XOR2_X1 ref_1_maj_145_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_145_n16) );
  OR2_X1 ref_1_maj_145_U6 ( .A1(ref_1_maj_145_n20), .A2(ref_1_maj_145_n19), 
        .ZN(ref_1_maj_145_n24) );
  NAND2_X1 ref_1_maj_145_U5 ( .A1(ref_1_maj_145_n24), .A2(ref_1_maj_145_n23), 
        .ZN(ref_1_maj_145_n25) );
  NAND2_X1 ref_1_maj_145_U4 ( .A1(ref_1_maj_145_n20), .A2(ref_1_maj_145_n19), 
        .ZN(ref_1_maj_145_n26) );
  NAND2_X1 ref_1_maj_145_U3 ( .A1(ref_1_maj_145_n26), .A2(ref_1_maj_145_n25), 
        .ZN(ref_1_maj_145_port_o) );
  XOR2_X1 ref_1_maj_145_U2 ( .A(ref_1_maj_145_n22), .B(ref_1_maj_145_n21), .Z(
        ref_1_maj_145_n23) );
  NAND2_X1 ref_1_maj_146_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_146_n18) );
  NAND2_X1 ref_1_maj_146_U14 ( .A1(ref_1_maj_146_n21), .A2(ref_1_maj_146_n22), 
        .ZN(ref_1_maj_146_n17) );
  NAND2_X1 ref_1_maj_146_U13 ( .A1(ref_1_maj_146_n18), .A2(ref_1_maj_146_n17), 
        .ZN(ref_1_maj_146_n19) );
  NAND2_X1 ref_1_maj_146_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_146_n16), .ZN(
        ref_1_maj_146_n14) );
  NAND2_X1 ref_1_maj_146_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_146_n15) );
  NAND2_X1 ref_1_maj_146_U10 ( .A1(ref_1_maj_146_n15), .A2(ref_1_maj_146_n14), 
        .ZN(ref_1_maj_146_n20) );
  XOR2_X1 ref_1_maj_146_U9 ( .A(ref_1_n36), .B(ref_1_maj_146_n16), .Z(
        ref_1_maj_146_n21) );
  XOR2_X1 ref_1_maj_146_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_146_n22) );
  XOR2_X1 ref_1_maj_146_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_146_n16) );
  OR2_X1 ref_1_maj_146_U6 ( .A1(ref_1_maj_146_n20), .A2(ref_1_maj_146_n19), 
        .ZN(ref_1_maj_146_n24) );
  NAND2_X1 ref_1_maj_146_U5 ( .A1(ref_1_maj_146_n24), .A2(ref_1_maj_146_n23), 
        .ZN(ref_1_maj_146_n25) );
  NAND2_X1 ref_1_maj_146_U4 ( .A1(ref_1_maj_146_n20), .A2(ref_1_maj_146_n19), 
        .ZN(ref_1_maj_146_n26) );
  NAND2_X1 ref_1_maj_146_U3 ( .A1(ref_1_maj_146_n26), .A2(ref_1_maj_146_n25), 
        .ZN(ref_1_maj_146_port_o) );
  XOR2_X1 ref_1_maj_146_U2 ( .A(ref_1_maj_146_n22), .B(ref_1_maj_146_n21), .Z(
        ref_1_maj_146_n23) );
  NAND2_X1 ref_1_maj_147_U15 ( .A1(ref_1_n38), .A2(ref_1_n40), .ZN(
        ref_1_maj_147_n18) );
  NAND2_X1 ref_1_maj_147_U14 ( .A1(ref_1_maj_147_n21), .A2(ref_1_maj_147_n22), 
        .ZN(ref_1_maj_147_n17) );
  NAND2_X1 ref_1_maj_147_U13 ( .A1(ref_1_maj_147_n18), .A2(ref_1_maj_147_n17), 
        .ZN(ref_1_maj_147_n19) );
  NAND2_X1 ref_1_maj_147_U12 ( .A1(ref_1_n36), .A2(ref_1_maj_147_n16), .ZN(
        ref_1_maj_147_n14) );
  NAND2_X1 ref_1_maj_147_U11 ( .A1(ref_1_n32), .A2(ref_1_n34), .ZN(
        ref_1_maj_147_n15) );
  NAND2_X1 ref_1_maj_147_U10 ( .A1(ref_1_maj_147_n15), .A2(ref_1_maj_147_n14), 
        .ZN(ref_1_maj_147_n20) );
  XOR2_X1 ref_1_maj_147_U9 ( .A(ref_1_n36), .B(ref_1_maj_147_n16), .Z(
        ref_1_maj_147_n21) );
  XOR2_X1 ref_1_maj_147_U8 ( .A(ref_1_n38), .B(ref_1_n40), .Z(
        ref_1_maj_147_n22) );
  XOR2_X1 ref_1_maj_147_U7 ( .A(ref_1_n32), .B(ref_1_n34), .Z(
        ref_1_maj_147_n16) );
  OR2_X1 ref_1_maj_147_U6 ( .A1(ref_1_maj_147_n20), .A2(ref_1_maj_147_n19), 
        .ZN(ref_1_maj_147_n24) );
  NAND2_X1 ref_1_maj_147_U5 ( .A1(ref_1_maj_147_n24), .A2(ref_1_maj_147_n23), 
        .ZN(ref_1_maj_147_n25) );
  NAND2_X1 ref_1_maj_147_U4 ( .A1(ref_1_maj_147_n20), .A2(ref_1_maj_147_n19), 
        .ZN(ref_1_maj_147_n26) );
  NAND2_X1 ref_1_maj_147_U3 ( .A1(ref_1_maj_147_n26), .A2(ref_1_maj_147_n25), 
        .ZN(ref_1_maj_147_port_o) );
  XOR2_X1 ref_1_maj_147_U2 ( .A(ref_1_maj_147_n22), .B(ref_1_maj_147_n21), .Z(
        ref_1_maj_147_n23) );
  NAND2_X1 ref_1_maj_148_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_148_n18) );
  NAND2_X1 ref_1_maj_148_U14 ( .A1(ref_1_maj_148_n21), .A2(ref_1_maj_148_n22), 
        .ZN(ref_1_maj_148_n17) );
  NAND2_X1 ref_1_maj_148_U13 ( .A1(ref_1_maj_148_n18), .A2(ref_1_maj_148_n17), 
        .ZN(ref_1_maj_148_n19) );
  NAND2_X1 ref_1_maj_148_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_148_n16), .ZN(
        ref_1_maj_148_n14) );
  NAND2_X1 ref_1_maj_148_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_148_n15) );
  NAND2_X1 ref_1_maj_148_U10 ( .A1(ref_1_maj_148_n15), .A2(ref_1_maj_148_n14), 
        .ZN(ref_1_maj_148_n20) );
  XOR2_X1 ref_1_maj_148_U9 ( .A(ref_1_n26), .B(ref_1_maj_148_n16), .Z(
        ref_1_maj_148_n21) );
  XOR2_X1 ref_1_maj_148_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_148_n22) );
  XOR2_X1 ref_1_maj_148_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_148_n16) );
  OR2_X1 ref_1_maj_148_U6 ( .A1(ref_1_maj_148_n20), .A2(ref_1_maj_148_n19), 
        .ZN(ref_1_maj_148_n24) );
  NAND2_X1 ref_1_maj_148_U5 ( .A1(ref_1_maj_148_n24), .A2(ref_1_maj_148_n23), 
        .ZN(ref_1_maj_148_n25) );
  NAND2_X1 ref_1_maj_148_U4 ( .A1(ref_1_maj_148_n20), .A2(ref_1_maj_148_n19), 
        .ZN(ref_1_maj_148_n26) );
  NAND2_X1 ref_1_maj_148_U3 ( .A1(ref_1_maj_148_n26), .A2(ref_1_maj_148_n25), 
        .ZN(ref_1_maj_148_port_o) );
  XOR2_X1 ref_1_maj_148_U2 ( .A(ref_1_maj_148_n22), .B(ref_1_maj_148_n21), .Z(
        ref_1_maj_148_n23) );
  NAND2_X1 ref_1_maj_149_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_149_n18) );
  NAND2_X1 ref_1_maj_149_U14 ( .A1(ref_1_maj_149_n21), .A2(ref_1_maj_149_n22), 
        .ZN(ref_1_maj_149_n17) );
  NAND2_X1 ref_1_maj_149_U13 ( .A1(ref_1_maj_149_n18), .A2(ref_1_maj_149_n17), 
        .ZN(ref_1_maj_149_n19) );
  NAND2_X1 ref_1_maj_149_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_149_n16), .ZN(
        ref_1_maj_149_n14) );
  NAND2_X1 ref_1_maj_149_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_149_n15) );
  NAND2_X1 ref_1_maj_149_U10 ( .A1(ref_1_maj_149_n15), .A2(ref_1_maj_149_n14), 
        .ZN(ref_1_maj_149_n20) );
  XOR2_X1 ref_1_maj_149_U9 ( .A(ref_1_n26), .B(ref_1_maj_149_n16), .Z(
        ref_1_maj_149_n21) );
  XOR2_X1 ref_1_maj_149_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_149_n22) );
  XOR2_X1 ref_1_maj_149_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_149_n16) );
  OR2_X1 ref_1_maj_149_U6 ( .A1(ref_1_maj_149_n20), .A2(ref_1_maj_149_n19), 
        .ZN(ref_1_maj_149_n24) );
  NAND2_X1 ref_1_maj_149_U5 ( .A1(ref_1_maj_149_n24), .A2(ref_1_maj_149_n23), 
        .ZN(ref_1_maj_149_n25) );
  NAND2_X1 ref_1_maj_149_U4 ( .A1(ref_1_maj_149_n20), .A2(ref_1_maj_149_n19), 
        .ZN(ref_1_maj_149_n26) );
  NAND2_X1 ref_1_maj_149_U3 ( .A1(ref_1_maj_149_n26), .A2(ref_1_maj_149_n25), 
        .ZN(ref_1_maj_149_port_o) );
  XOR2_X1 ref_1_maj_149_U2 ( .A(ref_1_maj_149_n22), .B(ref_1_maj_149_n21), .Z(
        ref_1_maj_149_n23) );
  NAND2_X1 ref_1_maj_150_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_150_n18) );
  NAND2_X1 ref_1_maj_150_U14 ( .A1(ref_1_maj_150_n21), .A2(ref_1_maj_150_n22), 
        .ZN(ref_1_maj_150_n17) );
  NAND2_X1 ref_1_maj_150_U13 ( .A1(ref_1_maj_150_n18), .A2(ref_1_maj_150_n17), 
        .ZN(ref_1_maj_150_n19) );
  NAND2_X1 ref_1_maj_150_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_150_n16), .ZN(
        ref_1_maj_150_n14) );
  NAND2_X1 ref_1_maj_150_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_150_n15) );
  NAND2_X1 ref_1_maj_150_U10 ( .A1(ref_1_maj_150_n15), .A2(ref_1_maj_150_n14), 
        .ZN(ref_1_maj_150_n20) );
  XOR2_X1 ref_1_maj_150_U9 ( .A(ref_1_n26), .B(ref_1_maj_150_n16), .Z(
        ref_1_maj_150_n21) );
  XOR2_X1 ref_1_maj_150_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_150_n22) );
  XOR2_X1 ref_1_maj_150_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_150_n16) );
  OR2_X1 ref_1_maj_150_U6 ( .A1(ref_1_maj_150_n20), .A2(ref_1_maj_150_n19), 
        .ZN(ref_1_maj_150_n24) );
  NAND2_X1 ref_1_maj_150_U5 ( .A1(ref_1_maj_150_n24), .A2(ref_1_maj_150_n23), 
        .ZN(ref_1_maj_150_n25) );
  NAND2_X1 ref_1_maj_150_U4 ( .A1(ref_1_maj_150_n20), .A2(ref_1_maj_150_n19), 
        .ZN(ref_1_maj_150_n26) );
  NAND2_X1 ref_1_maj_150_U3 ( .A1(ref_1_maj_150_n26), .A2(ref_1_maj_150_n25), 
        .ZN(ref_1_maj_150_port_o) );
  XOR2_X1 ref_1_maj_150_U2 ( .A(ref_1_maj_150_n22), .B(ref_1_maj_150_n21), .Z(
        ref_1_maj_150_n23) );
  NAND2_X1 ref_1_maj_151_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_151_n18) );
  NAND2_X1 ref_1_maj_151_U14 ( .A1(ref_1_maj_151_n21), .A2(ref_1_maj_151_n22), 
        .ZN(ref_1_maj_151_n17) );
  NAND2_X1 ref_1_maj_151_U13 ( .A1(ref_1_maj_151_n18), .A2(ref_1_maj_151_n17), 
        .ZN(ref_1_maj_151_n19) );
  NAND2_X1 ref_1_maj_151_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_151_n16), .ZN(
        ref_1_maj_151_n14) );
  NAND2_X1 ref_1_maj_151_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_151_n15) );
  NAND2_X1 ref_1_maj_151_U10 ( .A1(ref_1_maj_151_n15), .A2(ref_1_maj_151_n14), 
        .ZN(ref_1_maj_151_n20) );
  XOR2_X1 ref_1_maj_151_U9 ( .A(ref_1_n26), .B(ref_1_maj_151_n16), .Z(
        ref_1_maj_151_n21) );
  XOR2_X1 ref_1_maj_151_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(
        ref_1_maj_151_n22) );
  XOR2_X1 ref_1_maj_151_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(
        ref_1_maj_151_n16) );
  OR2_X1 ref_1_maj_151_U6 ( .A1(ref_1_maj_151_n20), .A2(ref_1_maj_151_n19), 
        .ZN(ref_1_maj_151_n24) );
  NAND2_X1 ref_1_maj_151_U5 ( .A1(ref_1_maj_151_n24), .A2(ref_1_maj_151_n23), 
        .ZN(ref_1_maj_151_n25) );
  NAND2_X1 ref_1_maj_151_U4 ( .A1(ref_1_maj_151_n20), .A2(ref_1_maj_151_n19), 
        .ZN(ref_1_maj_151_n26) );
  NAND2_X1 ref_1_maj_151_U3 ( .A1(ref_1_maj_151_n26), .A2(ref_1_maj_151_n25), 
        .ZN(ref_1_maj_151_port_o) );
  XOR2_X1 ref_1_maj_151_U2 ( .A(ref_1_maj_151_n22), .B(ref_1_maj_151_n21), .Z(
        ref_1_maj_151_n23) );
  NAND2_X1 ref_1_maj_152_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_152_n18) );
  NAND2_X1 ref_1_maj_152_U14 ( .A1(ref_1_maj_152_n21), .A2(ref_1_maj_152_n22), 
        .ZN(ref_1_maj_152_n17) );
  NAND2_X1 ref_1_maj_152_U13 ( .A1(ref_1_maj_152_n18), .A2(ref_1_maj_152_n17), 
        .ZN(ref_1_maj_152_n19) );
  NAND2_X1 ref_1_maj_152_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_152_n16), .ZN(
        ref_1_maj_152_n14) );
  NAND2_X1 ref_1_maj_152_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_152_n15) );
  NAND2_X1 ref_1_maj_152_U10 ( .A1(ref_1_maj_152_n15), .A2(ref_1_maj_152_n14), 
        .ZN(ref_1_maj_152_n20) );
  XOR2_X1 ref_1_maj_152_U9 ( .A(ref_1_n16), .B(ref_1_maj_152_n16), .Z(
        ref_1_maj_152_n21) );
  XOR2_X1 ref_1_maj_152_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_152_n22) );
  XOR2_X1 ref_1_maj_152_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_152_n16) );
  OR2_X1 ref_1_maj_152_U6 ( .A1(ref_1_maj_152_n20), .A2(ref_1_maj_152_n19), 
        .ZN(ref_1_maj_152_n24) );
  NAND2_X1 ref_1_maj_152_U5 ( .A1(ref_1_maj_152_n24), .A2(ref_1_maj_152_n23), 
        .ZN(ref_1_maj_152_n25) );
  NAND2_X1 ref_1_maj_152_U4 ( .A1(ref_1_maj_152_n20), .A2(ref_1_maj_152_n19), 
        .ZN(ref_1_maj_152_n26) );
  NAND2_X1 ref_1_maj_152_U3 ( .A1(ref_1_maj_152_n26), .A2(ref_1_maj_152_n25), 
        .ZN(ref_1_maj_152_port_o) );
  XOR2_X1 ref_1_maj_152_U2 ( .A(ref_1_maj_152_n22), .B(ref_1_maj_152_n21), .Z(
        ref_1_maj_152_n23) );
  NAND2_X1 ref_1_maj_153_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_153_n18) );
  NAND2_X1 ref_1_maj_153_U14 ( .A1(ref_1_maj_153_n21), .A2(ref_1_maj_153_n22), 
        .ZN(ref_1_maj_153_n17) );
  NAND2_X1 ref_1_maj_153_U13 ( .A1(ref_1_maj_153_n18), .A2(ref_1_maj_153_n17), 
        .ZN(ref_1_maj_153_n19) );
  NAND2_X1 ref_1_maj_153_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_153_n16), .ZN(
        ref_1_maj_153_n14) );
  NAND2_X1 ref_1_maj_153_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_153_n15) );
  NAND2_X1 ref_1_maj_153_U10 ( .A1(ref_1_maj_153_n15), .A2(ref_1_maj_153_n14), 
        .ZN(ref_1_maj_153_n20) );
  XOR2_X1 ref_1_maj_153_U9 ( .A(ref_1_n16), .B(ref_1_maj_153_n16), .Z(
        ref_1_maj_153_n21) );
  XOR2_X1 ref_1_maj_153_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_153_n22) );
  XOR2_X1 ref_1_maj_153_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_153_n16) );
  OR2_X1 ref_1_maj_153_U6 ( .A1(ref_1_maj_153_n20), .A2(ref_1_maj_153_n19), 
        .ZN(ref_1_maj_153_n24) );
  NAND2_X1 ref_1_maj_153_U5 ( .A1(ref_1_maj_153_n24), .A2(ref_1_maj_153_n23), 
        .ZN(ref_1_maj_153_n25) );
  NAND2_X1 ref_1_maj_153_U4 ( .A1(ref_1_maj_153_n20), .A2(ref_1_maj_153_n19), 
        .ZN(ref_1_maj_153_n26) );
  NAND2_X1 ref_1_maj_153_U3 ( .A1(ref_1_maj_153_n26), .A2(ref_1_maj_153_n25), 
        .ZN(ref_1_maj_153_port_o) );
  XOR2_X1 ref_1_maj_153_U2 ( .A(ref_1_maj_153_n22), .B(ref_1_maj_153_n21), .Z(
        ref_1_maj_153_n23) );
  NAND2_X1 ref_1_maj_154_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_154_n18) );
  NAND2_X1 ref_1_maj_154_U14 ( .A1(ref_1_maj_154_n21), .A2(ref_1_maj_154_n22), 
        .ZN(ref_1_maj_154_n17) );
  NAND2_X1 ref_1_maj_154_U13 ( .A1(ref_1_maj_154_n18), .A2(ref_1_maj_154_n17), 
        .ZN(ref_1_maj_154_n19) );
  NAND2_X1 ref_1_maj_154_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_154_n16), .ZN(
        ref_1_maj_154_n14) );
  NAND2_X1 ref_1_maj_154_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_154_n15) );
  NAND2_X1 ref_1_maj_154_U10 ( .A1(ref_1_maj_154_n15), .A2(ref_1_maj_154_n14), 
        .ZN(ref_1_maj_154_n20) );
  XOR2_X1 ref_1_maj_154_U9 ( .A(ref_1_n16), .B(ref_1_maj_154_n16), .Z(
        ref_1_maj_154_n21) );
  XOR2_X1 ref_1_maj_154_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_154_n22) );
  XOR2_X1 ref_1_maj_154_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_154_n16) );
  OR2_X1 ref_1_maj_154_U6 ( .A1(ref_1_maj_154_n20), .A2(ref_1_maj_154_n19), 
        .ZN(ref_1_maj_154_n24) );
  NAND2_X1 ref_1_maj_154_U5 ( .A1(ref_1_maj_154_n24), .A2(ref_1_maj_154_n23), 
        .ZN(ref_1_maj_154_n25) );
  NAND2_X1 ref_1_maj_154_U4 ( .A1(ref_1_maj_154_n20), .A2(ref_1_maj_154_n19), 
        .ZN(ref_1_maj_154_n26) );
  NAND2_X1 ref_1_maj_154_U3 ( .A1(ref_1_maj_154_n26), .A2(ref_1_maj_154_n25), 
        .ZN(ref_1_maj_154_port_o) );
  XOR2_X1 ref_1_maj_154_U2 ( .A(ref_1_maj_154_n22), .B(ref_1_maj_154_n21), .Z(
        ref_1_maj_154_n23) );
  NAND2_X1 ref_1_maj_155_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_155_n18) );
  NAND2_X1 ref_1_maj_155_U14 ( .A1(ref_1_maj_155_n21), .A2(ref_1_maj_155_n22), 
        .ZN(ref_1_maj_155_n17) );
  NAND2_X1 ref_1_maj_155_U13 ( .A1(ref_1_maj_155_n18), .A2(ref_1_maj_155_n17), 
        .ZN(ref_1_maj_155_n19) );
  NAND2_X1 ref_1_maj_155_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_155_n16), .ZN(
        ref_1_maj_155_n14) );
  NAND2_X1 ref_1_maj_155_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_155_n15) );
  NAND2_X1 ref_1_maj_155_U10 ( .A1(ref_1_maj_155_n15), .A2(ref_1_maj_155_n14), 
        .ZN(ref_1_maj_155_n20) );
  XOR2_X1 ref_1_maj_155_U9 ( .A(ref_1_n16), .B(ref_1_maj_155_n16), .Z(
        ref_1_maj_155_n21) );
  XOR2_X1 ref_1_maj_155_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(
        ref_1_maj_155_n22) );
  XOR2_X1 ref_1_maj_155_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(
        ref_1_maj_155_n16) );
  OR2_X1 ref_1_maj_155_U6 ( .A1(ref_1_maj_155_n20), .A2(ref_1_maj_155_n19), 
        .ZN(ref_1_maj_155_n24) );
  NAND2_X1 ref_1_maj_155_U5 ( .A1(ref_1_maj_155_n24), .A2(ref_1_maj_155_n23), 
        .ZN(ref_1_maj_155_n25) );
  NAND2_X1 ref_1_maj_155_U4 ( .A1(ref_1_maj_155_n20), .A2(ref_1_maj_155_n19), 
        .ZN(ref_1_maj_155_n26) );
  NAND2_X1 ref_1_maj_155_U3 ( .A1(ref_1_maj_155_n26), .A2(ref_1_maj_155_n25), 
        .ZN(ref_1_maj_155_port_o) );
  XOR2_X1 ref_1_maj_155_U2 ( .A(ref_1_maj_155_n22), .B(ref_1_maj_155_n21), .Z(
        ref_1_maj_155_n23) );
  NAND2_X1 ref_1_maj_156_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_156_n18) );
  NAND2_X1 ref_1_maj_156_U14 ( .A1(ref_1_maj_156_n21), .A2(ref_1_maj_156_n22), 
        .ZN(ref_1_maj_156_n17) );
  NAND2_X1 ref_1_maj_156_U13 ( .A1(ref_1_maj_156_n18), .A2(ref_1_maj_156_n17), 
        .ZN(ref_1_maj_156_n19) );
  NAND2_X1 ref_1_maj_156_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_156_n16), .ZN(
        ref_1_maj_156_n14) );
  NAND2_X1 ref_1_maj_156_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_156_n15) );
  NAND2_X1 ref_1_maj_156_U10 ( .A1(ref_1_maj_156_n15), .A2(ref_1_maj_156_n14), 
        .ZN(ref_1_maj_156_n20) );
  XOR2_X1 ref_1_maj_156_U9 ( .A(ref_1_n6), .B(ref_1_maj_156_n16), .Z(
        ref_1_maj_156_n21) );
  XOR2_X1 ref_1_maj_156_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_156_n22) );
  XOR2_X1 ref_1_maj_156_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_156_n16)
         );
  OR2_X1 ref_1_maj_156_U6 ( .A1(ref_1_maj_156_n20), .A2(ref_1_maj_156_n19), 
        .ZN(ref_1_maj_156_n24) );
  NAND2_X1 ref_1_maj_156_U5 ( .A1(ref_1_maj_156_n24), .A2(ref_1_maj_156_n23), 
        .ZN(ref_1_maj_156_n25) );
  NAND2_X1 ref_1_maj_156_U4 ( .A1(ref_1_maj_156_n20), .A2(ref_1_maj_156_n19), 
        .ZN(ref_1_maj_156_n26) );
  NAND2_X1 ref_1_maj_156_U3 ( .A1(ref_1_maj_156_n26), .A2(ref_1_maj_156_n25), 
        .ZN(ref_1_maj_156_port_o) );
  XOR2_X1 ref_1_maj_156_U2 ( .A(ref_1_maj_156_n22), .B(ref_1_maj_156_n21), .Z(
        ref_1_maj_156_n23) );
  NAND2_X1 ref_1_maj_157_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_157_n18) );
  NAND2_X1 ref_1_maj_157_U14 ( .A1(ref_1_maj_157_n21), .A2(ref_1_maj_157_n22), 
        .ZN(ref_1_maj_157_n17) );
  NAND2_X1 ref_1_maj_157_U13 ( .A1(ref_1_maj_157_n18), .A2(ref_1_maj_157_n17), 
        .ZN(ref_1_maj_157_n19) );
  NAND2_X1 ref_1_maj_157_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_157_n16), .ZN(
        ref_1_maj_157_n14) );
  NAND2_X1 ref_1_maj_157_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_157_n15) );
  NAND2_X1 ref_1_maj_157_U10 ( .A1(ref_1_maj_157_n15), .A2(ref_1_maj_157_n14), 
        .ZN(ref_1_maj_157_n20) );
  XOR2_X1 ref_1_maj_157_U9 ( .A(ref_1_n6), .B(ref_1_maj_157_n16), .Z(
        ref_1_maj_157_n21) );
  XOR2_X1 ref_1_maj_157_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_157_n22) );
  XOR2_X1 ref_1_maj_157_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_157_n16)
         );
  OR2_X1 ref_1_maj_157_U6 ( .A1(ref_1_maj_157_n20), .A2(ref_1_maj_157_n19), 
        .ZN(ref_1_maj_157_n24) );
  NAND2_X1 ref_1_maj_157_U5 ( .A1(ref_1_maj_157_n24), .A2(ref_1_maj_157_n23), 
        .ZN(ref_1_maj_157_n25) );
  NAND2_X1 ref_1_maj_157_U4 ( .A1(ref_1_maj_157_n20), .A2(ref_1_maj_157_n19), 
        .ZN(ref_1_maj_157_n26) );
  NAND2_X1 ref_1_maj_157_U3 ( .A1(ref_1_maj_157_n26), .A2(ref_1_maj_157_n25), 
        .ZN(ref_1_maj_157_port_o) );
  XOR2_X1 ref_1_maj_157_U2 ( .A(ref_1_maj_157_n22), .B(ref_1_maj_157_n21), .Z(
        ref_1_maj_157_n23) );
  NAND2_X1 ref_1_maj_158_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_158_n18) );
  NAND2_X1 ref_1_maj_158_U14 ( .A1(ref_1_maj_158_n21), .A2(ref_1_maj_158_n22), 
        .ZN(ref_1_maj_158_n17) );
  NAND2_X1 ref_1_maj_158_U13 ( .A1(ref_1_maj_158_n18), .A2(ref_1_maj_158_n17), 
        .ZN(ref_1_maj_158_n19) );
  NAND2_X1 ref_1_maj_158_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_158_n16), .ZN(
        ref_1_maj_158_n14) );
  NAND2_X1 ref_1_maj_158_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_158_n15) );
  NAND2_X1 ref_1_maj_158_U10 ( .A1(ref_1_maj_158_n15), .A2(ref_1_maj_158_n14), 
        .ZN(ref_1_maj_158_n20) );
  XOR2_X1 ref_1_maj_158_U9 ( .A(ref_1_n6), .B(ref_1_maj_158_n16), .Z(
        ref_1_maj_158_n21) );
  XOR2_X1 ref_1_maj_158_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_158_n22) );
  XOR2_X1 ref_1_maj_158_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_158_n16)
         );
  OR2_X1 ref_1_maj_158_U6 ( .A1(ref_1_maj_158_n20), .A2(ref_1_maj_158_n19), 
        .ZN(ref_1_maj_158_n24) );
  NAND2_X1 ref_1_maj_158_U5 ( .A1(ref_1_maj_158_n24), .A2(ref_1_maj_158_n23), 
        .ZN(ref_1_maj_158_n25) );
  NAND2_X1 ref_1_maj_158_U4 ( .A1(ref_1_maj_158_n20), .A2(ref_1_maj_158_n19), 
        .ZN(ref_1_maj_158_n26) );
  NAND2_X1 ref_1_maj_158_U3 ( .A1(ref_1_maj_158_n26), .A2(ref_1_maj_158_n25), 
        .ZN(ref_1_maj_158_port_o) );
  XOR2_X1 ref_1_maj_158_U2 ( .A(ref_1_maj_158_n22), .B(ref_1_maj_158_n21), .Z(
        ref_1_maj_158_n23) );
  NAND2_X1 ref_1_maj_159_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_159_n18) );
  NAND2_X1 ref_1_maj_159_U14 ( .A1(ref_1_maj_159_n21), .A2(ref_1_maj_159_n22), 
        .ZN(ref_1_maj_159_n17) );
  NAND2_X1 ref_1_maj_159_U13 ( .A1(ref_1_maj_159_n18), .A2(ref_1_maj_159_n17), 
        .ZN(ref_1_maj_159_n19) );
  NAND2_X1 ref_1_maj_159_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_159_n16), .ZN(
        ref_1_maj_159_n14) );
  NAND2_X1 ref_1_maj_159_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_159_n15) );
  NAND2_X1 ref_1_maj_159_U10 ( .A1(ref_1_maj_159_n15), .A2(ref_1_maj_159_n14), 
        .ZN(ref_1_maj_159_n20) );
  XOR2_X1 ref_1_maj_159_U9 ( .A(ref_1_n6), .B(ref_1_maj_159_n16), .Z(
        ref_1_maj_159_n21) );
  XOR2_X1 ref_1_maj_159_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_159_n22) );
  XOR2_X1 ref_1_maj_159_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_159_n16)
         );
  OR2_X1 ref_1_maj_159_U6 ( .A1(ref_1_maj_159_n20), .A2(ref_1_maj_159_n19), 
        .ZN(ref_1_maj_159_n24) );
  NAND2_X1 ref_1_maj_159_U5 ( .A1(ref_1_maj_159_n24), .A2(ref_1_maj_159_n23), 
        .ZN(ref_1_maj_159_n25) );
  NAND2_X1 ref_1_maj_159_U4 ( .A1(ref_1_maj_159_n20), .A2(ref_1_maj_159_n19), 
        .ZN(ref_1_maj_159_n26) );
  NAND2_X1 ref_1_maj_159_U3 ( .A1(ref_1_maj_159_n26), .A2(ref_1_maj_159_n25), 
        .ZN(ref_1_maj_159_port_o) );
  XOR2_X1 ref_1_maj_159_U2 ( .A(ref_1_maj_159_n22), .B(ref_1_maj_159_n21), .Z(
        ref_1_maj_159_n23) );
  XOR2_X1 simpleXor_240_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_240_port_a0), 
        .Z(simpleXor_240_port_z) );
  XOR2_X1 simpleXor_241_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_240_port_z), 
        .Z(simpleXor_241_port_z) );
  XOR2_X1 simpleXor_242_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_242_port_a0), 
        .Z(simpleXor_242_port_z) );
  XOR2_X1 simpleXor_243_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_242_port_z), 
        .Z(simpleXor_243_port_z) );
  XOR2_X1 simpleXor_244_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_244_port_a0), 
        .Z(simpleXor_244_port_z) );
  XOR2_X1 simpleXor_245_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_244_port_z), 
        .Z(simpleXor_245_port_z) );
  XOR2_X1 simpleXor_246_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_246_port_a0), 
        .Z(simpleXor_246_port_z) );
  XOR2_X1 simpleXor_247_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_246_port_z), 
        .Z(simpleXor_247_port_z) );
  XOR2_X1 simpleXor_248_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_248_port_a0), 
        .Z(simpleXor_248_port_z) );
  XOR2_X1 simpleXor_249_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_248_port_z), 
        .Z(simpleXor_249_port_z) );
  XOR2_X1 simpleXor_250_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_250_port_a0), 
        .Z(simpleXor_250_port_z) );
  XOR2_X1 simpleXor_251_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_250_port_z), 
        .Z(simpleXor_251_port_z) );
  XOR2_X1 simpleXor_252_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_252_port_a0), 
        .Z(simpleXor_252_port_z) );
  XOR2_X1 simpleXor_253_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_252_port_z), 
        .Z(simpleXor_253_port_z) );
  XOR2_X1 simpleXor_254_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_254_port_a0), 
        .Z(simpleXor_254_port_z) );
  XOR2_X1 simpleXor_255_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_254_port_z), 
        .Z(simpleXor_255_port_z) );
  XOR2_X1 simpleXor_256_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_256_port_a0), 
        .Z(simpleXor_256_port_z) );
  XOR2_X1 simpleXor_257_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_256_port_z), 
        .Z(simpleXor_257_port_z) );
  XOR2_X1 simpleXor_258_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_258_port_a0), 
        .Z(simpleXor_258_port_z) );
  XOR2_X1 simpleXor_259_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_258_port_z), 
        .Z(simpleXor_259_port_z) );
  XOR2_X1 simpleXor_260_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_260_port_a0), 
        .Z(simpleXor_260_port_z) );
  XOR2_X1 simpleXor_261_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_260_port_z), 
        .Z(simpleXor_261_port_z) );
  XOR2_X1 simpleXor_262_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_262_port_a0), 
        .Z(simpleXor_262_port_z) );
  XOR2_X1 simpleXor_263_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_262_port_z), 
        .Z(simpleXor_263_port_z) );
  XOR2_X1 simpleXor_264_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_264_port_a0), 
        .Z(simpleXor_264_port_z) );
  XOR2_X1 simpleXor_265_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_264_port_z), 
        .Z(simpleXor_265_port_z) );
  XOR2_X1 simpleXor_266_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_266_port_a0), 
        .Z(simpleXor_266_port_z) );
  XOR2_X1 simpleXor_267_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_266_port_z), 
        .Z(simpleXor_267_port_z) );
  XOR2_X1 simpleXor_268_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_268_port_a0), 
        .Z(simpleXor_268_port_z) );
  XOR2_X1 simpleXor_269_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_268_port_z), 
        .Z(simpleXor_269_port_z) );
  XOR2_X1 simpleXor_270_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_270_port_a0), 
        .Z(simpleXor_270_port_z) );
  XOR2_X1 simpleXor_271_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_270_port_z), 
        .Z(simpleXor_271_port_z) );
  XOR2_X1 simpleXor_272_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_272_port_a0), 
        .Z(simpleXor_272_port_z) );
  XOR2_X1 simpleXor_273_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_272_port_z), 
        .Z(simpleXor_273_port_z) );
  XOR2_X1 simpleXor_274_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_274_port_a0), 
        .Z(simpleXor_274_port_z) );
  XOR2_X1 simpleXor_275_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_274_port_z), 
        .Z(simpleXor_275_port_z) );
  XOR2_X1 simpleXor_276_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_276_port_a0), 
        .Z(simpleXor_276_port_z) );
  XOR2_X1 simpleXor_277_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_276_port_z), 
        .Z(simpleXor_277_port_z) );
  XOR2_X1 simpleXor_278_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_278_port_a0), 
        .Z(simpleXor_278_port_z) );
  XOR2_X1 simpleXor_279_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_278_port_z), 
        .Z(simpleXor_279_port_z) );
  XOR2_X1 simpleXor_280_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_280_port_a0), 
        .Z(simpleXor_280_port_z) );
  XOR2_X1 simpleXor_281_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_280_port_z), 
        .Z(simpleXor_281_port_z) );
  XOR2_X1 simpleXor_282_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_282_port_a0), 
        .Z(simpleXor_282_port_z) );
  XOR2_X1 simpleXor_283_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_282_port_z), 
        .Z(simpleXor_283_port_z) );
  XOR2_X1 simpleXor_284_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_284_port_a0), 
        .Z(simpleXor_284_port_z) );
  XOR2_X1 simpleXor_285_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_284_port_z), 
        .Z(simpleXor_285_port_z) );
  XOR2_X1 simpleXor_286_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_286_port_a0), 
        .Z(simpleXor_286_port_z) );
  XOR2_X1 simpleXor_287_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_286_port_z), 
        .Z(simpleXor_287_port_z) );
  XOR2_X1 simpleXor_288_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_288_port_a0), 
        .Z(simpleXor_288_port_z) );
  XOR2_X1 simpleXor_289_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_288_port_z), 
        .Z(simpleXor_289_port_z) );
  XOR2_X1 simpleXor_290_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_290_port_a0), 
        .Z(simpleXor_290_port_z) );
  XOR2_X1 simpleXor_291_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_290_port_z), 
        .Z(simpleXor_291_port_z) );
  XOR2_X1 simpleXor_292_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_292_port_a0), 
        .Z(simpleXor_292_port_z) );
  XOR2_X1 simpleXor_293_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_292_port_z), 
        .Z(simpleXor_293_port_z) );
  XOR2_X1 simpleXor_294_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_294_port_a0), 
        .Z(simpleXor_294_port_z) );
  XOR2_X1 simpleXor_295_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_294_port_z), 
        .Z(simpleXor_295_port_z) );
  XOR2_X1 simpleXor_296_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_296_port_a0), 
        .Z(simpleXor_296_port_z) );
  XOR2_X1 simpleXor_297_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_296_port_z), 
        .Z(simpleXor_297_port_z) );
  XOR2_X1 simpleXor_298_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_298_port_a0), 
        .Z(simpleXor_298_port_z) );
  XOR2_X1 simpleXor_299_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_298_port_z), 
        .Z(simpleXor_299_port_z) );
  XOR2_X1 simpleXor_300_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_300_port_a0), 
        .Z(simpleXor_300_port_z) );
  XOR2_X1 simpleXor_301_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_300_port_z), 
        .Z(simpleXor_301_port_z) );
  XOR2_X1 simpleXor_302_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_302_port_a0), 
        .Z(simpleXor_302_port_z) );
  XOR2_X1 simpleXor_303_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_302_port_z), 
        .Z(simpleXor_303_port_z) );
  XOR2_X1 simpleXor_304_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_304_port_a0), 
        .Z(simpleXor_304_port_z) );
  XOR2_X1 simpleXor_305_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_304_port_z), 
        .Z(simpleXor_305_port_z) );
  XOR2_X1 simpleXor_306_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_306_port_a0), 
        .Z(simpleXor_306_port_z) );
  XOR2_X1 simpleXor_307_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_306_port_z), 
        .Z(simpleXor_307_port_z) );
  XOR2_X1 simpleXor_308_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_308_port_a0), 
        .Z(simpleXor_308_port_z) );
  XOR2_X1 simpleXor_309_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_308_port_z), 
        .Z(simpleXor_309_port_z) );
  XOR2_X1 simpleXor_310_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_310_port_a0), 
        .Z(simpleXor_310_port_z) );
  XOR2_X1 simpleXor_311_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_310_port_z), 
        .Z(simpleXor_311_port_z) );
  XOR2_X1 simpleXor_312_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_312_port_a0), 
        .Z(simpleXor_312_port_z) );
  XOR2_X1 simpleXor_313_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_312_port_z), 
        .Z(simpleXor_313_port_z) );
  XOR2_X1 simpleXor_314_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_314_port_a0), 
        .Z(simpleXor_314_port_z) );
  XOR2_X1 simpleXor_315_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_314_port_z), 
        .Z(simpleXor_315_port_z) );
  XOR2_X1 simpleXor_316_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_316_port_a0), 
        .Z(simpleXor_316_port_z) );
  XOR2_X1 simpleXor_317_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_316_port_z), 
        .Z(simpleXor_317_port_z) );
  XOR2_X1 simpleXor_318_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_318_port_a0), 
        .Z(simpleXor_318_port_z) );
  XOR2_X1 simpleXor_319_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_318_port_z), 
        .Z(simpleXor_319_port_z) );
  XOR2_X1 simpleXor_320_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_320_port_a0), 
        .Z(simpleXor_320_port_z) );
  XOR2_X1 simpleXor_321_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_320_port_z), 
        .Z(simpleXor_321_port_z) );
  XOR2_X1 simpleXor_322_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_322_port_a0), 
        .Z(simpleXor_322_port_z) );
  XOR2_X1 simpleXor_323_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_322_port_z), 
        .Z(simpleXor_323_port_z) );
  XOR2_X1 simpleXor_324_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_324_port_a0), 
        .Z(simpleXor_324_port_z) );
  XOR2_X1 simpleXor_325_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_324_port_z), 
        .Z(simpleXor_325_port_z) );
  XOR2_X1 simpleXor_326_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_326_port_a0), 
        .Z(simpleXor_326_port_z) );
  XOR2_X1 simpleXor_327_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_326_port_z), 
        .Z(simpleXor_327_port_z) );
  XOR2_X1 simpleXor_328_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_328_port_a0), 
        .Z(simpleXor_328_port_z) );
  XOR2_X1 simpleXor_329_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_328_port_z), 
        .Z(simpleXor_329_port_z) );
  XOR2_X1 simpleXor_330_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_330_port_a0), 
        .Z(simpleXor_330_port_z) );
  XOR2_X1 simpleXor_331_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_330_port_z), 
        .Z(simpleXor_331_port_z) );
  XOR2_X1 simpleXor_332_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_332_port_a0), 
        .Z(simpleXor_332_port_z) );
  XOR2_X1 simpleXor_333_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_332_port_z), 
        .Z(simpleXor_333_port_z) );
  XOR2_X1 simpleXor_334_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_334_port_a0), 
        .Z(simpleXor_334_port_z) );
  XOR2_X1 simpleXor_335_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_334_port_z), 
        .Z(simpleXor_335_port_z) );
  XOR2_X1 simpleXor_336_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_336_port_a0), 
        .Z(simpleXor_336_port_z) );
  XOR2_X1 simpleXor_337_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_336_port_z), 
        .Z(simpleXor_337_port_z) );
  XOR2_X1 simpleXor_338_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_338_port_a0), 
        .Z(simpleXor_338_port_z) );
  XOR2_X1 simpleXor_339_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_338_port_z), 
        .Z(simpleXor_339_port_z) );
  XOR2_X1 simpleXor_340_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_340_port_a0), 
        .Z(simpleXor_340_port_z) );
  XOR2_X1 simpleXor_341_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_340_port_z), 
        .Z(simpleXor_341_port_z) );
  XOR2_X1 simpleXor_342_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_342_port_a0), 
        .Z(simpleXor_342_port_z) );
  XOR2_X1 simpleXor_343_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_342_port_z), 
        .Z(simpleXor_343_port_z) );
  XOR2_X1 simpleXor_344_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_344_port_a0), 
        .Z(simpleXor_344_port_z) );
  XOR2_X1 simpleXor_345_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_344_port_z), 
        .Z(simpleXor_345_port_z) );
  XOR2_X1 simpleXor_346_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_346_port_a0), 
        .Z(simpleXor_346_port_z) );
  XOR2_X1 simpleXor_347_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_346_port_z), 
        .Z(simpleXor_347_port_z) );
  XOR2_X1 simpleXor_348_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_348_port_a0), 
        .Z(simpleXor_348_port_z) );
  XOR2_X1 simpleXor_349_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_348_port_z), 
        .Z(simpleXor_349_port_z) );
  XOR2_X1 simpleXor_350_U1 ( .A(port_rand_mul_3[0]), .B(simpleXor_350_port_a0), 
        .Z(simpleXor_350_port_z) );
  XOR2_X1 simpleXor_351_U1 ( .A(port_rand_mul_3[1]), .B(simpleXor_350_port_z), 
        .Z(simpleXor_351_port_z) );
  XOR2_X1 simpleXor_352_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_352_port_a0), 
        .Z(simpleXor_352_port_z) );
  XOR2_X1 simpleXor_353_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_352_port_z), 
        .Z(simpleXor_353_port_z) );
  XOR2_X1 simpleXor_354_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_354_port_a0), 
        .Z(simpleXor_354_port_z) );
  XOR2_X1 simpleXor_355_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_354_port_z), 
        .Z(simpleXor_355_port_z) );
  XOR2_X1 simpleXor_356_U1 ( .A(port_rand_mul_4[0]), .B(simpleXor_356_port_a0), 
        .Z(simpleXor_356_port_z) );
  XOR2_X1 simpleXor_357_U1 ( .A(port_rand_mul_4[1]), .B(simpleXor_356_port_z), 
        .Z(simpleXor_357_port_z) );
  XOR2_X1 simpleXor_358_U1 ( .A(port_rand_mul_5[0]), .B(simpleXor_358_port_a0), 
        .Z(simpleXor_358_port_z) );
  XOR2_X1 simpleXor_359_U1 ( .A(port_rand_mul_5[1]), .B(simpleXor_358_port_z), 
        .Z(simpleXor_359_port_z) );
endmodule

