
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i0_s5, io_i0_s6, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, 
        io_i1_s4, io_i1_s5, io_i1_s6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, 
        p_rand_4, p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, 
        p_rand_11, p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16, 
        p_rand_17, p_rand_18, p_rand_19, p_rand_20, io_o0_s0, io_o0_s1, 
        io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5, io_o0_s6 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i0_s5, io_i0_s6, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4,
         io_i1_s5, io_i1_s6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4,
         p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10,
         p_rand_11, p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16,
         p_rand_17, p_rand_18, p_rand_19, p_rand_20;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5, io_o0_s6;
  wire   n_hpc2_0_n287, n_hpc2_0_n286, n_hpc2_0_n285, n_hpc2_0_n284,
         n_hpc2_0_n283, n_hpc2_0_n282, n_hpc2_0_n281, n_hpc2_0_n280,
         n_hpc2_0_n279, n_hpc2_0_n278, n_hpc2_0_n277, n_hpc2_0_n276,
         n_hpc2_0_n275, n_hpc2_0_n274, n_hpc2_0_n273, n_hpc2_0_n272,
         n_hpc2_0_n271, n_hpc2_0_n270, n_hpc2_0_n269, n_hpc2_0_n268,
         n_hpc2_0_n267, n_hpc2_0_n266, n_hpc2_0_n265, n_hpc2_0_n264,
         n_hpc2_0_n263, n_hpc2_0_n262, n_hpc2_0_n261, n_hpc2_0_n260,
         n_hpc2_0_n259, n_hpc2_0_n258, n_hpc2_0_n257, n_hpc2_0_n256,
         n_hpc2_0_n255, n_hpc2_0_n254, n_hpc2_0_n253, n_hpc2_0_n252,
         n_hpc2_0_n251, n_hpc2_0_n250, n_hpc2_0_n249, n_hpc2_0_n248,
         n_hpc2_0_n247, n_hpc2_0_n246, n_hpc2_0_n245, n_hpc2_0_n244,
         n_hpc2_0_n243, n_hpc2_0_n242, n_hpc2_0_n241, n_hpc2_0_n240,
         n_hpc2_0_n239, n_hpc2_0_n238, n_hpc2_0_n237, n_hpc2_0_n236,
         n_hpc2_0_n235, n_hpc2_0_n234, n_hpc2_0_n233, n_hpc2_0_n232,
         n_hpc2_0_n231, n_hpc2_0_n230, n_hpc2_0_n229, n_hpc2_0_n228,
         n_hpc2_0_n227, n_hpc2_0_n226, n_hpc2_0_n225, n_hpc2_0_n224,
         n_hpc2_0_n223, n_hpc2_0_n222, n_hpc2_0_n221, n_hpc2_0_n220,
         n_hpc2_0_n219, n_hpc2_0_n218, n_hpc2_0_n217, n_hpc2_0_n216,
         n_hpc2_0_n215, n_hpc2_0_n214, n_hpc2_0_n213, n_hpc2_0_n212,
         n_hpc2_0_n211, n_hpc2_0_n210, n_hpc2_0_n209, n_hpc2_0_n208,
         n_hpc2_0_n207, n_hpc2_0_n206, n_hpc2_0_n205, n_hpc2_0_n204,
         n_hpc2_0_n203, n_hpc2_0_n202, n_hpc2_0_n201, n_hpc2_0_n200,
         n_hpc2_0_n199, n_hpc2_0_n198, n_hpc2_0_n197, n_hpc2_0_n196,
         n_hpc2_0_n195, n_hpc2_0_n194, n_hpc2_0_n193, n_hpc2_0_n192,
         n_hpc2_0_n191, n_hpc2_0_n190, n_hpc2_0_n189, n_hpc2_0_n188,
         n_hpc2_0_n187, n_hpc2_0_n186, n_hpc2_0_n185, n_hpc2_0_n184,
         n_hpc2_0_n183, n_hpc2_0_n182, n_hpc2_0_n181, n_hpc2_0_n180,
         n_hpc2_0_n179, n_hpc2_0_n178, n_hpc2_0_n177, n_hpc2_0_n176,
         n_hpc2_0_n175, n_hpc2_0_n174, n_hpc2_0_n173, n_hpc2_0_n172,
         n_hpc2_0_n171, n_hpc2_0_n170, n_hpc2_0_n169, n_hpc2_0_n168,
         n_hpc2_0_n167, n_hpc2_0_n166, n_hpc2_0_n165, n_hpc2_0_n164,
         n_hpc2_0_n163, n_hpc2_0_n162, n_hpc2_0_n161, n_hpc2_0_n160,
         n_hpc2_0_n159, n_hpc2_0_n158, n_hpc2_0_n157, n_hpc2_0_n156,
         n_hpc2_0_n155, n_hpc2_0_n154, n_hpc2_0_n153, n_hpc2_0_n152,
         n_hpc2_0_n151, n_hpc2_0_n150, n_hpc2_0_n149, n_hpc2_0_n148,
         n_hpc2_0_n147, n_hpc2_0_n146, n_hpc2_0_n145, n_hpc2_0_n144,
         n_hpc2_0_n143, n_hpc2_0_n142, n_hpc2_0_n141, n_hpc2_0_n140,
         n_hpc2_0_n139, n_hpc2_0_n138, n_hpc2_0_n137, n_hpc2_0_n136,
         n_hpc2_0_n135, n_hpc2_0_n134, n_hpc2_0_n133, n_hpc2_0_n132,
         n_hpc2_0_n131, n_hpc2_0_n130, n_hpc2_0_n129, n_hpc2_0_n128,
         n_hpc2_0_n127, n_hpc2_0_n126, n_hpc2_0_n125, n_hpc2_0_n124,
         n_hpc2_0_n123, n_hpc2_0_n122, n_hpc2_0_n121, n_hpc2_0_n120,
         n_hpc2_0_n119, n_hpc2_0_n118, n_hpc2_0_n117, n_hpc2_0_n116,
         n_hpc2_0_n115, n_hpc2_0_n114, n_hpc2_0_n113, n_hpc2_0_n112,
         n_hpc2_0_n111, n_hpc2_0_n110, n_hpc2_0_n109, n_hpc2_0_n108,
         n_hpc2_0_n107, n_hpc2_0_n106, n_hpc2_0_n105, n_hpc2_0_n104,
         n_hpc2_0_n103, n_hpc2_0_n102, n_hpc2_0_n101, n_hpc2_0_n100,
         n_hpc2_0_n99, n_hpc2_0_n98, n_hpc2_0_n97, n_hpc2_0_n96, n_hpc2_0_n95,
         n_hpc2_0_n94, n_hpc2_0_n93, n_hpc2_0_n92, n_hpc2_0_n91, n_hpc2_0_n90,
         n_hpc2_0_n89, n_hpc2_0_n88, n_hpc2_0_n87, n_hpc2_0_n86, n_hpc2_0_n85,
         n_hpc2_0_n84, n_hpc2_0_n83, n_hpc2_0_n82, n_hpc2_0_n81, n_hpc2_0_n80,
         n_hpc2_0_n79, n_hpc2_0_n78, n_hpc2_0_n77, n_hpc2_0_n76, n_hpc2_0_n75,
         n_hpc2_0_n74, n_hpc2_0_n73, n_hpc2_0_n72, n_hpc2_0_n71, n_hpc2_0_n70,
         n_hpc2_0_n69, n_hpc2_0_n68, n_hpc2_0_n67, n_hpc2_0_n66, n_hpc2_0_n65,
         n_hpc2_0_n64, n_hpc2_0_n63, n_hpc2_0_n62, n_hpc2_0_n61, n_hpc2_0_n60,
         n_hpc2_0_n59, n_hpc2_0_n58, n_hpc2_0_n57, n_hpc2_0_n56, n_hpc2_0_n55,
         n_hpc2_0_n54, n_hpc2_0_n53, n_hpc2_0_n52, n_hpc2_0_n51, n_hpc2_0_n50,
         n_hpc2_0_n49, n_hpc2_0_n48, n_hpc2_0_n47, n_hpc2_0_n46, n_hpc2_0_n45,
         n_hpc2_0_n44, n_hpc2_0_n43, n_hpc2_0_n42, n_hpc2_0_n41, n_hpc2_0_n40,
         n_hpc2_0_n39, n_hpc2_0_n38, n_hpc2_0_n37, n_hpc2_0_n36, n_hpc2_0_n35,
         n_hpc2_0_n34, n_hpc2_0_n33, n_hpc2_0_n32, n_hpc2_0_n31, n_hpc2_0_n30,
         n_hpc2_0_n29, n_hpc2_0_n28, n_hpc2_0_n27, n_hpc2_0_n26, n_hpc2_0_n25,
         n_hpc2_0_n24, n_hpc2_0_n23, n_hpc2_0_n22, n_hpc2_0_n21, n_hpc2_0_n20,
         n_hpc2_0_n19, n_hpc2_0_n18, n_hpc2_0_n17, n_hpc2_0_n16, n_hpc2_0_n15,
         n_hpc2_0_n14, n_hpc2_0_n13, n_hpc2_0_n12, n_hpc2_0_n11, n_hpc2_0_n10,
         n_hpc2_0_n9, n_hpc2_0_n8, n_hpc2_0_n7, n_hpc2_0_n6, n_hpc2_0_n5,
         n_hpc2_0_n4, n_hpc2_0_n3, n_hpc2_0_n2, n_hpc2_0_n1, n_hpc2_0_N139,
         n_hpc2_0_N138, n_hpc2_0_N137, n_hpc2_0_N136, n_hpc2_0_N135,
         n_hpc2_0_N134, n_hpc2_0_N133, n_hpc2_0_N132, n_hpc2_0_N131,
         n_hpc2_0_N130, n_hpc2_0_N129, n_hpc2_0_N128, n_hpc2_0_N127,
         n_hpc2_0_N126, n_hpc2_0_N125, n_hpc2_0_N124, n_hpc2_0_N123,
         n_hpc2_0_N122, n_hpc2_0_N121, n_hpc2_0_N120, n_hpc2_0_N119,
         n_hpc2_0_N118, n_hpc2_0_N117, n_hpc2_0_N116, n_hpc2_0_N115,
         n_hpc2_0_N114, n_hpc2_0_N113, n_hpc2_0_N112, n_hpc2_0_N111,
         n_hpc2_0_N110, n_hpc2_0_N109, n_hpc2_0_N108, n_hpc2_0_N107,
         n_hpc2_0_N106, n_hpc2_0_N105, n_hpc2_0_N104, n_hpc2_0_N103,
         n_hpc2_0_N102, n_hpc2_0_N101, n_hpc2_0_N100, n_hpc2_0_N99,
         n_hpc2_0_N98, n_hpc2_0_N97, n_hpc2_0_N96, n_hpc2_0_N95, n_hpc2_0_N94,
         n_hpc2_0_N93, n_hpc2_0_N92, n_hpc2_0_N91, n_hpc2_0_N90, n_hpc2_0_N89,
         n_hpc2_0_N88, n_hpc2_0_N87, n_hpc2_0_N86, n_hpc2_0_N85, n_hpc2_0_N84,
         n_hpc2_0_N83, n_hpc2_0_N82, n_hpc2_0_N81, n_hpc2_0_N80, n_hpc2_0_N79,
         n_hpc2_0_N78, n_hpc2_0_N77, n_hpc2_0_N76, n_hpc2_0_N75, n_hpc2_0_N74,
         n_hpc2_0_N73, n_hpc2_0_N72, n_hpc2_0_N71, n_hpc2_0_N70, n_hpc2_0_N69,
         n_hpc2_0_N68, n_hpc2_0_N67, n_hpc2_0_N66, n_hpc2_0_N65, n_hpc2_0_N64,
         n_hpc2_0_N63, n_hpc2_0_N62, n_hpc2_0_N61, n_hpc2_0_N60, n_hpc2_0_N59,
         n_hpc2_0_N58, n_hpc2_0_N57, n_hpc2_0_N56, n_hpc2_0_N55, n_hpc2_0_N54,
         n_hpc2_0_N53, n_hpc2_0_N52, n_hpc2_0_N51, n_hpc2_0_N50, n_hpc2_0_N49,
         n_hpc2_0_N48, n_hpc2_0_N47, n_hpc2_0_N46, n_hpc2_0_N45, n_hpc2_0_N44,
         n_hpc2_0_N43, n_hpc2_0_N42, n_hpc2_0_N41, n_hpc2_0_N40, n_hpc2_0_N39,
         n_hpc2_0_N38, n_hpc2_0_N37, n_hpc2_0_N36, n_hpc2_0_N35, n_hpc2_0_N34,
         n_hpc2_0_N33, n_hpc2_0_N32, n_hpc2_0_N31, n_hpc2_0_N30, n_hpc2_0_N29,
         n_hpc2_0_N28, n_hpc2_0_N27, n_hpc2_0_N26, n_hpc2_0_N25, n_hpc2_0_N24,
         n_hpc2_0_N23, n_hpc2_0_N22, n_hpc2_0_N21, n_hpc2_0_N20, n_hpc2_0_N19,
         n_hpc2_0_N18, n_hpc2_0_N17, n_hpc2_0_N16, n_hpc2_0_N15, n_hpc2_0_N14,
         n_hpc2_0_N13, n_hpc2_0_N12, n_hpc2_0_N11, n_hpc2_0_N10, n_hpc2_0_N9,
         n_hpc2_0_N8, n_hpc2_0_N7, n_hpc2_0__hpc_av62, n_hpc2_0__hpc_av52,
         n_hpc2_0__hpc_av42, n_hpc2_0__hpc_av32, n_hpc2_0__hpc_av23,
         n_hpc2_0__hpc_av13, n_hpc2_0__hpc_av03;

  NOR2_X1 u_hpc2_0_U226 ( .A1(n_hpc2_0_n287), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N10) );
  XOR2_X1 u_hpc2_0_U225 ( .A(io_i1_s3), .B(p_rand_2), .Z(n_hpc2_0_N100) );
  XOR2_X1 u_hpc2_0_U224 ( .A(io_i1_s4), .B(p_rand_3), .Z(n_hpc2_0_N101) );
  XOR2_X1 u_hpc2_0_U223 ( .A(io_i1_s5), .B(p_rand_4), .Z(n_hpc2_0_N102) );
  XOR2_X1 u_hpc2_0_U222 ( .A(io_i1_s6), .B(p_rand_5), .Z(n_hpc2_0_N103) );
  XOR2_X1 u_hpc2_0_U221 ( .A(io_i1_s0), .B(p_rand_0), .Z(n_hpc2_0_N104) );
  XOR2_X1 u_hpc2_0_U220 ( .A(io_i1_s2), .B(p_rand_6), .Z(n_hpc2_0_N105) );
  XOR2_X1 u_hpc2_0_U219 ( .A(io_i1_s3), .B(p_rand_7), .Z(n_hpc2_0_N106) );
  XOR2_X1 u_hpc2_0_U218 ( .A(io_i1_s4), .B(p_rand_8), .Z(n_hpc2_0_N107) );
  XOR2_X1 u_hpc2_0_U217 ( .A(io_i1_s5), .B(p_rand_9), .Z(n_hpc2_0_N108) );
  XOR2_X1 u_hpc2_0_U216 ( .A(io_i1_s6), .B(p_rand_10), .Z(n_hpc2_0_N109) );
  NOR2_X1 u_hpc2_0_U215 ( .A1(n_hpc2_0_n286), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N11) );
  XOR2_X1 u_hpc2_0_U214 ( .A(io_i1_s0), .B(p_rand_1), .Z(n_hpc2_0_N110) );
  XOR2_X1 u_hpc2_0_U213 ( .A(io_i1_s1), .B(p_rand_6), .Z(n_hpc2_0_N111) );
  XOR2_X1 u_hpc2_0_U212 ( .A(io_i1_s3), .B(p_rand_11), .Z(n_hpc2_0_N112) );
  XOR2_X1 u_hpc2_0_U211 ( .A(io_i1_s4), .B(p_rand_12), .Z(n_hpc2_0_N113) );
  XOR2_X1 u_hpc2_0_U210 ( .A(io_i1_s5), .B(p_rand_13), .Z(n_hpc2_0_N114) );
  XOR2_X1 u_hpc2_0_U209 ( .A(io_i1_s6), .B(p_rand_14), .Z(n_hpc2_0_N115) );
  XOR2_X1 u_hpc2_0_U208 ( .A(io_i1_s0), .B(p_rand_2), .Z(n_hpc2_0_N116) );
  XOR2_X1 u_hpc2_0_U207 ( .A(io_i1_s1), .B(p_rand_7), .Z(n_hpc2_0_N117) );
  XOR2_X1 u_hpc2_0_U206 ( .A(io_i1_s2), .B(p_rand_11), .Z(n_hpc2_0_N118) );
  XOR2_X1 u_hpc2_0_U205 ( .A(io_i1_s4), .B(p_rand_15), .Z(n_hpc2_0_N119) );
  NOR2_X1 u_hpc2_0_U204 ( .A1(n_hpc2_0_n285), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N12) );
  XOR2_X1 u_hpc2_0_U203 ( .A(io_i1_s5), .B(p_rand_16), .Z(n_hpc2_0_N120) );
  XOR2_X1 u_hpc2_0_U202 ( .A(io_i1_s6), .B(p_rand_17), .Z(n_hpc2_0_N121) );
  XOR2_X1 u_hpc2_0_U201 ( .A(io_i1_s0), .B(p_rand_3), .Z(n_hpc2_0_N122) );
  XOR2_X1 u_hpc2_0_U200 ( .A(io_i1_s1), .B(p_rand_8), .Z(n_hpc2_0_N123) );
  XOR2_X1 u_hpc2_0_U199 ( .A(io_i1_s2), .B(p_rand_12), .Z(n_hpc2_0_N124) );
  XOR2_X1 u_hpc2_0_U198 ( .A(io_i1_s3), .B(p_rand_15), .Z(n_hpc2_0_N125) );
  XOR2_X1 u_hpc2_0_U197 ( .A(io_i1_s5), .B(p_rand_18), .Z(n_hpc2_0_N126) );
  XOR2_X1 u_hpc2_0_U196 ( .A(io_i1_s6), .B(p_rand_19), .Z(n_hpc2_0_N127) );
  XOR2_X1 u_hpc2_0_U195 ( .A(io_i1_s0), .B(p_rand_4), .Z(n_hpc2_0_N128) );
  XOR2_X1 u_hpc2_0_U194 ( .A(io_i1_s1), .B(p_rand_9), .Z(n_hpc2_0_N129) );
  NOR2_X1 u_hpc2_0_U193 ( .A1(n_hpc2_0_n284), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N13) );
  XOR2_X1 u_hpc2_0_U192 ( .A(io_i1_s2), .B(p_rand_13), .Z(n_hpc2_0_N130) );
  XOR2_X1 u_hpc2_0_U191 ( .A(io_i1_s3), .B(p_rand_16), .Z(n_hpc2_0_N131) );
  XOR2_X1 u_hpc2_0_U190 ( .A(io_i1_s4), .B(p_rand_18), .Z(n_hpc2_0_N132) );
  XOR2_X1 u_hpc2_0_U189 ( .A(io_i1_s6), .B(p_rand_20), .Z(n_hpc2_0_N133) );
  XOR2_X1 u_hpc2_0_U188 ( .A(io_i1_s0), .B(p_rand_5), .Z(n_hpc2_0_N134) );
  XOR2_X1 u_hpc2_0_U187 ( .A(io_i1_s1), .B(p_rand_10), .Z(n_hpc2_0_N135) );
  XOR2_X1 u_hpc2_0_U186 ( .A(io_i1_s2), .B(p_rand_14), .Z(n_hpc2_0_N136) );
  XOR2_X1 u_hpc2_0_U185 ( .A(io_i1_s3), .B(p_rand_17), .Z(n_hpc2_0_N137) );
  XOR2_X1 u_hpc2_0_U184 ( .A(io_i1_s4), .B(p_rand_19), .Z(n_hpc2_0_N138) );
  XOR2_X1 u_hpc2_0_U183 ( .A(io_i1_s5), .B(p_rand_20), .Z(n_hpc2_0_N139) );
  NOR2_X1 u_hpc2_0_U182 ( .A1(n_hpc2_0_n283), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N14) );
  NOR2_X1 u_hpc2_0_U181 ( .A1(n_hpc2_0_n282), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N15) );
  NOR2_X1 u_hpc2_0_U180 ( .A1(n_hpc2_0_n281), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N16) );
  NOR2_X1 u_hpc2_0_U179 ( .A1(n_hpc2_0_n280), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N17) );
  NOR2_X1 u_hpc2_0_U178 ( .A1(n_hpc2_0_n279), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N18) );
  NOR2_X1 u_hpc2_0_U177 ( .A1(n_hpc2_0_n278), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N19) );
  NOR2_X1 u_hpc2_0_U176 ( .A1(n_hpc2_0_n277), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N20) );
  NOR2_X1 u_hpc2_0_U175 ( .A1(n_hpc2_0_n276), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N21) );
  NOR2_X1 u_hpc2_0_U174 ( .A1(n_hpc2_0_n275), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N22) );
  NOR2_X1 u_hpc2_0_U173 ( .A1(n_hpc2_0_n274), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N23) );
  NOR2_X1 u_hpc2_0_U172 ( .A1(n_hpc2_0_n273), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N24) );
  NOR2_X1 u_hpc2_0_U171 ( .A1(n_hpc2_0_n272), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N25) );
  NOR2_X1 u_hpc2_0_U170 ( .A1(n_hpc2_0_n271), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N26) );
  NOR2_X1 u_hpc2_0_U169 ( .A1(n_hpc2_0_n270), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N27) );
  NOR2_X1 u_hpc2_0_U168 ( .A1(n_hpc2_0_n269), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N28) );
  NOR2_X1 u_hpc2_0_U167 ( .A1(n_hpc2_0_n268), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N29) );
  NOR2_X1 u_hpc2_0_U166 ( .A1(n_hpc2_0_n267), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N30) );
  NOR2_X1 u_hpc2_0_U165 ( .A1(n_hpc2_0_n266), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N31) );
  NOR2_X1 u_hpc2_0_U164 ( .A1(n_hpc2_0_n265), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N32) );
  NOR2_X1 u_hpc2_0_U163 ( .A1(n_hpc2_0_n264), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N33) );
  NOR2_X1 u_hpc2_0_U162 ( .A1(n_hpc2_0_n263), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N34) );
  NOR2_X1 u_hpc2_0_U161 ( .A1(n_hpc2_0_n262), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N35) );
  NOR2_X1 u_hpc2_0_U160 ( .A1(n_hpc2_0_n261), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N36) );
  NOR2_X1 u_hpc2_0_U159 ( .A1(n_hpc2_0_n260), .A2(n_hpc2_0_n14), .ZN(
        n_hpc2_0_N37) );
  NOR2_X1 u_hpc2_0_U158 ( .A1(n_hpc2_0_n259), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N38) );
  NOR2_X1 u_hpc2_0_U157 ( .A1(n_hpc2_0_n258), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N39) );
  NOR2_X1 u_hpc2_0_U156 ( .A1(n_hpc2_0_n257), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N40) );
  NOR2_X1 u_hpc2_0_U155 ( .A1(n_hpc2_0_n256), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N41) );
  NOR2_X1 u_hpc2_0_U154 ( .A1(n_hpc2_0_n255), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N42) );
  NOR2_X1 u_hpc2_0_U153 ( .A1(n_hpc2_0_n254), .A2(n_hpc2_0_n13), .ZN(
        n_hpc2_0_N43) );
  NOR2_X1 u_hpc2_0_U152 ( .A1(n_hpc2_0_n253), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N44) );
  NOR2_X1 u_hpc2_0_U151 ( .A1(n_hpc2_0_n252), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N45) );
  NOR2_X1 u_hpc2_0_U150 ( .A1(n_hpc2_0_n251), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N46) );
  NOR2_X1 u_hpc2_0_U149 ( .A1(n_hpc2_0_n250), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N47) );
  NOR2_X1 u_hpc2_0_U148 ( .A1(n_hpc2_0_n249), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N48) );
  NOR2_X1 u_hpc2_0_U147 ( .A1(n_hpc2_0_n248), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N49) );
  NOR2_X1 u_hpc2_0_U146 ( .A1(n_hpc2_0_n247), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N50) );
  NOR2_X1 u_hpc2_0_U145 ( .A1(n_hpc2_0_n246), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N51) );
  NOR2_X1 u_hpc2_0_U144 ( .A1(n_hpc2_0_n245), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N52) );
  NOR2_X1 u_hpc2_0_U143 ( .A1(n_hpc2_0_n244), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N53) );
  NOR2_X1 u_hpc2_0_U142 ( .A1(n_hpc2_0_n243), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N54) );
  NOR2_X1 u_hpc2_0_U141 ( .A1(n_hpc2_0_n242), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N55) );
  NOR2_X1 u_hpc2_0_U140 ( .A1(n_hpc2_0_n240), .A2(n_hpc2_0_n241), .ZN(
        n_hpc2_0_N56) );
  NOR2_X1 u_hpc2_0_U139 ( .A1(n_hpc2_0_n238), .A2(n_hpc2_0_n239), .ZN(
        n_hpc2_0_N57) );
  NOR2_X1 u_hpc2_0_U138 ( .A1(n_hpc2_0_n236), .A2(n_hpc2_0_n237), .ZN(
        n_hpc2_0_N58) );
  NOR2_X1 u_hpc2_0_U137 ( .A1(n_hpc2_0_n234), .A2(n_hpc2_0_n235), .ZN(
        n_hpc2_0_N59) );
  NOR2_X1 u_hpc2_0_U136 ( .A1(n_hpc2_0_n232), .A2(n_hpc2_0_n233), .ZN(
        n_hpc2_0_N60) );
  NOR2_X1 u_hpc2_0_U135 ( .A1(n_hpc2_0_n230), .A2(n_hpc2_0_n231), .ZN(
        n_hpc2_0_N61) );
  NOR2_X1 u_hpc2_0_U134 ( .A1(n_hpc2_0_n240), .A2(n_hpc2_0_n229), .ZN(
        n_hpc2_0_N62) );
  NOR2_X1 u_hpc2_0_U133 ( .A1(n_hpc2_0_n227), .A2(n_hpc2_0_n228), .ZN(
        n_hpc2_0_N63) );
  NOR2_X1 u_hpc2_0_U132 ( .A1(n_hpc2_0_n225), .A2(n_hpc2_0_n226), .ZN(
        n_hpc2_0_N64) );
  NOR2_X1 u_hpc2_0_U131 ( .A1(n_hpc2_0_n223), .A2(n_hpc2_0_n224), .ZN(
        n_hpc2_0_N65) );
  NOR2_X1 u_hpc2_0_U130 ( .A1(n_hpc2_0_n221), .A2(n_hpc2_0_n222), .ZN(
        n_hpc2_0_N66) );
  NOR2_X1 u_hpc2_0_U129 ( .A1(n_hpc2_0_n219), .A2(n_hpc2_0_n220), .ZN(
        n_hpc2_0_N67) );
  NOR2_X1 u_hpc2_0_U128 ( .A1(n_hpc2_0_n238), .A2(n_hpc2_0_n218), .ZN(
        n_hpc2_0_N68) );
  NOR2_X1 u_hpc2_0_U127 ( .A1(n_hpc2_0_n227), .A2(n_hpc2_0_n217), .ZN(
        n_hpc2_0_N69) );
  NOR2_X1 u_hpc2_0_U126 ( .A1(n_hpc2_0_n216), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N7) );
  NOR2_X1 u_hpc2_0_U125 ( .A1(n_hpc2_0_n214), .A2(n_hpc2_0_n215), .ZN(
        n_hpc2_0_N70) );
  NOR2_X1 u_hpc2_0_U124 ( .A1(n_hpc2_0_n212), .A2(n_hpc2_0_n213), .ZN(
        n_hpc2_0_N71) );
  NOR2_X1 u_hpc2_0_U123 ( .A1(n_hpc2_0_n210), .A2(n_hpc2_0_n211), .ZN(
        n_hpc2_0_N72) );
  NOR2_X1 u_hpc2_0_U122 ( .A1(n_hpc2_0_n208), .A2(n_hpc2_0_n209), .ZN(
        n_hpc2_0_N73) );
  NOR2_X1 u_hpc2_0_U121 ( .A1(n_hpc2_0_n236), .A2(n_hpc2_0_n207), .ZN(
        n_hpc2_0_N74) );
  NOR2_X1 u_hpc2_0_U120 ( .A1(n_hpc2_0_n225), .A2(n_hpc2_0_n206), .ZN(
        n_hpc2_0_N75) );
  NOR2_X1 u_hpc2_0_U119 ( .A1(n_hpc2_0_n214), .A2(n_hpc2_0_n205), .ZN(
        n_hpc2_0_N76) );
  NOR2_X1 u_hpc2_0_U118 ( .A1(n_hpc2_0_n203), .A2(n_hpc2_0_n204), .ZN(
        n_hpc2_0_N77) );
  NOR2_X1 u_hpc2_0_U117 ( .A1(n_hpc2_0_n201), .A2(n_hpc2_0_n202), .ZN(
        n_hpc2_0_N78) );
  NOR2_X1 u_hpc2_0_U116 ( .A1(n_hpc2_0_n199), .A2(n_hpc2_0_n200), .ZN(
        n_hpc2_0_N79) );
  NOR2_X1 u_hpc2_0_U115 ( .A1(n_hpc2_0_n198), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N8) );
  NOR2_X1 u_hpc2_0_U114 ( .A1(n_hpc2_0_n234), .A2(n_hpc2_0_n197), .ZN(
        n_hpc2_0_N80) );
  NOR2_X1 u_hpc2_0_U113 ( .A1(n_hpc2_0_n223), .A2(n_hpc2_0_n196), .ZN(
        n_hpc2_0_N81) );
  NOR2_X1 u_hpc2_0_U112 ( .A1(n_hpc2_0_n212), .A2(n_hpc2_0_n195), .ZN(
        n_hpc2_0_N82) );
  NOR2_X1 u_hpc2_0_U111 ( .A1(n_hpc2_0_n203), .A2(n_hpc2_0_n194), .ZN(
        n_hpc2_0_N83) );
  NOR2_X1 u_hpc2_0_U110 ( .A1(n_hpc2_0_n192), .A2(n_hpc2_0_n193), .ZN(
        n_hpc2_0_N84) );
  NOR2_X1 u_hpc2_0_U109 ( .A1(n_hpc2_0_n190), .A2(n_hpc2_0_n191), .ZN(
        n_hpc2_0_N85) );
  NOR2_X1 u_hpc2_0_U108 ( .A1(n_hpc2_0_n232), .A2(n_hpc2_0_n189), .ZN(
        n_hpc2_0_N86) );
  NOR2_X1 u_hpc2_0_U107 ( .A1(n_hpc2_0_n221), .A2(n_hpc2_0_n188), .ZN(
        n_hpc2_0_N87) );
  NOR2_X1 u_hpc2_0_U106 ( .A1(n_hpc2_0_n210), .A2(n_hpc2_0_n187), .ZN(
        n_hpc2_0_N88) );
  NOR2_X1 u_hpc2_0_U105 ( .A1(n_hpc2_0_n201), .A2(n_hpc2_0_n186), .ZN(
        n_hpc2_0_N89) );
  NOR2_X1 u_hpc2_0_U104 ( .A1(n_hpc2_0_n185), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N9) );
  NOR2_X1 u_hpc2_0_U103 ( .A1(n_hpc2_0_n192), .A2(n_hpc2_0_n184), .ZN(
        n_hpc2_0_N90) );
  NOR2_X1 u_hpc2_0_U102 ( .A1(n_hpc2_0_n182), .A2(n_hpc2_0_n183), .ZN(
        n_hpc2_0_N91) );
  NOR2_X1 u_hpc2_0_U101 ( .A1(n_hpc2_0_n230), .A2(n_hpc2_0_n181), .ZN(
        n_hpc2_0_N92) );
  NOR2_X1 u_hpc2_0_U100 ( .A1(n_hpc2_0_n219), .A2(n_hpc2_0_n180), .ZN(
        n_hpc2_0_N93) );
  NOR2_X1 u_hpc2_0_U99 ( .A1(n_hpc2_0_n208), .A2(n_hpc2_0_n179), .ZN(
        n_hpc2_0_N94) );
  NOR2_X1 u_hpc2_0_U98 ( .A1(n_hpc2_0_n199), .A2(n_hpc2_0_n178), .ZN(
        n_hpc2_0_N95) );
  NOR2_X1 u_hpc2_0_U97 ( .A1(n_hpc2_0_n190), .A2(n_hpc2_0_n177), .ZN(
        n_hpc2_0_N96) );
  NOR2_X1 u_hpc2_0_U96 ( .A1(n_hpc2_0_n182), .A2(n_hpc2_0_n176), .ZN(
        n_hpc2_0_N97) );
  XOR2_X1 u_hpc2_0_U95 ( .A(io_i1_s1), .B(p_rand_0), .Z(n_hpc2_0_N98) );
  XOR2_X1 u_hpc2_0_U94 ( .A(io_i1_s2), .B(p_rand_1), .Z(n_hpc2_0_N99) );
  INV_X1 u_hpc2_0_U93 ( .A(io_i0_s0), .ZN(n_hpc2_0_n1) );
  INV_X1 u_hpc2_0_U92 ( .A(io_i0_s1), .ZN(n_hpc2_0_n2) );
  INV_X1 u_hpc2_0_U91 ( .A(io_i0_s2), .ZN(n_hpc2_0_n3) );
  INV_X1 u_hpc2_0_U90 ( .A(io_i0_s3), .ZN(n_hpc2_0_n4) );
  INV_X1 u_hpc2_0_U89 ( .A(io_i0_s4), .ZN(n_hpc2_0_n5) );
  INV_X1 u_hpc2_0_U88 ( .A(io_i0_s5), .ZN(n_hpc2_0_n6) );
  INV_X1 u_hpc2_0_U87 ( .A(io_i0_s6), .ZN(n_hpc2_0_n7) );
  XOR2_X1 u_hpc2_0_U86 ( .A(n_hpc2_0__hpc_av03), .B(n_hpc2_0_n166), .Z(
        n_hpc2_0_n90) );
  XOR2_X1 u_hpc2_0_U85 ( .A(n_hpc2_0_n164), .B(n_hpc2_0_n165), .Z(n_hpc2_0_n91) );
  XOR2_X1 u_hpc2_0_U84 ( .A(n_hpc2_0_n90), .B(n_hpc2_0_n91), .Z(n_hpc2_0_n87)
         );
  XOR2_X1 u_hpc2_0_U83 ( .A(n_hpc2_0_n173), .B(n_hpc2_0_n174), .Z(n_hpc2_0_n89) );
  XOR2_X1 u_hpc2_0_U82 ( .A(n_hpc2_0_n175), .B(n_hpc2_0_n89), .Z(n_hpc2_0_n88)
         );
  XOR2_X1 u_hpc2_0_U81 ( .A(n_hpc2_0_n87), .B(n_hpc2_0_n88), .Z(n_hpc2_0_n85)
         );
  XOR2_X1 u_hpc2_0_U80 ( .A(n_hpc2_0_n171), .B(n_hpc2_0_n172), .Z(n_hpc2_0_n86) );
  XOR2_X1 u_hpc2_0_U79 ( .A(n_hpc2_0_n85), .B(n_hpc2_0_n86), .Z(n_hpc2_0_n81)
         );
  XOR2_X1 u_hpc2_0_U78 ( .A(n_hpc2_0_n167), .B(n_hpc2_0_n168), .Z(n_hpc2_0_n83) );
  XOR2_X1 u_hpc2_0_U77 ( .A(n_hpc2_0_n169), .B(n_hpc2_0_n170), .Z(n_hpc2_0_n84) );
  XOR2_X1 u_hpc2_0_U76 ( .A(n_hpc2_0_n83), .B(n_hpc2_0_n84), .Z(n_hpc2_0_n82)
         );
  XOR2_X1 u_hpc2_0_U75 ( .A(n_hpc2_0_n81), .B(n_hpc2_0_n82), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U74 ( .A(n_hpc2_0__hpc_av13), .B(n_hpc2_0_n154), .Z(
        n_hpc2_0_n79) );
  XOR2_X1 u_hpc2_0_U73 ( .A(n_hpc2_0_n152), .B(n_hpc2_0_n153), .Z(n_hpc2_0_n80) );
  XOR2_X1 u_hpc2_0_U72 ( .A(n_hpc2_0_n79), .B(n_hpc2_0_n80), .Z(n_hpc2_0_n76)
         );
  XOR2_X1 u_hpc2_0_U71 ( .A(n_hpc2_0_n161), .B(n_hpc2_0_n162), .Z(n_hpc2_0_n78) );
  XOR2_X1 u_hpc2_0_U70 ( .A(n_hpc2_0_n163), .B(n_hpc2_0_n78), .Z(n_hpc2_0_n77)
         );
  XOR2_X1 u_hpc2_0_U69 ( .A(n_hpc2_0_n76), .B(n_hpc2_0_n77), .Z(n_hpc2_0_n74)
         );
  XOR2_X1 u_hpc2_0_U68 ( .A(n_hpc2_0_n159), .B(n_hpc2_0_n160), .Z(n_hpc2_0_n75) );
  XOR2_X1 u_hpc2_0_U67 ( .A(n_hpc2_0_n74), .B(n_hpc2_0_n75), .Z(n_hpc2_0_n70)
         );
  XOR2_X1 u_hpc2_0_U66 ( .A(n_hpc2_0_n155), .B(n_hpc2_0_n156), .Z(n_hpc2_0_n72) );
  XOR2_X1 u_hpc2_0_U65 ( .A(n_hpc2_0_n157), .B(n_hpc2_0_n158), .Z(n_hpc2_0_n73) );
  XOR2_X1 u_hpc2_0_U64 ( .A(n_hpc2_0_n72), .B(n_hpc2_0_n73), .Z(n_hpc2_0_n71)
         );
  XOR2_X1 u_hpc2_0_U63 ( .A(n_hpc2_0_n70), .B(n_hpc2_0_n71), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U62 ( .A(n_hpc2_0__hpc_av23), .B(n_hpc2_0_n142), .Z(
        n_hpc2_0_n68) );
  XOR2_X1 u_hpc2_0_U61 ( .A(n_hpc2_0_n140), .B(n_hpc2_0_n141), .Z(n_hpc2_0_n69) );
  XOR2_X1 u_hpc2_0_U60 ( .A(n_hpc2_0_n68), .B(n_hpc2_0_n69), .Z(n_hpc2_0_n65)
         );
  XOR2_X1 u_hpc2_0_U59 ( .A(n_hpc2_0_n149), .B(n_hpc2_0_n150), .Z(n_hpc2_0_n67) );
  XOR2_X1 u_hpc2_0_U58 ( .A(n_hpc2_0_n151), .B(n_hpc2_0_n67), .Z(n_hpc2_0_n66)
         );
  XOR2_X1 u_hpc2_0_U57 ( .A(n_hpc2_0_n65), .B(n_hpc2_0_n66), .Z(n_hpc2_0_n63)
         );
  XOR2_X1 u_hpc2_0_U56 ( .A(n_hpc2_0_n147), .B(n_hpc2_0_n148), .Z(n_hpc2_0_n64) );
  XOR2_X1 u_hpc2_0_U55 ( .A(n_hpc2_0_n63), .B(n_hpc2_0_n64), .Z(n_hpc2_0_n59)
         );
  XOR2_X1 u_hpc2_0_U54 ( .A(n_hpc2_0_n143), .B(n_hpc2_0_n144), .Z(n_hpc2_0_n61) );
  XOR2_X1 u_hpc2_0_U53 ( .A(n_hpc2_0_n145), .B(n_hpc2_0_n146), .Z(n_hpc2_0_n62) );
  XOR2_X1 u_hpc2_0_U52 ( .A(n_hpc2_0_n61), .B(n_hpc2_0_n62), .Z(n_hpc2_0_n60)
         );
  XOR2_X1 u_hpc2_0_U51 ( .A(n_hpc2_0_n59), .B(n_hpc2_0_n60), .Z(io_o0_s2) );
  XOR2_X1 u_hpc2_0_U50 ( .A(n_hpc2_0__hpc_av32), .B(n_hpc2_0_n130), .Z(
        n_hpc2_0_n57) );
  XOR2_X1 u_hpc2_0_U49 ( .A(n_hpc2_0_n128), .B(n_hpc2_0_n129), .Z(n_hpc2_0_n58) );
  XOR2_X1 u_hpc2_0_U48 ( .A(n_hpc2_0_n57), .B(n_hpc2_0_n58), .Z(n_hpc2_0_n54)
         );
  XOR2_X1 u_hpc2_0_U47 ( .A(n_hpc2_0_n137), .B(n_hpc2_0_n138), .Z(n_hpc2_0_n56) );
  XOR2_X1 u_hpc2_0_U46 ( .A(n_hpc2_0_n139), .B(n_hpc2_0_n56), .Z(n_hpc2_0_n55)
         );
  XOR2_X1 u_hpc2_0_U45 ( .A(n_hpc2_0_n54), .B(n_hpc2_0_n55), .Z(n_hpc2_0_n52)
         );
  XOR2_X1 u_hpc2_0_U44 ( .A(n_hpc2_0_n135), .B(n_hpc2_0_n136), .Z(n_hpc2_0_n53) );
  XOR2_X1 u_hpc2_0_U43 ( .A(n_hpc2_0_n52), .B(n_hpc2_0_n53), .Z(n_hpc2_0_n48)
         );
  XOR2_X1 u_hpc2_0_U42 ( .A(n_hpc2_0_n131), .B(n_hpc2_0_n132), .Z(n_hpc2_0_n50) );
  XOR2_X1 u_hpc2_0_U41 ( .A(n_hpc2_0_n133), .B(n_hpc2_0_n134), .Z(n_hpc2_0_n51) );
  XOR2_X1 u_hpc2_0_U40 ( .A(n_hpc2_0_n50), .B(n_hpc2_0_n51), .Z(n_hpc2_0_n49)
         );
  XOR2_X1 u_hpc2_0_U39 ( .A(n_hpc2_0_n48), .B(n_hpc2_0_n49), .Z(io_o0_s3) );
  XOR2_X1 u_hpc2_0_U38 ( .A(n_hpc2_0__hpc_av42), .B(n_hpc2_0_n118), .Z(
        n_hpc2_0_n46) );
  XOR2_X1 u_hpc2_0_U37 ( .A(n_hpc2_0_n116), .B(n_hpc2_0_n117), .Z(n_hpc2_0_n47) );
  XOR2_X1 u_hpc2_0_U36 ( .A(n_hpc2_0_n46), .B(n_hpc2_0_n47), .Z(n_hpc2_0_n43)
         );
  XOR2_X1 u_hpc2_0_U35 ( .A(n_hpc2_0_n125), .B(n_hpc2_0_n126), .Z(n_hpc2_0_n45) );
  XOR2_X1 u_hpc2_0_U34 ( .A(n_hpc2_0_n127), .B(n_hpc2_0_n45), .Z(n_hpc2_0_n44)
         );
  XOR2_X1 u_hpc2_0_U33 ( .A(n_hpc2_0_n43), .B(n_hpc2_0_n44), .Z(n_hpc2_0_n41)
         );
  XOR2_X1 u_hpc2_0_U32 ( .A(n_hpc2_0_n123), .B(n_hpc2_0_n124), .Z(n_hpc2_0_n42) );
  XOR2_X1 u_hpc2_0_U31 ( .A(n_hpc2_0_n41), .B(n_hpc2_0_n42), .Z(n_hpc2_0_n37)
         );
  XOR2_X1 u_hpc2_0_U30 ( .A(n_hpc2_0_n119), .B(n_hpc2_0_n120), .Z(n_hpc2_0_n39) );
  XOR2_X1 u_hpc2_0_U29 ( .A(n_hpc2_0_n121), .B(n_hpc2_0_n122), .Z(n_hpc2_0_n40) );
  XOR2_X1 u_hpc2_0_U28 ( .A(n_hpc2_0_n39), .B(n_hpc2_0_n40), .Z(n_hpc2_0_n38)
         );
  XOR2_X1 u_hpc2_0_U27 ( .A(n_hpc2_0_n37), .B(n_hpc2_0_n38), .Z(io_o0_s4) );
  XOR2_X1 u_hpc2_0_U26 ( .A(n_hpc2_0__hpc_av52), .B(n_hpc2_0_n106), .Z(
        n_hpc2_0_n35) );
  XOR2_X1 u_hpc2_0_U25 ( .A(n_hpc2_0_n104), .B(n_hpc2_0_n105), .Z(n_hpc2_0_n36) );
  XOR2_X1 u_hpc2_0_U24 ( .A(n_hpc2_0_n35), .B(n_hpc2_0_n36), .Z(n_hpc2_0_n32)
         );
  XOR2_X1 u_hpc2_0_U23 ( .A(n_hpc2_0_n113), .B(n_hpc2_0_n114), .Z(n_hpc2_0_n34) );
  XOR2_X1 u_hpc2_0_U22 ( .A(n_hpc2_0_n115), .B(n_hpc2_0_n34), .Z(n_hpc2_0_n33)
         );
  XOR2_X1 u_hpc2_0_U21 ( .A(n_hpc2_0_n32), .B(n_hpc2_0_n33), .Z(n_hpc2_0_n30)
         );
  XOR2_X1 u_hpc2_0_U20 ( .A(n_hpc2_0_n111), .B(n_hpc2_0_n112), .Z(n_hpc2_0_n31) );
  XOR2_X1 u_hpc2_0_U19 ( .A(n_hpc2_0_n30), .B(n_hpc2_0_n31), .Z(n_hpc2_0_n26)
         );
  XOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0_n107), .B(n_hpc2_0_n108), .Z(n_hpc2_0_n28) );
  XOR2_X1 u_hpc2_0_U17 ( .A(n_hpc2_0_n109), .B(n_hpc2_0_n110), .Z(n_hpc2_0_n29) );
  XOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_n28), .B(n_hpc2_0_n29), .Z(n_hpc2_0_n27)
         );
  XOR2_X1 u_hpc2_0_U15 ( .A(n_hpc2_0_n26), .B(n_hpc2_0_n27), .Z(io_o0_s5) );
  XOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0__hpc_av62), .B(n_hpc2_0_n94), .Z(
        n_hpc2_0_n24) );
  XOR2_X1 u_hpc2_0_U13 ( .A(n_hpc2_0_n92), .B(n_hpc2_0_n93), .Z(n_hpc2_0_n25)
         );
  XOR2_X1 u_hpc2_0_U12 ( .A(n_hpc2_0_n24), .B(n_hpc2_0_n25), .Z(n_hpc2_0_n21)
         );
  XOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_n101), .B(n_hpc2_0_n102), .Z(n_hpc2_0_n23) );
  XOR2_X1 u_hpc2_0_U10 ( .A(n_hpc2_0_n103), .B(n_hpc2_0_n23), .Z(n_hpc2_0_n22)
         );
  XOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_n21), .B(n_hpc2_0_n22), .Z(n_hpc2_0_n19)
         );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0_n99), .B(n_hpc2_0_n100), .Z(n_hpc2_0_n20)
         );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0_n19), .B(n_hpc2_0_n20), .Z(n_hpc2_0_n15)
         );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0_n95), .B(n_hpc2_0_n96), .Z(n_hpc2_0_n17)
         );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0_n97), .B(n_hpc2_0_n98), .Z(n_hpc2_0_n18)
         );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0_n17), .B(n_hpc2_0_n18), .Z(n_hpc2_0_n16)
         );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n15), .B(n_hpc2_0_n16), .Z(io_o0_s6) );
  DFF_X1 u_hpc2_0__hpc_av65_reg ( .D(n_hpc2_0_N55), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n97) );
  DFF_X1 u_hpc2_0__hpc_v65_reg ( .D(n_hpc2_0_N139), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n242) );
  DFF_X1 u_hpc2_0__hpc_av64_reg ( .D(n_hpc2_0_N54), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n96) );
  DFF_X1 u_hpc2_0__hpc_v64_reg ( .D(n_hpc2_0_N138), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n243) );
  DFF_X1 u_hpc2_0__hpc_av63_reg ( .D(n_hpc2_0_N53), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n95) );
  DFF_X1 u_hpc2_0__hpc_v63_reg ( .D(n_hpc2_0_N137), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n244) );
  DFF_X1 u_hpc2_0__hpc_av62_reg ( .D(n_hpc2_0_N52), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av62), .QN() );
  DFF_X1 u_hpc2_0__hpc_v62_reg ( .D(n_hpc2_0_N136), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n245) );
  DFF_X1 u_hpc2_0__hpc_av61_reg ( .D(n_hpc2_0_N51), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n93) );
  DFF_X1 u_hpc2_0__hpc_v61_reg ( .D(n_hpc2_0_N135), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n246) );
  DFF_X1 u_hpc2_0__hpc_av60_reg ( .D(n_hpc2_0_N50), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n92) );
  DFF_X1 u_hpc2_0__hpc_v60_reg ( .D(n_hpc2_0_N134), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n247) );
  DFF_X1 u_hpc2_0__hpc_av56_reg ( .D(n_hpc2_0_N49), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n109) );
  DFF_X1 u_hpc2_0__hpc_v56_reg ( .D(n_hpc2_0_N133), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n248) );
  DFF_X1 u_hpc2_0__hpc_av54_reg ( .D(n_hpc2_0_N48), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n108) );
  DFF_X1 u_hpc2_0__hpc_v54_reg ( .D(n_hpc2_0_N132), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n249) );
  DFF_X1 u_hpc2_0__hpc_av53_reg ( .D(n_hpc2_0_N47), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n107) );
  DFF_X1 u_hpc2_0__hpc_v53_reg ( .D(n_hpc2_0_N131), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n250) );
  DFF_X1 u_hpc2_0__hpc_av52_reg ( .D(n_hpc2_0_N46), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av52), .QN() );
  DFF_X1 u_hpc2_0__hpc_v52_reg ( .D(n_hpc2_0_N130), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n251) );
  DFF_X1 u_hpc2_0__hpc_av51_reg ( .D(n_hpc2_0_N45), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n105) );
  DFF_X1 u_hpc2_0__hpc_v51_reg ( .D(n_hpc2_0_N129), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n252) );
  DFF_X1 u_hpc2_0__hpc_av50_reg ( .D(n_hpc2_0_N44), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n104) );
  DFF_X1 u_hpc2_0__hpc_v50_reg ( .D(n_hpc2_0_N128), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n253) );
  DFF_X1 u_hpc2_0__hpc_av46_reg ( .D(n_hpc2_0_N43), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n121) );
  DFF_X1 u_hpc2_0__hpc_v46_reg ( .D(n_hpc2_0_N127), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n254) );
  DFF_X1 u_hpc2_0__hpc_av45_reg ( .D(n_hpc2_0_N42), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n120) );
  DFF_X1 u_hpc2_0__hpc_v45_reg ( .D(n_hpc2_0_N126), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n255) );
  DFF_X1 u_hpc2_0__hpc_av43_reg ( .D(n_hpc2_0_N41), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n119) );
  DFF_X1 u_hpc2_0__hpc_v43_reg ( .D(n_hpc2_0_N125), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n256) );
  DFF_X1 u_hpc2_0__hpc_av42_reg ( .D(n_hpc2_0_N40), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av42), .QN() );
  DFF_X1 u_hpc2_0__hpc_v42_reg ( .D(n_hpc2_0_N124), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n257) );
  DFF_X1 u_hpc2_0__hpc_av41_reg ( .D(n_hpc2_0_N39), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n117) );
  DFF_X1 u_hpc2_0__hpc_v41_reg ( .D(n_hpc2_0_N123), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n258) );
  DFF_X1 u_hpc2_0__hpc_av40_reg ( .D(n_hpc2_0_N38), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n116) );
  DFF_X1 u_hpc2_0__hpc_v40_reg ( .D(n_hpc2_0_N122), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n259) );
  DFF_X1 u_hpc2_0__hpc_av36_reg ( .D(n_hpc2_0_N37), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n133) );
  DFF_X1 u_hpc2_0__hpc_v36_reg ( .D(n_hpc2_0_N121), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n260) );
  DFF_X1 u_hpc2_0__hpc_av35_reg ( .D(n_hpc2_0_N36), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n132) );
  DFF_X1 u_hpc2_0__hpc_v35_reg ( .D(n_hpc2_0_N120), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n261) );
  DFF_X1 u_hpc2_0__hpc_av34_reg ( .D(n_hpc2_0_N35), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n131) );
  DFF_X1 u_hpc2_0__hpc_v34_reg ( .D(n_hpc2_0_N119), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n262) );
  DFF_X1 u_hpc2_0__hpc_av32_reg ( .D(n_hpc2_0_N34), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av32), .QN() );
  DFF_X1 u_hpc2_0__hpc_v32_reg ( .D(n_hpc2_0_N118), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n263) );
  DFF_X1 u_hpc2_0__hpc_av31_reg ( .D(n_hpc2_0_N33), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n129) );
  DFF_X1 u_hpc2_0__hpc_v31_reg ( .D(n_hpc2_0_N117), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n264) );
  DFF_X1 u_hpc2_0__hpc_av30_reg ( .D(n_hpc2_0_N32), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n128) );
  DFF_X1 u_hpc2_0__hpc_v30_reg ( .D(n_hpc2_0_N116), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n265) );
  DFF_X1 u_hpc2_0__hpc_av26_reg ( .D(n_hpc2_0_N31), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n145) );
  DFF_X1 u_hpc2_0__hpc_v26_reg ( .D(n_hpc2_0_N115), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n266) );
  DFF_X1 u_hpc2_0__hpc_av25_reg ( .D(n_hpc2_0_N30), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n144) );
  DFF_X1 u_hpc2_0__hpc_v25_reg ( .D(n_hpc2_0_N114), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n267) );
  DFF_X1 u_hpc2_0__hpc_av24_reg ( .D(n_hpc2_0_N29), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n143) );
  DFF_X1 u_hpc2_0__hpc_v24_reg ( .D(n_hpc2_0_N113), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n268) );
  DFF_X1 u_hpc2_0__hpc_av23_reg ( .D(n_hpc2_0_N28), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av23), .QN() );
  DFF_X1 u_hpc2_0__hpc_v23_reg ( .D(n_hpc2_0_N112), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n269) );
  DFF_X1 u_hpc2_0__hpc_av21_reg ( .D(n_hpc2_0_N27), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n141) );
  DFF_X1 u_hpc2_0__hpc_v21_reg ( .D(n_hpc2_0_N111), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n270) );
  DFF_X1 u_hpc2_0__hpc_av20_reg ( .D(n_hpc2_0_N26), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n140) );
  DFF_X1 u_hpc2_0__hpc_v20_reg ( .D(n_hpc2_0_N110), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n271) );
  DFF_X1 u_hpc2_0__hpc_av16_reg ( .D(n_hpc2_0_N25), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n157) );
  DFF_X1 u_hpc2_0__hpc_v16_reg ( .D(n_hpc2_0_N109), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n272) );
  DFF_X1 u_hpc2_0__hpc_av15_reg ( .D(n_hpc2_0_N24), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n156) );
  DFF_X1 u_hpc2_0__hpc_v15_reg ( .D(n_hpc2_0_N108), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n273) );
  DFF_X1 u_hpc2_0__hpc_av14_reg ( .D(n_hpc2_0_N23), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n155) );
  DFF_X1 u_hpc2_0__hpc_v14_reg ( .D(n_hpc2_0_N107), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n274) );
  DFF_X1 u_hpc2_0__hpc_av13_reg ( .D(n_hpc2_0_N22), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av13), .QN() );
  DFF_X1 u_hpc2_0__hpc_v13_reg ( .D(n_hpc2_0_N106), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n275) );
  DFF_X1 u_hpc2_0__hpc_av12_reg ( .D(n_hpc2_0_N21), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n153) );
  DFF_X1 u_hpc2_0__hpc_v12_reg ( .D(n_hpc2_0_N105), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n276) );
  DFF_X1 u_hpc2_0__hpc_av10_reg ( .D(n_hpc2_0_N20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n152) );
  DFF_X1 u_hpc2_0__hpc_v10_reg ( .D(n_hpc2_0_N104), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n277) );
  DFF_X1 u_hpc2_0__hpc_av06_reg ( .D(n_hpc2_0_N19), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n169) );
  DFF_X1 u_hpc2_0__hpc_v06_reg ( .D(n_hpc2_0_N103), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n278) );
  DFF_X1 u_hpc2_0__hpc_av05_reg ( .D(n_hpc2_0_N18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n168) );
  DFF_X1 u_hpc2_0__hpc_v05_reg ( .D(n_hpc2_0_N102), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n279) );
  DFF_X1 u_hpc2_0__hpc_av04_reg ( .D(n_hpc2_0_N17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n167) );
  DFF_X1 u_hpc2_0__hpc_v04_reg ( .D(n_hpc2_0_N101), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n280) );
  DFF_X1 u_hpc2_0__hpc_av03_reg ( .D(n_hpc2_0_N16), .CK(clock_0), .Q(
        n_hpc2_0__hpc_av03), .QN() );
  DFF_X1 u_hpc2_0__hpc_v03_reg ( .D(n_hpc2_0_N100), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n281) );
  DFF_X1 u_hpc2_0__hpc_av02_reg ( .D(n_hpc2_0_N15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n165) );
  DFF_X1 u_hpc2_0__hpc_v02_reg ( .D(n_hpc2_0_N99), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n282) );
  DFF_X1 u_hpc2_0__hpc_av01_reg ( .D(n_hpc2_0_N14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n164) );
  DFF_X1 u_hpc2_0__hpc_v01_reg ( .D(n_hpc2_0_N98), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n283) );
  DFF_X1 u_hpc2_0__hpc_u65_reg ( .D(n_hpc2_0_N97), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n100) );
  DFF_X1 u_hpc2_0__hpc_u64_reg ( .D(n_hpc2_0_N96), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n99) );
  DFF_X1 u_hpc2_0__hpc_u63_reg ( .D(n_hpc2_0_N95), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n98) );
  DFF_X1 u_hpc2_0__hpc_u62_reg ( .D(n_hpc2_0_N94), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n103) );
  DFF_X1 u_hpc2_0__hpc_u61_reg ( .D(n_hpc2_0_N93), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n102) );
  DFF_X1 u_hpc2_0__hpc_u60_reg ( .D(n_hpc2_0_N92), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n101) );
  DFF_X1 u_hpc2_0__hpc_u56_reg ( .D(n_hpc2_0_N91), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n112) );
  DFF_X1 u_hpc2_0__hpc_u54_reg ( .D(n_hpc2_0_N90), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n111) );
  DFF_X1 u_hpc2_0__hpc_u53_reg ( .D(n_hpc2_0_N89), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n110) );
  DFF_X1 u_hpc2_0__hpc_u52_reg ( .D(n_hpc2_0_N88), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n115) );
  DFF_X1 u_hpc2_0__hpc_u51_reg ( .D(n_hpc2_0_N87), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n114) );
  DFF_X1 u_hpc2_0__hpc_u50_reg ( .D(n_hpc2_0_N86), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n113) );
  DFF_X1 u_hpc2_0__hpc_u46_reg ( .D(n_hpc2_0_N85), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n124) );
  DFF_X1 u_hpc2_0__hpc_u45_reg ( .D(n_hpc2_0_N84), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n123) );
  DFF_X1 u_hpc2_0__hpc_u43_reg ( .D(n_hpc2_0_N83), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n122) );
  DFF_X1 u_hpc2_0__hpc_u42_reg ( .D(n_hpc2_0_N82), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n127) );
  DFF_X1 u_hpc2_0__hpc_u41_reg ( .D(n_hpc2_0_N81), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n126) );
  DFF_X1 u_hpc2_0__hpc_u40_reg ( .D(n_hpc2_0_N80), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n125) );
  DFF_X1 u_hpc2_0__hpc_u36_reg ( .D(n_hpc2_0_N79), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n136) );
  DFF_X1 u_hpc2_0__hpc_u35_reg ( .D(n_hpc2_0_N78), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n135) );
  DFF_X1 u_hpc2_0__hpc_u34_reg ( .D(n_hpc2_0_N77), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n134) );
  DFF_X1 u_hpc2_0__hpc_u32_reg ( .D(n_hpc2_0_N76), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n139) );
  DFF_X1 u_hpc2_0__hpc_u31_reg ( .D(n_hpc2_0_N75), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n138) );
  DFF_X1 u_hpc2_0__hpc_u30_reg ( .D(n_hpc2_0_N74), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n137) );
  DFF_X1 u_hpc2_0__hpc_u26_reg ( .D(n_hpc2_0_N73), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n148) );
  DFF_X1 u_hpc2_0__hpc_u25_reg ( .D(n_hpc2_0_N72), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n147) );
  DFF_X1 u_hpc2_0__hpc_u24_reg ( .D(n_hpc2_0_N71), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n146) );
  DFF_X1 u_hpc2_0__hpc_u23_reg ( .D(n_hpc2_0_N70), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n151) );
  DFF_X1 u_hpc2_0__hpc_u21_reg ( .D(n_hpc2_0_N69), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n150) );
  DFF_X1 u_hpc2_0__hpc_u20_reg ( .D(n_hpc2_0_N68), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n149) );
  DFF_X1 u_hpc2_0__hpc_u16_reg ( .D(n_hpc2_0_N67), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n160) );
  DFF_X1 u_hpc2_0__hpc_u15_reg ( .D(n_hpc2_0_N66), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n159) );
  DFF_X1 u_hpc2_0__hpc_u14_reg ( .D(n_hpc2_0_N65), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n158) );
  DFF_X1 u_hpc2_0__hpc_u13_reg ( .D(n_hpc2_0_N64), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n163) );
  DFF_X1 u_hpc2_0__hpc_u12_reg ( .D(n_hpc2_0_N63), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n162) );
  DFF_X1 u_hpc2_0__hpc_u10_reg ( .D(n_hpc2_0_N62), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n161) );
  DFF_X1 u_hpc2_0__hpc_u06_reg ( .D(n_hpc2_0_N61), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n172) );
  DFF_X1 u_hpc2_0__hpc_u05_reg ( .D(n_hpc2_0_N60), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n171) );
  DFF_X1 u_hpc2_0__hpc_u04_reg ( .D(n_hpc2_0_N59), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n170) );
  DFF_X1 u_hpc2_0__hpc_u03_reg ( .D(n_hpc2_0_N58), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n175) );
  DFF_X1 u_hpc2_0__hpc_u02_reg ( .D(n_hpc2_0_N57), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n174) );
  DFF_X1 u_hpc2_0__hpc_u01_reg ( .D(n_hpc2_0_N56), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n173) );
  DFF_X1 u_hpc2_0__hpc_ab6_reg ( .D(n_hpc2_0_N13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n94) );
  DFF_X1 u_hpc2_0__hpc_b6_reg ( .D(io_i1_s6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n284) );
  DFF_X1 u_hpc2_0__hpc_ab5_reg ( .D(n_hpc2_0_N12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n106) );
  DFF_X1 u_hpc2_0__hpc_b5_reg ( .D(io_i1_s5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n285) );
  DFF_X1 u_hpc2_0__hpc_ab4_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n118) );
  DFF_X1 u_hpc2_0__hpc_b4_reg ( .D(io_i1_s4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n286) );
  DFF_X1 u_hpc2_0__hpc_ab3_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n130) );
  DFF_X1 u_hpc2_0__hpc_b3_reg ( .D(io_i1_s3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n287) );
  DFF_X1 u_hpc2_0__hpc_ab2_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n142) );
  DFF_X1 u_hpc2_0__hpc_b2_reg ( .D(io_i1_s2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n185) );
  DFF_X1 u_hpc2_0__hpc_ab1_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n154) );
  DFF_X1 u_hpc2_0__hpc_b1_reg ( .D(io_i1_s1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n198) );
  DFF_X1 u_hpc2_0__hpc_ab0_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n166) );
  DFF_X1 u_hpc2_0__hpc_b0_reg ( .D(io_i1_s0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n216) );
  DFF_X1 u_hpc2_0_reg_pipeline_34_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n229) );
  DFF_X1 u_hpc2_0_reg_pipeline_33_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n228) );
  DFF_X1 u_hpc2_0_reg_pipeline_36_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n233) );
  DFF_X1 u_hpc2_0_reg_pipeline_32_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n226) );
  DFF_X1 u_hpc2_0_reg_pipeline_37_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n235) );
  DFF_X1 u_hpc2_0_reg_pipeline_31_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n224) );
  DFF_X1 u_hpc2_0_reg_pipeline_38_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n237) );
  DFF_X1 u_hpc2_0_reg_pipeline_30_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n222) );
  DFF_X1 u_hpc2_0_reg_pipeline_39_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n239) );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(n_hpc2_0_n7), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n180) );
  DFF_X1 u_hpc2_0_reg_pipeline_27_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n217) );
  DFF_X1 u_hpc2_0_reg_pipeline_29_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n220) );
  DFF_X1 u_hpc2_0_reg_pipeline_35_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n231) );
  DFF_X1 u_hpc2_0_reg_pipeline_28_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n218) );
  DFF_X1 u_hpc2_0_reg_pipeline_46_reg ( .D(io_i0_s5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n12) );
  DFF_X1 u_hpc2_0_reg_pipeline_47_reg ( .D(io_i0_s6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n11) );
  DFF_X1 u_hpc2_0_reg_pipeline_9_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n188) );
  DFF_X1 u_hpc2_0_reg_pipeline_5_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n183) );
  DFF_X1 u_hpc2_0__hpc_r9_reg ( .D(p_rand_9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n221) );
  DFF_X1 u_hpc2_0__hpc_r5_reg ( .D(p_rand_5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n230) );
  DFF_X1 u_hpc2_0_reg_pipeline_6_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n184) );
  DFF_X1 u_hpc2_0__hpc_r8_reg ( .D(p_rand_8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n223) );
  DFF_X1 u_hpc2_0__hpc_r4_reg ( .D(p_rand_4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n232) );
  DFF_X1 u_hpc2_0__hpc_r2_reg ( .D(p_rand_2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n236) );
  DFF_X1 u_hpc2_0_reg_pipeline_7_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n186) );
  DFF_X1 u_hpc2_0__hpc_r7_reg ( .D(p_rand_7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n225) );
  DFF_X1 u_hpc2_0__hpc_r3_reg ( .D(p_rand_3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n234) );
  DFF_X1 u_hpc2_0__hpc_r19_reg ( .D(p_rand_19), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n190) );
  DFF_X1 u_hpc2_0__hpc_r17_reg ( .D(p_rand_17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n199) );
  DFF_X1 u_hpc2_0_reg_pipeline_8_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n187) );
  DFF_X1 u_hpc2_0__hpc_r6_reg ( .D(p_rand_6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n227) );
  DFF_X1 u_hpc2_0__hpc_r20_reg ( .D(p_rand_20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n182) );
  DFF_X1 u_hpc2_0__hpc_r18_reg ( .D(p_rand_18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n192) );
  DFF_X1 u_hpc2_0__hpc_r16_reg ( .D(p_rand_16), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n201) );
  DFF_X1 u_hpc2_0__hpc_r15_reg ( .D(p_rand_15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n203) );
  DFF_X1 u_hpc2_0_reg_pipeline_26_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n215) );
  DFF_X1 u_hpc2_0_reg_pipeline_25_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n213) );
  DFF_X1 u_hpc2_0_reg_pipeline_24_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n211) );
  DFF_X1 u_hpc2_0_reg_pipeline_23_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n209) );
  DFF_X1 u_hpc2_0_reg_pipeline_22_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n207) );
  DFF_X1 u_hpc2_0_reg_pipeline_21_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n206) );
  DFF_X1 u_hpc2_0_reg_pipeline_20_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n205) );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(n_hpc2_0_n7), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n179) );
  DFF_X1 u_hpc2_0_reg_pipeline_19_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n204) );
  DFF_X1 u_hpc2_0_reg_pipeline_18_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n202) );
  DFF_X1 u_hpc2_0_reg_pipeline_17_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n200) );
  DFF_X1 u_hpc2_0_reg_pipeline_16_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n197) );
  DFF_X1 u_hpc2_0_reg_pipeline_15_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n196) );
  DFF_X1 u_hpc2_0_reg_pipeline_14_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n195) );
  DFF_X1 u_hpc2_0_reg_pipeline_13_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n194) );
  DFF_X1 u_hpc2_0_reg_pipeline_12_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n193) );
  DFF_X1 u_hpc2_0_reg_pipeline_11_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n191) );
  DFF_X1 u_hpc2_0_reg_pipeline_10_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n189) );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(n_hpc2_0_n7), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n178) );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(n_hpc2_0_n7), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n177) );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(n_hpc2_0_n7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n176) );
  DFF_X1 u_hpc2_0_reg_pipeline_45_reg ( .D(io_i0_s4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n13) );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(n_hpc2_0_n7), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n181) );
  DFF_X1 u_hpc2_0_reg_pipeline_40_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n241) );
  DFF_X1 u_hpc2_0_reg_pipeline_41_reg ( .D(io_i0_s0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n10) );
  DFF_X1 u_hpc2_0_reg_pipeline_42_reg ( .D(io_i0_s1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n9) );
  DFF_X1 u_hpc2_0_reg_pipeline_43_reg ( .D(io_i0_s2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n8) );
  DFF_X1 u_hpc2_0_reg_pipeline_44_reg ( .D(io_i0_s3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n14) );
  DFF_X1 u_hpc2_0__hpc_r14_reg ( .D(p_rand_14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n208) );
  DFF_X1 u_hpc2_0__hpc_r13_reg ( .D(p_rand_13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n210) );
  DFF_X1 u_hpc2_0__hpc_r12_reg ( .D(p_rand_12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n212) );
  DFF_X1 u_hpc2_0__hpc_r11_reg ( .D(p_rand_11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n214) );
  DFF_X1 u_hpc2_0__hpc_r10_reg ( .D(p_rand_10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n219) );
  DFF_X1 u_hpc2_0__hpc_r1_reg ( .D(p_rand_1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n238) );
  DFF_X1 u_hpc2_0__hpc_r0_reg ( .D(p_rand_0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n240) );
endmodule

