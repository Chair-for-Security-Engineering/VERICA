
module ISW_SifaTest ( port_a_in, port_b_in, port_rand, port_det_out, clk, 
        reset );
  input [1:0] port_a_in;
  input [1:0] port_b_in;
  input [0:0] port_rand;
  output [1:0] port_det_out;
  input clk, reset;
  wire   isw_0__zz_port_a_3, isw_0__zz_port_b_1, isw_0__zz_port_a_1,
         isw_0_xor_12_port_z, isw_0_z_0, isw_0__zz_port_a_4,
         isw_0_and_12_port_z, isw_0_xor_11_port_z, isw_0__zz_port_b_2,
         isw_0__zz_port_a_2, isw_0_and_11_port_z, isw_0_xor_10_port_z,
         isw_0__zz_port_b, isw_0__zz_port_a, isw_0_and_10_port_z,
         isw_0_xor_9_port_z, isw_0_and_9_port_z, isw_1__zz_port_a_3,
         isw_1__zz_port_b_1, isw_1__zz_port_a_1, isw_1_xor_12_port_z,
         isw_1_z_0, isw_1__zz_port_a_4, isw_1_and_12_port_z,
         isw_1_xor_11_port_z, isw_1__zz_port_b_2, isw_1__zz_port_a_2,
         isw_1_and_11_port_z, isw_1_xor_10_port_z, isw_1__zz_port_b,
         isw_1__zz_port_a, isw_1_and_10_port_z, isw_1_xor_9_port_z,
         isw_1_and_9_port_z;
  wire   [1:0] n_zz_unequal_0;
  wire   [1:0] n_zz_unequal_0_1;
  wire port_a_in0, port_a_in1;

  BUF_X1 B00 ( .A(port_a_in[0]), .Z(port_a_in0) );
  BUF_X1 B01 ( .A(port_a_in[1]), .Z(port_a_in1) );

  XNOR2_X1 U3 ( .A(n_zz_unequal_0_1[0]), .B(n_zz_unequal_0[0]), .ZN(
        port_det_out[0]) );
  XNOR2_X1 U4 ( .A(n_zz_unequal_0_1[1]), .B(n_zz_unequal_0[1]), .ZN(
        port_det_out[1]) );
  DFF_X1 isw_0_result_1_reg ( .D(isw_0_xor_12_port_z), .CK(clk), .Q(
        n_zz_unequal_0[1]), .QN() );
  DFF_X1 isw_0__zz_port_a_4_reg ( .D(isw_0__zz_port_a_3), .CK(clk), .Q(
        isw_0__zz_port_a_4), .QN() );
  DFF_X1 isw_0_result_0_reg ( .D(isw_0_xor_11_port_z), .CK(clk), .Q(
        n_zz_unequal_0[0]), .QN() );
  DFF_X1 isw_0__zz_port_b_2_reg ( .D(isw_0__zz_port_b_1), .CK(clk), .Q(
        isw_0__zz_port_b_2), .QN() );
  DFF_X1 isw_0__zz_port_a_2_reg ( .D(isw_0__zz_port_a_1), .CK(clk), .Q(
        isw_0__zz_port_a_2), .QN() );
  DFF_X1 isw_0_z_0_reg ( .D(isw_0_xor_10_port_z), .CK(clk), .Q(isw_0_z_0), 
        .QN() );
  DFF_X1 isw_0__zz_port_b_reg ( .D(isw_0_and_10_port_z), .CK(clk), .Q(
        isw_0__zz_port_b), .QN() );
  DFF_X1 isw_0__zz_port_a_reg ( .D(isw_0_xor_9_port_z), .CK(clk), .Q(
        isw_0__zz_port_a), .QN() );
  DFF_X1 isw_0__zz_port_a_1_reg ( .D(isw_0_and_11_port_z), .CK(clk), .Q(
        isw_0__zz_port_a_1), .QN() );
  DFF_X1 isw_0__zz_port_b_1_reg ( .D(port_rand[0]), .CK(clk), .Q(
        isw_0__zz_port_b_1), .QN() );
  DFF_X1 isw_0__zz_port_a_3_reg ( .D(isw_0_and_12_port_z), .CK(clk), .Q(
        isw_0__zz_port_a_3), .QN() );
  AND2_X1 isw_0_and_9_U1 ( .A1(port_b_in[1]), .A2(port_a_in0), .ZN(
        isw_0_and_9_port_z) );
  XOR2_X1 isw_0_xor_9_U1 ( .A(isw_0_and_9_port_z), .B(port_rand[0]), .Z(
        isw_0_xor_9_port_z) );
  AND2_X1 isw_0_and_10_U1 ( .A1(port_b_in[0]), .A2(port_a_in1), .ZN(
        isw_0_and_10_port_z) );
  XOR2_X1 isw_0_xor_10_U1 ( .A(isw_0__zz_port_b), .B(isw_0__zz_port_a), .Z(
        isw_0_xor_10_port_z) );
  AND2_X1 isw_0_and_11_U1 ( .A1(port_b_in[0]), .A2(port_a_in0), .ZN(
        isw_0_and_11_port_z) );
  XOR2_X1 isw_0_xor_11_U1 ( .A(isw_0__zz_port_b_2), .B(isw_0__zz_port_a_2), 
        .Z(isw_0_xor_11_port_z) );
  AND2_X1 isw_0_and_12_U1 ( .A1(port_b_in[1]), .A2(port_a_in1), .ZN(
        isw_0_and_12_port_z) );
  XOR2_X1 isw_0_xor_12_U1 ( .A(isw_0_z_0), .B(isw_0__zz_port_a_4), .Z(
        isw_0_xor_12_port_z) );
  DFF_X1 isw_1_result_1_reg ( .D(isw_1_xor_12_port_z), .CK(clk), .Q(
        n_zz_unequal_0_1[1]), .QN() );
  DFF_X1 isw_1__zz_port_a_4_reg ( .D(isw_1__zz_port_a_3), .CK(clk), .Q(
        isw_1__zz_port_a_4), .QN() );
  DFF_X1 isw_1_result_0_reg ( .D(isw_1_xor_11_port_z), .CK(clk), .Q(
        n_zz_unequal_0_1[0]), .QN() );
  DFF_X1 isw_1__zz_port_b_2_reg ( .D(isw_1__zz_port_b_1), .CK(clk), .Q(
        isw_1__zz_port_b_2), .QN() );
  DFF_X1 isw_1__zz_port_a_2_reg ( .D(isw_1__zz_port_a_1), .CK(clk), .Q(
        isw_1__zz_port_a_2), .QN() );
  DFF_X1 isw_1_z_0_reg ( .D(isw_1_xor_10_port_z), .CK(clk), .Q(isw_1_z_0), 
        .QN() );
  DFF_X1 isw_1__zz_port_b_reg ( .D(isw_1_and_10_port_z), .CK(clk), .Q(
        isw_1__zz_port_b), .QN() );
  DFF_X1 isw_1__zz_port_a_reg ( .D(isw_1_xor_9_port_z), .CK(clk), .Q(
        isw_1__zz_port_a), .QN() );
  DFF_X1 isw_1__zz_port_a_1_reg ( .D(isw_1_and_11_port_z), .CK(clk), .Q(
        isw_1__zz_port_a_1), .QN() );
  DFF_X1 isw_1__zz_port_b_1_reg ( .D(port_rand[0]), .CK(clk), .Q(
        isw_1__zz_port_b_1), .QN() );
  DFF_X1 isw_1__zz_port_a_3_reg ( .D(isw_1_and_12_port_z), .CK(clk), .Q(
        isw_1__zz_port_a_3), .QN() );
  AND2_X1 isw_1_and_9_U1 ( .A1(port_b_in[1]), .A2(port_a_in[0]), .ZN(
        isw_1_and_9_port_z) );
  XOR2_X1 isw_1_xor_9_U1 ( .A(isw_1_and_9_port_z), .B(port_rand[0]), .Z(
        isw_1_xor_9_port_z) );
  AND2_X1 isw_1_and_10_U1 ( .A1(port_b_in[0]), .A2(port_a_in[1]), .ZN(
        isw_1_and_10_port_z) );
  XOR2_X1 isw_1_xor_10_U1 ( .A(isw_1__zz_port_b), .B(isw_1__zz_port_a), .Z(
        isw_1_xor_10_port_z) );
  AND2_X1 isw_1_and_11_U1 ( .A1(port_b_in[0]), .A2(port_a_in[0]), .ZN(
        isw_1_and_11_port_z) );
  XOR2_X1 isw_1_xor_11_U1 ( .A(isw_1__zz_port_b_2), .B(isw_1__zz_port_a_2), 
        .Z(isw_1_xor_11_port_z) );
  AND2_X1 isw_1_and_12_U1 ( .A1(port_b_in[1]), .A2(port_a_in[1]), .ZN(
        isw_1_and_12_port_z) );
  XOR2_X1 isw_1_xor_12_U1 ( .A(isw_1_z_0), .B(isw_1__zz_port_a_4), .Z(
        isw_1_xor_12_port_z) );
endmodule

