
module And_gate ( clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, 
        clock_6, reset_0, reset_1, reset_2, reset_3, reset_4, reset_5, reset_6, 
        io_i0_s0_d0, io_i0_s0_d1, io_i0_s0_d2, io_i0_s0_d3, io_i0_s0_d4, 
        io_i0_s0_d5, io_i0_s0_d6, io_i0_s1_d0, io_i0_s1_d1, io_i0_s1_d2, 
        io_i0_s1_d3, io_i0_s1_d4, io_i0_s1_d5, io_i0_s1_d6, io_i0_s2_d0, 
        io_i0_s2_d1, io_i0_s2_d2, io_i0_s2_d3, io_i0_s2_d4, io_i0_s2_d5, 
        io_i0_s2_d6, io_i0_s3_d0, io_i0_s3_d1, io_i0_s3_d2, io_i0_s3_d3, 
        io_i0_s3_d4, io_i0_s3_d5, io_i0_s3_d6, io_i1_s0_d0, io_i1_s0_d1, 
        io_i1_s0_d2, io_i1_s0_d3, io_i1_s0_d4, io_i1_s0_d5, io_i1_s0_d6, 
        io_i1_s1_d0, io_i1_s1_d1, io_i1_s1_d2, io_i1_s1_d3, io_i1_s1_d4, 
        io_i1_s1_d5, io_i1_s1_d6, io_i1_s2_d0, io_i1_s2_d1, io_i1_s2_d2, 
        io_i1_s2_d3, io_i1_s2_d4, io_i1_s2_d5, io_i1_s2_d6, io_i1_s3_d0, 
        io_i1_s3_d1, io_i1_s3_d2, io_i1_s3_d3, io_i1_s3_d4, io_i1_s3_d5, 
        io_i1_s3_d6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, 
        p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, 
        io_o0_s0_d0, io_o0_s0_d1, io_o0_s0_d2, io_o0_s0_d3, io_o0_s0_d4, 
        io_o0_s0_d5, io_o0_s0_d6, io_o0_s1_d0, io_o0_s1_d1, io_o0_s1_d2, 
        io_o0_s1_d3, io_o0_s1_d4, io_o0_s1_d5, io_o0_s1_d6, io_o0_s2_d0, 
        io_o0_s2_d1, io_o0_s2_d2, io_o0_s2_d3, io_o0_s2_d4, io_o0_s2_d5, 
        io_o0_s2_d6, io_o0_s3_d0, io_o0_s3_d1, io_o0_s3_d2, io_o0_s3_d3, 
        io_o0_s3_d4, io_o0_s3_d5, io_o0_s3_d6 );
  input clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, clock_6, reset_0,
         reset_1, reset_2, reset_3, reset_4, reset_5, reset_6, io_i0_s0_d0,
         io_i0_s0_d1, io_i0_s0_d2, io_i0_s0_d3, io_i0_s0_d4, io_i0_s0_d5,
         io_i0_s0_d6, io_i0_s1_d0, io_i0_s1_d1, io_i0_s1_d2, io_i0_s1_d3,
         io_i0_s1_d4, io_i0_s1_d5, io_i0_s1_d6, io_i0_s2_d0, io_i0_s2_d1,
         io_i0_s2_d2, io_i0_s2_d3, io_i0_s2_d4, io_i0_s2_d5, io_i0_s2_d6,
         io_i0_s3_d0, io_i0_s3_d1, io_i0_s3_d2, io_i0_s3_d3, io_i0_s3_d4,
         io_i0_s3_d5, io_i0_s3_d6, io_i1_s0_d0, io_i1_s0_d1, io_i1_s0_d2,
         io_i1_s0_d3, io_i1_s0_d4, io_i1_s0_d5, io_i1_s0_d6, io_i1_s1_d0,
         io_i1_s1_d1, io_i1_s1_d2, io_i1_s1_d3, io_i1_s1_d4, io_i1_s1_d5,
         io_i1_s1_d6, io_i1_s2_d0, io_i1_s2_d1, io_i1_s2_d2, io_i1_s2_d3,
         io_i1_s2_d4, io_i1_s2_d5, io_i1_s2_d6, io_i1_s3_d0, io_i1_s3_d1,
         io_i1_s3_d2, io_i1_s3_d3, io_i1_s3_d4, io_i1_s3_d5, io_i1_s3_d6,
         p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6,
         p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11;
  output io_o0_s0_d0, io_o0_s0_d1, io_o0_s0_d2, io_o0_s0_d3, io_o0_s0_d4,
         io_o0_s0_d5, io_o0_s0_d6, io_o0_s1_d0, io_o0_s1_d1, io_o0_s1_d2,
         io_o0_s1_d3, io_o0_s1_d4, io_o0_s1_d5, io_o0_s1_d6, io_o0_s2_d0,
         io_o0_s2_d1, io_o0_s2_d2, io_o0_s2_d3, io_o0_s2_d4, io_o0_s2_d5,
         io_o0_s2_d6, io_o0_s3_d0, io_o0_s3_d1, io_o0_s3_d2, io_o0_s3_d3,
         io_o0_s3_d4, io_o0_s3_d5, io_o0_s3_d6;
  wire   n_xor_module_1_res, n_xor_module_2_res, n_xor_module_3_res,
         n_xor_module_4_res, n_xor_module_5_res, n_xor_module_6_res,
         n_xor_module_7_res, n_xor_module_8_res, n_xor_module_9_res,
         n_xor_module_10_res, n_xor_module_11_res, n_xor_module_12_res,
         n_xor_module_13_res, n_xor_module_14_res, n_xor_module_15_res,
         n_xor_module_16_res, n_xor_module_17_res, n_xor_module_18_res,
         n_xor_module_19_res, n_xor_module_20_res, n_xor_module_21_res,
         n_xor_module_22_res, n_xor_module_23_res, n_xor_module_24_res,
         n_xor_module_25_res, n_xor_module_26_res, n_xor_module_27_res,
         n_xor_module_28_res, n_xor_module_29_res, n_xor_module_30_res,
         n_xor_module_31_res, n_xor_module_32_res, n_xor_module_33_res,
         n_xor_module_34_res, n_xor_module_35_res, n_xor_module_36_res,
         n_xor_module_37_res, n_xor_module_38_res, n_xor_module_39_res,
         n_xor_module_40_res, n_xor_module_41_res, n_xor_module_42_res,
         n_xor_module_43_res, n_xor_module_44_res, n_xor_module_45_res,
         n_xor_module_46_res, n_xor_module_47_res, n_xor_module_48_res,
         n_xor_module_49_res, n_xor_module_50_res, n_xor_module_51_res,
         n_xor_module_52_res, n_xor_module_53_res, n_xor_module_54_res,
         n_xor_module_55_res, n_xor_module_56_res, n_xor_module_57_res,
         n_xor_module_58_res, n_xor_module_59_res, n_xor_module_60_res,
         n_xor_module_61_res, n_xor_module_62_res, n_xor_module_63_res,
         n_xor_module_64_res, n_xor_module_65_res, n_xor_module_66_res,
         n_xor_module_67_res, n_xor_module_68_res, n_xor_module_69_res,
         n_xor_module_70_res, n_xor_module_71_res, n_xor_module_72_res,
         n_xor_module_73_res, n_xor_module_74_res, n_xor_module_75_res,
         n_xor_module_76_res, n_xor_module_77_res, n_xor_module_78_res,
         n_xor_module_79_res, n_xor_module_80_res, n_xor_module_81_res,
         n_xor_module_82_res, n_xor_module_83_res, n_xor_module_84_res,
         n_majority7_module_0_res, n_reg_module_1_res,
         n_majority7_module_1_res, n_reg_module_2_res,
         n_majority7_module_2_res, n_reg_module_3_res,
         n_majority7_module_3_res, n_reg_module_4_res,
         n_majority7_module_4_res, n_reg_module_5_res,
         n_majority7_module_5_res, n_reg_module_6_res,
         n_majority7_module_6_res, n_reg_module_7_res,
         n_majority7_module_7_res, n_reg_module_8_res,
         n_majority7_module_8_res, n_reg_module_9_res,
         n_majority7_module_9_res, n_reg_module_10_res,
         n_majority7_module_10_res, n_reg_module_11_res,
         n_majority7_module_11_res, n_reg_module_12_res,
         n_majority7_module_12_res, n_reg_module_13_res,
         n_majority7_module_13_res, n_reg_module_14_res,
         n_majority7_module_14_res, n_reg_module_15_res,
         n_majority7_module_15_res, n_reg_module_16_res,
         n_majority7_module_16_res, n_reg_module_17_res,
         n_majority7_module_17_res, n_reg_module_18_res,
         n_majority7_module_18_res, n_reg_module_19_res,
         n_majority7_module_19_res, n_reg_module_20_res,
         n_majority7_module_20_res, n_reg_module_21_res,
         n_majority7_module_21_res, n_reg_module_22_res,
         n_majority7_module_22_res, n_reg_module_23_res,
         n_majority7_module_23_res, n_reg_module_24_res,
         n_majority7_module_24_res, n_reg_module_25_res,
         n_majority7_module_25_res, n_reg_module_26_res,
         n_majority7_module_26_res, n_reg_module_27_res,
         n_majority7_module_27_res, n_reg_module_28_res,
         n_majority7_module_28_res, n_reg_module_29_res,
         n_majority7_module_29_res, n_reg_module_30_res,
         n_majority7_module_30_res, n_reg_module_31_res,
         n_majority7_module_31_res, n_reg_module_32_res,
         n_majority7_module_32_res, n_reg_module_33_res,
         n_majority7_module_33_res, n_reg_module_34_res,
         n_majority7_module_34_res, n_reg_module_35_res,
         n_majority7_module_35_res, n_reg_module_36_res,
         n_majority7_module_36_res, n_reg_module_37_res,
         n_majority7_module_37_res, n_reg_module_38_res,
         n_majority7_module_38_res, n_reg_module_39_res,
         n_majority7_module_39_res, n_reg_module_40_res,
         n_majority7_module_40_res, n_reg_module_41_res,
         n_majority7_module_41_res, n_reg_module_42_res,
         n_majority7_module_42_res, n_reg_module_43_res,
         n_majority7_module_43_res, n_reg_module_44_res,
         n_majority7_module_44_res, n_reg_module_45_res,
         n_majority7_module_45_res, n_reg_module_46_res,
         n_majority7_module_46_res, n_reg_module_47_res,
         n_majority7_module_47_res, n_reg_module_48_res,
         n_majority7_module_48_res, n_reg_module_49_res,
         n_majority7_module_49_res, n_reg_module_50_res,
         n_majority7_module_50_res, n_reg_module_51_res,
         n_majority7_module_51_res, n_reg_module_52_res,
         n_majority7_module_52_res, n_reg_module_53_res,
         n_majority7_module_53_res, n_reg_module_54_res,
         n_majority7_module_54_res, n_reg_module_55_res,
         n_majority7_module_55_res, n_reg_module_56_res,
         n_majority7_module_56_res, n_reg_module_57_res,
         n_majority7_module_57_res, n_reg_module_58_res,
         n_majority7_module_58_res, n_reg_module_59_res,
         n_majority7_module_59_res, n_reg_module_60_res,
         n_majority7_module_60_res, n_reg_module_61_res,
         n_majority7_module_61_res, n_reg_module_62_res,
         n_majority7_module_62_res, n_reg_module_63_res,
         n_majority7_module_63_res, n_reg_module_64_res,
         n_majority7_module_64_res, n_reg_module_65_res,
         n_majority7_module_65_res, n_reg_module_66_res,
         n_majority7_module_66_res, n_reg_module_67_res,
         n_majority7_module_67_res, n_reg_module_68_res,
         n_majority7_module_68_res, n_reg_module_69_res,
         n_majority7_module_69_res, n_reg_module_70_res,
         n_majority7_module_70_res, n_reg_module_71_res,
         n_majority7_module_71_res, n_reg_module_72_res,
         n_majority7_module_72_res, n_reg_module_73_res,
         n_majority7_module_73_res, n_reg_module_74_res,
         n_majority7_module_74_res, n_reg_module_75_res,
         n_majority7_module_75_res, n_reg_module_76_res,
         n_majority7_module_76_res, n_reg_module_77_res,
         n_majority7_module_77_res, n_reg_module_78_res,
         n_majority7_module_78_res, n_reg_module_79_res,
         n_majority7_module_79_res, n_reg_module_80_res,
         n_majority7_module_80_res, n_reg_module_81_res,
         n_majority7_module_81_res, n_reg_module_82_res,
         n_majority7_module_82_res, n_reg_module_83_res,
         n_majority7_module_83_res, n_reg_module_84_res,
         n_majority7_module_84_res, n_reg_module_85_res,
         n_majority7_module_85_res, n_reg_module_86_res,
         n_majority7_module_86_res, n_reg_module_87_res,
         n_majority7_module_87_res, n_reg_module_88_res,
         n_majority7_module_88_res, n_reg_module_89_res,
         n_majority7_module_89_res, n_reg_module_90_res,
         n_majority7_module_90_res, n_reg_module_91_res,
         n_majority7_module_91_res, n_reg_module_92_res,
         n_majority7_module_92_res, n_reg_module_93_res,
         n_majority7_module_93_res, n_reg_module_94_res,
         n_majority7_module_94_res, n_reg_module_95_res,
         n_majority7_module_95_res, n_reg_module_96_res,
         n_majority7_module_96_res, n_reg_module_97_res,
         n_majority7_module_97_res, n_reg_module_98_res,
         n_majority7_module_98_res, n_reg_module_99_res,
         n_majority7_module_99_res, n_reg_module_100_res,
         n_majority7_module_100_res, n_reg_module_101_res,
         n_majority7_module_101_res, n_reg_module_102_res,
         n_majority7_module_102_res, n_reg_module_103_res,
         n_majority7_module_103_res, n_reg_module_104_res,
         n_majority7_module_104_res, n_reg_module_105_res,
         n_majority7_module_105_res, n_reg_module_106_res,
         n_majority7_module_106_res, n_reg_module_107_res,
         n_majority7_module_107_res, n_reg_module_108_res,
         n_majority7_module_108_res, n_reg_module_109_res,
         n_majority7_module_109_res, n_reg_module_110_res,
         n_majority7_module_110_res, n_reg_module_111_res,
         n_majority7_module_111_res, n_reg_module_112_res, n_and_module_1_res,
         n_reg_module_113_res, n_and_module_2_res, n_xor_module_85_res,
         n_reg_module_114_res, n_and_module_3_res, n_xor_module_86_res,
         n_reg_module_115_res, n_and_module_4_res, n_xor_module_87_res,
         n_reg_module_116_res, n_and_module_5_res, n_xor_module_88_res,
         n_reg_module_117_res, n_and_module_6_res, n_reg_module_118_res,
         n_and_module_7_res, n_xor_module_89_res, n_reg_module_119_res,
         n_and_module_8_res, n_xor_module_90_res, n_reg_module_120_res,
         n_and_module_9_res, n_xor_module_91_res, n_reg_module_121_res,
         n_and_module_10_res, n_xor_module_92_res, n_reg_module_122_res,
         n_and_module_11_res, n_reg_module_123_res, n_and_module_12_res,
         n_xor_module_93_res, n_reg_module_124_res, n_and_module_13_res,
         n_xor_module_94_res, n_reg_module_125_res, n_and_module_14_res,
         n_xor_module_95_res, n_reg_module_126_res, n_and_module_15_res,
         n_xor_module_96_res, n_reg_module_127_res, n_and_module_16_res,
         n_reg_module_128_res, n_and_module_17_res, n_reg_module_129_res,
         n_and_module_18_res, n_xor_module_97_res, n_reg_module_130_res,
         n_and_module_19_res, n_xor_module_98_res, n_reg_module_131_res,
         n_and_module_20_res, n_xor_module_99_res, n_reg_module_132_res,
         n_and_module_21_res, n_xor_module_100_res, n_reg_module_133_res,
         n_and_module_22_res, n_reg_module_134_res, n_and_module_23_res,
         n_xor_module_101_res, n_reg_module_135_res, n_and_module_24_res,
         n_xor_module_102_res, n_reg_module_136_res, n_and_module_25_res,
         n_xor_module_103_res, n_reg_module_137_res, n_and_module_26_res,
         n_xor_module_104_res, n_reg_module_138_res, n_and_module_27_res,
         n_reg_module_139_res, n_and_module_28_res, n_xor_module_105_res,
         n_reg_module_140_res, n_and_module_29_res, n_xor_module_106_res,
         n_reg_module_141_res, n_and_module_30_res, n_xor_module_107_res,
         n_reg_module_142_res, n_and_module_31_res, n_xor_module_108_res,
         n_reg_module_143_res, n_and_module_32_res, n_reg_module_144_res,
         n_and_module_33_res, n_reg_module_145_res, n_and_module_34_res,
         n_xor_module_109_res, n_reg_module_146_res, n_and_module_35_res,
         n_xor_module_110_res, n_reg_module_147_res, n_and_module_36_res,
         n_xor_module_111_res, n_reg_module_148_res, n_and_module_37_res,
         n_xor_module_112_res, n_reg_module_149_res, n_and_module_38_res,
         n_reg_module_150_res, n_and_module_39_res, n_xor_module_113_res,
         n_reg_module_151_res, n_and_module_40_res, n_xor_module_114_res,
         n_reg_module_152_res, n_and_module_41_res, n_xor_module_115_res,
         n_reg_module_153_res, n_and_module_42_res, n_xor_module_116_res,
         n_reg_module_154_res, n_and_module_43_res, n_reg_module_155_res,
         n_and_module_44_res, n_xor_module_117_res, n_reg_module_156_res,
         n_and_module_45_res, n_xor_module_118_res, n_reg_module_157_res,
         n_and_module_46_res, n_xor_module_119_res, n_reg_module_158_res,
         n_and_module_47_res, n_xor_module_120_res, n_reg_module_159_res,
         n_and_module_48_res, n_reg_module_160_res, n_and_module_49_res,
         n_reg_module_161_res, n_and_module_50_res, n_xor_module_121_res,
         n_reg_module_162_res, n_and_module_51_res, n_xor_module_122_res,
         n_reg_module_163_res, n_and_module_52_res, n_xor_module_123_res,
         n_reg_module_164_res, n_and_module_53_res, n_xor_module_124_res,
         n_reg_module_165_res, n_and_module_54_res, n_reg_module_166_res,
         n_and_module_55_res, n_xor_module_125_res, n_reg_module_167_res,
         n_and_module_56_res, n_xor_module_126_res, n_reg_module_168_res,
         n_and_module_57_res, n_xor_module_127_res, n_reg_module_169_res,
         n_and_module_58_res, n_xor_module_128_res, n_reg_module_170_res,
         n_and_module_59_res, n_reg_module_171_res, n_and_module_60_res,
         n_xor_module_129_res, n_reg_module_172_res, n_and_module_61_res,
         n_xor_module_130_res, n_reg_module_173_res, n_and_module_62_res,
         n_xor_module_131_res, n_reg_module_174_res, n_and_module_63_res,
         n_xor_module_132_res, n_reg_module_175_res, n_and_module_64_res,
         n_reg_module_176_res, n_and_module_65_res, n_reg_module_177_res,
         n_and_module_66_res, n_xor_module_133_res, n_reg_module_178_res,
         n_and_module_67_res, n_xor_module_134_res, n_reg_module_179_res,
         n_and_module_68_res, n_xor_module_135_res, n_reg_module_180_res,
         n_and_module_69_res, n_xor_module_136_res, n_reg_module_181_res,
         n_and_module_70_res, n_reg_module_182_res, n_and_module_71_res,
         n_xor_module_137_res, n_reg_module_183_res, n_and_module_72_res,
         n_xor_module_138_res, n_reg_module_184_res, n_and_module_73_res,
         n_xor_module_139_res, n_reg_module_185_res, n_and_module_74_res,
         n_xor_module_140_res, n_reg_module_186_res, n_and_module_75_res,
         n_reg_module_187_res, n_and_module_76_res, n_xor_module_141_res,
         n_reg_module_188_res, n_and_module_77_res, n_xor_module_142_res,
         n_reg_module_189_res, n_and_module_78_res, n_xor_module_143_res,
         n_reg_module_190_res, n_and_module_79_res, n_xor_module_144_res,
         n_reg_module_191_res, n_and_module_80_res, n_reg_module_192_res,
         n_and_module_81_res, n_reg_module_193_res, n_and_module_82_res,
         n_xor_module_145_res, n_reg_module_194_res, n_and_module_83_res,
         n_xor_module_146_res, n_reg_module_195_res, n_and_module_84_res,
         n_xor_module_147_res, n_reg_module_196_res, n_and_module_85_res,
         n_xor_module_148_res, n_reg_module_197_res, n_and_module_86_res,
         n_reg_module_198_res, n_and_module_87_res, n_xor_module_149_res,
         n_reg_module_199_res, n_and_module_88_res, n_xor_module_150_res,
         n_reg_module_200_res, n_and_module_89_res, n_xor_module_151_res,
         n_reg_module_201_res, n_and_module_90_res, n_xor_module_152_res,
         n_reg_module_202_res, n_and_module_91_res, n_reg_module_203_res,
         n_and_module_92_res, n_xor_module_153_res, n_reg_module_204_res,
         n_and_module_93_res, n_xor_module_154_res, n_reg_module_205_res,
         n_and_module_94_res, n_xor_module_155_res, n_reg_module_206_res,
         n_and_module_95_res, n_xor_module_156_res, n_reg_module_207_res,
         n_and_module_96_res, n_reg_module_208_res, n_and_module_97_res,
         n_reg_module_209_res, n_and_module_98_res, n_xor_module_157_res,
         n_reg_module_210_res, n_and_module_99_res, n_xor_module_158_res,
         n_reg_module_211_res, n_and_module_100_res, n_xor_module_159_res,
         n_reg_module_212_res, n_and_module_101_res, n_xor_module_160_res,
         n_reg_module_213_res, n_and_module_102_res, n_reg_module_214_res,
         n_and_module_103_res, n_xor_module_161_res, n_reg_module_215_res,
         n_and_module_104_res, n_xor_module_162_res, n_reg_module_216_res,
         n_and_module_105_res, n_xor_module_163_res, n_reg_module_217_res,
         n_and_module_106_res, n_xor_module_164_res, n_reg_module_218_res,
         n_and_module_107_res, n_reg_module_219_res, n_and_module_108_res,
         n_xor_module_165_res, n_reg_module_220_res, n_and_module_109_res,
         n_xor_module_166_res, n_reg_module_221_res, n_and_module_110_res,
         n_xor_module_167_res, n_reg_module_222_res, n_and_module_111_res,
         n_xor_module_168_res, n_reg_module_223_res, n_and_module_112_res,
         n_reg_module_224_res, n_xor_module_169_res, n_xor_module_170_res,
         n_xor_module_172_res, n_xor_module_173_res, n_xor_module_175_res,
         n_xor_module_176_res, n_xor_module_178_res, n_xor_module_179_res,
         n_xor_module_181_res, n_xor_module_182_res, n_xor_module_184_res,
         n_xor_module_185_res, n_xor_module_187_res, n_xor_module_188_res,
         n_xor_module_190_res, n_xor_module_191_res, n_xor_module_193_res,
         n_xor_module_194_res, n_xor_module_196_res, n_xor_module_197_res,
         n_xor_module_199_res, n_xor_module_200_res, n_xor_module_202_res,
         n_xor_module_203_res, n_xor_module_205_res, n_xor_module_206_res,
         n_xor_module_208_res, n_xor_module_209_res, n_xor_module_211_res,
         n_xor_module_212_res, n_xor_module_214_res, n_xor_module_215_res,
         n_xor_module_217_res, n_xor_module_218_res, n_xor_module_220_res,
         n_xor_module_221_res, n_xor_module_223_res, n_xor_module_224_res,
         n_xor_module_226_res, n_xor_module_227_res, n_xor_module_229_res,
         n_xor_module_230_res, n_xor_module_232_res, n_xor_module_233_res,
         n_xor_module_235_res, n_xor_module_236_res, n_xor_module_238_res,
         n_xor_module_239_res, n_xor_module_241_res, n_xor_module_242_res,
         n_xor_module_244_res, n_xor_module_245_res, n_xor_module_247_res,
         n_xor_module_248_res, n_xor_module_250_res, n_xor_module_251_res,
         n_xor_module_3_n2, n_xor_module_6_n2, n_xor_module_9_n2,
         n_xor_module_12_n2, n_xor_module_15_n2, n_xor_module_18_n2,
         n_xor_module_21_n2, n_xor_module_24_n2, n_xor_module_27_n2,
         n_xor_module_30_n2, n_xor_module_33_n2, n_xor_module_36_n2,
         n_xor_module_39_n2, n_xor_module_42_n2, n_xor_module_45_n2,
         n_xor_module_48_n2, n_xor_module_51_n2, n_xor_module_54_n2,
         n_xor_module_57_n2, n_xor_module_60_n2, n_xor_module_63_n2,
         n_xor_module_66_n2, n_xor_module_69_n2, n_xor_module_72_n2,
         n_xor_module_75_n2, n_xor_module_78_n2, n_xor_module_81_n2,
         n_xor_module_84_n2, n_majority7_module_0_n7, n_majority7_module_0_n6,
         n_majority7_module_0_n5, n_majority7_module_0_n4,
         n_majority7_module_0_n3, n_majority7_module_0_n2,
         n_majority7_module_0_n1, n_majority7_module_0__and_module_10_res,
         n_majority7_module_0__or_module_11_res,
         n_majority7_module_0__and_module_9_res,
         n_majority7_module_0__or_module_10_res,
         n_majority7_module_0__or_module_9_res,
         n_majority7_module_0__and_module_8_res,
         n_majority7_module_0__or_module_8_res,
         n_majority7_module_0__and_module_7_res,
         n_majority7_module_0__or_module_7_res,
         n_majority7_module_0__or_module_6_res,
         n_majority7_module_0__and_module_6_res,
         n_majority7_module_0__or_module_5_res,
         n_majority7_module_0__and_module_5_res,
         n_majority7_module_0__or_module_4_res,
         n_majority7_module_0__and_module_4_res,
         n_majority7_module_0__or_module_3_res,
         n_majority7_module_0__and_module_3_res,
         n_majority7_module_0__or_module_2_res,
         n_majority7_module_0__and_module_2_res,
         n_majority7_module_0__or_module_1_res,
         n_majority7_module_0__and_module_1_res, n_majority7_module_1_n7,
         n_majority7_module_1_n6, n_majority7_module_1_n5,
         n_majority7_module_1_n4, n_majority7_module_1_n3,
         n_majority7_module_1_n2, n_majority7_module_1_n1,
         n_majority7_module_1__and_module_10_res,
         n_majority7_module_1__or_module_11_res,
         n_majority7_module_1__and_module_9_res,
         n_majority7_module_1__or_module_10_res,
         n_majority7_module_1__or_module_9_res,
         n_majority7_module_1__and_module_8_res,
         n_majority7_module_1__or_module_8_res,
         n_majority7_module_1__and_module_7_res,
         n_majority7_module_1__or_module_7_res,
         n_majority7_module_1__or_module_6_res,
         n_majority7_module_1__and_module_6_res,
         n_majority7_module_1__or_module_5_res,
         n_majority7_module_1__and_module_5_res,
         n_majority7_module_1__or_module_4_res,
         n_majority7_module_1__and_module_4_res,
         n_majority7_module_1__or_module_3_res,
         n_majority7_module_1__and_module_3_res,
         n_majority7_module_1__or_module_2_res,
         n_majority7_module_1__and_module_2_res,
         n_majority7_module_1__or_module_1_res,
         n_majority7_module_1__and_module_1_res, n_majority7_module_2_n7,
         n_majority7_module_2_n6, n_majority7_module_2_n5,
         n_majority7_module_2_n4, n_majority7_module_2_n3,
         n_majority7_module_2_n2, n_majority7_module_2_n1,
         n_majority7_module_2__and_module_10_res,
         n_majority7_module_2__or_module_11_res,
         n_majority7_module_2__and_module_9_res,
         n_majority7_module_2__or_module_10_res,
         n_majority7_module_2__or_module_9_res,
         n_majority7_module_2__and_module_8_res,
         n_majority7_module_2__or_module_8_res,
         n_majority7_module_2__and_module_7_res,
         n_majority7_module_2__or_module_7_res,
         n_majority7_module_2__or_module_6_res,
         n_majority7_module_2__and_module_6_res,
         n_majority7_module_2__or_module_5_res,
         n_majority7_module_2__and_module_5_res,
         n_majority7_module_2__or_module_4_res,
         n_majority7_module_2__and_module_4_res,
         n_majority7_module_2__or_module_3_res,
         n_majority7_module_2__and_module_3_res,
         n_majority7_module_2__or_module_2_res,
         n_majority7_module_2__and_module_2_res,
         n_majority7_module_2__or_module_1_res,
         n_majority7_module_2__and_module_1_res, n_majority7_module_3_n7,
         n_majority7_module_3_n6, n_majority7_module_3_n5,
         n_majority7_module_3_n4, n_majority7_module_3_n3,
         n_majority7_module_3_n2, n_majority7_module_3_n1,
         n_majority7_module_3__and_module_10_res,
         n_majority7_module_3__or_module_11_res,
         n_majority7_module_3__and_module_9_res,
         n_majority7_module_3__or_module_10_res,
         n_majority7_module_3__or_module_9_res,
         n_majority7_module_3__and_module_8_res,
         n_majority7_module_3__or_module_8_res,
         n_majority7_module_3__and_module_7_res,
         n_majority7_module_3__or_module_7_res,
         n_majority7_module_3__or_module_6_res,
         n_majority7_module_3__and_module_6_res,
         n_majority7_module_3__or_module_5_res,
         n_majority7_module_3__and_module_5_res,
         n_majority7_module_3__or_module_4_res,
         n_majority7_module_3__and_module_4_res,
         n_majority7_module_3__or_module_3_res,
         n_majority7_module_3__and_module_3_res,
         n_majority7_module_3__or_module_2_res,
         n_majority7_module_3__and_module_2_res,
         n_majority7_module_3__or_module_1_res,
         n_majority7_module_3__and_module_1_res, n_majority7_module_4_n7,
         n_majority7_module_4_n6, n_majority7_module_4_n5,
         n_majority7_module_4_n4, n_majority7_module_4_n3,
         n_majority7_module_4_n2, n_majority7_module_4_n1,
         n_majority7_module_4__and_module_10_res,
         n_majority7_module_4__or_module_11_res,
         n_majority7_module_4__and_module_9_res,
         n_majority7_module_4__or_module_10_res,
         n_majority7_module_4__or_module_9_res,
         n_majority7_module_4__and_module_8_res,
         n_majority7_module_4__or_module_8_res,
         n_majority7_module_4__and_module_7_res,
         n_majority7_module_4__or_module_7_res,
         n_majority7_module_4__or_module_6_res,
         n_majority7_module_4__and_module_6_res,
         n_majority7_module_4__or_module_5_res,
         n_majority7_module_4__and_module_5_res,
         n_majority7_module_4__or_module_4_res,
         n_majority7_module_4__and_module_4_res,
         n_majority7_module_4__or_module_3_res,
         n_majority7_module_4__and_module_3_res,
         n_majority7_module_4__or_module_2_res,
         n_majority7_module_4__and_module_2_res,
         n_majority7_module_4__or_module_1_res,
         n_majority7_module_4__and_module_1_res, n_majority7_module_5_n7,
         n_majority7_module_5_n6, n_majority7_module_5_n5,
         n_majority7_module_5_n4, n_majority7_module_5_n3,
         n_majority7_module_5_n2, n_majority7_module_5_n1,
         n_majority7_module_5__and_module_10_res,
         n_majority7_module_5__or_module_11_res,
         n_majority7_module_5__and_module_9_res,
         n_majority7_module_5__or_module_10_res,
         n_majority7_module_5__or_module_9_res,
         n_majority7_module_5__and_module_8_res,
         n_majority7_module_5__or_module_8_res,
         n_majority7_module_5__and_module_7_res,
         n_majority7_module_5__or_module_7_res,
         n_majority7_module_5__or_module_6_res,
         n_majority7_module_5__and_module_6_res,
         n_majority7_module_5__or_module_5_res,
         n_majority7_module_5__and_module_5_res,
         n_majority7_module_5__or_module_4_res,
         n_majority7_module_5__and_module_4_res,
         n_majority7_module_5__or_module_3_res,
         n_majority7_module_5__and_module_3_res,
         n_majority7_module_5__or_module_2_res,
         n_majority7_module_5__and_module_2_res,
         n_majority7_module_5__or_module_1_res,
         n_majority7_module_5__and_module_1_res, n_majority7_module_6_n7,
         n_majority7_module_6_n6, n_majority7_module_6_n5,
         n_majority7_module_6_n4, n_majority7_module_6_n3,
         n_majority7_module_6_n2, n_majority7_module_6_n1,
         n_majority7_module_6__and_module_10_res,
         n_majority7_module_6__or_module_11_res,
         n_majority7_module_6__and_module_9_res,
         n_majority7_module_6__or_module_10_res,
         n_majority7_module_6__or_module_9_res,
         n_majority7_module_6__and_module_8_res,
         n_majority7_module_6__or_module_8_res,
         n_majority7_module_6__and_module_7_res,
         n_majority7_module_6__or_module_7_res,
         n_majority7_module_6__or_module_6_res,
         n_majority7_module_6__and_module_6_res,
         n_majority7_module_6__or_module_5_res,
         n_majority7_module_6__and_module_5_res,
         n_majority7_module_6__or_module_4_res,
         n_majority7_module_6__and_module_4_res,
         n_majority7_module_6__or_module_3_res,
         n_majority7_module_6__and_module_3_res,
         n_majority7_module_6__or_module_2_res,
         n_majority7_module_6__and_module_2_res,
         n_majority7_module_6__or_module_1_res,
         n_majority7_module_6__and_module_1_res, n_majority7_module_7_n7,
         n_majority7_module_7_n6, n_majority7_module_7_n5,
         n_majority7_module_7_n4, n_majority7_module_7_n3,
         n_majority7_module_7_n2, n_majority7_module_7_n1,
         n_majority7_module_7__and_module_10_res,
         n_majority7_module_7__or_module_11_res,
         n_majority7_module_7__and_module_9_res,
         n_majority7_module_7__or_module_10_res,
         n_majority7_module_7__or_module_9_res,
         n_majority7_module_7__and_module_8_res,
         n_majority7_module_7__or_module_8_res,
         n_majority7_module_7__and_module_7_res,
         n_majority7_module_7__or_module_7_res,
         n_majority7_module_7__or_module_6_res,
         n_majority7_module_7__and_module_6_res,
         n_majority7_module_7__or_module_5_res,
         n_majority7_module_7__and_module_5_res,
         n_majority7_module_7__or_module_4_res,
         n_majority7_module_7__and_module_4_res,
         n_majority7_module_7__or_module_3_res,
         n_majority7_module_7__and_module_3_res,
         n_majority7_module_7__or_module_2_res,
         n_majority7_module_7__and_module_2_res,
         n_majority7_module_7__or_module_1_res,
         n_majority7_module_7__and_module_1_res, n_majority7_module_8_n7,
         n_majority7_module_8_n6, n_majority7_module_8_n5,
         n_majority7_module_8_n4, n_majority7_module_8_n3,
         n_majority7_module_8_n2, n_majority7_module_8_n1,
         n_majority7_module_8__and_module_10_res,
         n_majority7_module_8__or_module_11_res,
         n_majority7_module_8__and_module_9_res,
         n_majority7_module_8__or_module_10_res,
         n_majority7_module_8__or_module_9_res,
         n_majority7_module_8__and_module_8_res,
         n_majority7_module_8__or_module_8_res,
         n_majority7_module_8__and_module_7_res,
         n_majority7_module_8__or_module_7_res,
         n_majority7_module_8__or_module_6_res,
         n_majority7_module_8__and_module_6_res,
         n_majority7_module_8__or_module_5_res,
         n_majority7_module_8__and_module_5_res,
         n_majority7_module_8__or_module_4_res,
         n_majority7_module_8__and_module_4_res,
         n_majority7_module_8__or_module_3_res,
         n_majority7_module_8__and_module_3_res,
         n_majority7_module_8__or_module_2_res,
         n_majority7_module_8__and_module_2_res,
         n_majority7_module_8__or_module_1_res,
         n_majority7_module_8__and_module_1_res, n_majority7_module_9_n7,
         n_majority7_module_9_n6, n_majority7_module_9_n5,
         n_majority7_module_9_n4, n_majority7_module_9_n3,
         n_majority7_module_9_n2, n_majority7_module_9_n1,
         n_majority7_module_9__and_module_10_res,
         n_majority7_module_9__or_module_11_res,
         n_majority7_module_9__and_module_9_res,
         n_majority7_module_9__or_module_10_res,
         n_majority7_module_9__or_module_9_res,
         n_majority7_module_9__and_module_8_res,
         n_majority7_module_9__or_module_8_res,
         n_majority7_module_9__and_module_7_res,
         n_majority7_module_9__or_module_7_res,
         n_majority7_module_9__or_module_6_res,
         n_majority7_module_9__and_module_6_res,
         n_majority7_module_9__or_module_5_res,
         n_majority7_module_9__and_module_5_res,
         n_majority7_module_9__or_module_4_res,
         n_majority7_module_9__and_module_4_res,
         n_majority7_module_9__or_module_3_res,
         n_majority7_module_9__and_module_3_res,
         n_majority7_module_9__or_module_2_res,
         n_majority7_module_9__and_module_2_res,
         n_majority7_module_9__or_module_1_res,
         n_majority7_module_9__and_module_1_res, n_majority7_module_10_n7,
         n_majority7_module_10_n6, n_majority7_module_10_n5,
         n_majority7_module_10_n4, n_majority7_module_10_n3,
         n_majority7_module_10_n2, n_majority7_module_10_n1,
         n_majority7_module_10__and_module_10_res,
         n_majority7_module_10__or_module_11_res,
         n_majority7_module_10__and_module_9_res,
         n_majority7_module_10__or_module_10_res,
         n_majority7_module_10__or_module_9_res,
         n_majority7_module_10__and_module_8_res,
         n_majority7_module_10__or_module_8_res,
         n_majority7_module_10__and_module_7_res,
         n_majority7_module_10__or_module_7_res,
         n_majority7_module_10__or_module_6_res,
         n_majority7_module_10__and_module_6_res,
         n_majority7_module_10__or_module_5_res,
         n_majority7_module_10__and_module_5_res,
         n_majority7_module_10__or_module_4_res,
         n_majority7_module_10__and_module_4_res,
         n_majority7_module_10__or_module_3_res,
         n_majority7_module_10__and_module_3_res,
         n_majority7_module_10__or_module_2_res,
         n_majority7_module_10__and_module_2_res,
         n_majority7_module_10__or_module_1_res,
         n_majority7_module_10__and_module_1_res, n_majority7_module_11_n7,
         n_majority7_module_11_n6, n_majority7_module_11_n5,
         n_majority7_module_11_n4, n_majority7_module_11_n3,
         n_majority7_module_11_n2, n_majority7_module_11_n1,
         n_majority7_module_11__and_module_10_res,
         n_majority7_module_11__or_module_11_res,
         n_majority7_module_11__and_module_9_res,
         n_majority7_module_11__or_module_10_res,
         n_majority7_module_11__or_module_9_res,
         n_majority7_module_11__and_module_8_res,
         n_majority7_module_11__or_module_8_res,
         n_majority7_module_11__and_module_7_res,
         n_majority7_module_11__or_module_7_res,
         n_majority7_module_11__or_module_6_res,
         n_majority7_module_11__and_module_6_res,
         n_majority7_module_11__or_module_5_res,
         n_majority7_module_11__and_module_5_res,
         n_majority7_module_11__or_module_4_res,
         n_majority7_module_11__and_module_4_res,
         n_majority7_module_11__or_module_3_res,
         n_majority7_module_11__and_module_3_res,
         n_majority7_module_11__or_module_2_res,
         n_majority7_module_11__and_module_2_res,
         n_majority7_module_11__or_module_1_res,
         n_majority7_module_11__and_module_1_res, n_majority7_module_12_n7,
         n_majority7_module_12_n6, n_majority7_module_12_n5,
         n_majority7_module_12_n4, n_majority7_module_12_n3,
         n_majority7_module_12_n2, n_majority7_module_12_n1,
         n_majority7_module_12__and_module_10_res,
         n_majority7_module_12__or_module_11_res,
         n_majority7_module_12__and_module_9_res,
         n_majority7_module_12__or_module_10_res,
         n_majority7_module_12__or_module_9_res,
         n_majority7_module_12__and_module_8_res,
         n_majority7_module_12__or_module_8_res,
         n_majority7_module_12__and_module_7_res,
         n_majority7_module_12__or_module_7_res,
         n_majority7_module_12__or_module_6_res,
         n_majority7_module_12__and_module_6_res,
         n_majority7_module_12__or_module_5_res,
         n_majority7_module_12__and_module_5_res,
         n_majority7_module_12__or_module_4_res,
         n_majority7_module_12__and_module_4_res,
         n_majority7_module_12__or_module_3_res,
         n_majority7_module_12__and_module_3_res,
         n_majority7_module_12__or_module_2_res,
         n_majority7_module_12__and_module_2_res,
         n_majority7_module_12__or_module_1_res,
         n_majority7_module_12__and_module_1_res, n_majority7_module_13_n7,
         n_majority7_module_13_n6, n_majority7_module_13_n5,
         n_majority7_module_13_n4, n_majority7_module_13_n3,
         n_majority7_module_13_n2, n_majority7_module_13_n1,
         n_majority7_module_13__and_module_10_res,
         n_majority7_module_13__or_module_11_res,
         n_majority7_module_13__and_module_9_res,
         n_majority7_module_13__or_module_10_res,
         n_majority7_module_13__or_module_9_res,
         n_majority7_module_13__and_module_8_res,
         n_majority7_module_13__or_module_8_res,
         n_majority7_module_13__and_module_7_res,
         n_majority7_module_13__or_module_7_res,
         n_majority7_module_13__or_module_6_res,
         n_majority7_module_13__and_module_6_res,
         n_majority7_module_13__or_module_5_res,
         n_majority7_module_13__and_module_5_res,
         n_majority7_module_13__or_module_4_res,
         n_majority7_module_13__and_module_4_res,
         n_majority7_module_13__or_module_3_res,
         n_majority7_module_13__and_module_3_res,
         n_majority7_module_13__or_module_2_res,
         n_majority7_module_13__and_module_2_res,
         n_majority7_module_13__or_module_1_res,
         n_majority7_module_13__and_module_1_res, n_majority7_module_14_n7,
         n_majority7_module_14_n6, n_majority7_module_14_n5,
         n_majority7_module_14_n4, n_majority7_module_14_n3,
         n_majority7_module_14_n2, n_majority7_module_14_n1,
         n_majority7_module_14__and_module_10_res,
         n_majority7_module_14__or_module_11_res,
         n_majority7_module_14__and_module_9_res,
         n_majority7_module_14__or_module_10_res,
         n_majority7_module_14__or_module_9_res,
         n_majority7_module_14__and_module_8_res,
         n_majority7_module_14__or_module_8_res,
         n_majority7_module_14__and_module_7_res,
         n_majority7_module_14__or_module_7_res,
         n_majority7_module_14__or_module_6_res,
         n_majority7_module_14__and_module_6_res,
         n_majority7_module_14__or_module_5_res,
         n_majority7_module_14__and_module_5_res,
         n_majority7_module_14__or_module_4_res,
         n_majority7_module_14__and_module_4_res,
         n_majority7_module_14__or_module_3_res,
         n_majority7_module_14__and_module_3_res,
         n_majority7_module_14__or_module_2_res,
         n_majority7_module_14__and_module_2_res,
         n_majority7_module_14__or_module_1_res,
         n_majority7_module_14__and_module_1_res, n_majority7_module_15_n7,
         n_majority7_module_15_n6, n_majority7_module_15_n5,
         n_majority7_module_15_n4, n_majority7_module_15_n3,
         n_majority7_module_15_n2, n_majority7_module_15_n1,
         n_majority7_module_15__and_module_10_res,
         n_majority7_module_15__or_module_11_res,
         n_majority7_module_15__and_module_9_res,
         n_majority7_module_15__or_module_10_res,
         n_majority7_module_15__or_module_9_res,
         n_majority7_module_15__and_module_8_res,
         n_majority7_module_15__or_module_8_res,
         n_majority7_module_15__and_module_7_res,
         n_majority7_module_15__or_module_7_res,
         n_majority7_module_15__or_module_6_res,
         n_majority7_module_15__and_module_6_res,
         n_majority7_module_15__or_module_5_res,
         n_majority7_module_15__and_module_5_res,
         n_majority7_module_15__or_module_4_res,
         n_majority7_module_15__and_module_4_res,
         n_majority7_module_15__or_module_3_res,
         n_majority7_module_15__and_module_3_res,
         n_majority7_module_15__or_module_2_res,
         n_majority7_module_15__and_module_2_res,
         n_majority7_module_15__or_module_1_res,
         n_majority7_module_15__and_module_1_res, n_majority7_module_16_n7,
         n_majority7_module_16_n6, n_majority7_module_16_n5,
         n_majority7_module_16_n4, n_majority7_module_16_n3,
         n_majority7_module_16_n2, n_majority7_module_16_n1,
         n_majority7_module_16__and_module_10_res,
         n_majority7_module_16__or_module_11_res,
         n_majority7_module_16__and_module_9_res,
         n_majority7_module_16__or_module_10_res,
         n_majority7_module_16__or_module_9_res,
         n_majority7_module_16__and_module_8_res,
         n_majority7_module_16__or_module_8_res,
         n_majority7_module_16__and_module_7_res,
         n_majority7_module_16__or_module_7_res,
         n_majority7_module_16__or_module_6_res,
         n_majority7_module_16__and_module_6_res,
         n_majority7_module_16__or_module_5_res,
         n_majority7_module_16__and_module_5_res,
         n_majority7_module_16__or_module_4_res,
         n_majority7_module_16__and_module_4_res,
         n_majority7_module_16__or_module_3_res,
         n_majority7_module_16__and_module_3_res,
         n_majority7_module_16__or_module_2_res,
         n_majority7_module_16__and_module_2_res,
         n_majority7_module_16__or_module_1_res,
         n_majority7_module_16__and_module_1_res, n_majority7_module_17_n7,
         n_majority7_module_17_n6, n_majority7_module_17_n5,
         n_majority7_module_17_n4, n_majority7_module_17_n3,
         n_majority7_module_17_n2, n_majority7_module_17_n1,
         n_majority7_module_17__and_module_10_res,
         n_majority7_module_17__or_module_11_res,
         n_majority7_module_17__and_module_9_res,
         n_majority7_module_17__or_module_10_res,
         n_majority7_module_17__or_module_9_res,
         n_majority7_module_17__and_module_8_res,
         n_majority7_module_17__or_module_8_res,
         n_majority7_module_17__and_module_7_res,
         n_majority7_module_17__or_module_7_res,
         n_majority7_module_17__or_module_6_res,
         n_majority7_module_17__and_module_6_res,
         n_majority7_module_17__or_module_5_res,
         n_majority7_module_17__and_module_5_res,
         n_majority7_module_17__or_module_4_res,
         n_majority7_module_17__and_module_4_res,
         n_majority7_module_17__or_module_3_res,
         n_majority7_module_17__and_module_3_res,
         n_majority7_module_17__or_module_2_res,
         n_majority7_module_17__and_module_2_res,
         n_majority7_module_17__or_module_1_res,
         n_majority7_module_17__and_module_1_res, n_majority7_module_18_n7,
         n_majority7_module_18_n6, n_majority7_module_18_n5,
         n_majority7_module_18_n4, n_majority7_module_18_n3,
         n_majority7_module_18_n2, n_majority7_module_18_n1,
         n_majority7_module_18__and_module_10_res,
         n_majority7_module_18__or_module_11_res,
         n_majority7_module_18__and_module_9_res,
         n_majority7_module_18__or_module_10_res,
         n_majority7_module_18__or_module_9_res,
         n_majority7_module_18__and_module_8_res,
         n_majority7_module_18__or_module_8_res,
         n_majority7_module_18__and_module_7_res,
         n_majority7_module_18__or_module_7_res,
         n_majority7_module_18__or_module_6_res,
         n_majority7_module_18__and_module_6_res,
         n_majority7_module_18__or_module_5_res,
         n_majority7_module_18__and_module_5_res,
         n_majority7_module_18__or_module_4_res,
         n_majority7_module_18__and_module_4_res,
         n_majority7_module_18__or_module_3_res,
         n_majority7_module_18__and_module_3_res,
         n_majority7_module_18__or_module_2_res,
         n_majority7_module_18__and_module_2_res,
         n_majority7_module_18__or_module_1_res,
         n_majority7_module_18__and_module_1_res, n_majority7_module_19_n7,
         n_majority7_module_19_n6, n_majority7_module_19_n5,
         n_majority7_module_19_n4, n_majority7_module_19_n3,
         n_majority7_module_19_n2, n_majority7_module_19_n1,
         n_majority7_module_19__and_module_10_res,
         n_majority7_module_19__or_module_11_res,
         n_majority7_module_19__and_module_9_res,
         n_majority7_module_19__or_module_10_res,
         n_majority7_module_19__or_module_9_res,
         n_majority7_module_19__and_module_8_res,
         n_majority7_module_19__or_module_8_res,
         n_majority7_module_19__and_module_7_res,
         n_majority7_module_19__or_module_7_res,
         n_majority7_module_19__or_module_6_res,
         n_majority7_module_19__and_module_6_res,
         n_majority7_module_19__or_module_5_res,
         n_majority7_module_19__and_module_5_res,
         n_majority7_module_19__or_module_4_res,
         n_majority7_module_19__and_module_4_res,
         n_majority7_module_19__or_module_3_res,
         n_majority7_module_19__and_module_3_res,
         n_majority7_module_19__or_module_2_res,
         n_majority7_module_19__and_module_2_res,
         n_majority7_module_19__or_module_1_res,
         n_majority7_module_19__and_module_1_res, n_majority7_module_20_n7,
         n_majority7_module_20_n6, n_majority7_module_20_n5,
         n_majority7_module_20_n4, n_majority7_module_20_n3,
         n_majority7_module_20_n2, n_majority7_module_20_n1,
         n_majority7_module_20__and_module_10_res,
         n_majority7_module_20__or_module_11_res,
         n_majority7_module_20__and_module_9_res,
         n_majority7_module_20__or_module_10_res,
         n_majority7_module_20__or_module_9_res,
         n_majority7_module_20__and_module_8_res,
         n_majority7_module_20__or_module_8_res,
         n_majority7_module_20__and_module_7_res,
         n_majority7_module_20__or_module_7_res,
         n_majority7_module_20__or_module_6_res,
         n_majority7_module_20__and_module_6_res,
         n_majority7_module_20__or_module_5_res,
         n_majority7_module_20__and_module_5_res,
         n_majority7_module_20__or_module_4_res,
         n_majority7_module_20__and_module_4_res,
         n_majority7_module_20__or_module_3_res,
         n_majority7_module_20__and_module_3_res,
         n_majority7_module_20__or_module_2_res,
         n_majority7_module_20__and_module_2_res,
         n_majority7_module_20__or_module_1_res,
         n_majority7_module_20__and_module_1_res, n_majority7_module_21_n7,
         n_majority7_module_21_n6, n_majority7_module_21_n5,
         n_majority7_module_21_n4, n_majority7_module_21_n3,
         n_majority7_module_21_n2, n_majority7_module_21_n1,
         n_majority7_module_21__and_module_10_res,
         n_majority7_module_21__or_module_11_res,
         n_majority7_module_21__and_module_9_res,
         n_majority7_module_21__or_module_10_res,
         n_majority7_module_21__or_module_9_res,
         n_majority7_module_21__and_module_8_res,
         n_majority7_module_21__or_module_8_res,
         n_majority7_module_21__and_module_7_res,
         n_majority7_module_21__or_module_7_res,
         n_majority7_module_21__or_module_6_res,
         n_majority7_module_21__and_module_6_res,
         n_majority7_module_21__or_module_5_res,
         n_majority7_module_21__and_module_5_res,
         n_majority7_module_21__or_module_4_res,
         n_majority7_module_21__and_module_4_res,
         n_majority7_module_21__or_module_3_res,
         n_majority7_module_21__and_module_3_res,
         n_majority7_module_21__or_module_2_res,
         n_majority7_module_21__and_module_2_res,
         n_majority7_module_21__or_module_1_res,
         n_majority7_module_21__and_module_1_res, n_majority7_module_22_n7,
         n_majority7_module_22_n6, n_majority7_module_22_n5,
         n_majority7_module_22_n4, n_majority7_module_22_n3,
         n_majority7_module_22_n2, n_majority7_module_22_n1,
         n_majority7_module_22__and_module_10_res,
         n_majority7_module_22__or_module_11_res,
         n_majority7_module_22__and_module_9_res,
         n_majority7_module_22__or_module_10_res,
         n_majority7_module_22__or_module_9_res,
         n_majority7_module_22__and_module_8_res,
         n_majority7_module_22__or_module_8_res,
         n_majority7_module_22__and_module_7_res,
         n_majority7_module_22__or_module_7_res,
         n_majority7_module_22__or_module_6_res,
         n_majority7_module_22__and_module_6_res,
         n_majority7_module_22__or_module_5_res,
         n_majority7_module_22__and_module_5_res,
         n_majority7_module_22__or_module_4_res,
         n_majority7_module_22__and_module_4_res,
         n_majority7_module_22__or_module_3_res,
         n_majority7_module_22__and_module_3_res,
         n_majority7_module_22__or_module_2_res,
         n_majority7_module_22__and_module_2_res,
         n_majority7_module_22__or_module_1_res,
         n_majority7_module_22__and_module_1_res, n_majority7_module_23_n7,
         n_majority7_module_23_n6, n_majority7_module_23_n5,
         n_majority7_module_23_n4, n_majority7_module_23_n3,
         n_majority7_module_23_n2, n_majority7_module_23_n1,
         n_majority7_module_23__and_module_10_res,
         n_majority7_module_23__or_module_11_res,
         n_majority7_module_23__and_module_9_res,
         n_majority7_module_23__or_module_10_res,
         n_majority7_module_23__or_module_9_res,
         n_majority7_module_23__and_module_8_res,
         n_majority7_module_23__or_module_8_res,
         n_majority7_module_23__and_module_7_res,
         n_majority7_module_23__or_module_7_res,
         n_majority7_module_23__or_module_6_res,
         n_majority7_module_23__and_module_6_res,
         n_majority7_module_23__or_module_5_res,
         n_majority7_module_23__and_module_5_res,
         n_majority7_module_23__or_module_4_res,
         n_majority7_module_23__and_module_4_res,
         n_majority7_module_23__or_module_3_res,
         n_majority7_module_23__and_module_3_res,
         n_majority7_module_23__or_module_2_res,
         n_majority7_module_23__and_module_2_res,
         n_majority7_module_23__or_module_1_res,
         n_majority7_module_23__and_module_1_res, n_majority7_module_24_n7,
         n_majority7_module_24_n6, n_majority7_module_24_n5,
         n_majority7_module_24_n4, n_majority7_module_24_n3,
         n_majority7_module_24_n2, n_majority7_module_24_n1,
         n_majority7_module_24__and_module_10_res,
         n_majority7_module_24__or_module_11_res,
         n_majority7_module_24__and_module_9_res,
         n_majority7_module_24__or_module_10_res,
         n_majority7_module_24__or_module_9_res,
         n_majority7_module_24__and_module_8_res,
         n_majority7_module_24__or_module_8_res,
         n_majority7_module_24__and_module_7_res,
         n_majority7_module_24__or_module_7_res,
         n_majority7_module_24__or_module_6_res,
         n_majority7_module_24__and_module_6_res,
         n_majority7_module_24__or_module_5_res,
         n_majority7_module_24__and_module_5_res,
         n_majority7_module_24__or_module_4_res,
         n_majority7_module_24__and_module_4_res,
         n_majority7_module_24__or_module_3_res,
         n_majority7_module_24__and_module_3_res,
         n_majority7_module_24__or_module_2_res,
         n_majority7_module_24__and_module_2_res,
         n_majority7_module_24__or_module_1_res,
         n_majority7_module_24__and_module_1_res, n_majority7_module_25_n7,
         n_majority7_module_25_n6, n_majority7_module_25_n5,
         n_majority7_module_25_n4, n_majority7_module_25_n3,
         n_majority7_module_25_n2, n_majority7_module_25_n1,
         n_majority7_module_25__and_module_10_res,
         n_majority7_module_25__or_module_11_res,
         n_majority7_module_25__and_module_9_res,
         n_majority7_module_25__or_module_10_res,
         n_majority7_module_25__or_module_9_res,
         n_majority7_module_25__and_module_8_res,
         n_majority7_module_25__or_module_8_res,
         n_majority7_module_25__and_module_7_res,
         n_majority7_module_25__or_module_7_res,
         n_majority7_module_25__or_module_6_res,
         n_majority7_module_25__and_module_6_res,
         n_majority7_module_25__or_module_5_res,
         n_majority7_module_25__and_module_5_res,
         n_majority7_module_25__or_module_4_res,
         n_majority7_module_25__and_module_4_res,
         n_majority7_module_25__or_module_3_res,
         n_majority7_module_25__and_module_3_res,
         n_majority7_module_25__or_module_2_res,
         n_majority7_module_25__and_module_2_res,
         n_majority7_module_25__or_module_1_res,
         n_majority7_module_25__and_module_1_res, n_majority7_module_26_n7,
         n_majority7_module_26_n6, n_majority7_module_26_n5,
         n_majority7_module_26_n4, n_majority7_module_26_n3,
         n_majority7_module_26_n2, n_majority7_module_26_n1,
         n_majority7_module_26__and_module_10_res,
         n_majority7_module_26__or_module_11_res,
         n_majority7_module_26__and_module_9_res,
         n_majority7_module_26__or_module_10_res,
         n_majority7_module_26__or_module_9_res,
         n_majority7_module_26__and_module_8_res,
         n_majority7_module_26__or_module_8_res,
         n_majority7_module_26__and_module_7_res,
         n_majority7_module_26__or_module_7_res,
         n_majority7_module_26__or_module_6_res,
         n_majority7_module_26__and_module_6_res,
         n_majority7_module_26__or_module_5_res,
         n_majority7_module_26__and_module_5_res,
         n_majority7_module_26__or_module_4_res,
         n_majority7_module_26__and_module_4_res,
         n_majority7_module_26__or_module_3_res,
         n_majority7_module_26__and_module_3_res,
         n_majority7_module_26__or_module_2_res,
         n_majority7_module_26__and_module_2_res,
         n_majority7_module_26__or_module_1_res,
         n_majority7_module_26__and_module_1_res, n_majority7_module_27_n7,
         n_majority7_module_27_n6, n_majority7_module_27_n5,
         n_majority7_module_27_n4, n_majority7_module_27_n3,
         n_majority7_module_27_n2, n_majority7_module_27_n1,
         n_majority7_module_27__and_module_10_res,
         n_majority7_module_27__or_module_11_res,
         n_majority7_module_27__and_module_9_res,
         n_majority7_module_27__or_module_10_res,
         n_majority7_module_27__or_module_9_res,
         n_majority7_module_27__and_module_8_res,
         n_majority7_module_27__or_module_8_res,
         n_majority7_module_27__and_module_7_res,
         n_majority7_module_27__or_module_7_res,
         n_majority7_module_27__or_module_6_res,
         n_majority7_module_27__and_module_6_res,
         n_majority7_module_27__or_module_5_res,
         n_majority7_module_27__and_module_5_res,
         n_majority7_module_27__or_module_4_res,
         n_majority7_module_27__and_module_4_res,
         n_majority7_module_27__or_module_3_res,
         n_majority7_module_27__and_module_3_res,
         n_majority7_module_27__or_module_2_res,
         n_majority7_module_27__and_module_2_res,
         n_majority7_module_27__or_module_1_res,
         n_majority7_module_27__and_module_1_res, n_majority7_module_28_n7,
         n_majority7_module_28_n6, n_majority7_module_28_n5,
         n_majority7_module_28_n4, n_majority7_module_28_n3,
         n_majority7_module_28_n2, n_majority7_module_28_n1,
         n_majority7_module_28__and_module_10_res,
         n_majority7_module_28__or_module_11_res,
         n_majority7_module_28__and_module_9_res,
         n_majority7_module_28__or_module_10_res,
         n_majority7_module_28__or_module_9_res,
         n_majority7_module_28__and_module_8_res,
         n_majority7_module_28__or_module_8_res,
         n_majority7_module_28__and_module_7_res,
         n_majority7_module_28__or_module_7_res,
         n_majority7_module_28__or_module_6_res,
         n_majority7_module_28__and_module_6_res,
         n_majority7_module_28__or_module_5_res,
         n_majority7_module_28__and_module_5_res,
         n_majority7_module_28__or_module_4_res,
         n_majority7_module_28__and_module_4_res,
         n_majority7_module_28__or_module_3_res,
         n_majority7_module_28__and_module_3_res,
         n_majority7_module_28__or_module_2_res,
         n_majority7_module_28__and_module_2_res,
         n_majority7_module_28__or_module_1_res,
         n_majority7_module_28__and_module_1_res, n_majority7_module_29_n7,
         n_majority7_module_29_n6, n_majority7_module_29_n5,
         n_majority7_module_29_n4, n_majority7_module_29_n3,
         n_majority7_module_29_n2, n_majority7_module_29_n1,
         n_majority7_module_29__and_module_10_res,
         n_majority7_module_29__or_module_11_res,
         n_majority7_module_29__and_module_9_res,
         n_majority7_module_29__or_module_10_res,
         n_majority7_module_29__or_module_9_res,
         n_majority7_module_29__and_module_8_res,
         n_majority7_module_29__or_module_8_res,
         n_majority7_module_29__and_module_7_res,
         n_majority7_module_29__or_module_7_res,
         n_majority7_module_29__or_module_6_res,
         n_majority7_module_29__and_module_6_res,
         n_majority7_module_29__or_module_5_res,
         n_majority7_module_29__and_module_5_res,
         n_majority7_module_29__or_module_4_res,
         n_majority7_module_29__and_module_4_res,
         n_majority7_module_29__or_module_3_res,
         n_majority7_module_29__and_module_3_res,
         n_majority7_module_29__or_module_2_res,
         n_majority7_module_29__and_module_2_res,
         n_majority7_module_29__or_module_1_res,
         n_majority7_module_29__and_module_1_res, n_majority7_module_30_n7,
         n_majority7_module_30_n6, n_majority7_module_30_n5,
         n_majority7_module_30_n4, n_majority7_module_30_n3,
         n_majority7_module_30_n2, n_majority7_module_30_n1,
         n_majority7_module_30__and_module_10_res,
         n_majority7_module_30__or_module_11_res,
         n_majority7_module_30__and_module_9_res,
         n_majority7_module_30__or_module_10_res,
         n_majority7_module_30__or_module_9_res,
         n_majority7_module_30__and_module_8_res,
         n_majority7_module_30__or_module_8_res,
         n_majority7_module_30__and_module_7_res,
         n_majority7_module_30__or_module_7_res,
         n_majority7_module_30__or_module_6_res,
         n_majority7_module_30__and_module_6_res,
         n_majority7_module_30__or_module_5_res,
         n_majority7_module_30__and_module_5_res,
         n_majority7_module_30__or_module_4_res,
         n_majority7_module_30__and_module_4_res,
         n_majority7_module_30__or_module_3_res,
         n_majority7_module_30__and_module_3_res,
         n_majority7_module_30__or_module_2_res,
         n_majority7_module_30__and_module_2_res,
         n_majority7_module_30__or_module_1_res,
         n_majority7_module_30__and_module_1_res, n_majority7_module_31_n7,
         n_majority7_module_31_n6, n_majority7_module_31_n5,
         n_majority7_module_31_n4, n_majority7_module_31_n3,
         n_majority7_module_31_n2, n_majority7_module_31_n1,
         n_majority7_module_31__and_module_10_res,
         n_majority7_module_31__or_module_11_res,
         n_majority7_module_31__and_module_9_res,
         n_majority7_module_31__or_module_10_res,
         n_majority7_module_31__or_module_9_res,
         n_majority7_module_31__and_module_8_res,
         n_majority7_module_31__or_module_8_res,
         n_majority7_module_31__and_module_7_res,
         n_majority7_module_31__or_module_7_res,
         n_majority7_module_31__or_module_6_res,
         n_majority7_module_31__and_module_6_res,
         n_majority7_module_31__or_module_5_res,
         n_majority7_module_31__and_module_5_res,
         n_majority7_module_31__or_module_4_res,
         n_majority7_module_31__and_module_4_res,
         n_majority7_module_31__or_module_3_res,
         n_majority7_module_31__and_module_3_res,
         n_majority7_module_31__or_module_2_res,
         n_majority7_module_31__and_module_2_res,
         n_majority7_module_31__or_module_1_res,
         n_majority7_module_31__and_module_1_res, n_majority7_module_32_n7,
         n_majority7_module_32_n6, n_majority7_module_32_n5,
         n_majority7_module_32_n4, n_majority7_module_32_n3,
         n_majority7_module_32_n2, n_majority7_module_32_n1,
         n_majority7_module_32__and_module_10_res,
         n_majority7_module_32__or_module_11_res,
         n_majority7_module_32__and_module_9_res,
         n_majority7_module_32__or_module_10_res,
         n_majority7_module_32__or_module_9_res,
         n_majority7_module_32__and_module_8_res,
         n_majority7_module_32__or_module_8_res,
         n_majority7_module_32__and_module_7_res,
         n_majority7_module_32__or_module_7_res,
         n_majority7_module_32__or_module_6_res,
         n_majority7_module_32__and_module_6_res,
         n_majority7_module_32__or_module_5_res,
         n_majority7_module_32__and_module_5_res,
         n_majority7_module_32__or_module_4_res,
         n_majority7_module_32__and_module_4_res,
         n_majority7_module_32__or_module_3_res,
         n_majority7_module_32__and_module_3_res,
         n_majority7_module_32__or_module_2_res,
         n_majority7_module_32__and_module_2_res,
         n_majority7_module_32__or_module_1_res,
         n_majority7_module_32__and_module_1_res, n_majority7_module_33_n7,
         n_majority7_module_33_n6, n_majority7_module_33_n5,
         n_majority7_module_33_n4, n_majority7_module_33_n3,
         n_majority7_module_33_n2, n_majority7_module_33_n1,
         n_majority7_module_33__and_module_10_res,
         n_majority7_module_33__or_module_11_res,
         n_majority7_module_33__and_module_9_res,
         n_majority7_module_33__or_module_10_res,
         n_majority7_module_33__or_module_9_res,
         n_majority7_module_33__and_module_8_res,
         n_majority7_module_33__or_module_8_res,
         n_majority7_module_33__and_module_7_res,
         n_majority7_module_33__or_module_7_res,
         n_majority7_module_33__or_module_6_res,
         n_majority7_module_33__and_module_6_res,
         n_majority7_module_33__or_module_5_res,
         n_majority7_module_33__and_module_5_res,
         n_majority7_module_33__or_module_4_res,
         n_majority7_module_33__and_module_4_res,
         n_majority7_module_33__or_module_3_res,
         n_majority7_module_33__and_module_3_res,
         n_majority7_module_33__or_module_2_res,
         n_majority7_module_33__and_module_2_res,
         n_majority7_module_33__or_module_1_res,
         n_majority7_module_33__and_module_1_res, n_majority7_module_34_n7,
         n_majority7_module_34_n6, n_majority7_module_34_n5,
         n_majority7_module_34_n4, n_majority7_module_34_n3,
         n_majority7_module_34_n2, n_majority7_module_34_n1,
         n_majority7_module_34__and_module_10_res,
         n_majority7_module_34__or_module_11_res,
         n_majority7_module_34__and_module_9_res,
         n_majority7_module_34__or_module_10_res,
         n_majority7_module_34__or_module_9_res,
         n_majority7_module_34__and_module_8_res,
         n_majority7_module_34__or_module_8_res,
         n_majority7_module_34__and_module_7_res,
         n_majority7_module_34__or_module_7_res,
         n_majority7_module_34__or_module_6_res,
         n_majority7_module_34__and_module_6_res,
         n_majority7_module_34__or_module_5_res,
         n_majority7_module_34__and_module_5_res,
         n_majority7_module_34__or_module_4_res,
         n_majority7_module_34__and_module_4_res,
         n_majority7_module_34__or_module_3_res,
         n_majority7_module_34__and_module_3_res,
         n_majority7_module_34__or_module_2_res,
         n_majority7_module_34__and_module_2_res,
         n_majority7_module_34__or_module_1_res,
         n_majority7_module_34__and_module_1_res, n_majority7_module_35_n7,
         n_majority7_module_35_n6, n_majority7_module_35_n5,
         n_majority7_module_35_n4, n_majority7_module_35_n3,
         n_majority7_module_35_n2, n_majority7_module_35_n1,
         n_majority7_module_35__and_module_10_res,
         n_majority7_module_35__or_module_11_res,
         n_majority7_module_35__and_module_9_res,
         n_majority7_module_35__or_module_10_res,
         n_majority7_module_35__or_module_9_res,
         n_majority7_module_35__and_module_8_res,
         n_majority7_module_35__or_module_8_res,
         n_majority7_module_35__and_module_7_res,
         n_majority7_module_35__or_module_7_res,
         n_majority7_module_35__or_module_6_res,
         n_majority7_module_35__and_module_6_res,
         n_majority7_module_35__or_module_5_res,
         n_majority7_module_35__and_module_5_res,
         n_majority7_module_35__or_module_4_res,
         n_majority7_module_35__and_module_4_res,
         n_majority7_module_35__or_module_3_res,
         n_majority7_module_35__and_module_3_res,
         n_majority7_module_35__or_module_2_res,
         n_majority7_module_35__and_module_2_res,
         n_majority7_module_35__or_module_1_res,
         n_majority7_module_35__and_module_1_res, n_majority7_module_36_n7,
         n_majority7_module_36_n6, n_majority7_module_36_n5,
         n_majority7_module_36_n4, n_majority7_module_36_n3,
         n_majority7_module_36_n2, n_majority7_module_36_n1,
         n_majority7_module_36__and_module_10_res,
         n_majority7_module_36__or_module_11_res,
         n_majority7_module_36__and_module_9_res,
         n_majority7_module_36__or_module_10_res,
         n_majority7_module_36__or_module_9_res,
         n_majority7_module_36__and_module_8_res,
         n_majority7_module_36__or_module_8_res,
         n_majority7_module_36__and_module_7_res,
         n_majority7_module_36__or_module_7_res,
         n_majority7_module_36__or_module_6_res,
         n_majority7_module_36__and_module_6_res,
         n_majority7_module_36__or_module_5_res,
         n_majority7_module_36__and_module_5_res,
         n_majority7_module_36__or_module_4_res,
         n_majority7_module_36__and_module_4_res,
         n_majority7_module_36__or_module_3_res,
         n_majority7_module_36__and_module_3_res,
         n_majority7_module_36__or_module_2_res,
         n_majority7_module_36__and_module_2_res,
         n_majority7_module_36__or_module_1_res,
         n_majority7_module_36__and_module_1_res, n_majority7_module_37_n7,
         n_majority7_module_37_n6, n_majority7_module_37_n5,
         n_majority7_module_37_n4, n_majority7_module_37_n3,
         n_majority7_module_37_n2, n_majority7_module_37_n1,
         n_majority7_module_37__and_module_10_res,
         n_majority7_module_37__or_module_11_res,
         n_majority7_module_37__and_module_9_res,
         n_majority7_module_37__or_module_10_res,
         n_majority7_module_37__or_module_9_res,
         n_majority7_module_37__and_module_8_res,
         n_majority7_module_37__or_module_8_res,
         n_majority7_module_37__and_module_7_res,
         n_majority7_module_37__or_module_7_res,
         n_majority7_module_37__or_module_6_res,
         n_majority7_module_37__and_module_6_res,
         n_majority7_module_37__or_module_5_res,
         n_majority7_module_37__and_module_5_res,
         n_majority7_module_37__or_module_4_res,
         n_majority7_module_37__and_module_4_res,
         n_majority7_module_37__or_module_3_res,
         n_majority7_module_37__and_module_3_res,
         n_majority7_module_37__or_module_2_res,
         n_majority7_module_37__and_module_2_res,
         n_majority7_module_37__or_module_1_res,
         n_majority7_module_37__and_module_1_res, n_majority7_module_38_n7,
         n_majority7_module_38_n6, n_majority7_module_38_n5,
         n_majority7_module_38_n4, n_majority7_module_38_n3,
         n_majority7_module_38_n2, n_majority7_module_38_n1,
         n_majority7_module_38__and_module_10_res,
         n_majority7_module_38__or_module_11_res,
         n_majority7_module_38__and_module_9_res,
         n_majority7_module_38__or_module_10_res,
         n_majority7_module_38__or_module_9_res,
         n_majority7_module_38__and_module_8_res,
         n_majority7_module_38__or_module_8_res,
         n_majority7_module_38__and_module_7_res,
         n_majority7_module_38__or_module_7_res,
         n_majority7_module_38__or_module_6_res,
         n_majority7_module_38__and_module_6_res,
         n_majority7_module_38__or_module_5_res,
         n_majority7_module_38__and_module_5_res,
         n_majority7_module_38__or_module_4_res,
         n_majority7_module_38__and_module_4_res,
         n_majority7_module_38__or_module_3_res,
         n_majority7_module_38__and_module_3_res,
         n_majority7_module_38__or_module_2_res,
         n_majority7_module_38__and_module_2_res,
         n_majority7_module_38__or_module_1_res,
         n_majority7_module_38__and_module_1_res, n_majority7_module_39_n7,
         n_majority7_module_39_n6, n_majority7_module_39_n5,
         n_majority7_module_39_n4, n_majority7_module_39_n3,
         n_majority7_module_39_n2, n_majority7_module_39_n1,
         n_majority7_module_39__and_module_10_res,
         n_majority7_module_39__or_module_11_res,
         n_majority7_module_39__and_module_9_res,
         n_majority7_module_39__or_module_10_res,
         n_majority7_module_39__or_module_9_res,
         n_majority7_module_39__and_module_8_res,
         n_majority7_module_39__or_module_8_res,
         n_majority7_module_39__and_module_7_res,
         n_majority7_module_39__or_module_7_res,
         n_majority7_module_39__or_module_6_res,
         n_majority7_module_39__and_module_6_res,
         n_majority7_module_39__or_module_5_res,
         n_majority7_module_39__and_module_5_res,
         n_majority7_module_39__or_module_4_res,
         n_majority7_module_39__and_module_4_res,
         n_majority7_module_39__or_module_3_res,
         n_majority7_module_39__and_module_3_res,
         n_majority7_module_39__or_module_2_res,
         n_majority7_module_39__and_module_2_res,
         n_majority7_module_39__or_module_1_res,
         n_majority7_module_39__and_module_1_res, n_majority7_module_40_n7,
         n_majority7_module_40_n6, n_majority7_module_40_n5,
         n_majority7_module_40_n4, n_majority7_module_40_n3,
         n_majority7_module_40_n2, n_majority7_module_40_n1,
         n_majority7_module_40__and_module_10_res,
         n_majority7_module_40__or_module_11_res,
         n_majority7_module_40__and_module_9_res,
         n_majority7_module_40__or_module_10_res,
         n_majority7_module_40__or_module_9_res,
         n_majority7_module_40__and_module_8_res,
         n_majority7_module_40__or_module_8_res,
         n_majority7_module_40__and_module_7_res,
         n_majority7_module_40__or_module_7_res,
         n_majority7_module_40__or_module_6_res,
         n_majority7_module_40__and_module_6_res,
         n_majority7_module_40__or_module_5_res,
         n_majority7_module_40__and_module_5_res,
         n_majority7_module_40__or_module_4_res,
         n_majority7_module_40__and_module_4_res,
         n_majority7_module_40__or_module_3_res,
         n_majority7_module_40__and_module_3_res,
         n_majority7_module_40__or_module_2_res,
         n_majority7_module_40__and_module_2_res,
         n_majority7_module_40__or_module_1_res,
         n_majority7_module_40__and_module_1_res, n_majority7_module_41_n7,
         n_majority7_module_41_n6, n_majority7_module_41_n5,
         n_majority7_module_41_n4, n_majority7_module_41_n3,
         n_majority7_module_41_n2, n_majority7_module_41_n1,
         n_majority7_module_41__and_module_10_res,
         n_majority7_module_41__or_module_11_res,
         n_majority7_module_41__and_module_9_res,
         n_majority7_module_41__or_module_10_res,
         n_majority7_module_41__or_module_9_res,
         n_majority7_module_41__and_module_8_res,
         n_majority7_module_41__or_module_8_res,
         n_majority7_module_41__and_module_7_res,
         n_majority7_module_41__or_module_7_res,
         n_majority7_module_41__or_module_6_res,
         n_majority7_module_41__and_module_6_res,
         n_majority7_module_41__or_module_5_res,
         n_majority7_module_41__and_module_5_res,
         n_majority7_module_41__or_module_4_res,
         n_majority7_module_41__and_module_4_res,
         n_majority7_module_41__or_module_3_res,
         n_majority7_module_41__and_module_3_res,
         n_majority7_module_41__or_module_2_res,
         n_majority7_module_41__and_module_2_res,
         n_majority7_module_41__or_module_1_res,
         n_majority7_module_41__and_module_1_res, n_majority7_module_42_n7,
         n_majority7_module_42_n6, n_majority7_module_42_n5,
         n_majority7_module_42_n4, n_majority7_module_42_n3,
         n_majority7_module_42_n2, n_majority7_module_42_n1,
         n_majority7_module_42__and_module_10_res,
         n_majority7_module_42__or_module_11_res,
         n_majority7_module_42__and_module_9_res,
         n_majority7_module_42__or_module_10_res,
         n_majority7_module_42__or_module_9_res,
         n_majority7_module_42__and_module_8_res,
         n_majority7_module_42__or_module_8_res,
         n_majority7_module_42__and_module_7_res,
         n_majority7_module_42__or_module_7_res,
         n_majority7_module_42__or_module_6_res,
         n_majority7_module_42__and_module_6_res,
         n_majority7_module_42__or_module_5_res,
         n_majority7_module_42__and_module_5_res,
         n_majority7_module_42__or_module_4_res,
         n_majority7_module_42__and_module_4_res,
         n_majority7_module_42__or_module_3_res,
         n_majority7_module_42__and_module_3_res,
         n_majority7_module_42__or_module_2_res,
         n_majority7_module_42__and_module_2_res,
         n_majority7_module_42__or_module_1_res,
         n_majority7_module_42__and_module_1_res, n_majority7_module_43_n7,
         n_majority7_module_43_n6, n_majority7_module_43_n5,
         n_majority7_module_43_n4, n_majority7_module_43_n3,
         n_majority7_module_43_n2, n_majority7_module_43_n1,
         n_majority7_module_43__and_module_10_res,
         n_majority7_module_43__or_module_11_res,
         n_majority7_module_43__and_module_9_res,
         n_majority7_module_43__or_module_10_res,
         n_majority7_module_43__or_module_9_res,
         n_majority7_module_43__and_module_8_res,
         n_majority7_module_43__or_module_8_res,
         n_majority7_module_43__and_module_7_res,
         n_majority7_module_43__or_module_7_res,
         n_majority7_module_43__or_module_6_res,
         n_majority7_module_43__and_module_6_res,
         n_majority7_module_43__or_module_5_res,
         n_majority7_module_43__and_module_5_res,
         n_majority7_module_43__or_module_4_res,
         n_majority7_module_43__and_module_4_res,
         n_majority7_module_43__or_module_3_res,
         n_majority7_module_43__and_module_3_res,
         n_majority7_module_43__or_module_2_res,
         n_majority7_module_43__and_module_2_res,
         n_majority7_module_43__or_module_1_res,
         n_majority7_module_43__and_module_1_res, n_majority7_module_44_n7,
         n_majority7_module_44_n6, n_majority7_module_44_n5,
         n_majority7_module_44_n4, n_majority7_module_44_n3,
         n_majority7_module_44_n2, n_majority7_module_44_n1,
         n_majority7_module_44__and_module_10_res,
         n_majority7_module_44__or_module_11_res,
         n_majority7_module_44__and_module_9_res,
         n_majority7_module_44__or_module_10_res,
         n_majority7_module_44__or_module_9_res,
         n_majority7_module_44__and_module_8_res,
         n_majority7_module_44__or_module_8_res,
         n_majority7_module_44__and_module_7_res,
         n_majority7_module_44__or_module_7_res,
         n_majority7_module_44__or_module_6_res,
         n_majority7_module_44__and_module_6_res,
         n_majority7_module_44__or_module_5_res,
         n_majority7_module_44__and_module_5_res,
         n_majority7_module_44__or_module_4_res,
         n_majority7_module_44__and_module_4_res,
         n_majority7_module_44__or_module_3_res,
         n_majority7_module_44__and_module_3_res,
         n_majority7_module_44__or_module_2_res,
         n_majority7_module_44__and_module_2_res,
         n_majority7_module_44__or_module_1_res,
         n_majority7_module_44__and_module_1_res, n_majority7_module_45_n7,
         n_majority7_module_45_n6, n_majority7_module_45_n5,
         n_majority7_module_45_n4, n_majority7_module_45_n3,
         n_majority7_module_45_n2, n_majority7_module_45_n1,
         n_majority7_module_45__and_module_10_res,
         n_majority7_module_45__or_module_11_res,
         n_majority7_module_45__and_module_9_res,
         n_majority7_module_45__or_module_10_res,
         n_majority7_module_45__or_module_9_res,
         n_majority7_module_45__and_module_8_res,
         n_majority7_module_45__or_module_8_res,
         n_majority7_module_45__and_module_7_res,
         n_majority7_module_45__or_module_7_res,
         n_majority7_module_45__or_module_6_res,
         n_majority7_module_45__and_module_6_res,
         n_majority7_module_45__or_module_5_res,
         n_majority7_module_45__and_module_5_res,
         n_majority7_module_45__or_module_4_res,
         n_majority7_module_45__and_module_4_res,
         n_majority7_module_45__or_module_3_res,
         n_majority7_module_45__and_module_3_res,
         n_majority7_module_45__or_module_2_res,
         n_majority7_module_45__and_module_2_res,
         n_majority7_module_45__or_module_1_res,
         n_majority7_module_45__and_module_1_res, n_majority7_module_46_n7,
         n_majority7_module_46_n6, n_majority7_module_46_n5,
         n_majority7_module_46_n4, n_majority7_module_46_n3,
         n_majority7_module_46_n2, n_majority7_module_46_n1,
         n_majority7_module_46__and_module_10_res,
         n_majority7_module_46__or_module_11_res,
         n_majority7_module_46__and_module_9_res,
         n_majority7_module_46__or_module_10_res,
         n_majority7_module_46__or_module_9_res,
         n_majority7_module_46__and_module_8_res,
         n_majority7_module_46__or_module_8_res,
         n_majority7_module_46__and_module_7_res,
         n_majority7_module_46__or_module_7_res,
         n_majority7_module_46__or_module_6_res,
         n_majority7_module_46__and_module_6_res,
         n_majority7_module_46__or_module_5_res,
         n_majority7_module_46__and_module_5_res,
         n_majority7_module_46__or_module_4_res,
         n_majority7_module_46__and_module_4_res,
         n_majority7_module_46__or_module_3_res,
         n_majority7_module_46__and_module_3_res,
         n_majority7_module_46__or_module_2_res,
         n_majority7_module_46__and_module_2_res,
         n_majority7_module_46__or_module_1_res,
         n_majority7_module_46__and_module_1_res, n_majority7_module_47_n7,
         n_majority7_module_47_n6, n_majority7_module_47_n5,
         n_majority7_module_47_n4, n_majority7_module_47_n3,
         n_majority7_module_47_n2, n_majority7_module_47_n1,
         n_majority7_module_47__and_module_10_res,
         n_majority7_module_47__or_module_11_res,
         n_majority7_module_47__and_module_9_res,
         n_majority7_module_47__or_module_10_res,
         n_majority7_module_47__or_module_9_res,
         n_majority7_module_47__and_module_8_res,
         n_majority7_module_47__or_module_8_res,
         n_majority7_module_47__and_module_7_res,
         n_majority7_module_47__or_module_7_res,
         n_majority7_module_47__or_module_6_res,
         n_majority7_module_47__and_module_6_res,
         n_majority7_module_47__or_module_5_res,
         n_majority7_module_47__and_module_5_res,
         n_majority7_module_47__or_module_4_res,
         n_majority7_module_47__and_module_4_res,
         n_majority7_module_47__or_module_3_res,
         n_majority7_module_47__and_module_3_res,
         n_majority7_module_47__or_module_2_res,
         n_majority7_module_47__and_module_2_res,
         n_majority7_module_47__or_module_1_res,
         n_majority7_module_47__and_module_1_res, n_majority7_module_48_n7,
         n_majority7_module_48_n6, n_majority7_module_48_n5,
         n_majority7_module_48_n4, n_majority7_module_48_n3,
         n_majority7_module_48_n2, n_majority7_module_48_n1,
         n_majority7_module_48__and_module_10_res,
         n_majority7_module_48__or_module_11_res,
         n_majority7_module_48__and_module_9_res,
         n_majority7_module_48__or_module_10_res,
         n_majority7_module_48__or_module_9_res,
         n_majority7_module_48__and_module_8_res,
         n_majority7_module_48__or_module_8_res,
         n_majority7_module_48__and_module_7_res,
         n_majority7_module_48__or_module_7_res,
         n_majority7_module_48__or_module_6_res,
         n_majority7_module_48__and_module_6_res,
         n_majority7_module_48__or_module_5_res,
         n_majority7_module_48__and_module_5_res,
         n_majority7_module_48__or_module_4_res,
         n_majority7_module_48__and_module_4_res,
         n_majority7_module_48__or_module_3_res,
         n_majority7_module_48__and_module_3_res,
         n_majority7_module_48__or_module_2_res,
         n_majority7_module_48__and_module_2_res,
         n_majority7_module_48__or_module_1_res,
         n_majority7_module_48__and_module_1_res, n_majority7_module_49_n7,
         n_majority7_module_49_n6, n_majority7_module_49_n5,
         n_majority7_module_49_n4, n_majority7_module_49_n3,
         n_majority7_module_49_n2, n_majority7_module_49_n1,
         n_majority7_module_49__and_module_10_res,
         n_majority7_module_49__or_module_11_res,
         n_majority7_module_49__and_module_9_res,
         n_majority7_module_49__or_module_10_res,
         n_majority7_module_49__or_module_9_res,
         n_majority7_module_49__and_module_8_res,
         n_majority7_module_49__or_module_8_res,
         n_majority7_module_49__and_module_7_res,
         n_majority7_module_49__or_module_7_res,
         n_majority7_module_49__or_module_6_res,
         n_majority7_module_49__and_module_6_res,
         n_majority7_module_49__or_module_5_res,
         n_majority7_module_49__and_module_5_res,
         n_majority7_module_49__or_module_4_res,
         n_majority7_module_49__and_module_4_res,
         n_majority7_module_49__or_module_3_res,
         n_majority7_module_49__and_module_3_res,
         n_majority7_module_49__or_module_2_res,
         n_majority7_module_49__and_module_2_res,
         n_majority7_module_49__or_module_1_res,
         n_majority7_module_49__and_module_1_res, n_majority7_module_50_n7,
         n_majority7_module_50_n6, n_majority7_module_50_n5,
         n_majority7_module_50_n4, n_majority7_module_50_n3,
         n_majority7_module_50_n2, n_majority7_module_50_n1,
         n_majority7_module_50__and_module_10_res,
         n_majority7_module_50__or_module_11_res,
         n_majority7_module_50__and_module_9_res,
         n_majority7_module_50__or_module_10_res,
         n_majority7_module_50__or_module_9_res,
         n_majority7_module_50__and_module_8_res,
         n_majority7_module_50__or_module_8_res,
         n_majority7_module_50__and_module_7_res,
         n_majority7_module_50__or_module_7_res,
         n_majority7_module_50__or_module_6_res,
         n_majority7_module_50__and_module_6_res,
         n_majority7_module_50__or_module_5_res,
         n_majority7_module_50__and_module_5_res,
         n_majority7_module_50__or_module_4_res,
         n_majority7_module_50__and_module_4_res,
         n_majority7_module_50__or_module_3_res,
         n_majority7_module_50__and_module_3_res,
         n_majority7_module_50__or_module_2_res,
         n_majority7_module_50__and_module_2_res,
         n_majority7_module_50__or_module_1_res,
         n_majority7_module_50__and_module_1_res, n_majority7_module_51_n7,
         n_majority7_module_51_n6, n_majority7_module_51_n5,
         n_majority7_module_51_n4, n_majority7_module_51_n3,
         n_majority7_module_51_n2, n_majority7_module_51_n1,
         n_majority7_module_51__and_module_10_res,
         n_majority7_module_51__or_module_11_res,
         n_majority7_module_51__and_module_9_res,
         n_majority7_module_51__or_module_10_res,
         n_majority7_module_51__or_module_9_res,
         n_majority7_module_51__and_module_8_res,
         n_majority7_module_51__or_module_8_res,
         n_majority7_module_51__and_module_7_res,
         n_majority7_module_51__or_module_7_res,
         n_majority7_module_51__or_module_6_res,
         n_majority7_module_51__and_module_6_res,
         n_majority7_module_51__or_module_5_res,
         n_majority7_module_51__and_module_5_res,
         n_majority7_module_51__or_module_4_res,
         n_majority7_module_51__and_module_4_res,
         n_majority7_module_51__or_module_3_res,
         n_majority7_module_51__and_module_3_res,
         n_majority7_module_51__or_module_2_res,
         n_majority7_module_51__and_module_2_res,
         n_majority7_module_51__or_module_1_res,
         n_majority7_module_51__and_module_1_res, n_majority7_module_52_n7,
         n_majority7_module_52_n6, n_majority7_module_52_n5,
         n_majority7_module_52_n4, n_majority7_module_52_n3,
         n_majority7_module_52_n2, n_majority7_module_52_n1,
         n_majority7_module_52__and_module_10_res,
         n_majority7_module_52__or_module_11_res,
         n_majority7_module_52__and_module_9_res,
         n_majority7_module_52__or_module_10_res,
         n_majority7_module_52__or_module_9_res,
         n_majority7_module_52__and_module_8_res,
         n_majority7_module_52__or_module_8_res,
         n_majority7_module_52__and_module_7_res,
         n_majority7_module_52__or_module_7_res,
         n_majority7_module_52__or_module_6_res,
         n_majority7_module_52__and_module_6_res,
         n_majority7_module_52__or_module_5_res,
         n_majority7_module_52__and_module_5_res,
         n_majority7_module_52__or_module_4_res,
         n_majority7_module_52__and_module_4_res,
         n_majority7_module_52__or_module_3_res,
         n_majority7_module_52__and_module_3_res,
         n_majority7_module_52__or_module_2_res,
         n_majority7_module_52__and_module_2_res,
         n_majority7_module_52__or_module_1_res,
         n_majority7_module_52__and_module_1_res, n_majority7_module_53_n7,
         n_majority7_module_53_n6, n_majority7_module_53_n5,
         n_majority7_module_53_n4, n_majority7_module_53_n3,
         n_majority7_module_53_n2, n_majority7_module_53_n1,
         n_majority7_module_53__and_module_10_res,
         n_majority7_module_53__or_module_11_res,
         n_majority7_module_53__and_module_9_res,
         n_majority7_module_53__or_module_10_res,
         n_majority7_module_53__or_module_9_res,
         n_majority7_module_53__and_module_8_res,
         n_majority7_module_53__or_module_8_res,
         n_majority7_module_53__and_module_7_res,
         n_majority7_module_53__or_module_7_res,
         n_majority7_module_53__or_module_6_res,
         n_majority7_module_53__and_module_6_res,
         n_majority7_module_53__or_module_5_res,
         n_majority7_module_53__and_module_5_res,
         n_majority7_module_53__or_module_4_res,
         n_majority7_module_53__and_module_4_res,
         n_majority7_module_53__or_module_3_res,
         n_majority7_module_53__and_module_3_res,
         n_majority7_module_53__or_module_2_res,
         n_majority7_module_53__and_module_2_res,
         n_majority7_module_53__or_module_1_res,
         n_majority7_module_53__and_module_1_res, n_majority7_module_54_n7,
         n_majority7_module_54_n6, n_majority7_module_54_n5,
         n_majority7_module_54_n4, n_majority7_module_54_n3,
         n_majority7_module_54_n2, n_majority7_module_54_n1,
         n_majority7_module_54__and_module_10_res,
         n_majority7_module_54__or_module_11_res,
         n_majority7_module_54__and_module_9_res,
         n_majority7_module_54__or_module_10_res,
         n_majority7_module_54__or_module_9_res,
         n_majority7_module_54__and_module_8_res,
         n_majority7_module_54__or_module_8_res,
         n_majority7_module_54__and_module_7_res,
         n_majority7_module_54__or_module_7_res,
         n_majority7_module_54__or_module_6_res,
         n_majority7_module_54__and_module_6_res,
         n_majority7_module_54__or_module_5_res,
         n_majority7_module_54__and_module_5_res,
         n_majority7_module_54__or_module_4_res,
         n_majority7_module_54__and_module_4_res,
         n_majority7_module_54__or_module_3_res,
         n_majority7_module_54__and_module_3_res,
         n_majority7_module_54__or_module_2_res,
         n_majority7_module_54__and_module_2_res,
         n_majority7_module_54__or_module_1_res,
         n_majority7_module_54__and_module_1_res, n_majority7_module_55_n7,
         n_majority7_module_55_n6, n_majority7_module_55_n5,
         n_majority7_module_55_n4, n_majority7_module_55_n3,
         n_majority7_module_55_n2, n_majority7_module_55_n1,
         n_majority7_module_55__and_module_10_res,
         n_majority7_module_55__or_module_11_res,
         n_majority7_module_55__and_module_9_res,
         n_majority7_module_55__or_module_10_res,
         n_majority7_module_55__or_module_9_res,
         n_majority7_module_55__and_module_8_res,
         n_majority7_module_55__or_module_8_res,
         n_majority7_module_55__and_module_7_res,
         n_majority7_module_55__or_module_7_res,
         n_majority7_module_55__or_module_6_res,
         n_majority7_module_55__and_module_6_res,
         n_majority7_module_55__or_module_5_res,
         n_majority7_module_55__and_module_5_res,
         n_majority7_module_55__or_module_4_res,
         n_majority7_module_55__and_module_4_res,
         n_majority7_module_55__or_module_3_res,
         n_majority7_module_55__and_module_3_res,
         n_majority7_module_55__or_module_2_res,
         n_majority7_module_55__and_module_2_res,
         n_majority7_module_55__or_module_1_res,
         n_majority7_module_55__and_module_1_res, n_majority7_module_56_n7,
         n_majority7_module_56_n6, n_majority7_module_56_n5,
         n_majority7_module_56_n4, n_majority7_module_56_n3,
         n_majority7_module_56_n2, n_majority7_module_56_n1,
         n_majority7_module_56__and_module_10_res,
         n_majority7_module_56__or_module_11_res,
         n_majority7_module_56__and_module_9_res,
         n_majority7_module_56__or_module_10_res,
         n_majority7_module_56__or_module_9_res,
         n_majority7_module_56__and_module_8_res,
         n_majority7_module_56__or_module_8_res,
         n_majority7_module_56__and_module_7_res,
         n_majority7_module_56__or_module_7_res,
         n_majority7_module_56__or_module_6_res,
         n_majority7_module_56__and_module_6_res,
         n_majority7_module_56__or_module_5_res,
         n_majority7_module_56__and_module_5_res,
         n_majority7_module_56__or_module_4_res,
         n_majority7_module_56__and_module_4_res,
         n_majority7_module_56__or_module_3_res,
         n_majority7_module_56__and_module_3_res,
         n_majority7_module_56__or_module_2_res,
         n_majority7_module_56__and_module_2_res,
         n_majority7_module_56__or_module_1_res,
         n_majority7_module_56__and_module_1_res, n_majority7_module_57_n7,
         n_majority7_module_57_n6, n_majority7_module_57_n5,
         n_majority7_module_57_n4, n_majority7_module_57_n3,
         n_majority7_module_57_n2, n_majority7_module_57_n1,
         n_majority7_module_57__and_module_10_res,
         n_majority7_module_57__or_module_11_res,
         n_majority7_module_57__and_module_9_res,
         n_majority7_module_57__or_module_10_res,
         n_majority7_module_57__or_module_9_res,
         n_majority7_module_57__and_module_8_res,
         n_majority7_module_57__or_module_8_res,
         n_majority7_module_57__and_module_7_res,
         n_majority7_module_57__or_module_7_res,
         n_majority7_module_57__or_module_6_res,
         n_majority7_module_57__and_module_6_res,
         n_majority7_module_57__or_module_5_res,
         n_majority7_module_57__and_module_5_res,
         n_majority7_module_57__or_module_4_res,
         n_majority7_module_57__and_module_4_res,
         n_majority7_module_57__or_module_3_res,
         n_majority7_module_57__and_module_3_res,
         n_majority7_module_57__or_module_2_res,
         n_majority7_module_57__and_module_2_res,
         n_majority7_module_57__or_module_1_res,
         n_majority7_module_57__and_module_1_res, n_majority7_module_58_n7,
         n_majority7_module_58_n6, n_majority7_module_58_n5,
         n_majority7_module_58_n4, n_majority7_module_58_n3,
         n_majority7_module_58_n2, n_majority7_module_58_n1,
         n_majority7_module_58__and_module_10_res,
         n_majority7_module_58__or_module_11_res,
         n_majority7_module_58__and_module_9_res,
         n_majority7_module_58__or_module_10_res,
         n_majority7_module_58__or_module_9_res,
         n_majority7_module_58__and_module_8_res,
         n_majority7_module_58__or_module_8_res,
         n_majority7_module_58__and_module_7_res,
         n_majority7_module_58__or_module_7_res,
         n_majority7_module_58__or_module_6_res,
         n_majority7_module_58__and_module_6_res,
         n_majority7_module_58__or_module_5_res,
         n_majority7_module_58__and_module_5_res,
         n_majority7_module_58__or_module_4_res,
         n_majority7_module_58__and_module_4_res,
         n_majority7_module_58__or_module_3_res,
         n_majority7_module_58__and_module_3_res,
         n_majority7_module_58__or_module_2_res,
         n_majority7_module_58__and_module_2_res,
         n_majority7_module_58__or_module_1_res,
         n_majority7_module_58__and_module_1_res, n_majority7_module_59_n7,
         n_majority7_module_59_n6, n_majority7_module_59_n5,
         n_majority7_module_59_n4, n_majority7_module_59_n3,
         n_majority7_module_59_n2, n_majority7_module_59_n1,
         n_majority7_module_59__and_module_10_res,
         n_majority7_module_59__or_module_11_res,
         n_majority7_module_59__and_module_9_res,
         n_majority7_module_59__or_module_10_res,
         n_majority7_module_59__or_module_9_res,
         n_majority7_module_59__and_module_8_res,
         n_majority7_module_59__or_module_8_res,
         n_majority7_module_59__and_module_7_res,
         n_majority7_module_59__or_module_7_res,
         n_majority7_module_59__or_module_6_res,
         n_majority7_module_59__and_module_6_res,
         n_majority7_module_59__or_module_5_res,
         n_majority7_module_59__and_module_5_res,
         n_majority7_module_59__or_module_4_res,
         n_majority7_module_59__and_module_4_res,
         n_majority7_module_59__or_module_3_res,
         n_majority7_module_59__and_module_3_res,
         n_majority7_module_59__or_module_2_res,
         n_majority7_module_59__and_module_2_res,
         n_majority7_module_59__or_module_1_res,
         n_majority7_module_59__and_module_1_res, n_majority7_module_60_n7,
         n_majority7_module_60_n6, n_majority7_module_60_n5,
         n_majority7_module_60_n4, n_majority7_module_60_n3,
         n_majority7_module_60_n2, n_majority7_module_60_n1,
         n_majority7_module_60__and_module_10_res,
         n_majority7_module_60__or_module_11_res,
         n_majority7_module_60__and_module_9_res,
         n_majority7_module_60__or_module_10_res,
         n_majority7_module_60__or_module_9_res,
         n_majority7_module_60__and_module_8_res,
         n_majority7_module_60__or_module_8_res,
         n_majority7_module_60__and_module_7_res,
         n_majority7_module_60__or_module_7_res,
         n_majority7_module_60__or_module_6_res,
         n_majority7_module_60__and_module_6_res,
         n_majority7_module_60__or_module_5_res,
         n_majority7_module_60__and_module_5_res,
         n_majority7_module_60__or_module_4_res,
         n_majority7_module_60__and_module_4_res,
         n_majority7_module_60__or_module_3_res,
         n_majority7_module_60__and_module_3_res,
         n_majority7_module_60__or_module_2_res,
         n_majority7_module_60__and_module_2_res,
         n_majority7_module_60__or_module_1_res,
         n_majority7_module_60__and_module_1_res, n_majority7_module_61_n7,
         n_majority7_module_61_n6, n_majority7_module_61_n5,
         n_majority7_module_61_n4, n_majority7_module_61_n3,
         n_majority7_module_61_n2, n_majority7_module_61_n1,
         n_majority7_module_61__and_module_10_res,
         n_majority7_module_61__or_module_11_res,
         n_majority7_module_61__and_module_9_res,
         n_majority7_module_61__or_module_10_res,
         n_majority7_module_61__or_module_9_res,
         n_majority7_module_61__and_module_8_res,
         n_majority7_module_61__or_module_8_res,
         n_majority7_module_61__and_module_7_res,
         n_majority7_module_61__or_module_7_res,
         n_majority7_module_61__or_module_6_res,
         n_majority7_module_61__and_module_6_res,
         n_majority7_module_61__or_module_5_res,
         n_majority7_module_61__and_module_5_res,
         n_majority7_module_61__or_module_4_res,
         n_majority7_module_61__and_module_4_res,
         n_majority7_module_61__or_module_3_res,
         n_majority7_module_61__and_module_3_res,
         n_majority7_module_61__or_module_2_res,
         n_majority7_module_61__and_module_2_res,
         n_majority7_module_61__or_module_1_res,
         n_majority7_module_61__and_module_1_res, n_majority7_module_62_n7,
         n_majority7_module_62_n6, n_majority7_module_62_n5,
         n_majority7_module_62_n4, n_majority7_module_62_n3,
         n_majority7_module_62_n2, n_majority7_module_62_n1,
         n_majority7_module_62__and_module_10_res,
         n_majority7_module_62__or_module_11_res,
         n_majority7_module_62__and_module_9_res,
         n_majority7_module_62__or_module_10_res,
         n_majority7_module_62__or_module_9_res,
         n_majority7_module_62__and_module_8_res,
         n_majority7_module_62__or_module_8_res,
         n_majority7_module_62__and_module_7_res,
         n_majority7_module_62__or_module_7_res,
         n_majority7_module_62__or_module_6_res,
         n_majority7_module_62__and_module_6_res,
         n_majority7_module_62__or_module_5_res,
         n_majority7_module_62__and_module_5_res,
         n_majority7_module_62__or_module_4_res,
         n_majority7_module_62__and_module_4_res,
         n_majority7_module_62__or_module_3_res,
         n_majority7_module_62__and_module_3_res,
         n_majority7_module_62__or_module_2_res,
         n_majority7_module_62__and_module_2_res,
         n_majority7_module_62__or_module_1_res,
         n_majority7_module_62__and_module_1_res, n_majority7_module_63_n7,
         n_majority7_module_63_n6, n_majority7_module_63_n5,
         n_majority7_module_63_n4, n_majority7_module_63_n3,
         n_majority7_module_63_n2, n_majority7_module_63_n1,
         n_majority7_module_63__and_module_10_res,
         n_majority7_module_63__or_module_11_res,
         n_majority7_module_63__and_module_9_res,
         n_majority7_module_63__or_module_10_res,
         n_majority7_module_63__or_module_9_res,
         n_majority7_module_63__and_module_8_res,
         n_majority7_module_63__or_module_8_res,
         n_majority7_module_63__and_module_7_res,
         n_majority7_module_63__or_module_7_res,
         n_majority7_module_63__or_module_6_res,
         n_majority7_module_63__and_module_6_res,
         n_majority7_module_63__or_module_5_res,
         n_majority7_module_63__and_module_5_res,
         n_majority7_module_63__or_module_4_res,
         n_majority7_module_63__and_module_4_res,
         n_majority7_module_63__or_module_3_res,
         n_majority7_module_63__and_module_3_res,
         n_majority7_module_63__or_module_2_res,
         n_majority7_module_63__and_module_2_res,
         n_majority7_module_63__or_module_1_res,
         n_majority7_module_63__and_module_1_res, n_majority7_module_64_n7,
         n_majority7_module_64_n6, n_majority7_module_64_n5,
         n_majority7_module_64_n4, n_majority7_module_64_n3,
         n_majority7_module_64_n2, n_majority7_module_64_n1,
         n_majority7_module_64__and_module_10_res,
         n_majority7_module_64__or_module_11_res,
         n_majority7_module_64__and_module_9_res,
         n_majority7_module_64__or_module_10_res,
         n_majority7_module_64__or_module_9_res,
         n_majority7_module_64__and_module_8_res,
         n_majority7_module_64__or_module_8_res,
         n_majority7_module_64__and_module_7_res,
         n_majority7_module_64__or_module_7_res,
         n_majority7_module_64__or_module_6_res,
         n_majority7_module_64__and_module_6_res,
         n_majority7_module_64__or_module_5_res,
         n_majority7_module_64__and_module_5_res,
         n_majority7_module_64__or_module_4_res,
         n_majority7_module_64__and_module_4_res,
         n_majority7_module_64__or_module_3_res,
         n_majority7_module_64__and_module_3_res,
         n_majority7_module_64__or_module_2_res,
         n_majority7_module_64__and_module_2_res,
         n_majority7_module_64__or_module_1_res,
         n_majority7_module_64__and_module_1_res, n_majority7_module_65_n7,
         n_majority7_module_65_n6, n_majority7_module_65_n5,
         n_majority7_module_65_n4, n_majority7_module_65_n3,
         n_majority7_module_65_n2, n_majority7_module_65_n1,
         n_majority7_module_65__and_module_10_res,
         n_majority7_module_65__or_module_11_res,
         n_majority7_module_65__and_module_9_res,
         n_majority7_module_65__or_module_10_res,
         n_majority7_module_65__or_module_9_res,
         n_majority7_module_65__and_module_8_res,
         n_majority7_module_65__or_module_8_res,
         n_majority7_module_65__and_module_7_res,
         n_majority7_module_65__or_module_7_res,
         n_majority7_module_65__or_module_6_res,
         n_majority7_module_65__and_module_6_res,
         n_majority7_module_65__or_module_5_res,
         n_majority7_module_65__and_module_5_res,
         n_majority7_module_65__or_module_4_res,
         n_majority7_module_65__and_module_4_res,
         n_majority7_module_65__or_module_3_res,
         n_majority7_module_65__and_module_3_res,
         n_majority7_module_65__or_module_2_res,
         n_majority7_module_65__and_module_2_res,
         n_majority7_module_65__or_module_1_res,
         n_majority7_module_65__and_module_1_res, n_majority7_module_66_n7,
         n_majority7_module_66_n6, n_majority7_module_66_n5,
         n_majority7_module_66_n4, n_majority7_module_66_n3,
         n_majority7_module_66_n2, n_majority7_module_66_n1,
         n_majority7_module_66__and_module_10_res,
         n_majority7_module_66__or_module_11_res,
         n_majority7_module_66__and_module_9_res,
         n_majority7_module_66__or_module_10_res,
         n_majority7_module_66__or_module_9_res,
         n_majority7_module_66__and_module_8_res,
         n_majority7_module_66__or_module_8_res,
         n_majority7_module_66__and_module_7_res,
         n_majority7_module_66__or_module_7_res,
         n_majority7_module_66__or_module_6_res,
         n_majority7_module_66__and_module_6_res,
         n_majority7_module_66__or_module_5_res,
         n_majority7_module_66__and_module_5_res,
         n_majority7_module_66__or_module_4_res,
         n_majority7_module_66__and_module_4_res,
         n_majority7_module_66__or_module_3_res,
         n_majority7_module_66__and_module_3_res,
         n_majority7_module_66__or_module_2_res,
         n_majority7_module_66__and_module_2_res,
         n_majority7_module_66__or_module_1_res,
         n_majority7_module_66__and_module_1_res, n_majority7_module_67_n7,
         n_majority7_module_67_n6, n_majority7_module_67_n5,
         n_majority7_module_67_n4, n_majority7_module_67_n3,
         n_majority7_module_67_n2, n_majority7_module_67_n1,
         n_majority7_module_67__and_module_10_res,
         n_majority7_module_67__or_module_11_res,
         n_majority7_module_67__and_module_9_res,
         n_majority7_module_67__or_module_10_res,
         n_majority7_module_67__or_module_9_res,
         n_majority7_module_67__and_module_8_res,
         n_majority7_module_67__or_module_8_res,
         n_majority7_module_67__and_module_7_res,
         n_majority7_module_67__or_module_7_res,
         n_majority7_module_67__or_module_6_res,
         n_majority7_module_67__and_module_6_res,
         n_majority7_module_67__or_module_5_res,
         n_majority7_module_67__and_module_5_res,
         n_majority7_module_67__or_module_4_res,
         n_majority7_module_67__and_module_4_res,
         n_majority7_module_67__or_module_3_res,
         n_majority7_module_67__and_module_3_res,
         n_majority7_module_67__or_module_2_res,
         n_majority7_module_67__and_module_2_res,
         n_majority7_module_67__or_module_1_res,
         n_majority7_module_67__and_module_1_res, n_majority7_module_68_n7,
         n_majority7_module_68_n6, n_majority7_module_68_n5,
         n_majority7_module_68_n4, n_majority7_module_68_n3,
         n_majority7_module_68_n2, n_majority7_module_68_n1,
         n_majority7_module_68__and_module_10_res,
         n_majority7_module_68__or_module_11_res,
         n_majority7_module_68__and_module_9_res,
         n_majority7_module_68__or_module_10_res,
         n_majority7_module_68__or_module_9_res,
         n_majority7_module_68__and_module_8_res,
         n_majority7_module_68__or_module_8_res,
         n_majority7_module_68__and_module_7_res,
         n_majority7_module_68__or_module_7_res,
         n_majority7_module_68__or_module_6_res,
         n_majority7_module_68__and_module_6_res,
         n_majority7_module_68__or_module_5_res,
         n_majority7_module_68__and_module_5_res,
         n_majority7_module_68__or_module_4_res,
         n_majority7_module_68__and_module_4_res,
         n_majority7_module_68__or_module_3_res,
         n_majority7_module_68__and_module_3_res,
         n_majority7_module_68__or_module_2_res,
         n_majority7_module_68__and_module_2_res,
         n_majority7_module_68__or_module_1_res,
         n_majority7_module_68__and_module_1_res, n_majority7_module_69_n7,
         n_majority7_module_69_n6, n_majority7_module_69_n5,
         n_majority7_module_69_n4, n_majority7_module_69_n3,
         n_majority7_module_69_n2, n_majority7_module_69_n1,
         n_majority7_module_69__and_module_10_res,
         n_majority7_module_69__or_module_11_res,
         n_majority7_module_69__and_module_9_res,
         n_majority7_module_69__or_module_10_res,
         n_majority7_module_69__or_module_9_res,
         n_majority7_module_69__and_module_8_res,
         n_majority7_module_69__or_module_8_res,
         n_majority7_module_69__and_module_7_res,
         n_majority7_module_69__or_module_7_res,
         n_majority7_module_69__or_module_6_res,
         n_majority7_module_69__and_module_6_res,
         n_majority7_module_69__or_module_5_res,
         n_majority7_module_69__and_module_5_res,
         n_majority7_module_69__or_module_4_res,
         n_majority7_module_69__and_module_4_res,
         n_majority7_module_69__or_module_3_res,
         n_majority7_module_69__and_module_3_res,
         n_majority7_module_69__or_module_2_res,
         n_majority7_module_69__and_module_2_res,
         n_majority7_module_69__or_module_1_res,
         n_majority7_module_69__and_module_1_res, n_majority7_module_70_n7,
         n_majority7_module_70_n6, n_majority7_module_70_n5,
         n_majority7_module_70_n4, n_majority7_module_70_n3,
         n_majority7_module_70_n2, n_majority7_module_70_n1,
         n_majority7_module_70__and_module_10_res,
         n_majority7_module_70__or_module_11_res,
         n_majority7_module_70__and_module_9_res,
         n_majority7_module_70__or_module_10_res,
         n_majority7_module_70__or_module_9_res,
         n_majority7_module_70__and_module_8_res,
         n_majority7_module_70__or_module_8_res,
         n_majority7_module_70__and_module_7_res,
         n_majority7_module_70__or_module_7_res,
         n_majority7_module_70__or_module_6_res,
         n_majority7_module_70__and_module_6_res,
         n_majority7_module_70__or_module_5_res,
         n_majority7_module_70__and_module_5_res,
         n_majority7_module_70__or_module_4_res,
         n_majority7_module_70__and_module_4_res,
         n_majority7_module_70__or_module_3_res,
         n_majority7_module_70__and_module_3_res,
         n_majority7_module_70__or_module_2_res,
         n_majority7_module_70__and_module_2_res,
         n_majority7_module_70__or_module_1_res,
         n_majority7_module_70__and_module_1_res, n_majority7_module_71_n7,
         n_majority7_module_71_n6, n_majority7_module_71_n5,
         n_majority7_module_71_n4, n_majority7_module_71_n3,
         n_majority7_module_71_n2, n_majority7_module_71_n1,
         n_majority7_module_71__and_module_10_res,
         n_majority7_module_71__or_module_11_res,
         n_majority7_module_71__and_module_9_res,
         n_majority7_module_71__or_module_10_res,
         n_majority7_module_71__or_module_9_res,
         n_majority7_module_71__and_module_8_res,
         n_majority7_module_71__or_module_8_res,
         n_majority7_module_71__and_module_7_res,
         n_majority7_module_71__or_module_7_res,
         n_majority7_module_71__or_module_6_res,
         n_majority7_module_71__and_module_6_res,
         n_majority7_module_71__or_module_5_res,
         n_majority7_module_71__and_module_5_res,
         n_majority7_module_71__or_module_4_res,
         n_majority7_module_71__and_module_4_res,
         n_majority7_module_71__or_module_3_res,
         n_majority7_module_71__and_module_3_res,
         n_majority7_module_71__or_module_2_res,
         n_majority7_module_71__and_module_2_res,
         n_majority7_module_71__or_module_1_res,
         n_majority7_module_71__and_module_1_res, n_majority7_module_72_n7,
         n_majority7_module_72_n6, n_majority7_module_72_n5,
         n_majority7_module_72_n4, n_majority7_module_72_n3,
         n_majority7_module_72_n2, n_majority7_module_72_n1,
         n_majority7_module_72__and_module_10_res,
         n_majority7_module_72__or_module_11_res,
         n_majority7_module_72__and_module_9_res,
         n_majority7_module_72__or_module_10_res,
         n_majority7_module_72__or_module_9_res,
         n_majority7_module_72__and_module_8_res,
         n_majority7_module_72__or_module_8_res,
         n_majority7_module_72__and_module_7_res,
         n_majority7_module_72__or_module_7_res,
         n_majority7_module_72__or_module_6_res,
         n_majority7_module_72__and_module_6_res,
         n_majority7_module_72__or_module_5_res,
         n_majority7_module_72__and_module_5_res,
         n_majority7_module_72__or_module_4_res,
         n_majority7_module_72__and_module_4_res,
         n_majority7_module_72__or_module_3_res,
         n_majority7_module_72__and_module_3_res,
         n_majority7_module_72__or_module_2_res,
         n_majority7_module_72__and_module_2_res,
         n_majority7_module_72__or_module_1_res,
         n_majority7_module_72__and_module_1_res, n_majority7_module_73_n7,
         n_majority7_module_73_n6, n_majority7_module_73_n5,
         n_majority7_module_73_n4, n_majority7_module_73_n3,
         n_majority7_module_73_n2, n_majority7_module_73_n1,
         n_majority7_module_73__and_module_10_res,
         n_majority7_module_73__or_module_11_res,
         n_majority7_module_73__and_module_9_res,
         n_majority7_module_73__or_module_10_res,
         n_majority7_module_73__or_module_9_res,
         n_majority7_module_73__and_module_8_res,
         n_majority7_module_73__or_module_8_res,
         n_majority7_module_73__and_module_7_res,
         n_majority7_module_73__or_module_7_res,
         n_majority7_module_73__or_module_6_res,
         n_majority7_module_73__and_module_6_res,
         n_majority7_module_73__or_module_5_res,
         n_majority7_module_73__and_module_5_res,
         n_majority7_module_73__or_module_4_res,
         n_majority7_module_73__and_module_4_res,
         n_majority7_module_73__or_module_3_res,
         n_majority7_module_73__and_module_3_res,
         n_majority7_module_73__or_module_2_res,
         n_majority7_module_73__and_module_2_res,
         n_majority7_module_73__or_module_1_res,
         n_majority7_module_73__and_module_1_res, n_majority7_module_74_n7,
         n_majority7_module_74_n6, n_majority7_module_74_n5,
         n_majority7_module_74_n4, n_majority7_module_74_n3,
         n_majority7_module_74_n2, n_majority7_module_74_n1,
         n_majority7_module_74__and_module_10_res,
         n_majority7_module_74__or_module_11_res,
         n_majority7_module_74__and_module_9_res,
         n_majority7_module_74__or_module_10_res,
         n_majority7_module_74__or_module_9_res,
         n_majority7_module_74__and_module_8_res,
         n_majority7_module_74__or_module_8_res,
         n_majority7_module_74__and_module_7_res,
         n_majority7_module_74__or_module_7_res,
         n_majority7_module_74__or_module_6_res,
         n_majority7_module_74__and_module_6_res,
         n_majority7_module_74__or_module_5_res,
         n_majority7_module_74__and_module_5_res,
         n_majority7_module_74__or_module_4_res,
         n_majority7_module_74__and_module_4_res,
         n_majority7_module_74__or_module_3_res,
         n_majority7_module_74__and_module_3_res,
         n_majority7_module_74__or_module_2_res,
         n_majority7_module_74__and_module_2_res,
         n_majority7_module_74__or_module_1_res,
         n_majority7_module_74__and_module_1_res, n_majority7_module_75_n7,
         n_majority7_module_75_n6, n_majority7_module_75_n5,
         n_majority7_module_75_n4, n_majority7_module_75_n3,
         n_majority7_module_75_n2, n_majority7_module_75_n1,
         n_majority7_module_75__and_module_10_res,
         n_majority7_module_75__or_module_11_res,
         n_majority7_module_75__and_module_9_res,
         n_majority7_module_75__or_module_10_res,
         n_majority7_module_75__or_module_9_res,
         n_majority7_module_75__and_module_8_res,
         n_majority7_module_75__or_module_8_res,
         n_majority7_module_75__and_module_7_res,
         n_majority7_module_75__or_module_7_res,
         n_majority7_module_75__or_module_6_res,
         n_majority7_module_75__and_module_6_res,
         n_majority7_module_75__or_module_5_res,
         n_majority7_module_75__and_module_5_res,
         n_majority7_module_75__or_module_4_res,
         n_majority7_module_75__and_module_4_res,
         n_majority7_module_75__or_module_3_res,
         n_majority7_module_75__and_module_3_res,
         n_majority7_module_75__or_module_2_res,
         n_majority7_module_75__and_module_2_res,
         n_majority7_module_75__or_module_1_res,
         n_majority7_module_75__and_module_1_res, n_majority7_module_76_n7,
         n_majority7_module_76_n6, n_majority7_module_76_n5,
         n_majority7_module_76_n4, n_majority7_module_76_n3,
         n_majority7_module_76_n2, n_majority7_module_76_n1,
         n_majority7_module_76__and_module_10_res,
         n_majority7_module_76__or_module_11_res,
         n_majority7_module_76__and_module_9_res,
         n_majority7_module_76__or_module_10_res,
         n_majority7_module_76__or_module_9_res,
         n_majority7_module_76__and_module_8_res,
         n_majority7_module_76__or_module_8_res,
         n_majority7_module_76__and_module_7_res,
         n_majority7_module_76__or_module_7_res,
         n_majority7_module_76__or_module_6_res,
         n_majority7_module_76__and_module_6_res,
         n_majority7_module_76__or_module_5_res,
         n_majority7_module_76__and_module_5_res,
         n_majority7_module_76__or_module_4_res,
         n_majority7_module_76__and_module_4_res,
         n_majority7_module_76__or_module_3_res,
         n_majority7_module_76__and_module_3_res,
         n_majority7_module_76__or_module_2_res,
         n_majority7_module_76__and_module_2_res,
         n_majority7_module_76__or_module_1_res,
         n_majority7_module_76__and_module_1_res, n_majority7_module_77_n7,
         n_majority7_module_77_n6, n_majority7_module_77_n5,
         n_majority7_module_77_n4, n_majority7_module_77_n3,
         n_majority7_module_77_n2, n_majority7_module_77_n1,
         n_majority7_module_77__and_module_10_res,
         n_majority7_module_77__or_module_11_res,
         n_majority7_module_77__and_module_9_res,
         n_majority7_module_77__or_module_10_res,
         n_majority7_module_77__or_module_9_res,
         n_majority7_module_77__and_module_8_res,
         n_majority7_module_77__or_module_8_res,
         n_majority7_module_77__and_module_7_res,
         n_majority7_module_77__or_module_7_res,
         n_majority7_module_77__or_module_6_res,
         n_majority7_module_77__and_module_6_res,
         n_majority7_module_77__or_module_5_res,
         n_majority7_module_77__and_module_5_res,
         n_majority7_module_77__or_module_4_res,
         n_majority7_module_77__and_module_4_res,
         n_majority7_module_77__or_module_3_res,
         n_majority7_module_77__and_module_3_res,
         n_majority7_module_77__or_module_2_res,
         n_majority7_module_77__and_module_2_res,
         n_majority7_module_77__or_module_1_res,
         n_majority7_module_77__and_module_1_res, n_majority7_module_78_n7,
         n_majority7_module_78_n6, n_majority7_module_78_n5,
         n_majority7_module_78_n4, n_majority7_module_78_n3,
         n_majority7_module_78_n2, n_majority7_module_78_n1,
         n_majority7_module_78__and_module_10_res,
         n_majority7_module_78__or_module_11_res,
         n_majority7_module_78__and_module_9_res,
         n_majority7_module_78__or_module_10_res,
         n_majority7_module_78__or_module_9_res,
         n_majority7_module_78__and_module_8_res,
         n_majority7_module_78__or_module_8_res,
         n_majority7_module_78__and_module_7_res,
         n_majority7_module_78__or_module_7_res,
         n_majority7_module_78__or_module_6_res,
         n_majority7_module_78__and_module_6_res,
         n_majority7_module_78__or_module_5_res,
         n_majority7_module_78__and_module_5_res,
         n_majority7_module_78__or_module_4_res,
         n_majority7_module_78__and_module_4_res,
         n_majority7_module_78__or_module_3_res,
         n_majority7_module_78__and_module_3_res,
         n_majority7_module_78__or_module_2_res,
         n_majority7_module_78__and_module_2_res,
         n_majority7_module_78__or_module_1_res,
         n_majority7_module_78__and_module_1_res, n_majority7_module_79_n7,
         n_majority7_module_79_n6, n_majority7_module_79_n5,
         n_majority7_module_79_n4, n_majority7_module_79_n3,
         n_majority7_module_79_n2, n_majority7_module_79_n1,
         n_majority7_module_79__and_module_10_res,
         n_majority7_module_79__or_module_11_res,
         n_majority7_module_79__and_module_9_res,
         n_majority7_module_79__or_module_10_res,
         n_majority7_module_79__or_module_9_res,
         n_majority7_module_79__and_module_8_res,
         n_majority7_module_79__or_module_8_res,
         n_majority7_module_79__and_module_7_res,
         n_majority7_module_79__or_module_7_res,
         n_majority7_module_79__or_module_6_res,
         n_majority7_module_79__and_module_6_res,
         n_majority7_module_79__or_module_5_res,
         n_majority7_module_79__and_module_5_res,
         n_majority7_module_79__or_module_4_res,
         n_majority7_module_79__and_module_4_res,
         n_majority7_module_79__or_module_3_res,
         n_majority7_module_79__and_module_3_res,
         n_majority7_module_79__or_module_2_res,
         n_majority7_module_79__and_module_2_res,
         n_majority7_module_79__or_module_1_res,
         n_majority7_module_79__and_module_1_res, n_majority7_module_80_n7,
         n_majority7_module_80_n6, n_majority7_module_80_n5,
         n_majority7_module_80_n4, n_majority7_module_80_n3,
         n_majority7_module_80_n2, n_majority7_module_80_n1,
         n_majority7_module_80__and_module_10_res,
         n_majority7_module_80__or_module_11_res,
         n_majority7_module_80__and_module_9_res,
         n_majority7_module_80__or_module_10_res,
         n_majority7_module_80__or_module_9_res,
         n_majority7_module_80__and_module_8_res,
         n_majority7_module_80__or_module_8_res,
         n_majority7_module_80__and_module_7_res,
         n_majority7_module_80__or_module_7_res,
         n_majority7_module_80__or_module_6_res,
         n_majority7_module_80__and_module_6_res,
         n_majority7_module_80__or_module_5_res,
         n_majority7_module_80__and_module_5_res,
         n_majority7_module_80__or_module_4_res,
         n_majority7_module_80__and_module_4_res,
         n_majority7_module_80__or_module_3_res,
         n_majority7_module_80__and_module_3_res,
         n_majority7_module_80__or_module_2_res,
         n_majority7_module_80__and_module_2_res,
         n_majority7_module_80__or_module_1_res,
         n_majority7_module_80__and_module_1_res, n_majority7_module_81_n7,
         n_majority7_module_81_n6, n_majority7_module_81_n5,
         n_majority7_module_81_n4, n_majority7_module_81_n3,
         n_majority7_module_81_n2, n_majority7_module_81_n1,
         n_majority7_module_81__and_module_10_res,
         n_majority7_module_81__or_module_11_res,
         n_majority7_module_81__and_module_9_res,
         n_majority7_module_81__or_module_10_res,
         n_majority7_module_81__or_module_9_res,
         n_majority7_module_81__and_module_8_res,
         n_majority7_module_81__or_module_8_res,
         n_majority7_module_81__and_module_7_res,
         n_majority7_module_81__or_module_7_res,
         n_majority7_module_81__or_module_6_res,
         n_majority7_module_81__and_module_6_res,
         n_majority7_module_81__or_module_5_res,
         n_majority7_module_81__and_module_5_res,
         n_majority7_module_81__or_module_4_res,
         n_majority7_module_81__and_module_4_res,
         n_majority7_module_81__or_module_3_res,
         n_majority7_module_81__and_module_3_res,
         n_majority7_module_81__or_module_2_res,
         n_majority7_module_81__and_module_2_res,
         n_majority7_module_81__or_module_1_res,
         n_majority7_module_81__and_module_1_res, n_majority7_module_82_n7,
         n_majority7_module_82_n6, n_majority7_module_82_n5,
         n_majority7_module_82_n4, n_majority7_module_82_n3,
         n_majority7_module_82_n2, n_majority7_module_82_n1,
         n_majority7_module_82__and_module_10_res,
         n_majority7_module_82__or_module_11_res,
         n_majority7_module_82__and_module_9_res,
         n_majority7_module_82__or_module_10_res,
         n_majority7_module_82__or_module_9_res,
         n_majority7_module_82__and_module_8_res,
         n_majority7_module_82__or_module_8_res,
         n_majority7_module_82__and_module_7_res,
         n_majority7_module_82__or_module_7_res,
         n_majority7_module_82__or_module_6_res,
         n_majority7_module_82__and_module_6_res,
         n_majority7_module_82__or_module_5_res,
         n_majority7_module_82__and_module_5_res,
         n_majority7_module_82__or_module_4_res,
         n_majority7_module_82__and_module_4_res,
         n_majority7_module_82__or_module_3_res,
         n_majority7_module_82__and_module_3_res,
         n_majority7_module_82__or_module_2_res,
         n_majority7_module_82__and_module_2_res,
         n_majority7_module_82__or_module_1_res,
         n_majority7_module_82__and_module_1_res, n_majority7_module_83_n7,
         n_majority7_module_83_n6, n_majority7_module_83_n5,
         n_majority7_module_83_n4, n_majority7_module_83_n3,
         n_majority7_module_83_n2, n_majority7_module_83_n1,
         n_majority7_module_83__and_module_10_res,
         n_majority7_module_83__or_module_11_res,
         n_majority7_module_83__and_module_9_res,
         n_majority7_module_83__or_module_10_res,
         n_majority7_module_83__or_module_9_res,
         n_majority7_module_83__and_module_8_res,
         n_majority7_module_83__or_module_8_res,
         n_majority7_module_83__and_module_7_res,
         n_majority7_module_83__or_module_7_res,
         n_majority7_module_83__or_module_6_res,
         n_majority7_module_83__and_module_6_res,
         n_majority7_module_83__or_module_5_res,
         n_majority7_module_83__and_module_5_res,
         n_majority7_module_83__or_module_4_res,
         n_majority7_module_83__and_module_4_res,
         n_majority7_module_83__or_module_3_res,
         n_majority7_module_83__and_module_3_res,
         n_majority7_module_83__or_module_2_res,
         n_majority7_module_83__and_module_2_res,
         n_majority7_module_83__or_module_1_res,
         n_majority7_module_83__and_module_1_res, n_majority7_module_84_n7,
         n_majority7_module_84_n6, n_majority7_module_84_n5,
         n_majority7_module_84_n4, n_majority7_module_84_n3,
         n_majority7_module_84_n2, n_majority7_module_84_n1,
         n_majority7_module_84__and_module_10_res,
         n_majority7_module_84__or_module_11_res,
         n_majority7_module_84__and_module_9_res,
         n_majority7_module_84__or_module_10_res,
         n_majority7_module_84__or_module_9_res,
         n_majority7_module_84__and_module_8_res,
         n_majority7_module_84__or_module_8_res,
         n_majority7_module_84__and_module_7_res,
         n_majority7_module_84__or_module_7_res,
         n_majority7_module_84__or_module_6_res,
         n_majority7_module_84__and_module_6_res,
         n_majority7_module_84__or_module_5_res,
         n_majority7_module_84__and_module_5_res,
         n_majority7_module_84__or_module_4_res,
         n_majority7_module_84__and_module_4_res,
         n_majority7_module_84__or_module_3_res,
         n_majority7_module_84__and_module_3_res,
         n_majority7_module_84__or_module_2_res,
         n_majority7_module_84__and_module_2_res,
         n_majority7_module_84__or_module_1_res,
         n_majority7_module_84__and_module_1_res, n_majority7_module_85_n7,
         n_majority7_module_85_n6, n_majority7_module_85_n5,
         n_majority7_module_85_n4, n_majority7_module_85_n3,
         n_majority7_module_85_n2, n_majority7_module_85_n1,
         n_majority7_module_85__and_module_10_res,
         n_majority7_module_85__or_module_11_res,
         n_majority7_module_85__and_module_9_res,
         n_majority7_module_85__or_module_10_res,
         n_majority7_module_85__or_module_9_res,
         n_majority7_module_85__and_module_8_res,
         n_majority7_module_85__or_module_8_res,
         n_majority7_module_85__and_module_7_res,
         n_majority7_module_85__or_module_7_res,
         n_majority7_module_85__or_module_6_res,
         n_majority7_module_85__and_module_6_res,
         n_majority7_module_85__or_module_5_res,
         n_majority7_module_85__and_module_5_res,
         n_majority7_module_85__or_module_4_res,
         n_majority7_module_85__and_module_4_res,
         n_majority7_module_85__or_module_3_res,
         n_majority7_module_85__and_module_3_res,
         n_majority7_module_85__or_module_2_res,
         n_majority7_module_85__and_module_2_res,
         n_majority7_module_85__or_module_1_res,
         n_majority7_module_85__and_module_1_res, n_majority7_module_86_n7,
         n_majority7_module_86_n6, n_majority7_module_86_n5,
         n_majority7_module_86_n4, n_majority7_module_86_n3,
         n_majority7_module_86_n2, n_majority7_module_86_n1,
         n_majority7_module_86__and_module_10_res,
         n_majority7_module_86__or_module_11_res,
         n_majority7_module_86__and_module_9_res,
         n_majority7_module_86__or_module_10_res,
         n_majority7_module_86__or_module_9_res,
         n_majority7_module_86__and_module_8_res,
         n_majority7_module_86__or_module_8_res,
         n_majority7_module_86__and_module_7_res,
         n_majority7_module_86__or_module_7_res,
         n_majority7_module_86__or_module_6_res,
         n_majority7_module_86__and_module_6_res,
         n_majority7_module_86__or_module_5_res,
         n_majority7_module_86__and_module_5_res,
         n_majority7_module_86__or_module_4_res,
         n_majority7_module_86__and_module_4_res,
         n_majority7_module_86__or_module_3_res,
         n_majority7_module_86__and_module_3_res,
         n_majority7_module_86__or_module_2_res,
         n_majority7_module_86__and_module_2_res,
         n_majority7_module_86__or_module_1_res,
         n_majority7_module_86__and_module_1_res, n_majority7_module_87_n7,
         n_majority7_module_87_n6, n_majority7_module_87_n5,
         n_majority7_module_87_n4, n_majority7_module_87_n3,
         n_majority7_module_87_n2, n_majority7_module_87_n1,
         n_majority7_module_87__and_module_10_res,
         n_majority7_module_87__or_module_11_res,
         n_majority7_module_87__and_module_9_res,
         n_majority7_module_87__or_module_10_res,
         n_majority7_module_87__or_module_9_res,
         n_majority7_module_87__and_module_8_res,
         n_majority7_module_87__or_module_8_res,
         n_majority7_module_87__and_module_7_res,
         n_majority7_module_87__or_module_7_res,
         n_majority7_module_87__or_module_6_res,
         n_majority7_module_87__and_module_6_res,
         n_majority7_module_87__or_module_5_res,
         n_majority7_module_87__and_module_5_res,
         n_majority7_module_87__or_module_4_res,
         n_majority7_module_87__and_module_4_res,
         n_majority7_module_87__or_module_3_res,
         n_majority7_module_87__and_module_3_res,
         n_majority7_module_87__or_module_2_res,
         n_majority7_module_87__and_module_2_res,
         n_majority7_module_87__or_module_1_res,
         n_majority7_module_87__and_module_1_res, n_majority7_module_88_n7,
         n_majority7_module_88_n6, n_majority7_module_88_n5,
         n_majority7_module_88_n4, n_majority7_module_88_n3,
         n_majority7_module_88_n2, n_majority7_module_88_n1,
         n_majority7_module_88__and_module_10_res,
         n_majority7_module_88__or_module_11_res,
         n_majority7_module_88__and_module_9_res,
         n_majority7_module_88__or_module_10_res,
         n_majority7_module_88__or_module_9_res,
         n_majority7_module_88__and_module_8_res,
         n_majority7_module_88__or_module_8_res,
         n_majority7_module_88__and_module_7_res,
         n_majority7_module_88__or_module_7_res,
         n_majority7_module_88__or_module_6_res,
         n_majority7_module_88__and_module_6_res,
         n_majority7_module_88__or_module_5_res,
         n_majority7_module_88__and_module_5_res,
         n_majority7_module_88__or_module_4_res,
         n_majority7_module_88__and_module_4_res,
         n_majority7_module_88__or_module_3_res,
         n_majority7_module_88__and_module_3_res,
         n_majority7_module_88__or_module_2_res,
         n_majority7_module_88__and_module_2_res,
         n_majority7_module_88__or_module_1_res,
         n_majority7_module_88__and_module_1_res, n_majority7_module_89_n7,
         n_majority7_module_89_n6, n_majority7_module_89_n5,
         n_majority7_module_89_n4, n_majority7_module_89_n3,
         n_majority7_module_89_n2, n_majority7_module_89_n1,
         n_majority7_module_89__and_module_10_res,
         n_majority7_module_89__or_module_11_res,
         n_majority7_module_89__and_module_9_res,
         n_majority7_module_89__or_module_10_res,
         n_majority7_module_89__or_module_9_res,
         n_majority7_module_89__and_module_8_res,
         n_majority7_module_89__or_module_8_res,
         n_majority7_module_89__and_module_7_res,
         n_majority7_module_89__or_module_7_res,
         n_majority7_module_89__or_module_6_res,
         n_majority7_module_89__and_module_6_res,
         n_majority7_module_89__or_module_5_res,
         n_majority7_module_89__and_module_5_res,
         n_majority7_module_89__or_module_4_res,
         n_majority7_module_89__and_module_4_res,
         n_majority7_module_89__or_module_3_res,
         n_majority7_module_89__and_module_3_res,
         n_majority7_module_89__or_module_2_res,
         n_majority7_module_89__and_module_2_res,
         n_majority7_module_89__or_module_1_res,
         n_majority7_module_89__and_module_1_res, n_majority7_module_90_n7,
         n_majority7_module_90_n6, n_majority7_module_90_n5,
         n_majority7_module_90_n4, n_majority7_module_90_n3,
         n_majority7_module_90_n2, n_majority7_module_90_n1,
         n_majority7_module_90__and_module_10_res,
         n_majority7_module_90__or_module_11_res,
         n_majority7_module_90__and_module_9_res,
         n_majority7_module_90__or_module_10_res,
         n_majority7_module_90__or_module_9_res,
         n_majority7_module_90__and_module_8_res,
         n_majority7_module_90__or_module_8_res,
         n_majority7_module_90__and_module_7_res,
         n_majority7_module_90__or_module_7_res,
         n_majority7_module_90__or_module_6_res,
         n_majority7_module_90__and_module_6_res,
         n_majority7_module_90__or_module_5_res,
         n_majority7_module_90__and_module_5_res,
         n_majority7_module_90__or_module_4_res,
         n_majority7_module_90__and_module_4_res,
         n_majority7_module_90__or_module_3_res,
         n_majority7_module_90__and_module_3_res,
         n_majority7_module_90__or_module_2_res,
         n_majority7_module_90__and_module_2_res,
         n_majority7_module_90__or_module_1_res,
         n_majority7_module_90__and_module_1_res, n_majority7_module_91_n7,
         n_majority7_module_91_n6, n_majority7_module_91_n5,
         n_majority7_module_91_n4, n_majority7_module_91_n3,
         n_majority7_module_91_n2, n_majority7_module_91_n1,
         n_majority7_module_91__and_module_10_res,
         n_majority7_module_91__or_module_11_res,
         n_majority7_module_91__and_module_9_res,
         n_majority7_module_91__or_module_10_res,
         n_majority7_module_91__or_module_9_res,
         n_majority7_module_91__and_module_8_res,
         n_majority7_module_91__or_module_8_res,
         n_majority7_module_91__and_module_7_res,
         n_majority7_module_91__or_module_7_res,
         n_majority7_module_91__or_module_6_res,
         n_majority7_module_91__and_module_6_res,
         n_majority7_module_91__or_module_5_res,
         n_majority7_module_91__and_module_5_res,
         n_majority7_module_91__or_module_4_res,
         n_majority7_module_91__and_module_4_res,
         n_majority7_module_91__or_module_3_res,
         n_majority7_module_91__and_module_3_res,
         n_majority7_module_91__or_module_2_res,
         n_majority7_module_91__and_module_2_res,
         n_majority7_module_91__or_module_1_res,
         n_majority7_module_91__and_module_1_res, n_majority7_module_92_n7,
         n_majority7_module_92_n6, n_majority7_module_92_n5,
         n_majority7_module_92_n4, n_majority7_module_92_n3,
         n_majority7_module_92_n2, n_majority7_module_92_n1,
         n_majority7_module_92__and_module_10_res,
         n_majority7_module_92__or_module_11_res,
         n_majority7_module_92__and_module_9_res,
         n_majority7_module_92__or_module_10_res,
         n_majority7_module_92__or_module_9_res,
         n_majority7_module_92__and_module_8_res,
         n_majority7_module_92__or_module_8_res,
         n_majority7_module_92__and_module_7_res,
         n_majority7_module_92__or_module_7_res,
         n_majority7_module_92__or_module_6_res,
         n_majority7_module_92__and_module_6_res,
         n_majority7_module_92__or_module_5_res,
         n_majority7_module_92__and_module_5_res,
         n_majority7_module_92__or_module_4_res,
         n_majority7_module_92__and_module_4_res,
         n_majority7_module_92__or_module_3_res,
         n_majority7_module_92__and_module_3_res,
         n_majority7_module_92__or_module_2_res,
         n_majority7_module_92__and_module_2_res,
         n_majority7_module_92__or_module_1_res,
         n_majority7_module_92__and_module_1_res, n_majority7_module_93_n7,
         n_majority7_module_93_n6, n_majority7_module_93_n5,
         n_majority7_module_93_n4, n_majority7_module_93_n3,
         n_majority7_module_93_n2, n_majority7_module_93_n1,
         n_majority7_module_93__and_module_10_res,
         n_majority7_module_93__or_module_11_res,
         n_majority7_module_93__and_module_9_res,
         n_majority7_module_93__or_module_10_res,
         n_majority7_module_93__or_module_9_res,
         n_majority7_module_93__and_module_8_res,
         n_majority7_module_93__or_module_8_res,
         n_majority7_module_93__and_module_7_res,
         n_majority7_module_93__or_module_7_res,
         n_majority7_module_93__or_module_6_res,
         n_majority7_module_93__and_module_6_res,
         n_majority7_module_93__or_module_5_res,
         n_majority7_module_93__and_module_5_res,
         n_majority7_module_93__or_module_4_res,
         n_majority7_module_93__and_module_4_res,
         n_majority7_module_93__or_module_3_res,
         n_majority7_module_93__and_module_3_res,
         n_majority7_module_93__or_module_2_res,
         n_majority7_module_93__and_module_2_res,
         n_majority7_module_93__or_module_1_res,
         n_majority7_module_93__and_module_1_res, n_majority7_module_94_n7,
         n_majority7_module_94_n6, n_majority7_module_94_n5,
         n_majority7_module_94_n4, n_majority7_module_94_n3,
         n_majority7_module_94_n2, n_majority7_module_94_n1,
         n_majority7_module_94__and_module_10_res,
         n_majority7_module_94__or_module_11_res,
         n_majority7_module_94__and_module_9_res,
         n_majority7_module_94__or_module_10_res,
         n_majority7_module_94__or_module_9_res,
         n_majority7_module_94__and_module_8_res,
         n_majority7_module_94__or_module_8_res,
         n_majority7_module_94__and_module_7_res,
         n_majority7_module_94__or_module_7_res,
         n_majority7_module_94__or_module_6_res,
         n_majority7_module_94__and_module_6_res,
         n_majority7_module_94__or_module_5_res,
         n_majority7_module_94__and_module_5_res,
         n_majority7_module_94__or_module_4_res,
         n_majority7_module_94__and_module_4_res,
         n_majority7_module_94__or_module_3_res,
         n_majority7_module_94__and_module_3_res,
         n_majority7_module_94__or_module_2_res,
         n_majority7_module_94__and_module_2_res,
         n_majority7_module_94__or_module_1_res,
         n_majority7_module_94__and_module_1_res, n_majority7_module_95_n7,
         n_majority7_module_95_n6, n_majority7_module_95_n5,
         n_majority7_module_95_n4, n_majority7_module_95_n3,
         n_majority7_module_95_n2, n_majority7_module_95_n1,
         n_majority7_module_95__and_module_10_res,
         n_majority7_module_95__or_module_11_res,
         n_majority7_module_95__and_module_9_res,
         n_majority7_module_95__or_module_10_res,
         n_majority7_module_95__or_module_9_res,
         n_majority7_module_95__and_module_8_res,
         n_majority7_module_95__or_module_8_res,
         n_majority7_module_95__and_module_7_res,
         n_majority7_module_95__or_module_7_res,
         n_majority7_module_95__or_module_6_res,
         n_majority7_module_95__and_module_6_res,
         n_majority7_module_95__or_module_5_res,
         n_majority7_module_95__and_module_5_res,
         n_majority7_module_95__or_module_4_res,
         n_majority7_module_95__and_module_4_res,
         n_majority7_module_95__or_module_3_res,
         n_majority7_module_95__and_module_3_res,
         n_majority7_module_95__or_module_2_res,
         n_majority7_module_95__and_module_2_res,
         n_majority7_module_95__or_module_1_res,
         n_majority7_module_95__and_module_1_res, n_majority7_module_96_n7,
         n_majority7_module_96_n6, n_majority7_module_96_n5,
         n_majority7_module_96_n4, n_majority7_module_96_n3,
         n_majority7_module_96_n2, n_majority7_module_96_n1,
         n_majority7_module_96__and_module_10_res,
         n_majority7_module_96__or_module_11_res,
         n_majority7_module_96__and_module_9_res,
         n_majority7_module_96__or_module_10_res,
         n_majority7_module_96__or_module_9_res,
         n_majority7_module_96__and_module_8_res,
         n_majority7_module_96__or_module_8_res,
         n_majority7_module_96__and_module_7_res,
         n_majority7_module_96__or_module_7_res,
         n_majority7_module_96__or_module_6_res,
         n_majority7_module_96__and_module_6_res,
         n_majority7_module_96__or_module_5_res,
         n_majority7_module_96__and_module_5_res,
         n_majority7_module_96__or_module_4_res,
         n_majority7_module_96__and_module_4_res,
         n_majority7_module_96__or_module_3_res,
         n_majority7_module_96__and_module_3_res,
         n_majority7_module_96__or_module_2_res,
         n_majority7_module_96__and_module_2_res,
         n_majority7_module_96__or_module_1_res,
         n_majority7_module_96__and_module_1_res, n_majority7_module_97_n7,
         n_majority7_module_97_n6, n_majority7_module_97_n5,
         n_majority7_module_97_n4, n_majority7_module_97_n3,
         n_majority7_module_97_n2, n_majority7_module_97_n1,
         n_majority7_module_97__and_module_10_res,
         n_majority7_module_97__or_module_11_res,
         n_majority7_module_97__and_module_9_res,
         n_majority7_module_97__or_module_10_res,
         n_majority7_module_97__or_module_9_res,
         n_majority7_module_97__and_module_8_res,
         n_majority7_module_97__or_module_8_res,
         n_majority7_module_97__and_module_7_res,
         n_majority7_module_97__or_module_7_res,
         n_majority7_module_97__or_module_6_res,
         n_majority7_module_97__and_module_6_res,
         n_majority7_module_97__or_module_5_res,
         n_majority7_module_97__and_module_5_res,
         n_majority7_module_97__or_module_4_res,
         n_majority7_module_97__and_module_4_res,
         n_majority7_module_97__or_module_3_res,
         n_majority7_module_97__and_module_3_res,
         n_majority7_module_97__or_module_2_res,
         n_majority7_module_97__and_module_2_res,
         n_majority7_module_97__or_module_1_res,
         n_majority7_module_97__and_module_1_res, n_majority7_module_98_n7,
         n_majority7_module_98_n6, n_majority7_module_98_n5,
         n_majority7_module_98_n4, n_majority7_module_98_n3,
         n_majority7_module_98_n2, n_majority7_module_98_n1,
         n_majority7_module_98__and_module_10_res,
         n_majority7_module_98__or_module_11_res,
         n_majority7_module_98__and_module_9_res,
         n_majority7_module_98__or_module_10_res,
         n_majority7_module_98__or_module_9_res,
         n_majority7_module_98__and_module_8_res,
         n_majority7_module_98__or_module_8_res,
         n_majority7_module_98__and_module_7_res,
         n_majority7_module_98__or_module_7_res,
         n_majority7_module_98__or_module_6_res,
         n_majority7_module_98__and_module_6_res,
         n_majority7_module_98__or_module_5_res,
         n_majority7_module_98__and_module_5_res,
         n_majority7_module_98__or_module_4_res,
         n_majority7_module_98__and_module_4_res,
         n_majority7_module_98__or_module_3_res,
         n_majority7_module_98__and_module_3_res,
         n_majority7_module_98__or_module_2_res,
         n_majority7_module_98__and_module_2_res,
         n_majority7_module_98__or_module_1_res,
         n_majority7_module_98__and_module_1_res, n_majority7_module_99_n7,
         n_majority7_module_99_n6, n_majority7_module_99_n5,
         n_majority7_module_99_n4, n_majority7_module_99_n3,
         n_majority7_module_99_n2, n_majority7_module_99_n1,
         n_majority7_module_99__and_module_10_res,
         n_majority7_module_99__or_module_11_res,
         n_majority7_module_99__and_module_9_res,
         n_majority7_module_99__or_module_10_res,
         n_majority7_module_99__or_module_9_res,
         n_majority7_module_99__and_module_8_res,
         n_majority7_module_99__or_module_8_res,
         n_majority7_module_99__and_module_7_res,
         n_majority7_module_99__or_module_7_res,
         n_majority7_module_99__or_module_6_res,
         n_majority7_module_99__and_module_6_res,
         n_majority7_module_99__or_module_5_res,
         n_majority7_module_99__and_module_5_res,
         n_majority7_module_99__or_module_4_res,
         n_majority7_module_99__and_module_4_res,
         n_majority7_module_99__or_module_3_res,
         n_majority7_module_99__and_module_3_res,
         n_majority7_module_99__or_module_2_res,
         n_majority7_module_99__and_module_2_res,
         n_majority7_module_99__or_module_1_res,
         n_majority7_module_99__and_module_1_res, n_majority7_module_100_n7,
         n_majority7_module_100_n6, n_majority7_module_100_n5,
         n_majority7_module_100_n4, n_majority7_module_100_n3,
         n_majority7_module_100_n2, n_majority7_module_100_n1,
         n_majority7_module_100__and_module_10_res,
         n_majority7_module_100__or_module_11_res,
         n_majority7_module_100__and_module_9_res,
         n_majority7_module_100__or_module_10_res,
         n_majority7_module_100__or_module_9_res,
         n_majority7_module_100__and_module_8_res,
         n_majority7_module_100__or_module_8_res,
         n_majority7_module_100__and_module_7_res,
         n_majority7_module_100__or_module_7_res,
         n_majority7_module_100__or_module_6_res,
         n_majority7_module_100__and_module_6_res,
         n_majority7_module_100__or_module_5_res,
         n_majority7_module_100__and_module_5_res,
         n_majority7_module_100__or_module_4_res,
         n_majority7_module_100__and_module_4_res,
         n_majority7_module_100__or_module_3_res,
         n_majority7_module_100__and_module_3_res,
         n_majority7_module_100__or_module_2_res,
         n_majority7_module_100__and_module_2_res,
         n_majority7_module_100__or_module_1_res,
         n_majority7_module_100__and_module_1_res, n_majority7_module_101_n7,
         n_majority7_module_101_n6, n_majority7_module_101_n5,
         n_majority7_module_101_n4, n_majority7_module_101_n3,
         n_majority7_module_101_n2, n_majority7_module_101_n1,
         n_majority7_module_101__and_module_10_res,
         n_majority7_module_101__or_module_11_res,
         n_majority7_module_101__and_module_9_res,
         n_majority7_module_101__or_module_10_res,
         n_majority7_module_101__or_module_9_res,
         n_majority7_module_101__and_module_8_res,
         n_majority7_module_101__or_module_8_res,
         n_majority7_module_101__and_module_7_res,
         n_majority7_module_101__or_module_7_res,
         n_majority7_module_101__or_module_6_res,
         n_majority7_module_101__and_module_6_res,
         n_majority7_module_101__or_module_5_res,
         n_majority7_module_101__and_module_5_res,
         n_majority7_module_101__or_module_4_res,
         n_majority7_module_101__and_module_4_res,
         n_majority7_module_101__or_module_3_res,
         n_majority7_module_101__and_module_3_res,
         n_majority7_module_101__or_module_2_res,
         n_majority7_module_101__and_module_2_res,
         n_majority7_module_101__or_module_1_res,
         n_majority7_module_101__and_module_1_res, n_majority7_module_102_n7,
         n_majority7_module_102_n6, n_majority7_module_102_n5,
         n_majority7_module_102_n4, n_majority7_module_102_n3,
         n_majority7_module_102_n2, n_majority7_module_102_n1,
         n_majority7_module_102__and_module_10_res,
         n_majority7_module_102__or_module_11_res,
         n_majority7_module_102__and_module_9_res,
         n_majority7_module_102__or_module_10_res,
         n_majority7_module_102__or_module_9_res,
         n_majority7_module_102__and_module_8_res,
         n_majority7_module_102__or_module_8_res,
         n_majority7_module_102__and_module_7_res,
         n_majority7_module_102__or_module_7_res,
         n_majority7_module_102__or_module_6_res,
         n_majority7_module_102__and_module_6_res,
         n_majority7_module_102__or_module_5_res,
         n_majority7_module_102__and_module_5_res,
         n_majority7_module_102__or_module_4_res,
         n_majority7_module_102__and_module_4_res,
         n_majority7_module_102__or_module_3_res,
         n_majority7_module_102__and_module_3_res,
         n_majority7_module_102__or_module_2_res,
         n_majority7_module_102__and_module_2_res,
         n_majority7_module_102__or_module_1_res,
         n_majority7_module_102__and_module_1_res, n_majority7_module_103_n7,
         n_majority7_module_103_n6, n_majority7_module_103_n5,
         n_majority7_module_103_n4, n_majority7_module_103_n3,
         n_majority7_module_103_n2, n_majority7_module_103_n1,
         n_majority7_module_103__and_module_10_res,
         n_majority7_module_103__or_module_11_res,
         n_majority7_module_103__and_module_9_res,
         n_majority7_module_103__or_module_10_res,
         n_majority7_module_103__or_module_9_res,
         n_majority7_module_103__and_module_8_res,
         n_majority7_module_103__or_module_8_res,
         n_majority7_module_103__and_module_7_res,
         n_majority7_module_103__or_module_7_res,
         n_majority7_module_103__or_module_6_res,
         n_majority7_module_103__and_module_6_res,
         n_majority7_module_103__or_module_5_res,
         n_majority7_module_103__and_module_5_res,
         n_majority7_module_103__or_module_4_res,
         n_majority7_module_103__and_module_4_res,
         n_majority7_module_103__or_module_3_res,
         n_majority7_module_103__and_module_3_res,
         n_majority7_module_103__or_module_2_res,
         n_majority7_module_103__and_module_2_res,
         n_majority7_module_103__or_module_1_res,
         n_majority7_module_103__and_module_1_res, n_majority7_module_104_n7,
         n_majority7_module_104_n6, n_majority7_module_104_n5,
         n_majority7_module_104_n4, n_majority7_module_104_n3,
         n_majority7_module_104_n2, n_majority7_module_104_n1,
         n_majority7_module_104__and_module_10_res,
         n_majority7_module_104__or_module_11_res,
         n_majority7_module_104__and_module_9_res,
         n_majority7_module_104__or_module_10_res,
         n_majority7_module_104__or_module_9_res,
         n_majority7_module_104__and_module_8_res,
         n_majority7_module_104__or_module_8_res,
         n_majority7_module_104__and_module_7_res,
         n_majority7_module_104__or_module_7_res,
         n_majority7_module_104__or_module_6_res,
         n_majority7_module_104__and_module_6_res,
         n_majority7_module_104__or_module_5_res,
         n_majority7_module_104__and_module_5_res,
         n_majority7_module_104__or_module_4_res,
         n_majority7_module_104__and_module_4_res,
         n_majority7_module_104__or_module_3_res,
         n_majority7_module_104__and_module_3_res,
         n_majority7_module_104__or_module_2_res,
         n_majority7_module_104__and_module_2_res,
         n_majority7_module_104__or_module_1_res,
         n_majority7_module_104__and_module_1_res, n_majority7_module_105_n7,
         n_majority7_module_105_n6, n_majority7_module_105_n5,
         n_majority7_module_105_n4, n_majority7_module_105_n3,
         n_majority7_module_105_n2, n_majority7_module_105_n1,
         n_majority7_module_105__and_module_10_res,
         n_majority7_module_105__or_module_11_res,
         n_majority7_module_105__and_module_9_res,
         n_majority7_module_105__or_module_10_res,
         n_majority7_module_105__or_module_9_res,
         n_majority7_module_105__and_module_8_res,
         n_majority7_module_105__or_module_8_res,
         n_majority7_module_105__and_module_7_res,
         n_majority7_module_105__or_module_7_res,
         n_majority7_module_105__or_module_6_res,
         n_majority7_module_105__and_module_6_res,
         n_majority7_module_105__or_module_5_res,
         n_majority7_module_105__and_module_5_res,
         n_majority7_module_105__or_module_4_res,
         n_majority7_module_105__and_module_4_res,
         n_majority7_module_105__or_module_3_res,
         n_majority7_module_105__and_module_3_res,
         n_majority7_module_105__or_module_2_res,
         n_majority7_module_105__and_module_2_res,
         n_majority7_module_105__or_module_1_res,
         n_majority7_module_105__and_module_1_res, n_majority7_module_106_n7,
         n_majority7_module_106_n6, n_majority7_module_106_n5,
         n_majority7_module_106_n4, n_majority7_module_106_n3,
         n_majority7_module_106_n2, n_majority7_module_106_n1,
         n_majority7_module_106__and_module_10_res,
         n_majority7_module_106__or_module_11_res,
         n_majority7_module_106__and_module_9_res,
         n_majority7_module_106__or_module_10_res,
         n_majority7_module_106__or_module_9_res,
         n_majority7_module_106__and_module_8_res,
         n_majority7_module_106__or_module_8_res,
         n_majority7_module_106__and_module_7_res,
         n_majority7_module_106__or_module_7_res,
         n_majority7_module_106__or_module_6_res,
         n_majority7_module_106__and_module_6_res,
         n_majority7_module_106__or_module_5_res,
         n_majority7_module_106__and_module_5_res,
         n_majority7_module_106__or_module_4_res,
         n_majority7_module_106__and_module_4_res,
         n_majority7_module_106__or_module_3_res,
         n_majority7_module_106__and_module_3_res,
         n_majority7_module_106__or_module_2_res,
         n_majority7_module_106__and_module_2_res,
         n_majority7_module_106__or_module_1_res,
         n_majority7_module_106__and_module_1_res, n_majority7_module_107_n7,
         n_majority7_module_107_n6, n_majority7_module_107_n5,
         n_majority7_module_107_n4, n_majority7_module_107_n3,
         n_majority7_module_107_n2, n_majority7_module_107_n1,
         n_majority7_module_107__and_module_10_res,
         n_majority7_module_107__or_module_11_res,
         n_majority7_module_107__and_module_9_res,
         n_majority7_module_107__or_module_10_res,
         n_majority7_module_107__or_module_9_res,
         n_majority7_module_107__and_module_8_res,
         n_majority7_module_107__or_module_8_res,
         n_majority7_module_107__and_module_7_res,
         n_majority7_module_107__or_module_7_res,
         n_majority7_module_107__or_module_6_res,
         n_majority7_module_107__and_module_6_res,
         n_majority7_module_107__or_module_5_res,
         n_majority7_module_107__and_module_5_res,
         n_majority7_module_107__or_module_4_res,
         n_majority7_module_107__and_module_4_res,
         n_majority7_module_107__or_module_3_res,
         n_majority7_module_107__and_module_3_res,
         n_majority7_module_107__or_module_2_res,
         n_majority7_module_107__and_module_2_res,
         n_majority7_module_107__or_module_1_res,
         n_majority7_module_107__and_module_1_res, n_majority7_module_108_n7,
         n_majority7_module_108_n6, n_majority7_module_108_n5,
         n_majority7_module_108_n4, n_majority7_module_108_n3,
         n_majority7_module_108_n2, n_majority7_module_108_n1,
         n_majority7_module_108__and_module_10_res,
         n_majority7_module_108__or_module_11_res,
         n_majority7_module_108__and_module_9_res,
         n_majority7_module_108__or_module_10_res,
         n_majority7_module_108__or_module_9_res,
         n_majority7_module_108__and_module_8_res,
         n_majority7_module_108__or_module_8_res,
         n_majority7_module_108__and_module_7_res,
         n_majority7_module_108__or_module_7_res,
         n_majority7_module_108__or_module_6_res,
         n_majority7_module_108__and_module_6_res,
         n_majority7_module_108__or_module_5_res,
         n_majority7_module_108__and_module_5_res,
         n_majority7_module_108__or_module_4_res,
         n_majority7_module_108__and_module_4_res,
         n_majority7_module_108__or_module_3_res,
         n_majority7_module_108__and_module_3_res,
         n_majority7_module_108__or_module_2_res,
         n_majority7_module_108__and_module_2_res,
         n_majority7_module_108__or_module_1_res,
         n_majority7_module_108__and_module_1_res, n_majority7_module_109_n7,
         n_majority7_module_109_n6, n_majority7_module_109_n5,
         n_majority7_module_109_n4, n_majority7_module_109_n3,
         n_majority7_module_109_n2, n_majority7_module_109_n1,
         n_majority7_module_109__and_module_10_res,
         n_majority7_module_109__or_module_11_res,
         n_majority7_module_109__and_module_9_res,
         n_majority7_module_109__or_module_10_res,
         n_majority7_module_109__or_module_9_res,
         n_majority7_module_109__and_module_8_res,
         n_majority7_module_109__or_module_8_res,
         n_majority7_module_109__and_module_7_res,
         n_majority7_module_109__or_module_7_res,
         n_majority7_module_109__or_module_6_res,
         n_majority7_module_109__and_module_6_res,
         n_majority7_module_109__or_module_5_res,
         n_majority7_module_109__and_module_5_res,
         n_majority7_module_109__or_module_4_res,
         n_majority7_module_109__and_module_4_res,
         n_majority7_module_109__or_module_3_res,
         n_majority7_module_109__and_module_3_res,
         n_majority7_module_109__or_module_2_res,
         n_majority7_module_109__and_module_2_res,
         n_majority7_module_109__or_module_1_res,
         n_majority7_module_109__and_module_1_res, n_majority7_module_110_n7,
         n_majority7_module_110_n6, n_majority7_module_110_n5,
         n_majority7_module_110_n4, n_majority7_module_110_n3,
         n_majority7_module_110_n2, n_majority7_module_110_n1,
         n_majority7_module_110__and_module_10_res,
         n_majority7_module_110__or_module_11_res,
         n_majority7_module_110__and_module_9_res,
         n_majority7_module_110__or_module_10_res,
         n_majority7_module_110__or_module_9_res,
         n_majority7_module_110__and_module_8_res,
         n_majority7_module_110__or_module_8_res,
         n_majority7_module_110__and_module_7_res,
         n_majority7_module_110__or_module_7_res,
         n_majority7_module_110__or_module_6_res,
         n_majority7_module_110__and_module_6_res,
         n_majority7_module_110__or_module_5_res,
         n_majority7_module_110__and_module_5_res,
         n_majority7_module_110__or_module_4_res,
         n_majority7_module_110__and_module_4_res,
         n_majority7_module_110__or_module_3_res,
         n_majority7_module_110__and_module_3_res,
         n_majority7_module_110__or_module_2_res,
         n_majority7_module_110__and_module_2_res,
         n_majority7_module_110__or_module_1_res,
         n_majority7_module_110__and_module_1_res, n_majority7_module_111_n7,
         n_majority7_module_111_n6, n_majority7_module_111_n5,
         n_majority7_module_111_n4, n_majority7_module_111_n3,
         n_majority7_module_111_n2, n_majority7_module_111_n1,
         n_majority7_module_111__and_module_10_res,
         n_majority7_module_111__or_module_11_res,
         n_majority7_module_111__and_module_9_res,
         n_majority7_module_111__or_module_10_res,
         n_majority7_module_111__or_module_9_res,
         n_majority7_module_111__and_module_8_res,
         n_majority7_module_111__or_module_8_res,
         n_majority7_module_111__and_module_7_res,
         n_majority7_module_111__or_module_7_res,
         n_majority7_module_111__or_module_6_res,
         n_majority7_module_111__and_module_6_res,
         n_majority7_module_111__or_module_5_res,
         n_majority7_module_111__and_module_5_res,
         n_majority7_module_111__or_module_4_res,
         n_majority7_module_111__and_module_4_res,
         n_majority7_module_111__or_module_3_res,
         n_majority7_module_111__and_module_3_res,
         n_majority7_module_111__or_module_2_res,
         n_majority7_module_111__and_module_2_res,
         n_majority7_module_111__or_module_1_res,
         n_majority7_module_111__and_module_1_res;

  XOR2_X1 u_xor_module_1_U1 ( .A(p_rand_0), .B(io_i1_s0_d0), .Z(
        n_xor_module_1_res) );
  XOR2_X1 u_xor_module_2_U1 ( .A(p_rand_1), .B(n_xor_module_1_res), .Z(
        n_xor_module_2_res) );
  INV_X1 u_xor_module_3_U2 ( .A(n_xor_module_3_n2), .ZN(n_xor_module_3_res) );
  XNOR2_X1 u_xor_module_3_U1 ( .A(p_rand_2), .B(n_xor_module_2_res), .ZN(
        n_xor_module_3_n2) );
  XOR2_X1 u_xor_module_4_U1 ( .A(p_rand_0), .B(io_i1_s1_d0), .Z(
        n_xor_module_4_res) );
  XOR2_X1 u_xor_module_5_U1 ( .A(p_rand_3), .B(n_xor_module_4_res), .Z(
        n_xor_module_5_res) );
  INV_X1 u_xor_module_6_U2 ( .A(n_xor_module_6_n2), .ZN(n_xor_module_6_res) );
  XNOR2_X1 u_xor_module_6_U1 ( .A(p_rand_4), .B(n_xor_module_5_res), .ZN(
        n_xor_module_6_n2) );
  XOR2_X1 u_xor_module_7_U1 ( .A(p_rand_1), .B(io_i1_s2_d0), .Z(
        n_xor_module_7_res) );
  XOR2_X1 u_xor_module_8_U1 ( .A(p_rand_3), .B(n_xor_module_7_res), .Z(
        n_xor_module_8_res) );
  INV_X1 u_xor_module_9_U2 ( .A(n_xor_module_9_n2), .ZN(n_xor_module_9_res) );
  XNOR2_X1 u_xor_module_9_U1 ( .A(p_rand_5), .B(n_xor_module_8_res), .ZN(
        n_xor_module_9_n2) );
  XOR2_X1 u_xor_module_10_U1 ( .A(p_rand_2), .B(io_i1_s3_d0), .Z(
        n_xor_module_10_res) );
  XOR2_X1 u_xor_module_11_U1 ( .A(p_rand_4), .B(n_xor_module_10_res), .Z(
        n_xor_module_11_res) );
  INV_X1 u_xor_module_12_U2 ( .A(n_xor_module_12_n2), .ZN(n_xor_module_12_res)
         );
  XNOR2_X1 u_xor_module_12_U1 ( .A(p_rand_5), .B(n_xor_module_11_res), .ZN(
        n_xor_module_12_n2) );
  XOR2_X1 u_xor_module_13_U1 ( .A(p_rand_0), .B(io_i1_s0_d1), .Z(
        n_xor_module_13_res) );
  XOR2_X1 u_xor_module_14_U1 ( .A(p_rand_1), .B(n_xor_module_13_res), .Z(
        n_xor_module_14_res) );
  INV_X1 u_xor_module_15_U2 ( .A(n_xor_module_15_n2), .ZN(n_xor_module_15_res)
         );
  XNOR2_X1 u_xor_module_15_U1 ( .A(p_rand_2), .B(n_xor_module_14_res), .ZN(
        n_xor_module_15_n2) );
  XOR2_X1 u_xor_module_16_U1 ( .A(p_rand_0), .B(io_i1_s1_d1), .Z(
        n_xor_module_16_res) );
  XOR2_X1 u_xor_module_17_U1 ( .A(p_rand_3), .B(n_xor_module_16_res), .Z(
        n_xor_module_17_res) );
  INV_X1 u_xor_module_18_U2 ( .A(n_xor_module_18_n2), .ZN(n_xor_module_18_res)
         );
  XNOR2_X1 u_xor_module_18_U1 ( .A(p_rand_4), .B(n_xor_module_17_res), .ZN(
        n_xor_module_18_n2) );
  XOR2_X1 u_xor_module_19_U1 ( .A(p_rand_1), .B(io_i1_s2_d1), .Z(
        n_xor_module_19_res) );
  XOR2_X1 u_xor_module_20_U1 ( .A(p_rand_3), .B(n_xor_module_19_res), .Z(
        n_xor_module_20_res) );
  INV_X1 u_xor_module_21_U2 ( .A(n_xor_module_21_n2), .ZN(n_xor_module_21_res)
         );
  XNOR2_X1 u_xor_module_21_U1 ( .A(p_rand_5), .B(n_xor_module_20_res), .ZN(
        n_xor_module_21_n2) );
  XOR2_X1 u_xor_module_22_U1 ( .A(p_rand_2), .B(io_i1_s3_d1), .Z(
        n_xor_module_22_res) );
  XOR2_X1 u_xor_module_23_U1 ( .A(p_rand_4), .B(n_xor_module_22_res), .Z(
        n_xor_module_23_res) );
  INV_X1 u_xor_module_24_U2 ( .A(n_xor_module_24_n2), .ZN(n_xor_module_24_res)
         );
  XNOR2_X1 u_xor_module_24_U1 ( .A(p_rand_5), .B(n_xor_module_23_res), .ZN(
        n_xor_module_24_n2) );
  XOR2_X1 u_xor_module_25_U1 ( .A(p_rand_0), .B(io_i1_s0_d2), .Z(
        n_xor_module_25_res) );
  XOR2_X1 u_xor_module_26_U1 ( .A(p_rand_1), .B(n_xor_module_25_res), .Z(
        n_xor_module_26_res) );
  INV_X1 u_xor_module_27_U2 ( .A(n_xor_module_27_n2), .ZN(n_xor_module_27_res)
         );
  XNOR2_X1 u_xor_module_27_U1 ( .A(p_rand_2), .B(n_xor_module_26_res), .ZN(
        n_xor_module_27_n2) );
  XOR2_X1 u_xor_module_28_U1 ( .A(p_rand_0), .B(io_i1_s1_d2), .Z(
        n_xor_module_28_res) );
  XOR2_X1 u_xor_module_29_U1 ( .A(p_rand_3), .B(n_xor_module_28_res), .Z(
        n_xor_module_29_res) );
  INV_X1 u_xor_module_30_U2 ( .A(n_xor_module_30_n2), .ZN(n_xor_module_30_res)
         );
  XNOR2_X1 u_xor_module_30_U1 ( .A(p_rand_4), .B(n_xor_module_29_res), .ZN(
        n_xor_module_30_n2) );
  XOR2_X1 u_xor_module_31_U1 ( .A(p_rand_1), .B(io_i1_s2_d2), .Z(
        n_xor_module_31_res) );
  XOR2_X1 u_xor_module_32_U1 ( .A(p_rand_3), .B(n_xor_module_31_res), .Z(
        n_xor_module_32_res) );
  INV_X1 u_xor_module_33_U2 ( .A(n_xor_module_33_n2), .ZN(n_xor_module_33_res)
         );
  XNOR2_X1 u_xor_module_33_U1 ( .A(p_rand_5), .B(n_xor_module_32_res), .ZN(
        n_xor_module_33_n2) );
  XOR2_X1 u_xor_module_34_U1 ( .A(p_rand_2), .B(io_i1_s3_d2), .Z(
        n_xor_module_34_res) );
  XOR2_X1 u_xor_module_35_U1 ( .A(p_rand_4), .B(n_xor_module_34_res), .Z(
        n_xor_module_35_res) );
  INV_X1 u_xor_module_36_U2 ( .A(n_xor_module_36_n2), .ZN(n_xor_module_36_res)
         );
  XNOR2_X1 u_xor_module_36_U1 ( .A(p_rand_5), .B(n_xor_module_35_res), .ZN(
        n_xor_module_36_n2) );
  XOR2_X1 u_xor_module_37_U1 ( .A(p_rand_0), .B(io_i1_s0_d3), .Z(
        n_xor_module_37_res) );
  XOR2_X1 u_xor_module_38_U1 ( .A(p_rand_1), .B(n_xor_module_37_res), .Z(
        n_xor_module_38_res) );
  INV_X1 u_xor_module_39_U2 ( .A(n_xor_module_39_n2), .ZN(n_xor_module_39_res)
         );
  XNOR2_X1 u_xor_module_39_U1 ( .A(p_rand_2), .B(n_xor_module_38_res), .ZN(
        n_xor_module_39_n2) );
  XOR2_X1 u_xor_module_40_U1 ( .A(p_rand_0), .B(io_i1_s1_d3), .Z(
        n_xor_module_40_res) );
  XOR2_X1 u_xor_module_41_U1 ( .A(p_rand_3), .B(n_xor_module_40_res), .Z(
        n_xor_module_41_res) );
  INV_X1 u_xor_module_42_U2 ( .A(n_xor_module_42_n2), .ZN(n_xor_module_42_res)
         );
  XNOR2_X1 u_xor_module_42_U1 ( .A(p_rand_4), .B(n_xor_module_41_res), .ZN(
        n_xor_module_42_n2) );
  XOR2_X1 u_xor_module_43_U1 ( .A(p_rand_1), .B(io_i1_s2_d3), .Z(
        n_xor_module_43_res) );
  XOR2_X1 u_xor_module_44_U1 ( .A(p_rand_3), .B(n_xor_module_43_res), .Z(
        n_xor_module_44_res) );
  INV_X1 u_xor_module_45_U2 ( .A(n_xor_module_45_n2), .ZN(n_xor_module_45_res)
         );
  XNOR2_X1 u_xor_module_45_U1 ( .A(p_rand_5), .B(n_xor_module_44_res), .ZN(
        n_xor_module_45_n2) );
  XOR2_X1 u_xor_module_46_U1 ( .A(p_rand_2), .B(io_i1_s3_d3), .Z(
        n_xor_module_46_res) );
  XOR2_X1 u_xor_module_47_U1 ( .A(p_rand_4), .B(n_xor_module_46_res), .Z(
        n_xor_module_47_res) );
  INV_X1 u_xor_module_48_U2 ( .A(n_xor_module_48_n2), .ZN(n_xor_module_48_res)
         );
  XNOR2_X1 u_xor_module_48_U1 ( .A(p_rand_5), .B(n_xor_module_47_res), .ZN(
        n_xor_module_48_n2) );
  XOR2_X1 u_xor_module_49_U1 ( .A(p_rand_0), .B(io_i1_s0_d4), .Z(
        n_xor_module_49_res) );
  XOR2_X1 u_xor_module_50_U1 ( .A(p_rand_1), .B(n_xor_module_49_res), .Z(
        n_xor_module_50_res) );
  INV_X1 u_xor_module_51_U2 ( .A(n_xor_module_51_n2), .ZN(n_xor_module_51_res)
         );
  XNOR2_X1 u_xor_module_51_U1 ( .A(p_rand_2), .B(n_xor_module_50_res), .ZN(
        n_xor_module_51_n2) );
  XOR2_X1 u_xor_module_52_U1 ( .A(p_rand_0), .B(io_i1_s1_d4), .Z(
        n_xor_module_52_res) );
  XOR2_X1 u_xor_module_53_U1 ( .A(p_rand_3), .B(n_xor_module_52_res), .Z(
        n_xor_module_53_res) );
  INV_X1 u_xor_module_54_U2 ( .A(n_xor_module_54_n2), .ZN(n_xor_module_54_res)
         );
  XNOR2_X1 u_xor_module_54_U1 ( .A(p_rand_4), .B(n_xor_module_53_res), .ZN(
        n_xor_module_54_n2) );
  XOR2_X1 u_xor_module_55_U1 ( .A(p_rand_1), .B(io_i1_s2_d4), .Z(
        n_xor_module_55_res) );
  XOR2_X1 u_xor_module_56_U1 ( .A(p_rand_3), .B(n_xor_module_55_res), .Z(
        n_xor_module_56_res) );
  INV_X1 u_xor_module_57_U2 ( .A(n_xor_module_57_n2), .ZN(n_xor_module_57_res)
         );
  XNOR2_X1 u_xor_module_57_U1 ( .A(p_rand_5), .B(n_xor_module_56_res), .ZN(
        n_xor_module_57_n2) );
  XOR2_X1 u_xor_module_58_U1 ( .A(p_rand_2), .B(io_i1_s3_d4), .Z(
        n_xor_module_58_res) );
  XOR2_X1 u_xor_module_59_U1 ( .A(p_rand_4), .B(n_xor_module_58_res), .Z(
        n_xor_module_59_res) );
  INV_X1 u_xor_module_60_U2 ( .A(n_xor_module_60_n2), .ZN(n_xor_module_60_res)
         );
  XNOR2_X1 u_xor_module_60_U1 ( .A(p_rand_5), .B(n_xor_module_59_res), .ZN(
        n_xor_module_60_n2) );
  XOR2_X1 u_xor_module_61_U1 ( .A(p_rand_0), .B(io_i1_s0_d5), .Z(
        n_xor_module_61_res) );
  XOR2_X1 u_xor_module_62_U1 ( .A(p_rand_1), .B(n_xor_module_61_res), .Z(
        n_xor_module_62_res) );
  INV_X1 u_xor_module_63_U2 ( .A(n_xor_module_63_n2), .ZN(n_xor_module_63_res)
         );
  XNOR2_X1 u_xor_module_63_U1 ( .A(p_rand_2), .B(n_xor_module_62_res), .ZN(
        n_xor_module_63_n2) );
  XOR2_X1 u_xor_module_64_U1 ( .A(p_rand_0), .B(io_i1_s1_d5), .Z(
        n_xor_module_64_res) );
  XOR2_X1 u_xor_module_65_U1 ( .A(p_rand_3), .B(n_xor_module_64_res), .Z(
        n_xor_module_65_res) );
  INV_X1 u_xor_module_66_U2 ( .A(n_xor_module_66_n2), .ZN(n_xor_module_66_res)
         );
  XNOR2_X1 u_xor_module_66_U1 ( .A(p_rand_4), .B(n_xor_module_65_res), .ZN(
        n_xor_module_66_n2) );
  XOR2_X1 u_xor_module_67_U1 ( .A(p_rand_1), .B(io_i1_s2_d5), .Z(
        n_xor_module_67_res) );
  XOR2_X1 u_xor_module_68_U1 ( .A(p_rand_3), .B(n_xor_module_67_res), .Z(
        n_xor_module_68_res) );
  INV_X1 u_xor_module_69_U2 ( .A(n_xor_module_69_n2), .ZN(n_xor_module_69_res)
         );
  XNOR2_X1 u_xor_module_69_U1 ( .A(p_rand_5), .B(n_xor_module_68_res), .ZN(
        n_xor_module_69_n2) );
  XOR2_X1 u_xor_module_70_U1 ( .A(p_rand_2), .B(io_i1_s3_d5), .Z(
        n_xor_module_70_res) );
  XOR2_X1 u_xor_module_71_U1 ( .A(p_rand_4), .B(n_xor_module_70_res), .Z(
        n_xor_module_71_res) );
  INV_X1 u_xor_module_72_U2 ( .A(n_xor_module_72_n2), .ZN(n_xor_module_72_res)
         );
  XNOR2_X1 u_xor_module_72_U1 ( .A(p_rand_5), .B(n_xor_module_71_res), .ZN(
        n_xor_module_72_n2) );
  XOR2_X1 u_xor_module_73_U1 ( .A(p_rand_0), .B(io_i1_s0_d6), .Z(
        n_xor_module_73_res) );
  XOR2_X1 u_xor_module_74_U1 ( .A(p_rand_1), .B(n_xor_module_73_res), .Z(
        n_xor_module_74_res) );
  INV_X1 u_xor_module_75_U2 ( .A(n_xor_module_75_n2), .ZN(n_xor_module_75_res)
         );
  XNOR2_X1 u_xor_module_75_U1 ( .A(p_rand_2), .B(n_xor_module_74_res), .ZN(
        n_xor_module_75_n2) );
  XOR2_X1 u_xor_module_76_U1 ( .A(p_rand_0), .B(io_i1_s1_d6), .Z(
        n_xor_module_76_res) );
  XOR2_X1 u_xor_module_77_U1 ( .A(p_rand_3), .B(n_xor_module_76_res), .Z(
        n_xor_module_77_res) );
  INV_X1 u_xor_module_78_U2 ( .A(n_xor_module_78_n2), .ZN(n_xor_module_78_res)
         );
  XNOR2_X1 u_xor_module_78_U1 ( .A(p_rand_4), .B(n_xor_module_77_res), .ZN(
        n_xor_module_78_n2) );
  XOR2_X1 u_xor_module_79_U1 ( .A(p_rand_1), .B(io_i1_s2_d6), .Z(
        n_xor_module_79_res) );
  XOR2_X1 u_xor_module_80_U1 ( .A(p_rand_3), .B(n_xor_module_79_res), .Z(
        n_xor_module_80_res) );
  INV_X1 u_xor_module_81_U2 ( .A(n_xor_module_81_n2), .ZN(n_xor_module_81_res)
         );
  XNOR2_X1 u_xor_module_81_U1 ( .A(p_rand_5), .B(n_xor_module_80_res), .ZN(
        n_xor_module_81_n2) );
  XOR2_X1 u_xor_module_82_U1 ( .A(p_rand_2), .B(io_i1_s3_d6), .Z(
        n_xor_module_82_res) );
  XOR2_X1 u_xor_module_83_U1 ( .A(p_rand_4), .B(n_xor_module_82_res), .Z(
        n_xor_module_83_res) );
  INV_X1 u_xor_module_84_U2 ( .A(n_xor_module_84_n2), .ZN(n_xor_module_84_res)
         );
  XNOR2_X1 u_xor_module_84_U1 ( .A(p_rand_5), .B(n_xor_module_83_res), .ZN(
        n_xor_module_84_n2) );
  BUF_X1 u_majority7_module_0_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_0_n7) );
  BUF_X1 u_majority7_module_0_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_0_n6) );
  BUF_X1 u_majority7_module_0_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_0_n5) );
  BUF_X1 u_majority7_module_0_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_0_n4) );
  BUF_X1 u_majority7_module_0_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_0_n3) );
  BUF_X1 u_majority7_module_0_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_0_n2) );
  BUF_X1 u_majority7_module_0_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_0_n1) );
  AND2_X1 u_majority7_module_0__and_module_1_U1 ( .A1(n_majority7_module_0_n5), 
        .A2(n_majority7_module_0_n4), .ZN(
        n_majority7_module_0__and_module_1_res) );
  OR2_X1 u_majority7_module_0__or_module_1_U1 ( .A1(n_majority7_module_0_n4), 
        .A2(n_majority7_module_0_n5), .ZN(
        n_majority7_module_0__or_module_1_res) );
  AND2_X1 u_majority7_module_0__and_module_2_U1 ( .A1(n_majority7_module_0_n7), 
        .A2(n_majority7_module_0_n2), .ZN(
        n_majority7_module_0__and_module_2_res) );
  OR2_X1 u_majority7_module_0__or_module_2_U1 ( .A1(n_majority7_module_0_n2), 
        .A2(n_majority7_module_0_n7), .ZN(
        n_majority7_module_0__or_module_2_res) );
  AND2_X1 u_majority7_module_0__and_module_3_U1 ( .A1(n_majority7_module_0_n6), 
        .A2(n_majority7_module_0_n1), .ZN(
        n_majority7_module_0__and_module_3_res) );
  OR2_X1 u_majority7_module_0__or_module_3_U1 ( .A1(n_majority7_module_0_n1), 
        .A2(n_majority7_module_0_n6), .ZN(
        n_majority7_module_0__or_module_3_res) );
  AND2_X1 u_majority7_module_0__and_module_4_U1 ( .A1(
        n_majority7_module_0__and_module_2_res), .A2(
        n_majority7_module_0__and_module_1_res), .ZN(
        n_majority7_module_0__and_module_4_res) );
  OR2_X1 u_majority7_module_0__or_module_4_U1 ( .A1(
        n_majority7_module_0__and_module_1_res), .A2(
        n_majority7_module_0__and_module_2_res), .ZN(
        n_majority7_module_0__or_module_4_res) );
  AND2_X1 u_majority7_module_0__and_module_5_U1 ( .A1(
        n_majority7_module_0__and_module_3_res), .A2(n_majority7_module_0_n3), 
        .ZN(n_majority7_module_0__and_module_5_res) );
  OR2_X1 u_majority7_module_0__or_module_5_U1 ( .A1(n_majority7_module_0_n3), 
        .A2(n_majority7_module_0__and_module_3_res), .ZN(
        n_majority7_module_0__or_module_5_res) );
  AND2_X1 u_majority7_module_0__and_module_6_U1 ( .A1(
        n_majority7_module_0__or_module_1_res), .A2(
        n_majority7_module_0__or_module_2_res), .ZN(
        n_majority7_module_0__and_module_6_res) );
  OR2_X1 u_majority7_module_0__or_module_6_U1 ( .A1(
        n_majority7_module_0__or_module_2_res), .A2(
        n_majority7_module_0__or_module_1_res), .ZN(
        n_majority7_module_0__or_module_6_res) );
  OR2_X1 u_majority7_module_0__or_module_7_U1 ( .A1(
        n_majority7_module_0__and_module_4_res), .A2(
        n_majority7_module_0__and_module_5_res), .ZN(
        n_majority7_module_0__or_module_7_res) );
  AND2_X1 u_majority7_module_0__and_module_7_U1 ( .A1(
        n_majority7_module_0__or_module_3_res), .A2(
        n_majority7_module_0__or_module_4_res), .ZN(
        n_majority7_module_0__and_module_7_res) );
  OR2_X1 u_majority7_module_0__or_module_8_U1 ( .A1(
        n_majority7_module_0__or_module_4_res), .A2(
        n_majority7_module_0__or_module_3_res), .ZN(
        n_majority7_module_0__or_module_8_res) );
  AND2_X1 u_majority7_module_0__and_module_8_U1 ( .A1(
        n_majority7_module_0__or_module_5_res), .A2(
        n_majority7_module_0__and_module_6_res), .ZN(
        n_majority7_module_0__and_module_8_res) );
  OR2_X1 u_majority7_module_0__or_module_9_U1 ( .A1(
        n_majority7_module_0__and_module_6_res), .A2(
        n_majority7_module_0__or_module_5_res), .ZN(
        n_majority7_module_0__or_module_9_res) );
  OR2_X1 u_majority7_module_0__or_module_10_U1 ( .A1(
        n_majority7_module_0__or_module_7_res), .A2(
        n_majority7_module_0__and_module_7_res), .ZN(
        n_majority7_module_0__or_module_10_res) );
  AND2_X1 u_majority7_module_0__and_module_9_U1 ( .A1(
        n_majority7_module_0__or_module_6_res), .A2(
        n_majority7_module_0__or_module_9_res), .ZN(
        n_majority7_module_0__and_module_9_res) );
  OR2_X1 u_majority7_module_0__or_module_11_U1 ( .A1(
        n_majority7_module_0__or_module_10_res), .A2(
        n_majority7_module_0__and_module_8_res), .ZN(
        n_majority7_module_0__or_module_11_res) );
  AND2_X1 u_majority7_module_0__and_module_10_U1 ( .A1(
        n_majority7_module_0__or_module_8_res), .A2(
        n_majority7_module_0__and_module_9_res), .ZN(
        n_majority7_module_0__and_module_10_res) );
  AND2_X1 u_majority7_module_0__and_module_11_U1 ( .A1(
        n_majority7_module_0__and_module_10_res), .A2(
        n_majority7_module_0__or_module_11_res), .ZN(n_majority7_module_0_res)
         );
  DFF_X1 u_reg_module_1__cini_mul_v000_reg ( .D(n_majority7_module_0_res), 
        .CK(clock_0), .Q(n_reg_module_1_res), .QN() );
  BUF_X1 u_majority7_module_1_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_1_n7) );
  BUF_X1 u_majority7_module_1_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_1_n6) );
  BUF_X1 u_majority7_module_1_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_1_n5) );
  BUF_X1 u_majority7_module_1_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_1_n4) );
  BUF_X1 u_majority7_module_1_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_1_n3) );
  BUF_X1 u_majority7_module_1_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_1_n2) );
  BUF_X1 u_majority7_module_1_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_1_n1) );
  AND2_X1 u_majority7_module_1__and_module_1_U1 ( .A1(n_majority7_module_1_n5), 
        .A2(n_majority7_module_1_n4), .ZN(
        n_majority7_module_1__and_module_1_res) );
  OR2_X1 u_majority7_module_1__or_module_1_U1 ( .A1(n_majority7_module_1_n4), 
        .A2(n_majority7_module_1_n5), .ZN(
        n_majority7_module_1__or_module_1_res) );
  AND2_X1 u_majority7_module_1__and_module_2_U1 ( .A1(n_majority7_module_1_n7), 
        .A2(n_majority7_module_1_n2), .ZN(
        n_majority7_module_1__and_module_2_res) );
  OR2_X1 u_majority7_module_1__or_module_2_U1 ( .A1(n_majority7_module_1_n2), 
        .A2(n_majority7_module_1_n7), .ZN(
        n_majority7_module_1__or_module_2_res) );
  AND2_X1 u_majority7_module_1__and_module_3_U1 ( .A1(n_majority7_module_1_n6), 
        .A2(n_majority7_module_1_n1), .ZN(
        n_majority7_module_1__and_module_3_res) );
  OR2_X1 u_majority7_module_1__or_module_3_U1 ( .A1(n_majority7_module_1_n1), 
        .A2(n_majority7_module_1_n6), .ZN(
        n_majority7_module_1__or_module_3_res) );
  AND2_X1 u_majority7_module_1__and_module_4_U1 ( .A1(
        n_majority7_module_1__and_module_2_res), .A2(
        n_majority7_module_1__and_module_1_res), .ZN(
        n_majority7_module_1__and_module_4_res) );
  OR2_X1 u_majority7_module_1__or_module_4_U1 ( .A1(
        n_majority7_module_1__and_module_1_res), .A2(
        n_majority7_module_1__and_module_2_res), .ZN(
        n_majority7_module_1__or_module_4_res) );
  AND2_X1 u_majority7_module_1__and_module_5_U1 ( .A1(
        n_majority7_module_1__and_module_3_res), .A2(n_majority7_module_1_n3), 
        .ZN(n_majority7_module_1__and_module_5_res) );
  OR2_X1 u_majority7_module_1__or_module_5_U1 ( .A1(n_majority7_module_1_n3), 
        .A2(n_majority7_module_1__and_module_3_res), .ZN(
        n_majority7_module_1__or_module_5_res) );
  AND2_X1 u_majority7_module_1__and_module_6_U1 ( .A1(
        n_majority7_module_1__or_module_1_res), .A2(
        n_majority7_module_1__or_module_2_res), .ZN(
        n_majority7_module_1__and_module_6_res) );
  OR2_X1 u_majority7_module_1__or_module_6_U1 ( .A1(
        n_majority7_module_1__or_module_2_res), .A2(
        n_majority7_module_1__or_module_1_res), .ZN(
        n_majority7_module_1__or_module_6_res) );
  OR2_X1 u_majority7_module_1__or_module_7_U1 ( .A1(
        n_majority7_module_1__and_module_4_res), .A2(
        n_majority7_module_1__and_module_5_res), .ZN(
        n_majority7_module_1__or_module_7_res) );
  AND2_X1 u_majority7_module_1__and_module_7_U1 ( .A1(
        n_majority7_module_1__or_module_3_res), .A2(
        n_majority7_module_1__or_module_4_res), .ZN(
        n_majority7_module_1__and_module_7_res) );
  OR2_X1 u_majority7_module_1__or_module_8_U1 ( .A1(
        n_majority7_module_1__or_module_4_res), .A2(
        n_majority7_module_1__or_module_3_res), .ZN(
        n_majority7_module_1__or_module_8_res) );
  AND2_X1 u_majority7_module_1__and_module_8_U1 ( .A1(
        n_majority7_module_1__or_module_5_res), .A2(
        n_majority7_module_1__and_module_6_res), .ZN(
        n_majority7_module_1__and_module_8_res) );
  OR2_X1 u_majority7_module_1__or_module_9_U1 ( .A1(
        n_majority7_module_1__and_module_6_res), .A2(
        n_majority7_module_1__or_module_5_res), .ZN(
        n_majority7_module_1__or_module_9_res) );
  OR2_X1 u_majority7_module_1__or_module_10_U1 ( .A1(
        n_majority7_module_1__or_module_7_res), .A2(
        n_majority7_module_1__and_module_7_res), .ZN(
        n_majority7_module_1__or_module_10_res) );
  AND2_X1 u_majority7_module_1__and_module_9_U1 ( .A1(
        n_majority7_module_1__or_module_6_res), .A2(
        n_majority7_module_1__or_module_9_res), .ZN(
        n_majority7_module_1__and_module_9_res) );
  OR2_X1 u_majority7_module_1__or_module_11_U1 ( .A1(
        n_majority7_module_1__or_module_10_res), .A2(
        n_majority7_module_1__and_module_8_res), .ZN(
        n_majority7_module_1__or_module_11_res) );
  AND2_X1 u_majority7_module_1__and_module_10_U1 ( .A1(
        n_majority7_module_1__or_module_8_res), .A2(
        n_majority7_module_1__and_module_9_res), .ZN(
        n_majority7_module_1__and_module_10_res) );
  AND2_X1 u_majority7_module_1__and_module_11_U1 ( .A1(
        n_majority7_module_1__and_module_10_res), .A2(
        n_majority7_module_1__or_module_11_res), .ZN(n_majority7_module_1_res)
         );
  DFF_X1 u_reg_module_2__cini_mul_v000_reg ( .D(n_majority7_module_1_res), 
        .CK(clock_0), .Q(n_reg_module_2_res), .QN() );
  BUF_X1 u_majority7_module_2_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_2_n7) );
  BUF_X1 u_majority7_module_2_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_2_n6) );
  BUF_X1 u_majority7_module_2_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_2_n5) );
  BUF_X1 u_majority7_module_2_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_2_n4) );
  BUF_X1 u_majority7_module_2_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_2_n3) );
  BUF_X1 u_majority7_module_2_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_2_n2) );
  BUF_X1 u_majority7_module_2_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_2_n1) );
  AND2_X1 u_majority7_module_2__and_module_1_U1 ( .A1(n_majority7_module_2_n5), 
        .A2(n_majority7_module_2_n4), .ZN(
        n_majority7_module_2__and_module_1_res) );
  OR2_X1 u_majority7_module_2__or_module_1_U1 ( .A1(n_majority7_module_2_n4), 
        .A2(n_majority7_module_2_n5), .ZN(
        n_majority7_module_2__or_module_1_res) );
  AND2_X1 u_majority7_module_2__and_module_2_U1 ( .A1(n_majority7_module_2_n7), 
        .A2(n_majority7_module_2_n2), .ZN(
        n_majority7_module_2__and_module_2_res) );
  OR2_X1 u_majority7_module_2__or_module_2_U1 ( .A1(n_majority7_module_2_n2), 
        .A2(n_majority7_module_2_n7), .ZN(
        n_majority7_module_2__or_module_2_res) );
  AND2_X1 u_majority7_module_2__and_module_3_U1 ( .A1(n_majority7_module_2_n6), 
        .A2(n_majority7_module_2_n1), .ZN(
        n_majority7_module_2__and_module_3_res) );
  OR2_X1 u_majority7_module_2__or_module_3_U1 ( .A1(n_majority7_module_2_n1), 
        .A2(n_majority7_module_2_n6), .ZN(
        n_majority7_module_2__or_module_3_res) );
  AND2_X1 u_majority7_module_2__and_module_4_U1 ( .A1(
        n_majority7_module_2__and_module_2_res), .A2(
        n_majority7_module_2__and_module_1_res), .ZN(
        n_majority7_module_2__and_module_4_res) );
  OR2_X1 u_majority7_module_2__or_module_4_U1 ( .A1(
        n_majority7_module_2__and_module_1_res), .A2(
        n_majority7_module_2__and_module_2_res), .ZN(
        n_majority7_module_2__or_module_4_res) );
  AND2_X1 u_majority7_module_2__and_module_5_U1 ( .A1(
        n_majority7_module_2__and_module_3_res), .A2(n_majority7_module_2_n3), 
        .ZN(n_majority7_module_2__and_module_5_res) );
  OR2_X1 u_majority7_module_2__or_module_5_U1 ( .A1(n_majority7_module_2_n3), 
        .A2(n_majority7_module_2__and_module_3_res), .ZN(
        n_majority7_module_2__or_module_5_res) );
  AND2_X1 u_majority7_module_2__and_module_6_U1 ( .A1(
        n_majority7_module_2__or_module_1_res), .A2(
        n_majority7_module_2__or_module_2_res), .ZN(
        n_majority7_module_2__and_module_6_res) );
  OR2_X1 u_majority7_module_2__or_module_6_U1 ( .A1(
        n_majority7_module_2__or_module_2_res), .A2(
        n_majority7_module_2__or_module_1_res), .ZN(
        n_majority7_module_2__or_module_6_res) );
  OR2_X1 u_majority7_module_2__or_module_7_U1 ( .A1(
        n_majority7_module_2__and_module_4_res), .A2(
        n_majority7_module_2__and_module_5_res), .ZN(
        n_majority7_module_2__or_module_7_res) );
  AND2_X1 u_majority7_module_2__and_module_7_U1 ( .A1(
        n_majority7_module_2__or_module_3_res), .A2(
        n_majority7_module_2__or_module_4_res), .ZN(
        n_majority7_module_2__and_module_7_res) );
  OR2_X1 u_majority7_module_2__or_module_8_U1 ( .A1(
        n_majority7_module_2__or_module_4_res), .A2(
        n_majority7_module_2__or_module_3_res), .ZN(
        n_majority7_module_2__or_module_8_res) );
  AND2_X1 u_majority7_module_2__and_module_8_U1 ( .A1(
        n_majority7_module_2__or_module_5_res), .A2(
        n_majority7_module_2__and_module_6_res), .ZN(
        n_majority7_module_2__and_module_8_res) );
  OR2_X1 u_majority7_module_2__or_module_9_U1 ( .A1(
        n_majority7_module_2__and_module_6_res), .A2(
        n_majority7_module_2__or_module_5_res), .ZN(
        n_majority7_module_2__or_module_9_res) );
  OR2_X1 u_majority7_module_2__or_module_10_U1 ( .A1(
        n_majority7_module_2__or_module_7_res), .A2(
        n_majority7_module_2__and_module_7_res), .ZN(
        n_majority7_module_2__or_module_10_res) );
  AND2_X1 u_majority7_module_2__and_module_9_U1 ( .A1(
        n_majority7_module_2__or_module_6_res), .A2(
        n_majority7_module_2__or_module_9_res), .ZN(
        n_majority7_module_2__and_module_9_res) );
  OR2_X1 u_majority7_module_2__or_module_11_U1 ( .A1(
        n_majority7_module_2__or_module_10_res), .A2(
        n_majority7_module_2__and_module_8_res), .ZN(
        n_majority7_module_2__or_module_11_res) );
  AND2_X1 u_majority7_module_2__and_module_10_U1 ( .A1(
        n_majority7_module_2__or_module_8_res), .A2(
        n_majority7_module_2__and_module_9_res), .ZN(
        n_majority7_module_2__and_module_10_res) );
  AND2_X1 u_majority7_module_2__and_module_11_U1 ( .A1(
        n_majority7_module_2__and_module_10_res), .A2(
        n_majority7_module_2__or_module_11_res), .ZN(n_majority7_module_2_res)
         );
  DFF_X1 u_reg_module_3__cini_mul_v000_reg ( .D(n_majority7_module_2_res), 
        .CK(clock_0), .Q(n_reg_module_3_res), .QN() );
  BUF_X1 u_majority7_module_3_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_3_n7) );
  BUF_X1 u_majority7_module_3_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_3_n6) );
  BUF_X1 u_majority7_module_3_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_3_n5) );
  BUF_X1 u_majority7_module_3_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_3_n4) );
  BUF_X1 u_majority7_module_3_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_3_n3) );
  BUF_X1 u_majority7_module_3_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_3_n2) );
  BUF_X1 u_majority7_module_3_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_3_n1) );
  AND2_X1 u_majority7_module_3__and_module_1_U1 ( .A1(n_majority7_module_3_n5), 
        .A2(n_majority7_module_3_n4), .ZN(
        n_majority7_module_3__and_module_1_res) );
  OR2_X1 u_majority7_module_3__or_module_1_U1 ( .A1(n_majority7_module_3_n4), 
        .A2(n_majority7_module_3_n5), .ZN(
        n_majority7_module_3__or_module_1_res) );
  AND2_X1 u_majority7_module_3__and_module_2_U1 ( .A1(n_majority7_module_3_n7), 
        .A2(n_majority7_module_3_n2), .ZN(
        n_majority7_module_3__and_module_2_res) );
  OR2_X1 u_majority7_module_3__or_module_2_U1 ( .A1(n_majority7_module_3_n2), 
        .A2(n_majority7_module_3_n7), .ZN(
        n_majority7_module_3__or_module_2_res) );
  AND2_X1 u_majority7_module_3__and_module_3_U1 ( .A1(n_majority7_module_3_n6), 
        .A2(n_majority7_module_3_n1), .ZN(
        n_majority7_module_3__and_module_3_res) );
  OR2_X1 u_majority7_module_3__or_module_3_U1 ( .A1(n_majority7_module_3_n1), 
        .A2(n_majority7_module_3_n6), .ZN(
        n_majority7_module_3__or_module_3_res) );
  AND2_X1 u_majority7_module_3__and_module_4_U1 ( .A1(
        n_majority7_module_3__and_module_2_res), .A2(
        n_majority7_module_3__and_module_1_res), .ZN(
        n_majority7_module_3__and_module_4_res) );
  OR2_X1 u_majority7_module_3__or_module_4_U1 ( .A1(
        n_majority7_module_3__and_module_1_res), .A2(
        n_majority7_module_3__and_module_2_res), .ZN(
        n_majority7_module_3__or_module_4_res) );
  AND2_X1 u_majority7_module_3__and_module_5_U1 ( .A1(
        n_majority7_module_3__and_module_3_res), .A2(n_majority7_module_3_n3), 
        .ZN(n_majority7_module_3__and_module_5_res) );
  OR2_X1 u_majority7_module_3__or_module_5_U1 ( .A1(n_majority7_module_3_n3), 
        .A2(n_majority7_module_3__and_module_3_res), .ZN(
        n_majority7_module_3__or_module_5_res) );
  AND2_X1 u_majority7_module_3__and_module_6_U1 ( .A1(
        n_majority7_module_3__or_module_1_res), .A2(
        n_majority7_module_3__or_module_2_res), .ZN(
        n_majority7_module_3__and_module_6_res) );
  OR2_X1 u_majority7_module_3__or_module_6_U1 ( .A1(
        n_majority7_module_3__or_module_2_res), .A2(
        n_majority7_module_3__or_module_1_res), .ZN(
        n_majority7_module_3__or_module_6_res) );
  OR2_X1 u_majority7_module_3__or_module_7_U1 ( .A1(
        n_majority7_module_3__and_module_4_res), .A2(
        n_majority7_module_3__and_module_5_res), .ZN(
        n_majority7_module_3__or_module_7_res) );
  AND2_X1 u_majority7_module_3__and_module_7_U1 ( .A1(
        n_majority7_module_3__or_module_3_res), .A2(
        n_majority7_module_3__or_module_4_res), .ZN(
        n_majority7_module_3__and_module_7_res) );
  OR2_X1 u_majority7_module_3__or_module_8_U1 ( .A1(
        n_majority7_module_3__or_module_4_res), .A2(
        n_majority7_module_3__or_module_3_res), .ZN(
        n_majority7_module_3__or_module_8_res) );
  AND2_X1 u_majority7_module_3__and_module_8_U1 ( .A1(
        n_majority7_module_3__or_module_5_res), .A2(
        n_majority7_module_3__and_module_6_res), .ZN(
        n_majority7_module_3__and_module_8_res) );
  OR2_X1 u_majority7_module_3__or_module_9_U1 ( .A1(
        n_majority7_module_3__and_module_6_res), .A2(
        n_majority7_module_3__or_module_5_res), .ZN(
        n_majority7_module_3__or_module_9_res) );
  OR2_X1 u_majority7_module_3__or_module_10_U1 ( .A1(
        n_majority7_module_3__or_module_7_res), .A2(
        n_majority7_module_3__and_module_7_res), .ZN(
        n_majority7_module_3__or_module_10_res) );
  AND2_X1 u_majority7_module_3__and_module_9_U1 ( .A1(
        n_majority7_module_3__or_module_6_res), .A2(
        n_majority7_module_3__or_module_9_res), .ZN(
        n_majority7_module_3__and_module_9_res) );
  OR2_X1 u_majority7_module_3__or_module_11_U1 ( .A1(
        n_majority7_module_3__or_module_10_res), .A2(
        n_majority7_module_3__and_module_8_res), .ZN(
        n_majority7_module_3__or_module_11_res) );
  AND2_X1 u_majority7_module_3__and_module_10_U1 ( .A1(
        n_majority7_module_3__or_module_8_res), .A2(
        n_majority7_module_3__and_module_9_res), .ZN(
        n_majority7_module_3__and_module_10_res) );
  AND2_X1 u_majority7_module_3__and_module_11_U1 ( .A1(
        n_majority7_module_3__and_module_10_res), .A2(
        n_majority7_module_3__or_module_11_res), .ZN(n_majority7_module_3_res)
         );
  DFF_X1 u_reg_module_4__cini_mul_v000_reg ( .D(n_majority7_module_3_res), 
        .CK(clock_0), .Q(n_reg_module_4_res), .QN() );
  BUF_X1 u_majority7_module_4_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_4_n7) );
  BUF_X1 u_majority7_module_4_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_4_n6) );
  BUF_X1 u_majority7_module_4_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_4_n5) );
  BUF_X1 u_majority7_module_4_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_4_n4) );
  BUF_X1 u_majority7_module_4_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_4_n3) );
  BUF_X1 u_majority7_module_4_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_4_n2) );
  BUF_X1 u_majority7_module_4_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_4_n1) );
  AND2_X1 u_majority7_module_4__and_module_1_U1 ( .A1(n_majority7_module_4_n5), 
        .A2(n_majority7_module_4_n4), .ZN(
        n_majority7_module_4__and_module_1_res) );
  OR2_X1 u_majority7_module_4__or_module_1_U1 ( .A1(n_majority7_module_4_n4), 
        .A2(n_majority7_module_4_n5), .ZN(
        n_majority7_module_4__or_module_1_res) );
  AND2_X1 u_majority7_module_4__and_module_2_U1 ( .A1(n_majority7_module_4_n7), 
        .A2(n_majority7_module_4_n2), .ZN(
        n_majority7_module_4__and_module_2_res) );
  OR2_X1 u_majority7_module_4__or_module_2_U1 ( .A1(n_majority7_module_4_n2), 
        .A2(n_majority7_module_4_n7), .ZN(
        n_majority7_module_4__or_module_2_res) );
  AND2_X1 u_majority7_module_4__and_module_3_U1 ( .A1(n_majority7_module_4_n6), 
        .A2(n_majority7_module_4_n1), .ZN(
        n_majority7_module_4__and_module_3_res) );
  OR2_X1 u_majority7_module_4__or_module_3_U1 ( .A1(n_majority7_module_4_n1), 
        .A2(n_majority7_module_4_n6), .ZN(
        n_majority7_module_4__or_module_3_res) );
  AND2_X1 u_majority7_module_4__and_module_4_U1 ( .A1(
        n_majority7_module_4__and_module_2_res), .A2(
        n_majority7_module_4__and_module_1_res), .ZN(
        n_majority7_module_4__and_module_4_res) );
  OR2_X1 u_majority7_module_4__or_module_4_U1 ( .A1(
        n_majority7_module_4__and_module_1_res), .A2(
        n_majority7_module_4__and_module_2_res), .ZN(
        n_majority7_module_4__or_module_4_res) );
  AND2_X1 u_majority7_module_4__and_module_5_U1 ( .A1(
        n_majority7_module_4__and_module_3_res), .A2(n_majority7_module_4_n3), 
        .ZN(n_majority7_module_4__and_module_5_res) );
  OR2_X1 u_majority7_module_4__or_module_5_U1 ( .A1(n_majority7_module_4_n3), 
        .A2(n_majority7_module_4__and_module_3_res), .ZN(
        n_majority7_module_4__or_module_5_res) );
  AND2_X1 u_majority7_module_4__and_module_6_U1 ( .A1(
        n_majority7_module_4__or_module_1_res), .A2(
        n_majority7_module_4__or_module_2_res), .ZN(
        n_majority7_module_4__and_module_6_res) );
  OR2_X1 u_majority7_module_4__or_module_6_U1 ( .A1(
        n_majority7_module_4__or_module_2_res), .A2(
        n_majority7_module_4__or_module_1_res), .ZN(
        n_majority7_module_4__or_module_6_res) );
  OR2_X1 u_majority7_module_4__or_module_7_U1 ( .A1(
        n_majority7_module_4__and_module_4_res), .A2(
        n_majority7_module_4__and_module_5_res), .ZN(
        n_majority7_module_4__or_module_7_res) );
  AND2_X1 u_majority7_module_4__and_module_7_U1 ( .A1(
        n_majority7_module_4__or_module_3_res), .A2(
        n_majority7_module_4__or_module_4_res), .ZN(
        n_majority7_module_4__and_module_7_res) );
  OR2_X1 u_majority7_module_4__or_module_8_U1 ( .A1(
        n_majority7_module_4__or_module_4_res), .A2(
        n_majority7_module_4__or_module_3_res), .ZN(
        n_majority7_module_4__or_module_8_res) );
  AND2_X1 u_majority7_module_4__and_module_8_U1 ( .A1(
        n_majority7_module_4__or_module_5_res), .A2(
        n_majority7_module_4__and_module_6_res), .ZN(
        n_majority7_module_4__and_module_8_res) );
  OR2_X1 u_majority7_module_4__or_module_9_U1 ( .A1(
        n_majority7_module_4__and_module_6_res), .A2(
        n_majority7_module_4__or_module_5_res), .ZN(
        n_majority7_module_4__or_module_9_res) );
  OR2_X1 u_majority7_module_4__or_module_10_U1 ( .A1(
        n_majority7_module_4__or_module_7_res), .A2(
        n_majority7_module_4__and_module_7_res), .ZN(
        n_majority7_module_4__or_module_10_res) );
  AND2_X1 u_majority7_module_4__and_module_9_U1 ( .A1(
        n_majority7_module_4__or_module_6_res), .A2(
        n_majority7_module_4__or_module_9_res), .ZN(
        n_majority7_module_4__and_module_9_res) );
  OR2_X1 u_majority7_module_4__or_module_11_U1 ( .A1(
        n_majority7_module_4__or_module_10_res), .A2(
        n_majority7_module_4__and_module_8_res), .ZN(
        n_majority7_module_4__or_module_11_res) );
  AND2_X1 u_majority7_module_4__and_module_10_U1 ( .A1(
        n_majority7_module_4__or_module_8_res), .A2(
        n_majority7_module_4__and_module_9_res), .ZN(
        n_majority7_module_4__and_module_10_res) );
  AND2_X1 u_majority7_module_4__and_module_11_U1 ( .A1(
        n_majority7_module_4__and_module_10_res), .A2(
        n_majority7_module_4__or_module_11_res), .ZN(n_majority7_module_4_res)
         );
  DFF_X1 u_reg_module_5__cini_mul_v000_reg ( .D(n_majority7_module_4_res), 
        .CK(clock_0), .Q(n_reg_module_5_res), .QN() );
  BUF_X1 u_majority7_module_5_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_5_n7) );
  BUF_X1 u_majority7_module_5_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_5_n6) );
  BUF_X1 u_majority7_module_5_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_5_n5) );
  BUF_X1 u_majority7_module_5_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_5_n4) );
  BUF_X1 u_majority7_module_5_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_5_n3) );
  BUF_X1 u_majority7_module_5_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_5_n2) );
  BUF_X1 u_majority7_module_5_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_5_n1) );
  AND2_X1 u_majority7_module_5__and_module_1_U1 ( .A1(n_majority7_module_5_n5), 
        .A2(n_majority7_module_5_n4), .ZN(
        n_majority7_module_5__and_module_1_res) );
  OR2_X1 u_majority7_module_5__or_module_1_U1 ( .A1(n_majority7_module_5_n4), 
        .A2(n_majority7_module_5_n5), .ZN(
        n_majority7_module_5__or_module_1_res) );
  AND2_X1 u_majority7_module_5__and_module_2_U1 ( .A1(n_majority7_module_5_n7), 
        .A2(n_majority7_module_5_n2), .ZN(
        n_majority7_module_5__and_module_2_res) );
  OR2_X1 u_majority7_module_5__or_module_2_U1 ( .A1(n_majority7_module_5_n2), 
        .A2(n_majority7_module_5_n7), .ZN(
        n_majority7_module_5__or_module_2_res) );
  AND2_X1 u_majority7_module_5__and_module_3_U1 ( .A1(n_majority7_module_5_n6), 
        .A2(n_majority7_module_5_n1), .ZN(
        n_majority7_module_5__and_module_3_res) );
  OR2_X1 u_majority7_module_5__or_module_3_U1 ( .A1(n_majority7_module_5_n1), 
        .A2(n_majority7_module_5_n6), .ZN(
        n_majority7_module_5__or_module_3_res) );
  AND2_X1 u_majority7_module_5__and_module_4_U1 ( .A1(
        n_majority7_module_5__and_module_2_res), .A2(
        n_majority7_module_5__and_module_1_res), .ZN(
        n_majority7_module_5__and_module_4_res) );
  OR2_X1 u_majority7_module_5__or_module_4_U1 ( .A1(
        n_majority7_module_5__and_module_1_res), .A2(
        n_majority7_module_5__and_module_2_res), .ZN(
        n_majority7_module_5__or_module_4_res) );
  AND2_X1 u_majority7_module_5__and_module_5_U1 ( .A1(
        n_majority7_module_5__and_module_3_res), .A2(n_majority7_module_5_n3), 
        .ZN(n_majority7_module_5__and_module_5_res) );
  OR2_X1 u_majority7_module_5__or_module_5_U1 ( .A1(n_majority7_module_5_n3), 
        .A2(n_majority7_module_5__and_module_3_res), .ZN(
        n_majority7_module_5__or_module_5_res) );
  AND2_X1 u_majority7_module_5__and_module_6_U1 ( .A1(
        n_majority7_module_5__or_module_1_res), .A2(
        n_majority7_module_5__or_module_2_res), .ZN(
        n_majority7_module_5__and_module_6_res) );
  OR2_X1 u_majority7_module_5__or_module_6_U1 ( .A1(
        n_majority7_module_5__or_module_2_res), .A2(
        n_majority7_module_5__or_module_1_res), .ZN(
        n_majority7_module_5__or_module_6_res) );
  OR2_X1 u_majority7_module_5__or_module_7_U1 ( .A1(
        n_majority7_module_5__and_module_4_res), .A2(
        n_majority7_module_5__and_module_5_res), .ZN(
        n_majority7_module_5__or_module_7_res) );
  AND2_X1 u_majority7_module_5__and_module_7_U1 ( .A1(
        n_majority7_module_5__or_module_3_res), .A2(
        n_majority7_module_5__or_module_4_res), .ZN(
        n_majority7_module_5__and_module_7_res) );
  OR2_X1 u_majority7_module_5__or_module_8_U1 ( .A1(
        n_majority7_module_5__or_module_4_res), .A2(
        n_majority7_module_5__or_module_3_res), .ZN(
        n_majority7_module_5__or_module_8_res) );
  AND2_X1 u_majority7_module_5__and_module_8_U1 ( .A1(
        n_majority7_module_5__or_module_5_res), .A2(
        n_majority7_module_5__and_module_6_res), .ZN(
        n_majority7_module_5__and_module_8_res) );
  OR2_X1 u_majority7_module_5__or_module_9_U1 ( .A1(
        n_majority7_module_5__and_module_6_res), .A2(
        n_majority7_module_5__or_module_5_res), .ZN(
        n_majority7_module_5__or_module_9_res) );
  OR2_X1 u_majority7_module_5__or_module_10_U1 ( .A1(
        n_majority7_module_5__or_module_7_res), .A2(
        n_majority7_module_5__and_module_7_res), .ZN(
        n_majority7_module_5__or_module_10_res) );
  AND2_X1 u_majority7_module_5__and_module_9_U1 ( .A1(
        n_majority7_module_5__or_module_6_res), .A2(
        n_majority7_module_5__or_module_9_res), .ZN(
        n_majority7_module_5__and_module_9_res) );
  OR2_X1 u_majority7_module_5__or_module_11_U1 ( .A1(
        n_majority7_module_5__or_module_10_res), .A2(
        n_majority7_module_5__and_module_8_res), .ZN(
        n_majority7_module_5__or_module_11_res) );
  AND2_X1 u_majority7_module_5__and_module_10_U1 ( .A1(
        n_majority7_module_5__or_module_8_res), .A2(
        n_majority7_module_5__and_module_9_res), .ZN(
        n_majority7_module_5__and_module_10_res) );
  AND2_X1 u_majority7_module_5__and_module_11_U1 ( .A1(
        n_majority7_module_5__and_module_10_res), .A2(
        n_majority7_module_5__or_module_11_res), .ZN(n_majority7_module_5_res)
         );
  DFF_X1 u_reg_module_6__cini_mul_v000_reg ( .D(n_majority7_module_5_res), 
        .CK(clock_0), .Q(n_reg_module_6_res), .QN() );
  BUF_X1 u_majority7_module_6_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_6_n7) );
  BUF_X1 u_majority7_module_6_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_6_n6) );
  BUF_X1 u_majority7_module_6_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_6_n5) );
  BUF_X1 u_majority7_module_6_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_6_n4) );
  BUF_X1 u_majority7_module_6_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_6_n3) );
  BUF_X1 u_majority7_module_6_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_6_n2) );
  BUF_X1 u_majority7_module_6_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_6_n1) );
  AND2_X1 u_majority7_module_6__and_module_1_U1 ( .A1(n_majority7_module_6_n5), 
        .A2(n_majority7_module_6_n4), .ZN(
        n_majority7_module_6__and_module_1_res) );
  OR2_X1 u_majority7_module_6__or_module_1_U1 ( .A1(n_majority7_module_6_n4), 
        .A2(n_majority7_module_6_n5), .ZN(
        n_majority7_module_6__or_module_1_res) );
  AND2_X1 u_majority7_module_6__and_module_2_U1 ( .A1(n_majority7_module_6_n7), 
        .A2(n_majority7_module_6_n2), .ZN(
        n_majority7_module_6__and_module_2_res) );
  OR2_X1 u_majority7_module_6__or_module_2_U1 ( .A1(n_majority7_module_6_n2), 
        .A2(n_majority7_module_6_n7), .ZN(
        n_majority7_module_6__or_module_2_res) );
  AND2_X1 u_majority7_module_6__and_module_3_U1 ( .A1(n_majority7_module_6_n6), 
        .A2(n_majority7_module_6_n1), .ZN(
        n_majority7_module_6__and_module_3_res) );
  OR2_X1 u_majority7_module_6__or_module_3_U1 ( .A1(n_majority7_module_6_n1), 
        .A2(n_majority7_module_6_n6), .ZN(
        n_majority7_module_6__or_module_3_res) );
  AND2_X1 u_majority7_module_6__and_module_4_U1 ( .A1(
        n_majority7_module_6__and_module_2_res), .A2(
        n_majority7_module_6__and_module_1_res), .ZN(
        n_majority7_module_6__and_module_4_res) );
  OR2_X1 u_majority7_module_6__or_module_4_U1 ( .A1(
        n_majority7_module_6__and_module_1_res), .A2(
        n_majority7_module_6__and_module_2_res), .ZN(
        n_majority7_module_6__or_module_4_res) );
  AND2_X1 u_majority7_module_6__and_module_5_U1 ( .A1(
        n_majority7_module_6__and_module_3_res), .A2(n_majority7_module_6_n3), 
        .ZN(n_majority7_module_6__and_module_5_res) );
  OR2_X1 u_majority7_module_6__or_module_5_U1 ( .A1(n_majority7_module_6_n3), 
        .A2(n_majority7_module_6__and_module_3_res), .ZN(
        n_majority7_module_6__or_module_5_res) );
  AND2_X1 u_majority7_module_6__and_module_6_U1 ( .A1(
        n_majority7_module_6__or_module_1_res), .A2(
        n_majority7_module_6__or_module_2_res), .ZN(
        n_majority7_module_6__and_module_6_res) );
  OR2_X1 u_majority7_module_6__or_module_6_U1 ( .A1(
        n_majority7_module_6__or_module_2_res), .A2(
        n_majority7_module_6__or_module_1_res), .ZN(
        n_majority7_module_6__or_module_6_res) );
  OR2_X1 u_majority7_module_6__or_module_7_U1 ( .A1(
        n_majority7_module_6__and_module_4_res), .A2(
        n_majority7_module_6__and_module_5_res), .ZN(
        n_majority7_module_6__or_module_7_res) );
  AND2_X1 u_majority7_module_6__and_module_7_U1 ( .A1(
        n_majority7_module_6__or_module_3_res), .A2(
        n_majority7_module_6__or_module_4_res), .ZN(
        n_majority7_module_6__and_module_7_res) );
  OR2_X1 u_majority7_module_6__or_module_8_U1 ( .A1(
        n_majority7_module_6__or_module_4_res), .A2(
        n_majority7_module_6__or_module_3_res), .ZN(
        n_majority7_module_6__or_module_8_res) );
  AND2_X1 u_majority7_module_6__and_module_8_U1 ( .A1(
        n_majority7_module_6__or_module_5_res), .A2(
        n_majority7_module_6__and_module_6_res), .ZN(
        n_majority7_module_6__and_module_8_res) );
  OR2_X1 u_majority7_module_6__or_module_9_U1 ( .A1(
        n_majority7_module_6__and_module_6_res), .A2(
        n_majority7_module_6__or_module_5_res), .ZN(
        n_majority7_module_6__or_module_9_res) );
  OR2_X1 u_majority7_module_6__or_module_10_U1 ( .A1(
        n_majority7_module_6__or_module_7_res), .A2(
        n_majority7_module_6__and_module_7_res), .ZN(
        n_majority7_module_6__or_module_10_res) );
  AND2_X1 u_majority7_module_6__and_module_9_U1 ( .A1(
        n_majority7_module_6__or_module_6_res), .A2(
        n_majority7_module_6__or_module_9_res), .ZN(
        n_majority7_module_6__and_module_9_res) );
  OR2_X1 u_majority7_module_6__or_module_11_U1 ( .A1(
        n_majority7_module_6__or_module_10_res), .A2(
        n_majority7_module_6__and_module_8_res), .ZN(
        n_majority7_module_6__or_module_11_res) );
  AND2_X1 u_majority7_module_6__and_module_10_U1 ( .A1(
        n_majority7_module_6__or_module_8_res), .A2(
        n_majority7_module_6__and_module_9_res), .ZN(
        n_majority7_module_6__and_module_10_res) );
  AND2_X1 u_majority7_module_6__and_module_11_U1 ( .A1(
        n_majority7_module_6__and_module_10_res), .A2(
        n_majority7_module_6__or_module_11_res), .ZN(n_majority7_module_6_res)
         );
  DFF_X1 u_reg_module_7__cini_mul_v000_reg ( .D(n_majority7_module_6_res), 
        .CK(clock_0), .Q(n_reg_module_7_res), .QN() );
  BUF_X1 u_majority7_module_7_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_7_n7) );
  BUF_X1 u_majority7_module_7_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_7_n6) );
  BUF_X1 u_majority7_module_7_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_7_n5) );
  BUF_X1 u_majority7_module_7_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_7_n4) );
  BUF_X1 u_majority7_module_7_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_7_n3) );
  BUF_X1 u_majority7_module_7_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_7_n2) );
  BUF_X1 u_majority7_module_7_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_7_n1) );
  AND2_X1 u_majority7_module_7__and_module_1_U1 ( .A1(n_majority7_module_7_n5), 
        .A2(n_majority7_module_7_n4), .ZN(
        n_majority7_module_7__and_module_1_res) );
  OR2_X1 u_majority7_module_7__or_module_1_U1 ( .A1(n_majority7_module_7_n4), 
        .A2(n_majority7_module_7_n5), .ZN(
        n_majority7_module_7__or_module_1_res) );
  AND2_X1 u_majority7_module_7__and_module_2_U1 ( .A1(n_majority7_module_7_n7), 
        .A2(n_majority7_module_7_n2), .ZN(
        n_majority7_module_7__and_module_2_res) );
  OR2_X1 u_majority7_module_7__or_module_2_U1 ( .A1(n_majority7_module_7_n2), 
        .A2(n_majority7_module_7_n7), .ZN(
        n_majority7_module_7__or_module_2_res) );
  AND2_X1 u_majority7_module_7__and_module_3_U1 ( .A1(n_majority7_module_7_n6), 
        .A2(n_majority7_module_7_n1), .ZN(
        n_majority7_module_7__and_module_3_res) );
  OR2_X1 u_majority7_module_7__or_module_3_U1 ( .A1(n_majority7_module_7_n1), 
        .A2(n_majority7_module_7_n6), .ZN(
        n_majority7_module_7__or_module_3_res) );
  AND2_X1 u_majority7_module_7__and_module_4_U1 ( .A1(
        n_majority7_module_7__and_module_2_res), .A2(
        n_majority7_module_7__and_module_1_res), .ZN(
        n_majority7_module_7__and_module_4_res) );
  OR2_X1 u_majority7_module_7__or_module_4_U1 ( .A1(
        n_majority7_module_7__and_module_1_res), .A2(
        n_majority7_module_7__and_module_2_res), .ZN(
        n_majority7_module_7__or_module_4_res) );
  AND2_X1 u_majority7_module_7__and_module_5_U1 ( .A1(
        n_majority7_module_7__and_module_3_res), .A2(n_majority7_module_7_n3), 
        .ZN(n_majority7_module_7__and_module_5_res) );
  OR2_X1 u_majority7_module_7__or_module_5_U1 ( .A1(n_majority7_module_7_n3), 
        .A2(n_majority7_module_7__and_module_3_res), .ZN(
        n_majority7_module_7__or_module_5_res) );
  AND2_X1 u_majority7_module_7__and_module_6_U1 ( .A1(
        n_majority7_module_7__or_module_1_res), .A2(
        n_majority7_module_7__or_module_2_res), .ZN(
        n_majority7_module_7__and_module_6_res) );
  OR2_X1 u_majority7_module_7__or_module_6_U1 ( .A1(
        n_majority7_module_7__or_module_2_res), .A2(
        n_majority7_module_7__or_module_1_res), .ZN(
        n_majority7_module_7__or_module_6_res) );
  OR2_X1 u_majority7_module_7__or_module_7_U1 ( .A1(
        n_majority7_module_7__and_module_4_res), .A2(
        n_majority7_module_7__and_module_5_res), .ZN(
        n_majority7_module_7__or_module_7_res) );
  AND2_X1 u_majority7_module_7__and_module_7_U1 ( .A1(
        n_majority7_module_7__or_module_3_res), .A2(
        n_majority7_module_7__or_module_4_res), .ZN(
        n_majority7_module_7__and_module_7_res) );
  OR2_X1 u_majority7_module_7__or_module_8_U1 ( .A1(
        n_majority7_module_7__or_module_4_res), .A2(
        n_majority7_module_7__or_module_3_res), .ZN(
        n_majority7_module_7__or_module_8_res) );
  AND2_X1 u_majority7_module_7__and_module_8_U1 ( .A1(
        n_majority7_module_7__or_module_5_res), .A2(
        n_majority7_module_7__and_module_6_res), .ZN(
        n_majority7_module_7__and_module_8_res) );
  OR2_X1 u_majority7_module_7__or_module_9_U1 ( .A1(
        n_majority7_module_7__and_module_6_res), .A2(
        n_majority7_module_7__or_module_5_res), .ZN(
        n_majority7_module_7__or_module_9_res) );
  OR2_X1 u_majority7_module_7__or_module_10_U1 ( .A1(
        n_majority7_module_7__or_module_7_res), .A2(
        n_majority7_module_7__and_module_7_res), .ZN(
        n_majority7_module_7__or_module_10_res) );
  AND2_X1 u_majority7_module_7__and_module_9_U1 ( .A1(
        n_majority7_module_7__or_module_6_res), .A2(
        n_majority7_module_7__or_module_9_res), .ZN(
        n_majority7_module_7__and_module_9_res) );
  OR2_X1 u_majority7_module_7__or_module_11_U1 ( .A1(
        n_majority7_module_7__or_module_10_res), .A2(
        n_majority7_module_7__and_module_8_res), .ZN(
        n_majority7_module_7__or_module_11_res) );
  AND2_X1 u_majority7_module_7__and_module_10_U1 ( .A1(
        n_majority7_module_7__or_module_8_res), .A2(
        n_majority7_module_7__and_module_9_res), .ZN(
        n_majority7_module_7__and_module_10_res) );
  AND2_X1 u_majority7_module_7__and_module_11_U1 ( .A1(
        n_majority7_module_7__and_module_10_res), .A2(
        n_majority7_module_7__or_module_11_res), .ZN(n_majority7_module_7_res)
         );
  DFF_X1 u_reg_module_8__cini_mul_v000_reg ( .D(n_majority7_module_7_res), 
        .CK(clock_0), .Q(n_reg_module_8_res), .QN() );
  BUF_X1 u_majority7_module_8_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_8_n7) );
  BUF_X1 u_majority7_module_8_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_8_n6) );
  BUF_X1 u_majority7_module_8_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_8_n5) );
  BUF_X1 u_majority7_module_8_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_8_n4) );
  BUF_X1 u_majority7_module_8_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_8_n3) );
  BUF_X1 u_majority7_module_8_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_8_n2) );
  BUF_X1 u_majority7_module_8_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_8_n1) );
  AND2_X1 u_majority7_module_8__and_module_1_U1 ( .A1(n_majority7_module_8_n5), 
        .A2(n_majority7_module_8_n4), .ZN(
        n_majority7_module_8__and_module_1_res) );
  OR2_X1 u_majority7_module_8__or_module_1_U1 ( .A1(n_majority7_module_8_n4), 
        .A2(n_majority7_module_8_n5), .ZN(
        n_majority7_module_8__or_module_1_res) );
  AND2_X1 u_majority7_module_8__and_module_2_U1 ( .A1(n_majority7_module_8_n7), 
        .A2(n_majority7_module_8_n2), .ZN(
        n_majority7_module_8__and_module_2_res) );
  OR2_X1 u_majority7_module_8__or_module_2_U1 ( .A1(n_majority7_module_8_n2), 
        .A2(n_majority7_module_8_n7), .ZN(
        n_majority7_module_8__or_module_2_res) );
  AND2_X1 u_majority7_module_8__and_module_3_U1 ( .A1(n_majority7_module_8_n6), 
        .A2(n_majority7_module_8_n1), .ZN(
        n_majority7_module_8__and_module_3_res) );
  OR2_X1 u_majority7_module_8__or_module_3_U1 ( .A1(n_majority7_module_8_n1), 
        .A2(n_majority7_module_8_n6), .ZN(
        n_majority7_module_8__or_module_3_res) );
  AND2_X1 u_majority7_module_8__and_module_4_U1 ( .A1(
        n_majority7_module_8__and_module_2_res), .A2(
        n_majority7_module_8__and_module_1_res), .ZN(
        n_majority7_module_8__and_module_4_res) );
  OR2_X1 u_majority7_module_8__or_module_4_U1 ( .A1(
        n_majority7_module_8__and_module_1_res), .A2(
        n_majority7_module_8__and_module_2_res), .ZN(
        n_majority7_module_8__or_module_4_res) );
  AND2_X1 u_majority7_module_8__and_module_5_U1 ( .A1(
        n_majority7_module_8__and_module_3_res), .A2(n_majority7_module_8_n3), 
        .ZN(n_majority7_module_8__and_module_5_res) );
  OR2_X1 u_majority7_module_8__or_module_5_U1 ( .A1(n_majority7_module_8_n3), 
        .A2(n_majority7_module_8__and_module_3_res), .ZN(
        n_majority7_module_8__or_module_5_res) );
  AND2_X1 u_majority7_module_8__and_module_6_U1 ( .A1(
        n_majority7_module_8__or_module_1_res), .A2(
        n_majority7_module_8__or_module_2_res), .ZN(
        n_majority7_module_8__and_module_6_res) );
  OR2_X1 u_majority7_module_8__or_module_6_U1 ( .A1(
        n_majority7_module_8__or_module_2_res), .A2(
        n_majority7_module_8__or_module_1_res), .ZN(
        n_majority7_module_8__or_module_6_res) );
  OR2_X1 u_majority7_module_8__or_module_7_U1 ( .A1(
        n_majority7_module_8__and_module_4_res), .A2(
        n_majority7_module_8__and_module_5_res), .ZN(
        n_majority7_module_8__or_module_7_res) );
  AND2_X1 u_majority7_module_8__and_module_7_U1 ( .A1(
        n_majority7_module_8__or_module_3_res), .A2(
        n_majority7_module_8__or_module_4_res), .ZN(
        n_majority7_module_8__and_module_7_res) );
  OR2_X1 u_majority7_module_8__or_module_8_U1 ( .A1(
        n_majority7_module_8__or_module_4_res), .A2(
        n_majority7_module_8__or_module_3_res), .ZN(
        n_majority7_module_8__or_module_8_res) );
  AND2_X1 u_majority7_module_8__and_module_8_U1 ( .A1(
        n_majority7_module_8__or_module_5_res), .A2(
        n_majority7_module_8__and_module_6_res), .ZN(
        n_majority7_module_8__and_module_8_res) );
  OR2_X1 u_majority7_module_8__or_module_9_U1 ( .A1(
        n_majority7_module_8__and_module_6_res), .A2(
        n_majority7_module_8__or_module_5_res), .ZN(
        n_majority7_module_8__or_module_9_res) );
  OR2_X1 u_majority7_module_8__or_module_10_U1 ( .A1(
        n_majority7_module_8__or_module_7_res), .A2(
        n_majority7_module_8__and_module_7_res), .ZN(
        n_majority7_module_8__or_module_10_res) );
  AND2_X1 u_majority7_module_8__and_module_9_U1 ( .A1(
        n_majority7_module_8__or_module_6_res), .A2(
        n_majority7_module_8__or_module_9_res), .ZN(
        n_majority7_module_8__and_module_9_res) );
  OR2_X1 u_majority7_module_8__or_module_11_U1 ( .A1(
        n_majority7_module_8__or_module_10_res), .A2(
        n_majority7_module_8__and_module_8_res), .ZN(
        n_majority7_module_8__or_module_11_res) );
  AND2_X1 u_majority7_module_8__and_module_10_U1 ( .A1(
        n_majority7_module_8__or_module_8_res), .A2(
        n_majority7_module_8__and_module_9_res), .ZN(
        n_majority7_module_8__and_module_10_res) );
  AND2_X1 u_majority7_module_8__and_module_11_U1 ( .A1(
        n_majority7_module_8__and_module_10_res), .A2(
        n_majority7_module_8__or_module_11_res), .ZN(n_majority7_module_8_res)
         );
  DFF_X1 u_reg_module_9__cini_mul_v000_reg ( .D(n_majority7_module_8_res), 
        .CK(clock_0), .Q(n_reg_module_9_res), .QN() );
  BUF_X1 u_majority7_module_9_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_9_n7) );
  BUF_X1 u_majority7_module_9_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_9_n6) );
  BUF_X1 u_majority7_module_9_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_9_n5) );
  BUF_X1 u_majority7_module_9_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_9_n4) );
  BUF_X1 u_majority7_module_9_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_9_n3) );
  BUF_X1 u_majority7_module_9_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_9_n2) );
  BUF_X1 u_majority7_module_9_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_9_n1) );
  AND2_X1 u_majority7_module_9__and_module_1_U1 ( .A1(n_majority7_module_9_n5), 
        .A2(n_majority7_module_9_n4), .ZN(
        n_majority7_module_9__and_module_1_res) );
  OR2_X1 u_majority7_module_9__or_module_1_U1 ( .A1(n_majority7_module_9_n4), 
        .A2(n_majority7_module_9_n5), .ZN(
        n_majority7_module_9__or_module_1_res) );
  AND2_X1 u_majority7_module_9__and_module_2_U1 ( .A1(n_majority7_module_9_n7), 
        .A2(n_majority7_module_9_n2), .ZN(
        n_majority7_module_9__and_module_2_res) );
  OR2_X1 u_majority7_module_9__or_module_2_U1 ( .A1(n_majority7_module_9_n2), 
        .A2(n_majority7_module_9_n7), .ZN(
        n_majority7_module_9__or_module_2_res) );
  AND2_X1 u_majority7_module_9__and_module_3_U1 ( .A1(n_majority7_module_9_n6), 
        .A2(n_majority7_module_9_n1), .ZN(
        n_majority7_module_9__and_module_3_res) );
  OR2_X1 u_majority7_module_9__or_module_3_U1 ( .A1(n_majority7_module_9_n1), 
        .A2(n_majority7_module_9_n6), .ZN(
        n_majority7_module_9__or_module_3_res) );
  AND2_X1 u_majority7_module_9__and_module_4_U1 ( .A1(
        n_majority7_module_9__and_module_2_res), .A2(
        n_majority7_module_9__and_module_1_res), .ZN(
        n_majority7_module_9__and_module_4_res) );
  OR2_X1 u_majority7_module_9__or_module_4_U1 ( .A1(
        n_majority7_module_9__and_module_1_res), .A2(
        n_majority7_module_9__and_module_2_res), .ZN(
        n_majority7_module_9__or_module_4_res) );
  AND2_X1 u_majority7_module_9__and_module_5_U1 ( .A1(
        n_majority7_module_9__and_module_3_res), .A2(n_majority7_module_9_n3), 
        .ZN(n_majority7_module_9__and_module_5_res) );
  OR2_X1 u_majority7_module_9__or_module_5_U1 ( .A1(n_majority7_module_9_n3), 
        .A2(n_majority7_module_9__and_module_3_res), .ZN(
        n_majority7_module_9__or_module_5_res) );
  AND2_X1 u_majority7_module_9__and_module_6_U1 ( .A1(
        n_majority7_module_9__or_module_1_res), .A2(
        n_majority7_module_9__or_module_2_res), .ZN(
        n_majority7_module_9__and_module_6_res) );
  OR2_X1 u_majority7_module_9__or_module_6_U1 ( .A1(
        n_majority7_module_9__or_module_2_res), .A2(
        n_majority7_module_9__or_module_1_res), .ZN(
        n_majority7_module_9__or_module_6_res) );
  OR2_X1 u_majority7_module_9__or_module_7_U1 ( .A1(
        n_majority7_module_9__and_module_4_res), .A2(
        n_majority7_module_9__and_module_5_res), .ZN(
        n_majority7_module_9__or_module_7_res) );
  AND2_X1 u_majority7_module_9__and_module_7_U1 ( .A1(
        n_majority7_module_9__or_module_3_res), .A2(
        n_majority7_module_9__or_module_4_res), .ZN(
        n_majority7_module_9__and_module_7_res) );
  OR2_X1 u_majority7_module_9__or_module_8_U1 ( .A1(
        n_majority7_module_9__or_module_4_res), .A2(
        n_majority7_module_9__or_module_3_res), .ZN(
        n_majority7_module_9__or_module_8_res) );
  AND2_X1 u_majority7_module_9__and_module_8_U1 ( .A1(
        n_majority7_module_9__or_module_5_res), .A2(
        n_majority7_module_9__and_module_6_res), .ZN(
        n_majority7_module_9__and_module_8_res) );
  OR2_X1 u_majority7_module_9__or_module_9_U1 ( .A1(
        n_majority7_module_9__and_module_6_res), .A2(
        n_majority7_module_9__or_module_5_res), .ZN(
        n_majority7_module_9__or_module_9_res) );
  OR2_X1 u_majority7_module_9__or_module_10_U1 ( .A1(
        n_majority7_module_9__or_module_7_res), .A2(
        n_majority7_module_9__and_module_7_res), .ZN(
        n_majority7_module_9__or_module_10_res) );
  AND2_X1 u_majority7_module_9__and_module_9_U1 ( .A1(
        n_majority7_module_9__or_module_6_res), .A2(
        n_majority7_module_9__or_module_9_res), .ZN(
        n_majority7_module_9__and_module_9_res) );
  OR2_X1 u_majority7_module_9__or_module_11_U1 ( .A1(
        n_majority7_module_9__or_module_10_res), .A2(
        n_majority7_module_9__and_module_8_res), .ZN(
        n_majority7_module_9__or_module_11_res) );
  AND2_X1 u_majority7_module_9__and_module_10_U1 ( .A1(
        n_majority7_module_9__or_module_8_res), .A2(
        n_majority7_module_9__and_module_9_res), .ZN(
        n_majority7_module_9__and_module_10_res) );
  AND2_X1 u_majority7_module_9__and_module_11_U1 ( .A1(
        n_majority7_module_9__and_module_10_res), .A2(
        n_majority7_module_9__or_module_11_res), .ZN(n_majority7_module_9_res)
         );
  DFF_X1 u_reg_module_10__cini_mul_v000_reg ( .D(n_majority7_module_9_res), 
        .CK(clock_0), .Q(n_reg_module_10_res), .QN() );
  BUF_X1 u_majority7_module_10_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_10_n7) );
  BUF_X1 u_majority7_module_10_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_10_n6) );
  BUF_X1 u_majority7_module_10_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_10_n5) );
  BUF_X1 u_majority7_module_10_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_10_n4) );
  BUF_X1 u_majority7_module_10_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_10_n3) );
  BUF_X1 u_majority7_module_10_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_10_n2) );
  BUF_X1 u_majority7_module_10_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_10_n1) );
  AND2_X1 u_majority7_module_10__and_module_1_U1 ( .A1(
        n_majority7_module_10_n5), .A2(n_majority7_module_10_n4), .ZN(
        n_majority7_module_10__and_module_1_res) );
  OR2_X1 u_majority7_module_10__or_module_1_U1 ( .A1(n_majority7_module_10_n4), 
        .A2(n_majority7_module_10_n5), .ZN(
        n_majority7_module_10__or_module_1_res) );
  AND2_X1 u_majority7_module_10__and_module_2_U1 ( .A1(
        n_majority7_module_10_n7), .A2(n_majority7_module_10_n2), .ZN(
        n_majority7_module_10__and_module_2_res) );
  OR2_X1 u_majority7_module_10__or_module_2_U1 ( .A1(n_majority7_module_10_n2), 
        .A2(n_majority7_module_10_n7), .ZN(
        n_majority7_module_10__or_module_2_res) );
  AND2_X1 u_majority7_module_10__and_module_3_U1 ( .A1(
        n_majority7_module_10_n6), .A2(n_majority7_module_10_n1), .ZN(
        n_majority7_module_10__and_module_3_res) );
  OR2_X1 u_majority7_module_10__or_module_3_U1 ( .A1(n_majority7_module_10_n1), 
        .A2(n_majority7_module_10_n6), .ZN(
        n_majority7_module_10__or_module_3_res) );
  AND2_X1 u_majority7_module_10__and_module_4_U1 ( .A1(
        n_majority7_module_10__and_module_2_res), .A2(
        n_majority7_module_10__and_module_1_res), .ZN(
        n_majority7_module_10__and_module_4_res) );
  OR2_X1 u_majority7_module_10__or_module_4_U1 ( .A1(
        n_majority7_module_10__and_module_1_res), .A2(
        n_majority7_module_10__and_module_2_res), .ZN(
        n_majority7_module_10__or_module_4_res) );
  AND2_X1 u_majority7_module_10__and_module_5_U1 ( .A1(
        n_majority7_module_10__and_module_3_res), .A2(n_majority7_module_10_n3), .ZN(n_majority7_module_10__and_module_5_res) );
  OR2_X1 u_majority7_module_10__or_module_5_U1 ( .A1(n_majority7_module_10_n3), 
        .A2(n_majority7_module_10__and_module_3_res), .ZN(
        n_majority7_module_10__or_module_5_res) );
  AND2_X1 u_majority7_module_10__and_module_6_U1 ( .A1(
        n_majority7_module_10__or_module_1_res), .A2(
        n_majority7_module_10__or_module_2_res), .ZN(
        n_majority7_module_10__and_module_6_res) );
  OR2_X1 u_majority7_module_10__or_module_6_U1 ( .A1(
        n_majority7_module_10__or_module_2_res), .A2(
        n_majority7_module_10__or_module_1_res), .ZN(
        n_majority7_module_10__or_module_6_res) );
  OR2_X1 u_majority7_module_10__or_module_7_U1 ( .A1(
        n_majority7_module_10__and_module_4_res), .A2(
        n_majority7_module_10__and_module_5_res), .ZN(
        n_majority7_module_10__or_module_7_res) );
  AND2_X1 u_majority7_module_10__and_module_7_U1 ( .A1(
        n_majority7_module_10__or_module_3_res), .A2(
        n_majority7_module_10__or_module_4_res), .ZN(
        n_majority7_module_10__and_module_7_res) );
  OR2_X1 u_majority7_module_10__or_module_8_U1 ( .A1(
        n_majority7_module_10__or_module_4_res), .A2(
        n_majority7_module_10__or_module_3_res), .ZN(
        n_majority7_module_10__or_module_8_res) );
  AND2_X1 u_majority7_module_10__and_module_8_U1 ( .A1(
        n_majority7_module_10__or_module_5_res), .A2(
        n_majority7_module_10__and_module_6_res), .ZN(
        n_majority7_module_10__and_module_8_res) );
  OR2_X1 u_majority7_module_10__or_module_9_U1 ( .A1(
        n_majority7_module_10__and_module_6_res), .A2(
        n_majority7_module_10__or_module_5_res), .ZN(
        n_majority7_module_10__or_module_9_res) );
  OR2_X1 u_majority7_module_10__or_module_10_U1 ( .A1(
        n_majority7_module_10__or_module_7_res), .A2(
        n_majority7_module_10__and_module_7_res), .ZN(
        n_majority7_module_10__or_module_10_res) );
  AND2_X1 u_majority7_module_10__and_module_9_U1 ( .A1(
        n_majority7_module_10__or_module_6_res), .A2(
        n_majority7_module_10__or_module_9_res), .ZN(
        n_majority7_module_10__and_module_9_res) );
  OR2_X1 u_majority7_module_10__or_module_11_U1 ( .A1(
        n_majority7_module_10__or_module_10_res), .A2(
        n_majority7_module_10__and_module_8_res), .ZN(
        n_majority7_module_10__or_module_11_res) );
  AND2_X1 u_majority7_module_10__and_module_10_U1 ( .A1(
        n_majority7_module_10__or_module_8_res), .A2(
        n_majority7_module_10__and_module_9_res), .ZN(
        n_majority7_module_10__and_module_10_res) );
  AND2_X1 u_majority7_module_10__and_module_11_U1 ( .A1(
        n_majority7_module_10__and_module_10_res), .A2(
        n_majority7_module_10__or_module_11_res), .ZN(
        n_majority7_module_10_res) );
  DFF_X1 u_reg_module_11__cini_mul_v000_reg ( .D(n_majority7_module_10_res), 
        .CK(clock_0), .Q(n_reg_module_11_res), .QN() );
  BUF_X1 u_majority7_module_11_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_11_n7) );
  BUF_X1 u_majority7_module_11_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_11_n6) );
  BUF_X1 u_majority7_module_11_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_11_n5) );
  BUF_X1 u_majority7_module_11_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_11_n4) );
  BUF_X1 u_majority7_module_11_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_11_n3) );
  BUF_X1 u_majority7_module_11_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_11_n2) );
  BUF_X1 u_majority7_module_11_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_11_n1) );
  AND2_X1 u_majority7_module_11__and_module_1_U1 ( .A1(
        n_majority7_module_11_n5), .A2(n_majority7_module_11_n4), .ZN(
        n_majority7_module_11__and_module_1_res) );
  OR2_X1 u_majority7_module_11__or_module_1_U1 ( .A1(n_majority7_module_11_n4), 
        .A2(n_majority7_module_11_n5), .ZN(
        n_majority7_module_11__or_module_1_res) );
  AND2_X1 u_majority7_module_11__and_module_2_U1 ( .A1(
        n_majority7_module_11_n7), .A2(n_majority7_module_11_n2), .ZN(
        n_majority7_module_11__and_module_2_res) );
  OR2_X1 u_majority7_module_11__or_module_2_U1 ( .A1(n_majority7_module_11_n2), 
        .A2(n_majority7_module_11_n7), .ZN(
        n_majority7_module_11__or_module_2_res) );
  AND2_X1 u_majority7_module_11__and_module_3_U1 ( .A1(
        n_majority7_module_11_n6), .A2(n_majority7_module_11_n1), .ZN(
        n_majority7_module_11__and_module_3_res) );
  OR2_X1 u_majority7_module_11__or_module_3_U1 ( .A1(n_majority7_module_11_n1), 
        .A2(n_majority7_module_11_n6), .ZN(
        n_majority7_module_11__or_module_3_res) );
  AND2_X1 u_majority7_module_11__and_module_4_U1 ( .A1(
        n_majority7_module_11__and_module_2_res), .A2(
        n_majority7_module_11__and_module_1_res), .ZN(
        n_majority7_module_11__and_module_4_res) );
  OR2_X1 u_majority7_module_11__or_module_4_U1 ( .A1(
        n_majority7_module_11__and_module_1_res), .A2(
        n_majority7_module_11__and_module_2_res), .ZN(
        n_majority7_module_11__or_module_4_res) );
  AND2_X1 u_majority7_module_11__and_module_5_U1 ( .A1(
        n_majority7_module_11__and_module_3_res), .A2(n_majority7_module_11_n3), .ZN(n_majority7_module_11__and_module_5_res) );
  OR2_X1 u_majority7_module_11__or_module_5_U1 ( .A1(n_majority7_module_11_n3), 
        .A2(n_majority7_module_11__and_module_3_res), .ZN(
        n_majority7_module_11__or_module_5_res) );
  AND2_X1 u_majority7_module_11__and_module_6_U1 ( .A1(
        n_majority7_module_11__or_module_1_res), .A2(
        n_majority7_module_11__or_module_2_res), .ZN(
        n_majority7_module_11__and_module_6_res) );
  OR2_X1 u_majority7_module_11__or_module_6_U1 ( .A1(
        n_majority7_module_11__or_module_2_res), .A2(
        n_majority7_module_11__or_module_1_res), .ZN(
        n_majority7_module_11__or_module_6_res) );
  OR2_X1 u_majority7_module_11__or_module_7_U1 ( .A1(
        n_majority7_module_11__and_module_4_res), .A2(
        n_majority7_module_11__and_module_5_res), .ZN(
        n_majority7_module_11__or_module_7_res) );
  AND2_X1 u_majority7_module_11__and_module_7_U1 ( .A1(
        n_majority7_module_11__or_module_3_res), .A2(
        n_majority7_module_11__or_module_4_res), .ZN(
        n_majority7_module_11__and_module_7_res) );
  OR2_X1 u_majority7_module_11__or_module_8_U1 ( .A1(
        n_majority7_module_11__or_module_4_res), .A2(
        n_majority7_module_11__or_module_3_res), .ZN(
        n_majority7_module_11__or_module_8_res) );
  AND2_X1 u_majority7_module_11__and_module_8_U1 ( .A1(
        n_majority7_module_11__or_module_5_res), .A2(
        n_majority7_module_11__and_module_6_res), .ZN(
        n_majority7_module_11__and_module_8_res) );
  OR2_X1 u_majority7_module_11__or_module_9_U1 ( .A1(
        n_majority7_module_11__and_module_6_res), .A2(
        n_majority7_module_11__or_module_5_res), .ZN(
        n_majority7_module_11__or_module_9_res) );
  OR2_X1 u_majority7_module_11__or_module_10_U1 ( .A1(
        n_majority7_module_11__or_module_7_res), .A2(
        n_majority7_module_11__and_module_7_res), .ZN(
        n_majority7_module_11__or_module_10_res) );
  AND2_X1 u_majority7_module_11__and_module_9_U1 ( .A1(
        n_majority7_module_11__or_module_6_res), .A2(
        n_majority7_module_11__or_module_9_res), .ZN(
        n_majority7_module_11__and_module_9_res) );
  OR2_X1 u_majority7_module_11__or_module_11_U1 ( .A1(
        n_majority7_module_11__or_module_10_res), .A2(
        n_majority7_module_11__and_module_8_res), .ZN(
        n_majority7_module_11__or_module_11_res) );
  AND2_X1 u_majority7_module_11__and_module_10_U1 ( .A1(
        n_majority7_module_11__or_module_8_res), .A2(
        n_majority7_module_11__and_module_9_res), .ZN(
        n_majority7_module_11__and_module_10_res) );
  AND2_X1 u_majority7_module_11__and_module_11_U1 ( .A1(
        n_majority7_module_11__and_module_10_res), .A2(
        n_majority7_module_11__or_module_11_res), .ZN(
        n_majority7_module_11_res) );
  DFF_X1 u_reg_module_12__cini_mul_v000_reg ( .D(n_majority7_module_11_res), 
        .CK(clock_0), .Q(n_reg_module_12_res), .QN() );
  BUF_X1 u_majority7_module_12_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_12_n7) );
  BUF_X1 u_majority7_module_12_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_12_n6) );
  BUF_X1 u_majority7_module_12_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_12_n5) );
  BUF_X1 u_majority7_module_12_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_12_n4) );
  BUF_X1 u_majority7_module_12_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_12_n3) );
  BUF_X1 u_majority7_module_12_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_12_n2) );
  BUF_X1 u_majority7_module_12_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_12_n1) );
  AND2_X1 u_majority7_module_12__and_module_1_U1 ( .A1(
        n_majority7_module_12_n1), .A2(n_majority7_module_12_n5), .ZN(
        n_majority7_module_12__and_module_1_res) );
  OR2_X1 u_majority7_module_12__or_module_1_U1 ( .A1(n_majority7_module_12_n5), 
        .A2(n_majority7_module_12_n1), .ZN(
        n_majority7_module_12__or_module_1_res) );
  AND2_X1 u_majority7_module_12__and_module_2_U1 ( .A1(
        n_majority7_module_12_n7), .A2(n_majority7_module_12_n3), .ZN(
        n_majority7_module_12__and_module_2_res) );
  OR2_X1 u_majority7_module_12__or_module_2_U1 ( .A1(n_majority7_module_12_n3), 
        .A2(n_majority7_module_12_n7), .ZN(
        n_majority7_module_12__or_module_2_res) );
  AND2_X1 u_majority7_module_12__and_module_3_U1 ( .A1(
        n_majority7_module_12_n6), .A2(n_majority7_module_12_n2), .ZN(
        n_majority7_module_12__and_module_3_res) );
  OR2_X1 u_majority7_module_12__or_module_3_U1 ( .A1(n_majority7_module_12_n2), 
        .A2(n_majority7_module_12_n6), .ZN(
        n_majority7_module_12__or_module_3_res) );
  AND2_X1 u_majority7_module_12__and_module_4_U1 ( .A1(
        n_majority7_module_12__and_module_2_res), .A2(
        n_majority7_module_12__and_module_1_res), .ZN(
        n_majority7_module_12__and_module_4_res) );
  OR2_X1 u_majority7_module_12__or_module_4_U1 ( .A1(
        n_majority7_module_12__and_module_1_res), .A2(
        n_majority7_module_12__and_module_2_res), .ZN(
        n_majority7_module_12__or_module_4_res) );
  AND2_X1 u_majority7_module_12__and_module_5_U1 ( .A1(
        n_majority7_module_12__and_module_3_res), .A2(n_majority7_module_12_n4), .ZN(n_majority7_module_12__and_module_5_res) );
  OR2_X1 u_majority7_module_12__or_module_5_U1 ( .A1(n_majority7_module_12_n4), 
        .A2(n_majority7_module_12__and_module_3_res), .ZN(
        n_majority7_module_12__or_module_5_res) );
  AND2_X1 u_majority7_module_12__and_module_6_U1 ( .A1(
        n_majority7_module_12__or_module_1_res), .A2(
        n_majority7_module_12__or_module_2_res), .ZN(
        n_majority7_module_12__and_module_6_res) );
  OR2_X1 u_majority7_module_12__or_module_6_U1 ( .A1(
        n_majority7_module_12__or_module_2_res), .A2(
        n_majority7_module_12__or_module_1_res), .ZN(
        n_majority7_module_12__or_module_6_res) );
  OR2_X1 u_majority7_module_12__or_module_7_U1 ( .A1(
        n_majority7_module_12__and_module_4_res), .A2(
        n_majority7_module_12__and_module_5_res), .ZN(
        n_majority7_module_12__or_module_7_res) );
  AND2_X1 u_majority7_module_12__and_module_7_U1 ( .A1(
        n_majority7_module_12__or_module_3_res), .A2(
        n_majority7_module_12__or_module_4_res), .ZN(
        n_majority7_module_12__and_module_7_res) );
  OR2_X1 u_majority7_module_12__or_module_8_U1 ( .A1(
        n_majority7_module_12__or_module_4_res), .A2(
        n_majority7_module_12__or_module_3_res), .ZN(
        n_majority7_module_12__or_module_8_res) );
  AND2_X1 u_majority7_module_12__and_module_8_U1 ( .A1(
        n_majority7_module_12__or_module_5_res), .A2(
        n_majority7_module_12__and_module_6_res), .ZN(
        n_majority7_module_12__and_module_8_res) );
  OR2_X1 u_majority7_module_12__or_module_9_U1 ( .A1(
        n_majority7_module_12__and_module_6_res), .A2(
        n_majority7_module_12__or_module_5_res), .ZN(
        n_majority7_module_12__or_module_9_res) );
  OR2_X1 u_majority7_module_12__or_module_10_U1 ( .A1(
        n_majority7_module_12__or_module_7_res), .A2(
        n_majority7_module_12__and_module_7_res), .ZN(
        n_majority7_module_12__or_module_10_res) );
  AND2_X1 u_majority7_module_12__and_module_9_U1 ( .A1(
        n_majority7_module_12__or_module_6_res), .A2(
        n_majority7_module_12__or_module_9_res), .ZN(
        n_majority7_module_12__and_module_9_res) );
  OR2_X1 u_majority7_module_12__or_module_11_U1 ( .A1(
        n_majority7_module_12__or_module_10_res), .A2(
        n_majority7_module_12__and_module_8_res), .ZN(
        n_majority7_module_12__or_module_11_res) );
  AND2_X1 u_majority7_module_12__and_module_10_U1 ( .A1(
        n_majority7_module_12__or_module_8_res), .A2(
        n_majority7_module_12__and_module_9_res), .ZN(
        n_majority7_module_12__and_module_10_res) );
  AND2_X1 u_majority7_module_12__and_module_11_U1 ( .A1(
        n_majority7_module_12__and_module_10_res), .A2(
        n_majority7_module_12__or_module_11_res), .ZN(
        n_majority7_module_12_res) );
  DFF_X1 u_reg_module_13__cini_mul_v000_reg ( .D(n_majority7_module_12_res), 
        .CK(clock_0), .Q(n_reg_module_13_res), .QN() );
  BUF_X1 u_majority7_module_13_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_13_n7) );
  BUF_X1 u_majority7_module_13_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_13_n6) );
  BUF_X1 u_majority7_module_13_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_13_n5) );
  BUF_X1 u_majority7_module_13_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_13_n4) );
  BUF_X1 u_majority7_module_13_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_13_n3) );
  BUF_X1 u_majority7_module_13_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_13_n2) );
  BUF_X1 u_majority7_module_13_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_13_n1) );
  AND2_X1 u_majority7_module_13__and_module_1_U1 ( .A1(
        n_majority7_module_13_n1), .A2(n_majority7_module_13_n5), .ZN(
        n_majority7_module_13__and_module_1_res) );
  OR2_X1 u_majority7_module_13__or_module_1_U1 ( .A1(n_majority7_module_13_n5), 
        .A2(n_majority7_module_13_n1), .ZN(
        n_majority7_module_13__or_module_1_res) );
  AND2_X1 u_majority7_module_13__and_module_2_U1 ( .A1(
        n_majority7_module_13_n7), .A2(n_majority7_module_13_n3), .ZN(
        n_majority7_module_13__and_module_2_res) );
  OR2_X1 u_majority7_module_13__or_module_2_U1 ( .A1(n_majority7_module_13_n3), 
        .A2(n_majority7_module_13_n7), .ZN(
        n_majority7_module_13__or_module_2_res) );
  AND2_X1 u_majority7_module_13__and_module_3_U1 ( .A1(
        n_majority7_module_13_n6), .A2(n_majority7_module_13_n2), .ZN(
        n_majority7_module_13__and_module_3_res) );
  OR2_X1 u_majority7_module_13__or_module_3_U1 ( .A1(n_majority7_module_13_n2), 
        .A2(n_majority7_module_13_n6), .ZN(
        n_majority7_module_13__or_module_3_res) );
  AND2_X1 u_majority7_module_13__and_module_4_U1 ( .A1(
        n_majority7_module_13__and_module_2_res), .A2(
        n_majority7_module_13__and_module_1_res), .ZN(
        n_majority7_module_13__and_module_4_res) );
  OR2_X1 u_majority7_module_13__or_module_4_U1 ( .A1(
        n_majority7_module_13__and_module_1_res), .A2(
        n_majority7_module_13__and_module_2_res), .ZN(
        n_majority7_module_13__or_module_4_res) );
  AND2_X1 u_majority7_module_13__and_module_5_U1 ( .A1(
        n_majority7_module_13__and_module_3_res), .A2(n_majority7_module_13_n4), .ZN(n_majority7_module_13__and_module_5_res) );
  OR2_X1 u_majority7_module_13__or_module_5_U1 ( .A1(n_majority7_module_13_n4), 
        .A2(n_majority7_module_13__and_module_3_res), .ZN(
        n_majority7_module_13__or_module_5_res) );
  AND2_X1 u_majority7_module_13__and_module_6_U1 ( .A1(
        n_majority7_module_13__or_module_1_res), .A2(
        n_majority7_module_13__or_module_2_res), .ZN(
        n_majority7_module_13__and_module_6_res) );
  OR2_X1 u_majority7_module_13__or_module_6_U1 ( .A1(
        n_majority7_module_13__or_module_2_res), .A2(
        n_majority7_module_13__or_module_1_res), .ZN(
        n_majority7_module_13__or_module_6_res) );
  OR2_X1 u_majority7_module_13__or_module_7_U1 ( .A1(
        n_majority7_module_13__and_module_4_res), .A2(
        n_majority7_module_13__and_module_5_res), .ZN(
        n_majority7_module_13__or_module_7_res) );
  AND2_X1 u_majority7_module_13__and_module_7_U1 ( .A1(
        n_majority7_module_13__or_module_3_res), .A2(
        n_majority7_module_13__or_module_4_res), .ZN(
        n_majority7_module_13__and_module_7_res) );
  OR2_X1 u_majority7_module_13__or_module_8_U1 ( .A1(
        n_majority7_module_13__or_module_4_res), .A2(
        n_majority7_module_13__or_module_3_res), .ZN(
        n_majority7_module_13__or_module_8_res) );
  AND2_X1 u_majority7_module_13__and_module_8_U1 ( .A1(
        n_majority7_module_13__or_module_5_res), .A2(
        n_majority7_module_13__and_module_6_res), .ZN(
        n_majority7_module_13__and_module_8_res) );
  OR2_X1 u_majority7_module_13__or_module_9_U1 ( .A1(
        n_majority7_module_13__and_module_6_res), .A2(
        n_majority7_module_13__or_module_5_res), .ZN(
        n_majority7_module_13__or_module_9_res) );
  OR2_X1 u_majority7_module_13__or_module_10_U1 ( .A1(
        n_majority7_module_13__or_module_7_res), .A2(
        n_majority7_module_13__and_module_7_res), .ZN(
        n_majority7_module_13__or_module_10_res) );
  AND2_X1 u_majority7_module_13__and_module_9_U1 ( .A1(
        n_majority7_module_13__or_module_6_res), .A2(
        n_majority7_module_13__or_module_9_res), .ZN(
        n_majority7_module_13__and_module_9_res) );
  OR2_X1 u_majority7_module_13__or_module_11_U1 ( .A1(
        n_majority7_module_13__or_module_10_res), .A2(
        n_majority7_module_13__and_module_8_res), .ZN(
        n_majority7_module_13__or_module_11_res) );
  AND2_X1 u_majority7_module_13__and_module_10_U1 ( .A1(
        n_majority7_module_13__or_module_8_res), .A2(
        n_majority7_module_13__and_module_9_res), .ZN(
        n_majority7_module_13__and_module_10_res) );
  AND2_X1 u_majority7_module_13__and_module_11_U1 ( .A1(
        n_majority7_module_13__and_module_10_res), .A2(
        n_majority7_module_13__or_module_11_res), .ZN(
        n_majority7_module_13_res) );
  DFF_X1 u_reg_module_14__cini_mul_v000_reg ( .D(n_majority7_module_13_res), 
        .CK(clock_0), .Q(n_reg_module_14_res), .QN() );
  BUF_X1 u_majority7_module_14_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_14_n7) );
  BUF_X1 u_majority7_module_14_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_14_n6) );
  BUF_X1 u_majority7_module_14_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_14_n5) );
  BUF_X1 u_majority7_module_14_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_14_n4) );
  BUF_X1 u_majority7_module_14_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_14_n3) );
  BUF_X1 u_majority7_module_14_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_14_n2) );
  BUF_X1 u_majority7_module_14_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_14_n1) );
  AND2_X1 u_majority7_module_14__and_module_1_U1 ( .A1(
        n_majority7_module_14_n1), .A2(n_majority7_module_14_n5), .ZN(
        n_majority7_module_14__and_module_1_res) );
  OR2_X1 u_majority7_module_14__or_module_1_U1 ( .A1(n_majority7_module_14_n5), 
        .A2(n_majority7_module_14_n1), .ZN(
        n_majority7_module_14__or_module_1_res) );
  AND2_X1 u_majority7_module_14__and_module_2_U1 ( .A1(
        n_majority7_module_14_n7), .A2(n_majority7_module_14_n3), .ZN(
        n_majority7_module_14__and_module_2_res) );
  OR2_X1 u_majority7_module_14__or_module_2_U1 ( .A1(n_majority7_module_14_n3), 
        .A2(n_majority7_module_14_n7), .ZN(
        n_majority7_module_14__or_module_2_res) );
  AND2_X1 u_majority7_module_14__and_module_3_U1 ( .A1(
        n_majority7_module_14_n6), .A2(n_majority7_module_14_n2), .ZN(
        n_majority7_module_14__and_module_3_res) );
  OR2_X1 u_majority7_module_14__or_module_3_U1 ( .A1(n_majority7_module_14_n2), 
        .A2(n_majority7_module_14_n6), .ZN(
        n_majority7_module_14__or_module_3_res) );
  AND2_X1 u_majority7_module_14__and_module_4_U1 ( .A1(
        n_majority7_module_14__and_module_2_res), .A2(
        n_majority7_module_14__and_module_1_res), .ZN(
        n_majority7_module_14__and_module_4_res) );
  OR2_X1 u_majority7_module_14__or_module_4_U1 ( .A1(
        n_majority7_module_14__and_module_1_res), .A2(
        n_majority7_module_14__and_module_2_res), .ZN(
        n_majority7_module_14__or_module_4_res) );
  AND2_X1 u_majority7_module_14__and_module_5_U1 ( .A1(
        n_majority7_module_14__and_module_3_res), .A2(n_majority7_module_14_n4), .ZN(n_majority7_module_14__and_module_5_res) );
  OR2_X1 u_majority7_module_14__or_module_5_U1 ( .A1(n_majority7_module_14_n4), 
        .A2(n_majority7_module_14__and_module_3_res), .ZN(
        n_majority7_module_14__or_module_5_res) );
  AND2_X1 u_majority7_module_14__and_module_6_U1 ( .A1(
        n_majority7_module_14__or_module_1_res), .A2(
        n_majority7_module_14__or_module_2_res), .ZN(
        n_majority7_module_14__and_module_6_res) );
  OR2_X1 u_majority7_module_14__or_module_6_U1 ( .A1(
        n_majority7_module_14__or_module_2_res), .A2(
        n_majority7_module_14__or_module_1_res), .ZN(
        n_majority7_module_14__or_module_6_res) );
  OR2_X1 u_majority7_module_14__or_module_7_U1 ( .A1(
        n_majority7_module_14__and_module_4_res), .A2(
        n_majority7_module_14__and_module_5_res), .ZN(
        n_majority7_module_14__or_module_7_res) );
  AND2_X1 u_majority7_module_14__and_module_7_U1 ( .A1(
        n_majority7_module_14__or_module_3_res), .A2(
        n_majority7_module_14__or_module_4_res), .ZN(
        n_majority7_module_14__and_module_7_res) );
  OR2_X1 u_majority7_module_14__or_module_8_U1 ( .A1(
        n_majority7_module_14__or_module_4_res), .A2(
        n_majority7_module_14__or_module_3_res), .ZN(
        n_majority7_module_14__or_module_8_res) );
  AND2_X1 u_majority7_module_14__and_module_8_U1 ( .A1(
        n_majority7_module_14__or_module_5_res), .A2(
        n_majority7_module_14__and_module_6_res), .ZN(
        n_majority7_module_14__and_module_8_res) );
  OR2_X1 u_majority7_module_14__or_module_9_U1 ( .A1(
        n_majority7_module_14__and_module_6_res), .A2(
        n_majority7_module_14__or_module_5_res), .ZN(
        n_majority7_module_14__or_module_9_res) );
  OR2_X1 u_majority7_module_14__or_module_10_U1 ( .A1(
        n_majority7_module_14__or_module_7_res), .A2(
        n_majority7_module_14__and_module_7_res), .ZN(
        n_majority7_module_14__or_module_10_res) );
  AND2_X1 u_majority7_module_14__and_module_9_U1 ( .A1(
        n_majority7_module_14__or_module_6_res), .A2(
        n_majority7_module_14__or_module_9_res), .ZN(
        n_majority7_module_14__and_module_9_res) );
  OR2_X1 u_majority7_module_14__or_module_11_U1 ( .A1(
        n_majority7_module_14__or_module_10_res), .A2(
        n_majority7_module_14__and_module_8_res), .ZN(
        n_majority7_module_14__or_module_11_res) );
  AND2_X1 u_majority7_module_14__and_module_10_U1 ( .A1(
        n_majority7_module_14__or_module_8_res), .A2(
        n_majority7_module_14__and_module_9_res), .ZN(
        n_majority7_module_14__and_module_10_res) );
  AND2_X1 u_majority7_module_14__and_module_11_U1 ( .A1(
        n_majority7_module_14__and_module_10_res), .A2(
        n_majority7_module_14__or_module_11_res), .ZN(
        n_majority7_module_14_res) );
  DFF_X1 u_reg_module_15__cini_mul_v000_reg ( .D(n_majority7_module_14_res), 
        .CK(clock_0), .Q(n_reg_module_15_res), .QN() );
  BUF_X1 u_majority7_module_15_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_15_n7) );
  BUF_X1 u_majority7_module_15_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_15_n6) );
  BUF_X1 u_majority7_module_15_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_15_n5) );
  BUF_X1 u_majority7_module_15_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_15_n4) );
  BUF_X1 u_majority7_module_15_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_15_n3) );
  BUF_X1 u_majority7_module_15_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_15_n2) );
  BUF_X1 u_majority7_module_15_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_15_n1) );
  AND2_X1 u_majority7_module_15__and_module_1_U1 ( .A1(
        n_majority7_module_15_n1), .A2(n_majority7_module_15_n5), .ZN(
        n_majority7_module_15__and_module_1_res) );
  OR2_X1 u_majority7_module_15__or_module_1_U1 ( .A1(n_majority7_module_15_n5), 
        .A2(n_majority7_module_15_n1), .ZN(
        n_majority7_module_15__or_module_1_res) );
  AND2_X1 u_majority7_module_15__and_module_2_U1 ( .A1(
        n_majority7_module_15_n7), .A2(n_majority7_module_15_n3), .ZN(
        n_majority7_module_15__and_module_2_res) );
  OR2_X1 u_majority7_module_15__or_module_2_U1 ( .A1(n_majority7_module_15_n3), 
        .A2(n_majority7_module_15_n7), .ZN(
        n_majority7_module_15__or_module_2_res) );
  AND2_X1 u_majority7_module_15__and_module_3_U1 ( .A1(
        n_majority7_module_15_n6), .A2(n_majority7_module_15_n2), .ZN(
        n_majority7_module_15__and_module_3_res) );
  OR2_X1 u_majority7_module_15__or_module_3_U1 ( .A1(n_majority7_module_15_n2), 
        .A2(n_majority7_module_15_n6), .ZN(
        n_majority7_module_15__or_module_3_res) );
  AND2_X1 u_majority7_module_15__and_module_4_U1 ( .A1(
        n_majority7_module_15__and_module_2_res), .A2(
        n_majority7_module_15__and_module_1_res), .ZN(
        n_majority7_module_15__and_module_4_res) );
  OR2_X1 u_majority7_module_15__or_module_4_U1 ( .A1(
        n_majority7_module_15__and_module_1_res), .A2(
        n_majority7_module_15__and_module_2_res), .ZN(
        n_majority7_module_15__or_module_4_res) );
  AND2_X1 u_majority7_module_15__and_module_5_U1 ( .A1(
        n_majority7_module_15__and_module_3_res), .A2(n_majority7_module_15_n4), .ZN(n_majority7_module_15__and_module_5_res) );
  OR2_X1 u_majority7_module_15__or_module_5_U1 ( .A1(n_majority7_module_15_n4), 
        .A2(n_majority7_module_15__and_module_3_res), .ZN(
        n_majority7_module_15__or_module_5_res) );
  AND2_X1 u_majority7_module_15__and_module_6_U1 ( .A1(
        n_majority7_module_15__or_module_1_res), .A2(
        n_majority7_module_15__or_module_2_res), .ZN(
        n_majority7_module_15__and_module_6_res) );
  OR2_X1 u_majority7_module_15__or_module_6_U1 ( .A1(
        n_majority7_module_15__or_module_2_res), .A2(
        n_majority7_module_15__or_module_1_res), .ZN(
        n_majority7_module_15__or_module_6_res) );
  OR2_X1 u_majority7_module_15__or_module_7_U1 ( .A1(
        n_majority7_module_15__and_module_4_res), .A2(
        n_majority7_module_15__and_module_5_res), .ZN(
        n_majority7_module_15__or_module_7_res) );
  AND2_X1 u_majority7_module_15__and_module_7_U1 ( .A1(
        n_majority7_module_15__or_module_3_res), .A2(
        n_majority7_module_15__or_module_4_res), .ZN(
        n_majority7_module_15__and_module_7_res) );
  OR2_X1 u_majority7_module_15__or_module_8_U1 ( .A1(
        n_majority7_module_15__or_module_4_res), .A2(
        n_majority7_module_15__or_module_3_res), .ZN(
        n_majority7_module_15__or_module_8_res) );
  AND2_X1 u_majority7_module_15__and_module_8_U1 ( .A1(
        n_majority7_module_15__or_module_5_res), .A2(
        n_majority7_module_15__and_module_6_res), .ZN(
        n_majority7_module_15__and_module_8_res) );
  OR2_X1 u_majority7_module_15__or_module_9_U1 ( .A1(
        n_majority7_module_15__and_module_6_res), .A2(
        n_majority7_module_15__or_module_5_res), .ZN(
        n_majority7_module_15__or_module_9_res) );
  OR2_X1 u_majority7_module_15__or_module_10_U1 ( .A1(
        n_majority7_module_15__or_module_7_res), .A2(
        n_majority7_module_15__and_module_7_res), .ZN(
        n_majority7_module_15__or_module_10_res) );
  AND2_X1 u_majority7_module_15__and_module_9_U1 ( .A1(
        n_majority7_module_15__or_module_6_res), .A2(
        n_majority7_module_15__or_module_9_res), .ZN(
        n_majority7_module_15__and_module_9_res) );
  OR2_X1 u_majority7_module_15__or_module_11_U1 ( .A1(
        n_majority7_module_15__or_module_10_res), .A2(
        n_majority7_module_15__and_module_8_res), .ZN(
        n_majority7_module_15__or_module_11_res) );
  AND2_X1 u_majority7_module_15__and_module_10_U1 ( .A1(
        n_majority7_module_15__or_module_8_res), .A2(
        n_majority7_module_15__and_module_9_res), .ZN(
        n_majority7_module_15__and_module_10_res) );
  AND2_X1 u_majority7_module_15__and_module_11_U1 ( .A1(
        n_majority7_module_15__and_module_10_res), .A2(
        n_majority7_module_15__or_module_11_res), .ZN(
        n_majority7_module_15_res) );
  DFF_X1 u_reg_module_16__cini_mul_v000_reg ( .D(n_majority7_module_15_res), 
        .CK(clock_0), .Q(n_reg_module_16_res), .QN() );
  BUF_X1 u_majority7_module_16_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_16_n7) );
  BUF_X1 u_majority7_module_16_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_16_n6) );
  BUF_X1 u_majority7_module_16_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_16_n5) );
  BUF_X1 u_majority7_module_16_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_16_n4) );
  BUF_X1 u_majority7_module_16_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_16_n3) );
  BUF_X1 u_majority7_module_16_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_16_n2) );
  BUF_X1 u_majority7_module_16_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_16_n1) );
  AND2_X1 u_majority7_module_16__and_module_1_U1 ( .A1(
        n_majority7_module_16_n5), .A2(n_majority7_module_16_n4), .ZN(
        n_majority7_module_16__and_module_1_res) );
  OR2_X1 u_majority7_module_16__or_module_1_U1 ( .A1(n_majority7_module_16_n4), 
        .A2(n_majority7_module_16_n5), .ZN(
        n_majority7_module_16__or_module_1_res) );
  AND2_X1 u_majority7_module_16__and_module_2_U1 ( .A1(
        n_majority7_module_16_n7), .A2(n_majority7_module_16_n2), .ZN(
        n_majority7_module_16__and_module_2_res) );
  OR2_X1 u_majority7_module_16__or_module_2_U1 ( .A1(n_majority7_module_16_n2), 
        .A2(n_majority7_module_16_n7), .ZN(
        n_majority7_module_16__or_module_2_res) );
  AND2_X1 u_majority7_module_16__and_module_3_U1 ( .A1(
        n_majority7_module_16_n6), .A2(n_majority7_module_16_n1), .ZN(
        n_majority7_module_16__and_module_3_res) );
  OR2_X1 u_majority7_module_16__or_module_3_U1 ( .A1(n_majority7_module_16_n1), 
        .A2(n_majority7_module_16_n6), .ZN(
        n_majority7_module_16__or_module_3_res) );
  AND2_X1 u_majority7_module_16__and_module_4_U1 ( .A1(
        n_majority7_module_16__and_module_2_res), .A2(
        n_majority7_module_16__and_module_1_res), .ZN(
        n_majority7_module_16__and_module_4_res) );
  OR2_X1 u_majority7_module_16__or_module_4_U1 ( .A1(
        n_majority7_module_16__and_module_1_res), .A2(
        n_majority7_module_16__and_module_2_res), .ZN(
        n_majority7_module_16__or_module_4_res) );
  AND2_X1 u_majority7_module_16__and_module_5_U1 ( .A1(
        n_majority7_module_16__and_module_3_res), .A2(n_majority7_module_16_n3), .ZN(n_majority7_module_16__and_module_5_res) );
  OR2_X1 u_majority7_module_16__or_module_5_U1 ( .A1(n_majority7_module_16_n3), 
        .A2(n_majority7_module_16__and_module_3_res), .ZN(
        n_majority7_module_16__or_module_5_res) );
  AND2_X1 u_majority7_module_16__and_module_6_U1 ( .A1(
        n_majority7_module_16__or_module_1_res), .A2(
        n_majority7_module_16__or_module_2_res), .ZN(
        n_majority7_module_16__and_module_6_res) );
  OR2_X1 u_majority7_module_16__or_module_6_U1 ( .A1(
        n_majority7_module_16__or_module_2_res), .A2(
        n_majority7_module_16__or_module_1_res), .ZN(
        n_majority7_module_16__or_module_6_res) );
  OR2_X1 u_majority7_module_16__or_module_7_U1 ( .A1(
        n_majority7_module_16__and_module_4_res), .A2(
        n_majority7_module_16__and_module_5_res), .ZN(
        n_majority7_module_16__or_module_7_res) );
  AND2_X1 u_majority7_module_16__and_module_7_U1 ( .A1(
        n_majority7_module_16__or_module_3_res), .A2(
        n_majority7_module_16__or_module_4_res), .ZN(
        n_majority7_module_16__and_module_7_res) );
  OR2_X1 u_majority7_module_16__or_module_8_U1 ( .A1(
        n_majority7_module_16__or_module_4_res), .A2(
        n_majority7_module_16__or_module_3_res), .ZN(
        n_majority7_module_16__or_module_8_res) );
  AND2_X1 u_majority7_module_16__and_module_8_U1 ( .A1(
        n_majority7_module_16__or_module_5_res), .A2(
        n_majority7_module_16__and_module_6_res), .ZN(
        n_majority7_module_16__and_module_8_res) );
  OR2_X1 u_majority7_module_16__or_module_9_U1 ( .A1(
        n_majority7_module_16__and_module_6_res), .A2(
        n_majority7_module_16__or_module_5_res), .ZN(
        n_majority7_module_16__or_module_9_res) );
  OR2_X1 u_majority7_module_16__or_module_10_U1 ( .A1(
        n_majority7_module_16__or_module_7_res), .A2(
        n_majority7_module_16__and_module_7_res), .ZN(
        n_majority7_module_16__or_module_10_res) );
  AND2_X1 u_majority7_module_16__and_module_9_U1 ( .A1(
        n_majority7_module_16__or_module_6_res), .A2(
        n_majority7_module_16__or_module_9_res), .ZN(
        n_majority7_module_16__and_module_9_res) );
  OR2_X1 u_majority7_module_16__or_module_11_U1 ( .A1(
        n_majority7_module_16__or_module_10_res), .A2(
        n_majority7_module_16__and_module_8_res), .ZN(
        n_majority7_module_16__or_module_11_res) );
  AND2_X1 u_majority7_module_16__and_module_10_U1 ( .A1(
        n_majority7_module_16__or_module_8_res), .A2(
        n_majority7_module_16__and_module_9_res), .ZN(
        n_majority7_module_16__and_module_10_res) );
  AND2_X1 u_majority7_module_16__and_module_11_U1 ( .A1(
        n_majority7_module_16__and_module_10_res), .A2(
        n_majority7_module_16__or_module_11_res), .ZN(
        n_majority7_module_16_res) );
  DFF_X1 u_reg_module_17__cini_mul_v000_reg ( .D(n_majority7_module_16_res), 
        .CK(clock_1), .Q(n_reg_module_17_res), .QN() );
  BUF_X1 u_majority7_module_17_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_17_n7) );
  BUF_X1 u_majority7_module_17_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_17_n6) );
  BUF_X1 u_majority7_module_17_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_17_n5) );
  BUF_X1 u_majority7_module_17_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_17_n4) );
  BUF_X1 u_majority7_module_17_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_17_n3) );
  BUF_X1 u_majority7_module_17_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_17_n2) );
  BUF_X1 u_majority7_module_17_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_17_n1) );
  AND2_X1 u_majority7_module_17__and_module_1_U1 ( .A1(
        n_majority7_module_17_n5), .A2(n_majority7_module_17_n4), .ZN(
        n_majority7_module_17__and_module_1_res) );
  OR2_X1 u_majority7_module_17__or_module_1_U1 ( .A1(n_majority7_module_17_n4), 
        .A2(n_majority7_module_17_n5), .ZN(
        n_majority7_module_17__or_module_1_res) );
  AND2_X1 u_majority7_module_17__and_module_2_U1 ( .A1(
        n_majority7_module_17_n7), .A2(n_majority7_module_17_n2), .ZN(
        n_majority7_module_17__and_module_2_res) );
  OR2_X1 u_majority7_module_17__or_module_2_U1 ( .A1(n_majority7_module_17_n2), 
        .A2(n_majority7_module_17_n7), .ZN(
        n_majority7_module_17__or_module_2_res) );
  AND2_X1 u_majority7_module_17__and_module_3_U1 ( .A1(
        n_majority7_module_17_n6), .A2(n_majority7_module_17_n1), .ZN(
        n_majority7_module_17__and_module_3_res) );
  OR2_X1 u_majority7_module_17__or_module_3_U1 ( .A1(n_majority7_module_17_n1), 
        .A2(n_majority7_module_17_n6), .ZN(
        n_majority7_module_17__or_module_3_res) );
  AND2_X1 u_majority7_module_17__and_module_4_U1 ( .A1(
        n_majority7_module_17__and_module_2_res), .A2(
        n_majority7_module_17__and_module_1_res), .ZN(
        n_majority7_module_17__and_module_4_res) );
  OR2_X1 u_majority7_module_17__or_module_4_U1 ( .A1(
        n_majority7_module_17__and_module_1_res), .A2(
        n_majority7_module_17__and_module_2_res), .ZN(
        n_majority7_module_17__or_module_4_res) );
  AND2_X1 u_majority7_module_17__and_module_5_U1 ( .A1(
        n_majority7_module_17__and_module_3_res), .A2(n_majority7_module_17_n3), .ZN(n_majority7_module_17__and_module_5_res) );
  OR2_X1 u_majority7_module_17__or_module_5_U1 ( .A1(n_majority7_module_17_n3), 
        .A2(n_majority7_module_17__and_module_3_res), .ZN(
        n_majority7_module_17__or_module_5_res) );
  AND2_X1 u_majority7_module_17__and_module_6_U1 ( .A1(
        n_majority7_module_17__or_module_1_res), .A2(
        n_majority7_module_17__or_module_2_res), .ZN(
        n_majority7_module_17__and_module_6_res) );
  OR2_X1 u_majority7_module_17__or_module_6_U1 ( .A1(
        n_majority7_module_17__or_module_2_res), .A2(
        n_majority7_module_17__or_module_1_res), .ZN(
        n_majority7_module_17__or_module_6_res) );
  OR2_X1 u_majority7_module_17__or_module_7_U1 ( .A1(
        n_majority7_module_17__and_module_4_res), .A2(
        n_majority7_module_17__and_module_5_res), .ZN(
        n_majority7_module_17__or_module_7_res) );
  AND2_X1 u_majority7_module_17__and_module_7_U1 ( .A1(
        n_majority7_module_17__or_module_3_res), .A2(
        n_majority7_module_17__or_module_4_res), .ZN(
        n_majority7_module_17__and_module_7_res) );
  OR2_X1 u_majority7_module_17__or_module_8_U1 ( .A1(
        n_majority7_module_17__or_module_4_res), .A2(
        n_majority7_module_17__or_module_3_res), .ZN(
        n_majority7_module_17__or_module_8_res) );
  AND2_X1 u_majority7_module_17__and_module_8_U1 ( .A1(
        n_majority7_module_17__or_module_5_res), .A2(
        n_majority7_module_17__and_module_6_res), .ZN(
        n_majority7_module_17__and_module_8_res) );
  OR2_X1 u_majority7_module_17__or_module_9_U1 ( .A1(
        n_majority7_module_17__and_module_6_res), .A2(
        n_majority7_module_17__or_module_5_res), .ZN(
        n_majority7_module_17__or_module_9_res) );
  OR2_X1 u_majority7_module_17__or_module_10_U1 ( .A1(
        n_majority7_module_17__or_module_7_res), .A2(
        n_majority7_module_17__and_module_7_res), .ZN(
        n_majority7_module_17__or_module_10_res) );
  AND2_X1 u_majority7_module_17__and_module_9_U1 ( .A1(
        n_majority7_module_17__or_module_6_res), .A2(
        n_majority7_module_17__or_module_9_res), .ZN(
        n_majority7_module_17__and_module_9_res) );
  OR2_X1 u_majority7_module_17__or_module_11_U1 ( .A1(
        n_majority7_module_17__or_module_10_res), .A2(
        n_majority7_module_17__and_module_8_res), .ZN(
        n_majority7_module_17__or_module_11_res) );
  AND2_X1 u_majority7_module_17__and_module_10_U1 ( .A1(
        n_majority7_module_17__or_module_8_res), .A2(
        n_majority7_module_17__and_module_9_res), .ZN(
        n_majority7_module_17__and_module_10_res) );
  AND2_X1 u_majority7_module_17__and_module_11_U1 ( .A1(
        n_majority7_module_17__and_module_10_res), .A2(
        n_majority7_module_17__or_module_11_res), .ZN(
        n_majority7_module_17_res) );
  DFF_X1 u_reg_module_18__cini_mul_v000_reg ( .D(n_majority7_module_17_res), 
        .CK(clock_1), .Q(n_reg_module_18_res), .QN() );
  BUF_X1 u_majority7_module_18_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_18_n7) );
  BUF_X1 u_majority7_module_18_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_18_n6) );
  BUF_X1 u_majority7_module_18_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_18_n5) );
  BUF_X1 u_majority7_module_18_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_18_n4) );
  BUF_X1 u_majority7_module_18_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_18_n3) );
  BUF_X1 u_majority7_module_18_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_18_n2) );
  BUF_X1 u_majority7_module_18_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_18_n1) );
  AND2_X1 u_majority7_module_18__and_module_1_U1 ( .A1(
        n_majority7_module_18_n5), .A2(n_majority7_module_18_n4), .ZN(
        n_majority7_module_18__and_module_1_res) );
  OR2_X1 u_majority7_module_18__or_module_1_U1 ( .A1(n_majority7_module_18_n4), 
        .A2(n_majority7_module_18_n5), .ZN(
        n_majority7_module_18__or_module_1_res) );
  AND2_X1 u_majority7_module_18__and_module_2_U1 ( .A1(
        n_majority7_module_18_n7), .A2(n_majority7_module_18_n2), .ZN(
        n_majority7_module_18__and_module_2_res) );
  OR2_X1 u_majority7_module_18__or_module_2_U1 ( .A1(n_majority7_module_18_n2), 
        .A2(n_majority7_module_18_n7), .ZN(
        n_majority7_module_18__or_module_2_res) );
  AND2_X1 u_majority7_module_18__and_module_3_U1 ( .A1(
        n_majority7_module_18_n6), .A2(n_majority7_module_18_n1), .ZN(
        n_majority7_module_18__and_module_3_res) );
  OR2_X1 u_majority7_module_18__or_module_3_U1 ( .A1(n_majority7_module_18_n1), 
        .A2(n_majority7_module_18_n6), .ZN(
        n_majority7_module_18__or_module_3_res) );
  AND2_X1 u_majority7_module_18__and_module_4_U1 ( .A1(
        n_majority7_module_18__and_module_2_res), .A2(
        n_majority7_module_18__and_module_1_res), .ZN(
        n_majority7_module_18__and_module_4_res) );
  OR2_X1 u_majority7_module_18__or_module_4_U1 ( .A1(
        n_majority7_module_18__and_module_1_res), .A2(
        n_majority7_module_18__and_module_2_res), .ZN(
        n_majority7_module_18__or_module_4_res) );
  AND2_X1 u_majority7_module_18__and_module_5_U1 ( .A1(
        n_majority7_module_18__and_module_3_res), .A2(n_majority7_module_18_n3), .ZN(n_majority7_module_18__and_module_5_res) );
  OR2_X1 u_majority7_module_18__or_module_5_U1 ( .A1(n_majority7_module_18_n3), 
        .A2(n_majority7_module_18__and_module_3_res), .ZN(
        n_majority7_module_18__or_module_5_res) );
  AND2_X1 u_majority7_module_18__and_module_6_U1 ( .A1(
        n_majority7_module_18__or_module_1_res), .A2(
        n_majority7_module_18__or_module_2_res), .ZN(
        n_majority7_module_18__and_module_6_res) );
  OR2_X1 u_majority7_module_18__or_module_6_U1 ( .A1(
        n_majority7_module_18__or_module_2_res), .A2(
        n_majority7_module_18__or_module_1_res), .ZN(
        n_majority7_module_18__or_module_6_res) );
  OR2_X1 u_majority7_module_18__or_module_7_U1 ( .A1(
        n_majority7_module_18__and_module_4_res), .A2(
        n_majority7_module_18__and_module_5_res), .ZN(
        n_majority7_module_18__or_module_7_res) );
  AND2_X1 u_majority7_module_18__and_module_7_U1 ( .A1(
        n_majority7_module_18__or_module_3_res), .A2(
        n_majority7_module_18__or_module_4_res), .ZN(
        n_majority7_module_18__and_module_7_res) );
  OR2_X1 u_majority7_module_18__or_module_8_U1 ( .A1(
        n_majority7_module_18__or_module_4_res), .A2(
        n_majority7_module_18__or_module_3_res), .ZN(
        n_majority7_module_18__or_module_8_res) );
  AND2_X1 u_majority7_module_18__and_module_8_U1 ( .A1(
        n_majority7_module_18__or_module_5_res), .A2(
        n_majority7_module_18__and_module_6_res), .ZN(
        n_majority7_module_18__and_module_8_res) );
  OR2_X1 u_majority7_module_18__or_module_9_U1 ( .A1(
        n_majority7_module_18__and_module_6_res), .A2(
        n_majority7_module_18__or_module_5_res), .ZN(
        n_majority7_module_18__or_module_9_res) );
  OR2_X1 u_majority7_module_18__or_module_10_U1 ( .A1(
        n_majority7_module_18__or_module_7_res), .A2(
        n_majority7_module_18__and_module_7_res), .ZN(
        n_majority7_module_18__or_module_10_res) );
  AND2_X1 u_majority7_module_18__and_module_9_U1 ( .A1(
        n_majority7_module_18__or_module_6_res), .A2(
        n_majority7_module_18__or_module_9_res), .ZN(
        n_majority7_module_18__and_module_9_res) );
  OR2_X1 u_majority7_module_18__or_module_11_U1 ( .A1(
        n_majority7_module_18__or_module_10_res), .A2(
        n_majority7_module_18__and_module_8_res), .ZN(
        n_majority7_module_18__or_module_11_res) );
  AND2_X1 u_majority7_module_18__and_module_10_U1 ( .A1(
        n_majority7_module_18__or_module_8_res), .A2(
        n_majority7_module_18__and_module_9_res), .ZN(
        n_majority7_module_18__and_module_10_res) );
  AND2_X1 u_majority7_module_18__and_module_11_U1 ( .A1(
        n_majority7_module_18__and_module_10_res), .A2(
        n_majority7_module_18__or_module_11_res), .ZN(
        n_majority7_module_18_res) );
  DFF_X1 u_reg_module_19__cini_mul_v000_reg ( .D(n_majority7_module_18_res), 
        .CK(clock_1), .Q(n_reg_module_19_res), .QN() );
  BUF_X1 u_majority7_module_19_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_19_n7) );
  BUF_X1 u_majority7_module_19_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_19_n6) );
  BUF_X1 u_majority7_module_19_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_19_n5) );
  BUF_X1 u_majority7_module_19_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_19_n4) );
  BUF_X1 u_majority7_module_19_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_19_n3) );
  BUF_X1 u_majority7_module_19_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_19_n2) );
  BUF_X1 u_majority7_module_19_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_19_n1) );
  AND2_X1 u_majority7_module_19__and_module_1_U1 ( .A1(
        n_majority7_module_19_n5), .A2(n_majority7_module_19_n4), .ZN(
        n_majority7_module_19__and_module_1_res) );
  OR2_X1 u_majority7_module_19__or_module_1_U1 ( .A1(n_majority7_module_19_n4), 
        .A2(n_majority7_module_19_n5), .ZN(
        n_majority7_module_19__or_module_1_res) );
  AND2_X1 u_majority7_module_19__and_module_2_U1 ( .A1(
        n_majority7_module_19_n7), .A2(n_majority7_module_19_n2), .ZN(
        n_majority7_module_19__and_module_2_res) );
  OR2_X1 u_majority7_module_19__or_module_2_U1 ( .A1(n_majority7_module_19_n2), 
        .A2(n_majority7_module_19_n7), .ZN(
        n_majority7_module_19__or_module_2_res) );
  AND2_X1 u_majority7_module_19__and_module_3_U1 ( .A1(
        n_majority7_module_19_n6), .A2(n_majority7_module_19_n1), .ZN(
        n_majority7_module_19__and_module_3_res) );
  OR2_X1 u_majority7_module_19__or_module_3_U1 ( .A1(n_majority7_module_19_n1), 
        .A2(n_majority7_module_19_n6), .ZN(
        n_majority7_module_19__or_module_3_res) );
  AND2_X1 u_majority7_module_19__and_module_4_U1 ( .A1(
        n_majority7_module_19__and_module_2_res), .A2(
        n_majority7_module_19__and_module_1_res), .ZN(
        n_majority7_module_19__and_module_4_res) );
  OR2_X1 u_majority7_module_19__or_module_4_U1 ( .A1(
        n_majority7_module_19__and_module_1_res), .A2(
        n_majority7_module_19__and_module_2_res), .ZN(
        n_majority7_module_19__or_module_4_res) );
  AND2_X1 u_majority7_module_19__and_module_5_U1 ( .A1(
        n_majority7_module_19__and_module_3_res), .A2(n_majority7_module_19_n3), .ZN(n_majority7_module_19__and_module_5_res) );
  OR2_X1 u_majority7_module_19__or_module_5_U1 ( .A1(n_majority7_module_19_n3), 
        .A2(n_majority7_module_19__and_module_3_res), .ZN(
        n_majority7_module_19__or_module_5_res) );
  AND2_X1 u_majority7_module_19__and_module_6_U1 ( .A1(
        n_majority7_module_19__or_module_1_res), .A2(
        n_majority7_module_19__or_module_2_res), .ZN(
        n_majority7_module_19__and_module_6_res) );
  OR2_X1 u_majority7_module_19__or_module_6_U1 ( .A1(
        n_majority7_module_19__or_module_2_res), .A2(
        n_majority7_module_19__or_module_1_res), .ZN(
        n_majority7_module_19__or_module_6_res) );
  OR2_X1 u_majority7_module_19__or_module_7_U1 ( .A1(
        n_majority7_module_19__and_module_4_res), .A2(
        n_majority7_module_19__and_module_5_res), .ZN(
        n_majority7_module_19__or_module_7_res) );
  AND2_X1 u_majority7_module_19__and_module_7_U1 ( .A1(
        n_majority7_module_19__or_module_3_res), .A2(
        n_majority7_module_19__or_module_4_res), .ZN(
        n_majority7_module_19__and_module_7_res) );
  OR2_X1 u_majority7_module_19__or_module_8_U1 ( .A1(
        n_majority7_module_19__or_module_4_res), .A2(
        n_majority7_module_19__or_module_3_res), .ZN(
        n_majority7_module_19__or_module_8_res) );
  AND2_X1 u_majority7_module_19__and_module_8_U1 ( .A1(
        n_majority7_module_19__or_module_5_res), .A2(
        n_majority7_module_19__and_module_6_res), .ZN(
        n_majority7_module_19__and_module_8_res) );
  OR2_X1 u_majority7_module_19__or_module_9_U1 ( .A1(
        n_majority7_module_19__and_module_6_res), .A2(
        n_majority7_module_19__or_module_5_res), .ZN(
        n_majority7_module_19__or_module_9_res) );
  OR2_X1 u_majority7_module_19__or_module_10_U1 ( .A1(
        n_majority7_module_19__or_module_7_res), .A2(
        n_majority7_module_19__and_module_7_res), .ZN(
        n_majority7_module_19__or_module_10_res) );
  AND2_X1 u_majority7_module_19__and_module_9_U1 ( .A1(
        n_majority7_module_19__or_module_6_res), .A2(
        n_majority7_module_19__or_module_9_res), .ZN(
        n_majority7_module_19__and_module_9_res) );
  OR2_X1 u_majority7_module_19__or_module_11_U1 ( .A1(
        n_majority7_module_19__or_module_10_res), .A2(
        n_majority7_module_19__and_module_8_res), .ZN(
        n_majority7_module_19__or_module_11_res) );
  AND2_X1 u_majority7_module_19__and_module_10_U1 ( .A1(
        n_majority7_module_19__or_module_8_res), .A2(
        n_majority7_module_19__and_module_9_res), .ZN(
        n_majority7_module_19__and_module_10_res) );
  AND2_X1 u_majority7_module_19__and_module_11_U1 ( .A1(
        n_majority7_module_19__and_module_10_res), .A2(
        n_majority7_module_19__or_module_11_res), .ZN(
        n_majority7_module_19_res) );
  DFF_X1 u_reg_module_20__cini_mul_v000_reg ( .D(n_majority7_module_19_res), 
        .CK(clock_1), .Q(n_reg_module_20_res), .QN() );
  BUF_X1 u_majority7_module_20_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_20_n7) );
  BUF_X1 u_majority7_module_20_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_20_n6) );
  BUF_X1 u_majority7_module_20_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_20_n5) );
  BUF_X1 u_majority7_module_20_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_20_n4) );
  BUF_X1 u_majority7_module_20_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_20_n3) );
  BUF_X1 u_majority7_module_20_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_20_n2) );
  BUF_X1 u_majority7_module_20_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_20_n1) );
  AND2_X1 u_majority7_module_20__and_module_1_U1 ( .A1(
        n_majority7_module_20_n5), .A2(n_majority7_module_20_n4), .ZN(
        n_majority7_module_20__and_module_1_res) );
  OR2_X1 u_majority7_module_20__or_module_1_U1 ( .A1(n_majority7_module_20_n4), 
        .A2(n_majority7_module_20_n5), .ZN(
        n_majority7_module_20__or_module_1_res) );
  AND2_X1 u_majority7_module_20__and_module_2_U1 ( .A1(
        n_majority7_module_20_n7), .A2(n_majority7_module_20_n2), .ZN(
        n_majority7_module_20__and_module_2_res) );
  OR2_X1 u_majority7_module_20__or_module_2_U1 ( .A1(n_majority7_module_20_n2), 
        .A2(n_majority7_module_20_n7), .ZN(
        n_majority7_module_20__or_module_2_res) );
  AND2_X1 u_majority7_module_20__and_module_3_U1 ( .A1(
        n_majority7_module_20_n6), .A2(n_majority7_module_20_n1), .ZN(
        n_majority7_module_20__and_module_3_res) );
  OR2_X1 u_majority7_module_20__or_module_3_U1 ( .A1(n_majority7_module_20_n1), 
        .A2(n_majority7_module_20_n6), .ZN(
        n_majority7_module_20__or_module_3_res) );
  AND2_X1 u_majority7_module_20__and_module_4_U1 ( .A1(
        n_majority7_module_20__and_module_2_res), .A2(
        n_majority7_module_20__and_module_1_res), .ZN(
        n_majority7_module_20__and_module_4_res) );
  OR2_X1 u_majority7_module_20__or_module_4_U1 ( .A1(
        n_majority7_module_20__and_module_1_res), .A2(
        n_majority7_module_20__and_module_2_res), .ZN(
        n_majority7_module_20__or_module_4_res) );
  AND2_X1 u_majority7_module_20__and_module_5_U1 ( .A1(
        n_majority7_module_20__and_module_3_res), .A2(n_majority7_module_20_n3), .ZN(n_majority7_module_20__and_module_5_res) );
  OR2_X1 u_majority7_module_20__or_module_5_U1 ( .A1(n_majority7_module_20_n3), 
        .A2(n_majority7_module_20__and_module_3_res), .ZN(
        n_majority7_module_20__or_module_5_res) );
  AND2_X1 u_majority7_module_20__and_module_6_U1 ( .A1(
        n_majority7_module_20__or_module_1_res), .A2(
        n_majority7_module_20__or_module_2_res), .ZN(
        n_majority7_module_20__and_module_6_res) );
  OR2_X1 u_majority7_module_20__or_module_6_U1 ( .A1(
        n_majority7_module_20__or_module_2_res), .A2(
        n_majority7_module_20__or_module_1_res), .ZN(
        n_majority7_module_20__or_module_6_res) );
  OR2_X1 u_majority7_module_20__or_module_7_U1 ( .A1(
        n_majority7_module_20__and_module_4_res), .A2(
        n_majority7_module_20__and_module_5_res), .ZN(
        n_majority7_module_20__or_module_7_res) );
  AND2_X1 u_majority7_module_20__and_module_7_U1 ( .A1(
        n_majority7_module_20__or_module_3_res), .A2(
        n_majority7_module_20__or_module_4_res), .ZN(
        n_majority7_module_20__and_module_7_res) );
  OR2_X1 u_majority7_module_20__or_module_8_U1 ( .A1(
        n_majority7_module_20__or_module_4_res), .A2(
        n_majority7_module_20__or_module_3_res), .ZN(
        n_majority7_module_20__or_module_8_res) );
  AND2_X1 u_majority7_module_20__and_module_8_U1 ( .A1(
        n_majority7_module_20__or_module_5_res), .A2(
        n_majority7_module_20__and_module_6_res), .ZN(
        n_majority7_module_20__and_module_8_res) );
  OR2_X1 u_majority7_module_20__or_module_9_U1 ( .A1(
        n_majority7_module_20__and_module_6_res), .A2(
        n_majority7_module_20__or_module_5_res), .ZN(
        n_majority7_module_20__or_module_9_res) );
  OR2_X1 u_majority7_module_20__or_module_10_U1 ( .A1(
        n_majority7_module_20__or_module_7_res), .A2(
        n_majority7_module_20__and_module_7_res), .ZN(
        n_majority7_module_20__or_module_10_res) );
  AND2_X1 u_majority7_module_20__and_module_9_U1 ( .A1(
        n_majority7_module_20__or_module_6_res), .A2(
        n_majority7_module_20__or_module_9_res), .ZN(
        n_majority7_module_20__and_module_9_res) );
  OR2_X1 u_majority7_module_20__or_module_11_U1 ( .A1(
        n_majority7_module_20__or_module_10_res), .A2(
        n_majority7_module_20__and_module_8_res), .ZN(
        n_majority7_module_20__or_module_11_res) );
  AND2_X1 u_majority7_module_20__and_module_10_U1 ( .A1(
        n_majority7_module_20__or_module_8_res), .A2(
        n_majority7_module_20__and_module_9_res), .ZN(
        n_majority7_module_20__and_module_10_res) );
  AND2_X1 u_majority7_module_20__and_module_11_U1 ( .A1(
        n_majority7_module_20__and_module_10_res), .A2(
        n_majority7_module_20__or_module_11_res), .ZN(
        n_majority7_module_20_res) );
  DFF_X1 u_reg_module_21__cini_mul_v000_reg ( .D(n_majority7_module_20_res), 
        .CK(clock_1), .Q(n_reg_module_21_res), .QN() );
  BUF_X1 u_majority7_module_21_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_21_n7) );
  BUF_X1 u_majority7_module_21_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_21_n6) );
  BUF_X1 u_majority7_module_21_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_21_n5) );
  BUF_X1 u_majority7_module_21_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_21_n4) );
  BUF_X1 u_majority7_module_21_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_21_n3) );
  BUF_X1 u_majority7_module_21_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_21_n2) );
  BUF_X1 u_majority7_module_21_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_21_n1) );
  AND2_X1 u_majority7_module_21__and_module_1_U1 ( .A1(
        n_majority7_module_21_n5), .A2(n_majority7_module_21_n4), .ZN(
        n_majority7_module_21__and_module_1_res) );
  OR2_X1 u_majority7_module_21__or_module_1_U1 ( .A1(n_majority7_module_21_n4), 
        .A2(n_majority7_module_21_n5), .ZN(
        n_majority7_module_21__or_module_1_res) );
  AND2_X1 u_majority7_module_21__and_module_2_U1 ( .A1(
        n_majority7_module_21_n7), .A2(n_majority7_module_21_n2), .ZN(
        n_majority7_module_21__and_module_2_res) );
  OR2_X1 u_majority7_module_21__or_module_2_U1 ( .A1(n_majority7_module_21_n2), 
        .A2(n_majority7_module_21_n7), .ZN(
        n_majority7_module_21__or_module_2_res) );
  AND2_X1 u_majority7_module_21__and_module_3_U1 ( .A1(
        n_majority7_module_21_n6), .A2(n_majority7_module_21_n1), .ZN(
        n_majority7_module_21__and_module_3_res) );
  OR2_X1 u_majority7_module_21__or_module_3_U1 ( .A1(n_majority7_module_21_n1), 
        .A2(n_majority7_module_21_n6), .ZN(
        n_majority7_module_21__or_module_3_res) );
  AND2_X1 u_majority7_module_21__and_module_4_U1 ( .A1(
        n_majority7_module_21__and_module_2_res), .A2(
        n_majority7_module_21__and_module_1_res), .ZN(
        n_majority7_module_21__and_module_4_res) );
  OR2_X1 u_majority7_module_21__or_module_4_U1 ( .A1(
        n_majority7_module_21__and_module_1_res), .A2(
        n_majority7_module_21__and_module_2_res), .ZN(
        n_majority7_module_21__or_module_4_res) );
  AND2_X1 u_majority7_module_21__and_module_5_U1 ( .A1(
        n_majority7_module_21__and_module_3_res), .A2(n_majority7_module_21_n3), .ZN(n_majority7_module_21__and_module_5_res) );
  OR2_X1 u_majority7_module_21__or_module_5_U1 ( .A1(n_majority7_module_21_n3), 
        .A2(n_majority7_module_21__and_module_3_res), .ZN(
        n_majority7_module_21__or_module_5_res) );
  AND2_X1 u_majority7_module_21__and_module_6_U1 ( .A1(
        n_majority7_module_21__or_module_1_res), .A2(
        n_majority7_module_21__or_module_2_res), .ZN(
        n_majority7_module_21__and_module_6_res) );
  OR2_X1 u_majority7_module_21__or_module_6_U1 ( .A1(
        n_majority7_module_21__or_module_2_res), .A2(
        n_majority7_module_21__or_module_1_res), .ZN(
        n_majority7_module_21__or_module_6_res) );
  OR2_X1 u_majority7_module_21__or_module_7_U1 ( .A1(
        n_majority7_module_21__and_module_4_res), .A2(
        n_majority7_module_21__and_module_5_res), .ZN(
        n_majority7_module_21__or_module_7_res) );
  AND2_X1 u_majority7_module_21__and_module_7_U1 ( .A1(
        n_majority7_module_21__or_module_3_res), .A2(
        n_majority7_module_21__or_module_4_res), .ZN(
        n_majority7_module_21__and_module_7_res) );
  OR2_X1 u_majority7_module_21__or_module_8_U1 ( .A1(
        n_majority7_module_21__or_module_4_res), .A2(
        n_majority7_module_21__or_module_3_res), .ZN(
        n_majority7_module_21__or_module_8_res) );
  AND2_X1 u_majority7_module_21__and_module_8_U1 ( .A1(
        n_majority7_module_21__or_module_5_res), .A2(
        n_majority7_module_21__and_module_6_res), .ZN(
        n_majority7_module_21__and_module_8_res) );
  OR2_X1 u_majority7_module_21__or_module_9_U1 ( .A1(
        n_majority7_module_21__and_module_6_res), .A2(
        n_majority7_module_21__or_module_5_res), .ZN(
        n_majority7_module_21__or_module_9_res) );
  OR2_X1 u_majority7_module_21__or_module_10_U1 ( .A1(
        n_majority7_module_21__or_module_7_res), .A2(
        n_majority7_module_21__and_module_7_res), .ZN(
        n_majority7_module_21__or_module_10_res) );
  AND2_X1 u_majority7_module_21__and_module_9_U1 ( .A1(
        n_majority7_module_21__or_module_6_res), .A2(
        n_majority7_module_21__or_module_9_res), .ZN(
        n_majority7_module_21__and_module_9_res) );
  OR2_X1 u_majority7_module_21__or_module_11_U1 ( .A1(
        n_majority7_module_21__or_module_10_res), .A2(
        n_majority7_module_21__and_module_8_res), .ZN(
        n_majority7_module_21__or_module_11_res) );
  AND2_X1 u_majority7_module_21__and_module_10_U1 ( .A1(
        n_majority7_module_21__or_module_8_res), .A2(
        n_majority7_module_21__and_module_9_res), .ZN(
        n_majority7_module_21__and_module_10_res) );
  AND2_X1 u_majority7_module_21__and_module_11_U1 ( .A1(
        n_majority7_module_21__and_module_10_res), .A2(
        n_majority7_module_21__or_module_11_res), .ZN(
        n_majority7_module_21_res) );
  DFF_X1 u_reg_module_22__cini_mul_v000_reg ( .D(n_majority7_module_21_res), 
        .CK(clock_1), .Q(n_reg_module_22_res), .QN() );
  BUF_X1 u_majority7_module_22_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_22_n7) );
  BUF_X1 u_majority7_module_22_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_22_n6) );
  BUF_X1 u_majority7_module_22_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_22_n5) );
  BUF_X1 u_majority7_module_22_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_22_n4) );
  BUF_X1 u_majority7_module_22_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_22_n3) );
  BUF_X1 u_majority7_module_22_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_22_n2) );
  BUF_X1 u_majority7_module_22_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_22_n1) );
  AND2_X1 u_majority7_module_22__and_module_1_U1 ( .A1(
        n_majority7_module_22_n5), .A2(n_majority7_module_22_n4), .ZN(
        n_majority7_module_22__and_module_1_res) );
  OR2_X1 u_majority7_module_22__or_module_1_U1 ( .A1(n_majority7_module_22_n4), 
        .A2(n_majority7_module_22_n5), .ZN(
        n_majority7_module_22__or_module_1_res) );
  AND2_X1 u_majority7_module_22__and_module_2_U1 ( .A1(
        n_majority7_module_22_n7), .A2(n_majority7_module_22_n2), .ZN(
        n_majority7_module_22__and_module_2_res) );
  OR2_X1 u_majority7_module_22__or_module_2_U1 ( .A1(n_majority7_module_22_n2), 
        .A2(n_majority7_module_22_n7), .ZN(
        n_majority7_module_22__or_module_2_res) );
  AND2_X1 u_majority7_module_22__and_module_3_U1 ( .A1(
        n_majority7_module_22_n6), .A2(n_majority7_module_22_n1), .ZN(
        n_majority7_module_22__and_module_3_res) );
  OR2_X1 u_majority7_module_22__or_module_3_U1 ( .A1(n_majority7_module_22_n1), 
        .A2(n_majority7_module_22_n6), .ZN(
        n_majority7_module_22__or_module_3_res) );
  AND2_X1 u_majority7_module_22__and_module_4_U1 ( .A1(
        n_majority7_module_22__and_module_2_res), .A2(
        n_majority7_module_22__and_module_1_res), .ZN(
        n_majority7_module_22__and_module_4_res) );
  OR2_X1 u_majority7_module_22__or_module_4_U1 ( .A1(
        n_majority7_module_22__and_module_1_res), .A2(
        n_majority7_module_22__and_module_2_res), .ZN(
        n_majority7_module_22__or_module_4_res) );
  AND2_X1 u_majority7_module_22__and_module_5_U1 ( .A1(
        n_majority7_module_22__and_module_3_res), .A2(n_majority7_module_22_n3), .ZN(n_majority7_module_22__and_module_5_res) );
  OR2_X1 u_majority7_module_22__or_module_5_U1 ( .A1(n_majority7_module_22_n3), 
        .A2(n_majority7_module_22__and_module_3_res), .ZN(
        n_majority7_module_22__or_module_5_res) );
  AND2_X1 u_majority7_module_22__and_module_6_U1 ( .A1(
        n_majority7_module_22__or_module_1_res), .A2(
        n_majority7_module_22__or_module_2_res), .ZN(
        n_majority7_module_22__and_module_6_res) );
  OR2_X1 u_majority7_module_22__or_module_6_U1 ( .A1(
        n_majority7_module_22__or_module_2_res), .A2(
        n_majority7_module_22__or_module_1_res), .ZN(
        n_majority7_module_22__or_module_6_res) );
  OR2_X1 u_majority7_module_22__or_module_7_U1 ( .A1(
        n_majority7_module_22__and_module_4_res), .A2(
        n_majority7_module_22__and_module_5_res), .ZN(
        n_majority7_module_22__or_module_7_res) );
  AND2_X1 u_majority7_module_22__and_module_7_U1 ( .A1(
        n_majority7_module_22__or_module_3_res), .A2(
        n_majority7_module_22__or_module_4_res), .ZN(
        n_majority7_module_22__and_module_7_res) );
  OR2_X1 u_majority7_module_22__or_module_8_U1 ( .A1(
        n_majority7_module_22__or_module_4_res), .A2(
        n_majority7_module_22__or_module_3_res), .ZN(
        n_majority7_module_22__or_module_8_res) );
  AND2_X1 u_majority7_module_22__and_module_8_U1 ( .A1(
        n_majority7_module_22__or_module_5_res), .A2(
        n_majority7_module_22__and_module_6_res), .ZN(
        n_majority7_module_22__and_module_8_res) );
  OR2_X1 u_majority7_module_22__or_module_9_U1 ( .A1(
        n_majority7_module_22__and_module_6_res), .A2(
        n_majority7_module_22__or_module_5_res), .ZN(
        n_majority7_module_22__or_module_9_res) );
  OR2_X1 u_majority7_module_22__or_module_10_U1 ( .A1(
        n_majority7_module_22__or_module_7_res), .A2(
        n_majority7_module_22__and_module_7_res), .ZN(
        n_majority7_module_22__or_module_10_res) );
  AND2_X1 u_majority7_module_22__and_module_9_U1 ( .A1(
        n_majority7_module_22__or_module_6_res), .A2(
        n_majority7_module_22__or_module_9_res), .ZN(
        n_majority7_module_22__and_module_9_res) );
  OR2_X1 u_majority7_module_22__or_module_11_U1 ( .A1(
        n_majority7_module_22__or_module_10_res), .A2(
        n_majority7_module_22__and_module_8_res), .ZN(
        n_majority7_module_22__or_module_11_res) );
  AND2_X1 u_majority7_module_22__and_module_10_U1 ( .A1(
        n_majority7_module_22__or_module_8_res), .A2(
        n_majority7_module_22__and_module_9_res), .ZN(
        n_majority7_module_22__and_module_10_res) );
  AND2_X1 u_majority7_module_22__and_module_11_U1 ( .A1(
        n_majority7_module_22__and_module_10_res), .A2(
        n_majority7_module_22__or_module_11_res), .ZN(
        n_majority7_module_22_res) );
  DFF_X1 u_reg_module_23__cini_mul_v000_reg ( .D(n_majority7_module_22_res), 
        .CK(clock_1), .Q(n_reg_module_23_res), .QN() );
  BUF_X1 u_majority7_module_23_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_23_n7) );
  BUF_X1 u_majority7_module_23_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_23_n6) );
  BUF_X1 u_majority7_module_23_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_23_n5) );
  BUF_X1 u_majority7_module_23_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_23_n4) );
  BUF_X1 u_majority7_module_23_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_23_n3) );
  BUF_X1 u_majority7_module_23_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_23_n2) );
  BUF_X1 u_majority7_module_23_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_23_n1) );
  AND2_X1 u_majority7_module_23__and_module_1_U1 ( .A1(
        n_majority7_module_23_n5), .A2(n_majority7_module_23_n4), .ZN(
        n_majority7_module_23__and_module_1_res) );
  OR2_X1 u_majority7_module_23__or_module_1_U1 ( .A1(n_majority7_module_23_n4), 
        .A2(n_majority7_module_23_n5), .ZN(
        n_majority7_module_23__or_module_1_res) );
  AND2_X1 u_majority7_module_23__and_module_2_U1 ( .A1(
        n_majority7_module_23_n7), .A2(n_majority7_module_23_n2), .ZN(
        n_majority7_module_23__and_module_2_res) );
  OR2_X1 u_majority7_module_23__or_module_2_U1 ( .A1(n_majority7_module_23_n2), 
        .A2(n_majority7_module_23_n7), .ZN(
        n_majority7_module_23__or_module_2_res) );
  AND2_X1 u_majority7_module_23__and_module_3_U1 ( .A1(
        n_majority7_module_23_n6), .A2(n_majority7_module_23_n1), .ZN(
        n_majority7_module_23__and_module_3_res) );
  OR2_X1 u_majority7_module_23__or_module_3_U1 ( .A1(n_majority7_module_23_n1), 
        .A2(n_majority7_module_23_n6), .ZN(
        n_majority7_module_23__or_module_3_res) );
  AND2_X1 u_majority7_module_23__and_module_4_U1 ( .A1(
        n_majority7_module_23__and_module_2_res), .A2(
        n_majority7_module_23__and_module_1_res), .ZN(
        n_majority7_module_23__and_module_4_res) );
  OR2_X1 u_majority7_module_23__or_module_4_U1 ( .A1(
        n_majority7_module_23__and_module_1_res), .A2(
        n_majority7_module_23__and_module_2_res), .ZN(
        n_majority7_module_23__or_module_4_res) );
  AND2_X1 u_majority7_module_23__and_module_5_U1 ( .A1(
        n_majority7_module_23__and_module_3_res), .A2(n_majority7_module_23_n3), .ZN(n_majority7_module_23__and_module_5_res) );
  OR2_X1 u_majority7_module_23__or_module_5_U1 ( .A1(n_majority7_module_23_n3), 
        .A2(n_majority7_module_23__and_module_3_res), .ZN(
        n_majority7_module_23__or_module_5_res) );
  AND2_X1 u_majority7_module_23__and_module_6_U1 ( .A1(
        n_majority7_module_23__or_module_1_res), .A2(
        n_majority7_module_23__or_module_2_res), .ZN(
        n_majority7_module_23__and_module_6_res) );
  OR2_X1 u_majority7_module_23__or_module_6_U1 ( .A1(
        n_majority7_module_23__or_module_2_res), .A2(
        n_majority7_module_23__or_module_1_res), .ZN(
        n_majority7_module_23__or_module_6_res) );
  OR2_X1 u_majority7_module_23__or_module_7_U1 ( .A1(
        n_majority7_module_23__and_module_4_res), .A2(
        n_majority7_module_23__and_module_5_res), .ZN(
        n_majority7_module_23__or_module_7_res) );
  AND2_X1 u_majority7_module_23__and_module_7_U1 ( .A1(
        n_majority7_module_23__or_module_3_res), .A2(
        n_majority7_module_23__or_module_4_res), .ZN(
        n_majority7_module_23__and_module_7_res) );
  OR2_X1 u_majority7_module_23__or_module_8_U1 ( .A1(
        n_majority7_module_23__or_module_4_res), .A2(
        n_majority7_module_23__or_module_3_res), .ZN(
        n_majority7_module_23__or_module_8_res) );
  AND2_X1 u_majority7_module_23__and_module_8_U1 ( .A1(
        n_majority7_module_23__or_module_5_res), .A2(
        n_majority7_module_23__and_module_6_res), .ZN(
        n_majority7_module_23__and_module_8_res) );
  OR2_X1 u_majority7_module_23__or_module_9_U1 ( .A1(
        n_majority7_module_23__and_module_6_res), .A2(
        n_majority7_module_23__or_module_5_res), .ZN(
        n_majority7_module_23__or_module_9_res) );
  OR2_X1 u_majority7_module_23__or_module_10_U1 ( .A1(
        n_majority7_module_23__or_module_7_res), .A2(
        n_majority7_module_23__and_module_7_res), .ZN(
        n_majority7_module_23__or_module_10_res) );
  AND2_X1 u_majority7_module_23__and_module_9_U1 ( .A1(
        n_majority7_module_23__or_module_6_res), .A2(
        n_majority7_module_23__or_module_9_res), .ZN(
        n_majority7_module_23__and_module_9_res) );
  OR2_X1 u_majority7_module_23__or_module_11_U1 ( .A1(
        n_majority7_module_23__or_module_10_res), .A2(
        n_majority7_module_23__and_module_8_res), .ZN(
        n_majority7_module_23__or_module_11_res) );
  AND2_X1 u_majority7_module_23__and_module_10_U1 ( .A1(
        n_majority7_module_23__or_module_8_res), .A2(
        n_majority7_module_23__and_module_9_res), .ZN(
        n_majority7_module_23__and_module_10_res) );
  AND2_X1 u_majority7_module_23__and_module_11_U1 ( .A1(
        n_majority7_module_23__and_module_10_res), .A2(
        n_majority7_module_23__or_module_11_res), .ZN(
        n_majority7_module_23_res) );
  DFF_X1 u_reg_module_24__cini_mul_v000_reg ( .D(n_majority7_module_23_res), 
        .CK(clock_1), .Q(n_reg_module_24_res), .QN() );
  BUF_X1 u_majority7_module_24_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_24_n7) );
  BUF_X1 u_majority7_module_24_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_24_n6) );
  BUF_X1 u_majority7_module_24_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_24_n5) );
  BUF_X1 u_majority7_module_24_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_24_n4) );
  BUF_X1 u_majority7_module_24_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_24_n3) );
  BUF_X1 u_majority7_module_24_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_24_n2) );
  BUF_X1 u_majority7_module_24_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_24_n1) );
  AND2_X1 u_majority7_module_24__and_module_1_U1 ( .A1(
        n_majority7_module_24_n5), .A2(n_majority7_module_24_n4), .ZN(
        n_majority7_module_24__and_module_1_res) );
  OR2_X1 u_majority7_module_24__or_module_1_U1 ( .A1(n_majority7_module_24_n4), 
        .A2(n_majority7_module_24_n5), .ZN(
        n_majority7_module_24__or_module_1_res) );
  AND2_X1 u_majority7_module_24__and_module_2_U1 ( .A1(
        n_majority7_module_24_n7), .A2(n_majority7_module_24_n2), .ZN(
        n_majority7_module_24__and_module_2_res) );
  OR2_X1 u_majority7_module_24__or_module_2_U1 ( .A1(n_majority7_module_24_n2), 
        .A2(n_majority7_module_24_n7), .ZN(
        n_majority7_module_24__or_module_2_res) );
  AND2_X1 u_majority7_module_24__and_module_3_U1 ( .A1(
        n_majority7_module_24_n6), .A2(n_majority7_module_24_n1), .ZN(
        n_majority7_module_24__and_module_3_res) );
  OR2_X1 u_majority7_module_24__or_module_3_U1 ( .A1(n_majority7_module_24_n1), 
        .A2(n_majority7_module_24_n6), .ZN(
        n_majority7_module_24__or_module_3_res) );
  AND2_X1 u_majority7_module_24__and_module_4_U1 ( .A1(
        n_majority7_module_24__and_module_2_res), .A2(
        n_majority7_module_24__and_module_1_res), .ZN(
        n_majority7_module_24__and_module_4_res) );
  OR2_X1 u_majority7_module_24__or_module_4_U1 ( .A1(
        n_majority7_module_24__and_module_1_res), .A2(
        n_majority7_module_24__and_module_2_res), .ZN(
        n_majority7_module_24__or_module_4_res) );
  AND2_X1 u_majority7_module_24__and_module_5_U1 ( .A1(
        n_majority7_module_24__and_module_3_res), .A2(n_majority7_module_24_n3), .ZN(n_majority7_module_24__and_module_5_res) );
  OR2_X1 u_majority7_module_24__or_module_5_U1 ( .A1(n_majority7_module_24_n3), 
        .A2(n_majority7_module_24__and_module_3_res), .ZN(
        n_majority7_module_24__or_module_5_res) );
  AND2_X1 u_majority7_module_24__and_module_6_U1 ( .A1(
        n_majority7_module_24__or_module_1_res), .A2(
        n_majority7_module_24__or_module_2_res), .ZN(
        n_majority7_module_24__and_module_6_res) );
  OR2_X1 u_majority7_module_24__or_module_6_U1 ( .A1(
        n_majority7_module_24__or_module_2_res), .A2(
        n_majority7_module_24__or_module_1_res), .ZN(
        n_majority7_module_24__or_module_6_res) );
  OR2_X1 u_majority7_module_24__or_module_7_U1 ( .A1(
        n_majority7_module_24__and_module_4_res), .A2(
        n_majority7_module_24__and_module_5_res), .ZN(
        n_majority7_module_24__or_module_7_res) );
  AND2_X1 u_majority7_module_24__and_module_7_U1 ( .A1(
        n_majority7_module_24__or_module_3_res), .A2(
        n_majority7_module_24__or_module_4_res), .ZN(
        n_majority7_module_24__and_module_7_res) );
  OR2_X1 u_majority7_module_24__or_module_8_U1 ( .A1(
        n_majority7_module_24__or_module_4_res), .A2(
        n_majority7_module_24__or_module_3_res), .ZN(
        n_majority7_module_24__or_module_8_res) );
  AND2_X1 u_majority7_module_24__and_module_8_U1 ( .A1(
        n_majority7_module_24__or_module_5_res), .A2(
        n_majority7_module_24__and_module_6_res), .ZN(
        n_majority7_module_24__and_module_8_res) );
  OR2_X1 u_majority7_module_24__or_module_9_U1 ( .A1(
        n_majority7_module_24__and_module_6_res), .A2(
        n_majority7_module_24__or_module_5_res), .ZN(
        n_majority7_module_24__or_module_9_res) );
  OR2_X1 u_majority7_module_24__or_module_10_U1 ( .A1(
        n_majority7_module_24__or_module_7_res), .A2(
        n_majority7_module_24__and_module_7_res), .ZN(
        n_majority7_module_24__or_module_10_res) );
  AND2_X1 u_majority7_module_24__and_module_9_U1 ( .A1(
        n_majority7_module_24__or_module_6_res), .A2(
        n_majority7_module_24__or_module_9_res), .ZN(
        n_majority7_module_24__and_module_9_res) );
  OR2_X1 u_majority7_module_24__or_module_11_U1 ( .A1(
        n_majority7_module_24__or_module_10_res), .A2(
        n_majority7_module_24__and_module_8_res), .ZN(
        n_majority7_module_24__or_module_11_res) );
  AND2_X1 u_majority7_module_24__and_module_10_U1 ( .A1(
        n_majority7_module_24__or_module_8_res), .A2(
        n_majority7_module_24__and_module_9_res), .ZN(
        n_majority7_module_24__and_module_10_res) );
  AND2_X1 u_majority7_module_24__and_module_11_U1 ( .A1(
        n_majority7_module_24__and_module_10_res), .A2(
        n_majority7_module_24__or_module_11_res), .ZN(
        n_majority7_module_24_res) );
  DFF_X1 u_reg_module_25__cini_mul_v000_reg ( .D(n_majority7_module_24_res), 
        .CK(clock_1), .Q(n_reg_module_25_res), .QN() );
  BUF_X1 u_majority7_module_25_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_25_n7) );
  BUF_X1 u_majority7_module_25_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_25_n6) );
  BUF_X1 u_majority7_module_25_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_25_n5) );
  BUF_X1 u_majority7_module_25_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_25_n4) );
  BUF_X1 u_majority7_module_25_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_25_n3) );
  BUF_X1 u_majority7_module_25_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_25_n2) );
  BUF_X1 u_majority7_module_25_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_25_n1) );
  AND2_X1 u_majority7_module_25__and_module_1_U1 ( .A1(
        n_majority7_module_25_n5), .A2(n_majority7_module_25_n4), .ZN(
        n_majority7_module_25__and_module_1_res) );
  OR2_X1 u_majority7_module_25__or_module_1_U1 ( .A1(n_majority7_module_25_n4), 
        .A2(n_majority7_module_25_n5), .ZN(
        n_majority7_module_25__or_module_1_res) );
  AND2_X1 u_majority7_module_25__and_module_2_U1 ( .A1(
        n_majority7_module_25_n7), .A2(n_majority7_module_25_n2), .ZN(
        n_majority7_module_25__and_module_2_res) );
  OR2_X1 u_majority7_module_25__or_module_2_U1 ( .A1(n_majority7_module_25_n2), 
        .A2(n_majority7_module_25_n7), .ZN(
        n_majority7_module_25__or_module_2_res) );
  AND2_X1 u_majority7_module_25__and_module_3_U1 ( .A1(
        n_majority7_module_25_n6), .A2(n_majority7_module_25_n1), .ZN(
        n_majority7_module_25__and_module_3_res) );
  OR2_X1 u_majority7_module_25__or_module_3_U1 ( .A1(n_majority7_module_25_n1), 
        .A2(n_majority7_module_25_n6), .ZN(
        n_majority7_module_25__or_module_3_res) );
  AND2_X1 u_majority7_module_25__and_module_4_U1 ( .A1(
        n_majority7_module_25__and_module_2_res), .A2(
        n_majority7_module_25__and_module_1_res), .ZN(
        n_majority7_module_25__and_module_4_res) );
  OR2_X1 u_majority7_module_25__or_module_4_U1 ( .A1(
        n_majority7_module_25__and_module_1_res), .A2(
        n_majority7_module_25__and_module_2_res), .ZN(
        n_majority7_module_25__or_module_4_res) );
  AND2_X1 u_majority7_module_25__and_module_5_U1 ( .A1(
        n_majority7_module_25__and_module_3_res), .A2(n_majority7_module_25_n3), .ZN(n_majority7_module_25__and_module_5_res) );
  OR2_X1 u_majority7_module_25__or_module_5_U1 ( .A1(n_majority7_module_25_n3), 
        .A2(n_majority7_module_25__and_module_3_res), .ZN(
        n_majority7_module_25__or_module_5_res) );
  AND2_X1 u_majority7_module_25__and_module_6_U1 ( .A1(
        n_majority7_module_25__or_module_1_res), .A2(
        n_majority7_module_25__or_module_2_res), .ZN(
        n_majority7_module_25__and_module_6_res) );
  OR2_X1 u_majority7_module_25__or_module_6_U1 ( .A1(
        n_majority7_module_25__or_module_2_res), .A2(
        n_majority7_module_25__or_module_1_res), .ZN(
        n_majority7_module_25__or_module_6_res) );
  OR2_X1 u_majority7_module_25__or_module_7_U1 ( .A1(
        n_majority7_module_25__and_module_4_res), .A2(
        n_majority7_module_25__and_module_5_res), .ZN(
        n_majority7_module_25__or_module_7_res) );
  AND2_X1 u_majority7_module_25__and_module_7_U1 ( .A1(
        n_majority7_module_25__or_module_3_res), .A2(
        n_majority7_module_25__or_module_4_res), .ZN(
        n_majority7_module_25__and_module_7_res) );
  OR2_X1 u_majority7_module_25__or_module_8_U1 ( .A1(
        n_majority7_module_25__or_module_4_res), .A2(
        n_majority7_module_25__or_module_3_res), .ZN(
        n_majority7_module_25__or_module_8_res) );
  AND2_X1 u_majority7_module_25__and_module_8_U1 ( .A1(
        n_majority7_module_25__or_module_5_res), .A2(
        n_majority7_module_25__and_module_6_res), .ZN(
        n_majority7_module_25__and_module_8_res) );
  OR2_X1 u_majority7_module_25__or_module_9_U1 ( .A1(
        n_majority7_module_25__and_module_6_res), .A2(
        n_majority7_module_25__or_module_5_res), .ZN(
        n_majority7_module_25__or_module_9_res) );
  OR2_X1 u_majority7_module_25__or_module_10_U1 ( .A1(
        n_majority7_module_25__or_module_7_res), .A2(
        n_majority7_module_25__and_module_7_res), .ZN(
        n_majority7_module_25__or_module_10_res) );
  AND2_X1 u_majority7_module_25__and_module_9_U1 ( .A1(
        n_majority7_module_25__or_module_6_res), .A2(
        n_majority7_module_25__or_module_9_res), .ZN(
        n_majority7_module_25__and_module_9_res) );
  OR2_X1 u_majority7_module_25__or_module_11_U1 ( .A1(
        n_majority7_module_25__or_module_10_res), .A2(
        n_majority7_module_25__and_module_8_res), .ZN(
        n_majority7_module_25__or_module_11_res) );
  AND2_X1 u_majority7_module_25__and_module_10_U1 ( .A1(
        n_majority7_module_25__or_module_8_res), .A2(
        n_majority7_module_25__and_module_9_res), .ZN(
        n_majority7_module_25__and_module_10_res) );
  AND2_X1 u_majority7_module_25__and_module_11_U1 ( .A1(
        n_majority7_module_25__and_module_10_res), .A2(
        n_majority7_module_25__or_module_11_res), .ZN(
        n_majority7_module_25_res) );
  DFF_X1 u_reg_module_26__cini_mul_v000_reg ( .D(n_majority7_module_25_res), 
        .CK(clock_1), .Q(n_reg_module_26_res), .QN() );
  BUF_X1 u_majority7_module_26_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_26_n7) );
  BUF_X1 u_majority7_module_26_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_26_n6) );
  BUF_X1 u_majority7_module_26_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_26_n5) );
  BUF_X1 u_majority7_module_26_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_26_n4) );
  BUF_X1 u_majority7_module_26_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_26_n3) );
  BUF_X1 u_majority7_module_26_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_26_n2) );
  BUF_X1 u_majority7_module_26_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_26_n1) );
  AND2_X1 u_majority7_module_26__and_module_1_U1 ( .A1(
        n_majority7_module_26_n5), .A2(n_majority7_module_26_n4), .ZN(
        n_majority7_module_26__and_module_1_res) );
  OR2_X1 u_majority7_module_26__or_module_1_U1 ( .A1(n_majority7_module_26_n4), 
        .A2(n_majority7_module_26_n5), .ZN(
        n_majority7_module_26__or_module_1_res) );
  AND2_X1 u_majority7_module_26__and_module_2_U1 ( .A1(
        n_majority7_module_26_n7), .A2(n_majority7_module_26_n2), .ZN(
        n_majority7_module_26__and_module_2_res) );
  OR2_X1 u_majority7_module_26__or_module_2_U1 ( .A1(n_majority7_module_26_n2), 
        .A2(n_majority7_module_26_n7), .ZN(
        n_majority7_module_26__or_module_2_res) );
  AND2_X1 u_majority7_module_26__and_module_3_U1 ( .A1(
        n_majority7_module_26_n6), .A2(n_majority7_module_26_n1), .ZN(
        n_majority7_module_26__and_module_3_res) );
  OR2_X1 u_majority7_module_26__or_module_3_U1 ( .A1(n_majority7_module_26_n1), 
        .A2(n_majority7_module_26_n6), .ZN(
        n_majority7_module_26__or_module_3_res) );
  AND2_X1 u_majority7_module_26__and_module_4_U1 ( .A1(
        n_majority7_module_26__and_module_2_res), .A2(
        n_majority7_module_26__and_module_1_res), .ZN(
        n_majority7_module_26__and_module_4_res) );
  OR2_X1 u_majority7_module_26__or_module_4_U1 ( .A1(
        n_majority7_module_26__and_module_1_res), .A2(
        n_majority7_module_26__and_module_2_res), .ZN(
        n_majority7_module_26__or_module_4_res) );
  AND2_X1 u_majority7_module_26__and_module_5_U1 ( .A1(
        n_majority7_module_26__and_module_3_res), .A2(n_majority7_module_26_n3), .ZN(n_majority7_module_26__and_module_5_res) );
  OR2_X1 u_majority7_module_26__or_module_5_U1 ( .A1(n_majority7_module_26_n3), 
        .A2(n_majority7_module_26__and_module_3_res), .ZN(
        n_majority7_module_26__or_module_5_res) );
  AND2_X1 u_majority7_module_26__and_module_6_U1 ( .A1(
        n_majority7_module_26__or_module_1_res), .A2(
        n_majority7_module_26__or_module_2_res), .ZN(
        n_majority7_module_26__and_module_6_res) );
  OR2_X1 u_majority7_module_26__or_module_6_U1 ( .A1(
        n_majority7_module_26__or_module_2_res), .A2(
        n_majority7_module_26__or_module_1_res), .ZN(
        n_majority7_module_26__or_module_6_res) );
  OR2_X1 u_majority7_module_26__or_module_7_U1 ( .A1(
        n_majority7_module_26__and_module_4_res), .A2(
        n_majority7_module_26__and_module_5_res), .ZN(
        n_majority7_module_26__or_module_7_res) );
  AND2_X1 u_majority7_module_26__and_module_7_U1 ( .A1(
        n_majority7_module_26__or_module_3_res), .A2(
        n_majority7_module_26__or_module_4_res), .ZN(
        n_majority7_module_26__and_module_7_res) );
  OR2_X1 u_majority7_module_26__or_module_8_U1 ( .A1(
        n_majority7_module_26__or_module_4_res), .A2(
        n_majority7_module_26__or_module_3_res), .ZN(
        n_majority7_module_26__or_module_8_res) );
  AND2_X1 u_majority7_module_26__and_module_8_U1 ( .A1(
        n_majority7_module_26__or_module_5_res), .A2(
        n_majority7_module_26__and_module_6_res), .ZN(
        n_majority7_module_26__and_module_8_res) );
  OR2_X1 u_majority7_module_26__or_module_9_U1 ( .A1(
        n_majority7_module_26__and_module_6_res), .A2(
        n_majority7_module_26__or_module_5_res), .ZN(
        n_majority7_module_26__or_module_9_res) );
  OR2_X1 u_majority7_module_26__or_module_10_U1 ( .A1(
        n_majority7_module_26__or_module_7_res), .A2(
        n_majority7_module_26__and_module_7_res), .ZN(
        n_majority7_module_26__or_module_10_res) );
  AND2_X1 u_majority7_module_26__and_module_9_U1 ( .A1(
        n_majority7_module_26__or_module_6_res), .A2(
        n_majority7_module_26__or_module_9_res), .ZN(
        n_majority7_module_26__and_module_9_res) );
  OR2_X1 u_majority7_module_26__or_module_11_U1 ( .A1(
        n_majority7_module_26__or_module_10_res), .A2(
        n_majority7_module_26__and_module_8_res), .ZN(
        n_majority7_module_26__or_module_11_res) );
  AND2_X1 u_majority7_module_26__and_module_10_U1 ( .A1(
        n_majority7_module_26__or_module_8_res), .A2(
        n_majority7_module_26__and_module_9_res), .ZN(
        n_majority7_module_26__and_module_10_res) );
  AND2_X1 u_majority7_module_26__and_module_11_U1 ( .A1(
        n_majority7_module_26__and_module_10_res), .A2(
        n_majority7_module_26__or_module_11_res), .ZN(
        n_majority7_module_26_res) );
  DFF_X1 u_reg_module_27__cini_mul_v000_reg ( .D(n_majority7_module_26_res), 
        .CK(clock_1), .Q(n_reg_module_27_res), .QN() );
  BUF_X1 u_majority7_module_27_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_27_n7) );
  BUF_X1 u_majority7_module_27_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_27_n6) );
  BUF_X1 u_majority7_module_27_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_27_n5) );
  BUF_X1 u_majority7_module_27_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_27_n4) );
  BUF_X1 u_majority7_module_27_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_27_n3) );
  BUF_X1 u_majority7_module_27_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_27_n2) );
  BUF_X1 u_majority7_module_27_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_27_n1) );
  AND2_X1 u_majority7_module_27__and_module_1_U1 ( .A1(
        n_majority7_module_27_n5), .A2(n_majority7_module_27_n4), .ZN(
        n_majority7_module_27__and_module_1_res) );
  OR2_X1 u_majority7_module_27__or_module_1_U1 ( .A1(n_majority7_module_27_n4), 
        .A2(n_majority7_module_27_n5), .ZN(
        n_majority7_module_27__or_module_1_res) );
  AND2_X1 u_majority7_module_27__and_module_2_U1 ( .A1(
        n_majority7_module_27_n7), .A2(n_majority7_module_27_n2), .ZN(
        n_majority7_module_27__and_module_2_res) );
  OR2_X1 u_majority7_module_27__or_module_2_U1 ( .A1(n_majority7_module_27_n2), 
        .A2(n_majority7_module_27_n7), .ZN(
        n_majority7_module_27__or_module_2_res) );
  AND2_X1 u_majority7_module_27__and_module_3_U1 ( .A1(
        n_majority7_module_27_n6), .A2(n_majority7_module_27_n1), .ZN(
        n_majority7_module_27__and_module_3_res) );
  OR2_X1 u_majority7_module_27__or_module_3_U1 ( .A1(n_majority7_module_27_n1), 
        .A2(n_majority7_module_27_n6), .ZN(
        n_majority7_module_27__or_module_3_res) );
  AND2_X1 u_majority7_module_27__and_module_4_U1 ( .A1(
        n_majority7_module_27__and_module_2_res), .A2(
        n_majority7_module_27__and_module_1_res), .ZN(
        n_majority7_module_27__and_module_4_res) );
  OR2_X1 u_majority7_module_27__or_module_4_U1 ( .A1(
        n_majority7_module_27__and_module_1_res), .A2(
        n_majority7_module_27__and_module_2_res), .ZN(
        n_majority7_module_27__or_module_4_res) );
  AND2_X1 u_majority7_module_27__and_module_5_U1 ( .A1(
        n_majority7_module_27__and_module_3_res), .A2(n_majority7_module_27_n3), .ZN(n_majority7_module_27__and_module_5_res) );
  OR2_X1 u_majority7_module_27__or_module_5_U1 ( .A1(n_majority7_module_27_n3), 
        .A2(n_majority7_module_27__and_module_3_res), .ZN(
        n_majority7_module_27__or_module_5_res) );
  AND2_X1 u_majority7_module_27__and_module_6_U1 ( .A1(
        n_majority7_module_27__or_module_1_res), .A2(
        n_majority7_module_27__or_module_2_res), .ZN(
        n_majority7_module_27__and_module_6_res) );
  OR2_X1 u_majority7_module_27__or_module_6_U1 ( .A1(
        n_majority7_module_27__or_module_2_res), .A2(
        n_majority7_module_27__or_module_1_res), .ZN(
        n_majority7_module_27__or_module_6_res) );
  OR2_X1 u_majority7_module_27__or_module_7_U1 ( .A1(
        n_majority7_module_27__and_module_4_res), .A2(
        n_majority7_module_27__and_module_5_res), .ZN(
        n_majority7_module_27__or_module_7_res) );
  AND2_X1 u_majority7_module_27__and_module_7_U1 ( .A1(
        n_majority7_module_27__or_module_3_res), .A2(
        n_majority7_module_27__or_module_4_res), .ZN(
        n_majority7_module_27__and_module_7_res) );
  OR2_X1 u_majority7_module_27__or_module_8_U1 ( .A1(
        n_majority7_module_27__or_module_4_res), .A2(
        n_majority7_module_27__or_module_3_res), .ZN(
        n_majority7_module_27__or_module_8_res) );
  AND2_X1 u_majority7_module_27__and_module_8_U1 ( .A1(
        n_majority7_module_27__or_module_5_res), .A2(
        n_majority7_module_27__and_module_6_res), .ZN(
        n_majority7_module_27__and_module_8_res) );
  OR2_X1 u_majority7_module_27__or_module_9_U1 ( .A1(
        n_majority7_module_27__and_module_6_res), .A2(
        n_majority7_module_27__or_module_5_res), .ZN(
        n_majority7_module_27__or_module_9_res) );
  OR2_X1 u_majority7_module_27__or_module_10_U1 ( .A1(
        n_majority7_module_27__or_module_7_res), .A2(
        n_majority7_module_27__and_module_7_res), .ZN(
        n_majority7_module_27__or_module_10_res) );
  AND2_X1 u_majority7_module_27__and_module_9_U1 ( .A1(
        n_majority7_module_27__or_module_6_res), .A2(
        n_majority7_module_27__or_module_9_res), .ZN(
        n_majority7_module_27__and_module_9_res) );
  OR2_X1 u_majority7_module_27__or_module_11_U1 ( .A1(
        n_majority7_module_27__or_module_10_res), .A2(
        n_majority7_module_27__and_module_8_res), .ZN(
        n_majority7_module_27__or_module_11_res) );
  AND2_X1 u_majority7_module_27__and_module_10_U1 ( .A1(
        n_majority7_module_27__or_module_8_res), .A2(
        n_majority7_module_27__and_module_9_res), .ZN(
        n_majority7_module_27__and_module_10_res) );
  AND2_X1 u_majority7_module_27__and_module_11_U1 ( .A1(
        n_majority7_module_27__and_module_10_res), .A2(
        n_majority7_module_27__or_module_11_res), .ZN(
        n_majority7_module_27_res) );
  DFF_X1 u_reg_module_28__cini_mul_v000_reg ( .D(n_majority7_module_27_res), 
        .CK(clock_1), .Q(n_reg_module_28_res), .QN() );
  BUF_X1 u_majority7_module_28_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_28_n7) );
  BUF_X1 u_majority7_module_28_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_28_n6) );
  BUF_X1 u_majority7_module_28_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_28_n5) );
  BUF_X1 u_majority7_module_28_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_28_n4) );
  BUF_X1 u_majority7_module_28_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_28_n3) );
  BUF_X1 u_majority7_module_28_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_28_n2) );
  BUF_X1 u_majority7_module_28_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_28_n1) );
  AND2_X1 u_majority7_module_28__and_module_1_U1 ( .A1(
        n_majority7_module_28_n1), .A2(n_majority7_module_28_n5), .ZN(
        n_majority7_module_28__and_module_1_res) );
  OR2_X1 u_majority7_module_28__or_module_1_U1 ( .A1(n_majority7_module_28_n5), 
        .A2(n_majority7_module_28_n1), .ZN(
        n_majority7_module_28__or_module_1_res) );
  AND2_X1 u_majority7_module_28__and_module_2_U1 ( .A1(
        n_majority7_module_28_n7), .A2(n_majority7_module_28_n3), .ZN(
        n_majority7_module_28__and_module_2_res) );
  OR2_X1 u_majority7_module_28__or_module_2_U1 ( .A1(n_majority7_module_28_n3), 
        .A2(n_majority7_module_28_n7), .ZN(
        n_majority7_module_28__or_module_2_res) );
  AND2_X1 u_majority7_module_28__and_module_3_U1 ( .A1(
        n_majority7_module_28_n6), .A2(n_majority7_module_28_n2), .ZN(
        n_majority7_module_28__and_module_3_res) );
  OR2_X1 u_majority7_module_28__or_module_3_U1 ( .A1(n_majority7_module_28_n2), 
        .A2(n_majority7_module_28_n6), .ZN(
        n_majority7_module_28__or_module_3_res) );
  AND2_X1 u_majority7_module_28__and_module_4_U1 ( .A1(
        n_majority7_module_28__and_module_2_res), .A2(
        n_majority7_module_28__and_module_1_res), .ZN(
        n_majority7_module_28__and_module_4_res) );
  OR2_X1 u_majority7_module_28__or_module_4_U1 ( .A1(
        n_majority7_module_28__and_module_1_res), .A2(
        n_majority7_module_28__and_module_2_res), .ZN(
        n_majority7_module_28__or_module_4_res) );
  AND2_X1 u_majority7_module_28__and_module_5_U1 ( .A1(
        n_majority7_module_28__and_module_3_res), .A2(n_majority7_module_28_n4), .ZN(n_majority7_module_28__and_module_5_res) );
  OR2_X1 u_majority7_module_28__or_module_5_U1 ( .A1(n_majority7_module_28_n4), 
        .A2(n_majority7_module_28__and_module_3_res), .ZN(
        n_majority7_module_28__or_module_5_res) );
  AND2_X1 u_majority7_module_28__and_module_6_U1 ( .A1(
        n_majority7_module_28__or_module_1_res), .A2(
        n_majority7_module_28__or_module_2_res), .ZN(
        n_majority7_module_28__and_module_6_res) );
  OR2_X1 u_majority7_module_28__or_module_6_U1 ( .A1(
        n_majority7_module_28__or_module_2_res), .A2(
        n_majority7_module_28__or_module_1_res), .ZN(
        n_majority7_module_28__or_module_6_res) );
  OR2_X1 u_majority7_module_28__or_module_7_U1 ( .A1(
        n_majority7_module_28__and_module_4_res), .A2(
        n_majority7_module_28__and_module_5_res), .ZN(
        n_majority7_module_28__or_module_7_res) );
  AND2_X1 u_majority7_module_28__and_module_7_U1 ( .A1(
        n_majority7_module_28__or_module_3_res), .A2(
        n_majority7_module_28__or_module_4_res), .ZN(
        n_majority7_module_28__and_module_7_res) );
  OR2_X1 u_majority7_module_28__or_module_8_U1 ( .A1(
        n_majority7_module_28__or_module_4_res), .A2(
        n_majority7_module_28__or_module_3_res), .ZN(
        n_majority7_module_28__or_module_8_res) );
  AND2_X1 u_majority7_module_28__and_module_8_U1 ( .A1(
        n_majority7_module_28__or_module_5_res), .A2(
        n_majority7_module_28__and_module_6_res), .ZN(
        n_majority7_module_28__and_module_8_res) );
  OR2_X1 u_majority7_module_28__or_module_9_U1 ( .A1(
        n_majority7_module_28__and_module_6_res), .A2(
        n_majority7_module_28__or_module_5_res), .ZN(
        n_majority7_module_28__or_module_9_res) );
  OR2_X1 u_majority7_module_28__or_module_10_U1 ( .A1(
        n_majority7_module_28__or_module_7_res), .A2(
        n_majority7_module_28__and_module_7_res), .ZN(
        n_majority7_module_28__or_module_10_res) );
  AND2_X1 u_majority7_module_28__and_module_9_U1 ( .A1(
        n_majority7_module_28__or_module_6_res), .A2(
        n_majority7_module_28__or_module_9_res), .ZN(
        n_majority7_module_28__and_module_9_res) );
  OR2_X1 u_majority7_module_28__or_module_11_U1 ( .A1(
        n_majority7_module_28__or_module_10_res), .A2(
        n_majority7_module_28__and_module_8_res), .ZN(
        n_majority7_module_28__or_module_11_res) );
  AND2_X1 u_majority7_module_28__and_module_10_U1 ( .A1(
        n_majority7_module_28__or_module_8_res), .A2(
        n_majority7_module_28__and_module_9_res), .ZN(
        n_majority7_module_28__and_module_10_res) );
  AND2_X1 u_majority7_module_28__and_module_11_U1 ( .A1(
        n_majority7_module_28__and_module_10_res), .A2(
        n_majority7_module_28__or_module_11_res), .ZN(
        n_majority7_module_28_res) );
  DFF_X1 u_reg_module_29__cini_mul_v000_reg ( .D(n_majority7_module_28_res), 
        .CK(clock_1), .Q(n_reg_module_29_res), .QN() );
  BUF_X1 u_majority7_module_29_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_29_n7) );
  BUF_X1 u_majority7_module_29_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_29_n6) );
  BUF_X1 u_majority7_module_29_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_29_n5) );
  BUF_X1 u_majority7_module_29_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_29_n4) );
  BUF_X1 u_majority7_module_29_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_29_n3) );
  BUF_X1 u_majority7_module_29_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_29_n2) );
  BUF_X1 u_majority7_module_29_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_29_n1) );
  AND2_X1 u_majority7_module_29__and_module_1_U1 ( .A1(
        n_majority7_module_29_n1), .A2(n_majority7_module_29_n5), .ZN(
        n_majority7_module_29__and_module_1_res) );
  OR2_X1 u_majority7_module_29__or_module_1_U1 ( .A1(n_majority7_module_29_n5), 
        .A2(n_majority7_module_29_n1), .ZN(
        n_majority7_module_29__or_module_1_res) );
  AND2_X1 u_majority7_module_29__and_module_2_U1 ( .A1(
        n_majority7_module_29_n7), .A2(n_majority7_module_29_n3), .ZN(
        n_majority7_module_29__and_module_2_res) );
  OR2_X1 u_majority7_module_29__or_module_2_U1 ( .A1(n_majority7_module_29_n3), 
        .A2(n_majority7_module_29_n7), .ZN(
        n_majority7_module_29__or_module_2_res) );
  AND2_X1 u_majority7_module_29__and_module_3_U1 ( .A1(
        n_majority7_module_29_n6), .A2(n_majority7_module_29_n2), .ZN(
        n_majority7_module_29__and_module_3_res) );
  OR2_X1 u_majority7_module_29__or_module_3_U1 ( .A1(n_majority7_module_29_n2), 
        .A2(n_majority7_module_29_n6), .ZN(
        n_majority7_module_29__or_module_3_res) );
  AND2_X1 u_majority7_module_29__and_module_4_U1 ( .A1(
        n_majority7_module_29__and_module_2_res), .A2(
        n_majority7_module_29__and_module_1_res), .ZN(
        n_majority7_module_29__and_module_4_res) );
  OR2_X1 u_majority7_module_29__or_module_4_U1 ( .A1(
        n_majority7_module_29__and_module_1_res), .A2(
        n_majority7_module_29__and_module_2_res), .ZN(
        n_majority7_module_29__or_module_4_res) );
  AND2_X1 u_majority7_module_29__and_module_5_U1 ( .A1(
        n_majority7_module_29__and_module_3_res), .A2(n_majority7_module_29_n4), .ZN(n_majority7_module_29__and_module_5_res) );
  OR2_X1 u_majority7_module_29__or_module_5_U1 ( .A1(n_majority7_module_29_n4), 
        .A2(n_majority7_module_29__and_module_3_res), .ZN(
        n_majority7_module_29__or_module_5_res) );
  AND2_X1 u_majority7_module_29__and_module_6_U1 ( .A1(
        n_majority7_module_29__or_module_1_res), .A2(
        n_majority7_module_29__or_module_2_res), .ZN(
        n_majority7_module_29__and_module_6_res) );
  OR2_X1 u_majority7_module_29__or_module_6_U1 ( .A1(
        n_majority7_module_29__or_module_2_res), .A2(
        n_majority7_module_29__or_module_1_res), .ZN(
        n_majority7_module_29__or_module_6_res) );
  OR2_X1 u_majority7_module_29__or_module_7_U1 ( .A1(
        n_majority7_module_29__and_module_4_res), .A2(
        n_majority7_module_29__and_module_5_res), .ZN(
        n_majority7_module_29__or_module_7_res) );
  AND2_X1 u_majority7_module_29__and_module_7_U1 ( .A1(
        n_majority7_module_29__or_module_3_res), .A2(
        n_majority7_module_29__or_module_4_res), .ZN(
        n_majority7_module_29__and_module_7_res) );
  OR2_X1 u_majority7_module_29__or_module_8_U1 ( .A1(
        n_majority7_module_29__or_module_4_res), .A2(
        n_majority7_module_29__or_module_3_res), .ZN(
        n_majority7_module_29__or_module_8_res) );
  AND2_X1 u_majority7_module_29__and_module_8_U1 ( .A1(
        n_majority7_module_29__or_module_5_res), .A2(
        n_majority7_module_29__and_module_6_res), .ZN(
        n_majority7_module_29__and_module_8_res) );
  OR2_X1 u_majority7_module_29__or_module_9_U1 ( .A1(
        n_majority7_module_29__and_module_6_res), .A2(
        n_majority7_module_29__or_module_5_res), .ZN(
        n_majority7_module_29__or_module_9_res) );
  OR2_X1 u_majority7_module_29__or_module_10_U1 ( .A1(
        n_majority7_module_29__or_module_7_res), .A2(
        n_majority7_module_29__and_module_7_res), .ZN(
        n_majority7_module_29__or_module_10_res) );
  AND2_X1 u_majority7_module_29__and_module_9_U1 ( .A1(
        n_majority7_module_29__or_module_6_res), .A2(
        n_majority7_module_29__or_module_9_res), .ZN(
        n_majority7_module_29__and_module_9_res) );
  OR2_X1 u_majority7_module_29__or_module_11_U1 ( .A1(
        n_majority7_module_29__or_module_10_res), .A2(
        n_majority7_module_29__and_module_8_res), .ZN(
        n_majority7_module_29__or_module_11_res) );
  AND2_X1 u_majority7_module_29__and_module_10_U1 ( .A1(
        n_majority7_module_29__or_module_8_res), .A2(
        n_majority7_module_29__and_module_9_res), .ZN(
        n_majority7_module_29__and_module_10_res) );
  AND2_X1 u_majority7_module_29__and_module_11_U1 ( .A1(
        n_majority7_module_29__and_module_10_res), .A2(
        n_majority7_module_29__or_module_11_res), .ZN(
        n_majority7_module_29_res) );
  DFF_X1 u_reg_module_30__cini_mul_v000_reg ( .D(n_majority7_module_29_res), 
        .CK(clock_1), .Q(n_reg_module_30_res), .QN() );
  BUF_X1 u_majority7_module_30_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_30_n7) );
  BUF_X1 u_majority7_module_30_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_30_n6) );
  BUF_X1 u_majority7_module_30_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_30_n5) );
  BUF_X1 u_majority7_module_30_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_30_n4) );
  BUF_X1 u_majority7_module_30_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_30_n3) );
  BUF_X1 u_majority7_module_30_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_30_n2) );
  BUF_X1 u_majority7_module_30_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_30_n1) );
  AND2_X1 u_majority7_module_30__and_module_1_U1 ( .A1(
        n_majority7_module_30_n1), .A2(n_majority7_module_30_n5), .ZN(
        n_majority7_module_30__and_module_1_res) );
  OR2_X1 u_majority7_module_30__or_module_1_U1 ( .A1(n_majority7_module_30_n5), 
        .A2(n_majority7_module_30_n1), .ZN(
        n_majority7_module_30__or_module_1_res) );
  AND2_X1 u_majority7_module_30__and_module_2_U1 ( .A1(
        n_majority7_module_30_n7), .A2(n_majority7_module_30_n3), .ZN(
        n_majority7_module_30__and_module_2_res) );
  OR2_X1 u_majority7_module_30__or_module_2_U1 ( .A1(n_majority7_module_30_n3), 
        .A2(n_majority7_module_30_n7), .ZN(
        n_majority7_module_30__or_module_2_res) );
  AND2_X1 u_majority7_module_30__and_module_3_U1 ( .A1(
        n_majority7_module_30_n6), .A2(n_majority7_module_30_n2), .ZN(
        n_majority7_module_30__and_module_3_res) );
  OR2_X1 u_majority7_module_30__or_module_3_U1 ( .A1(n_majority7_module_30_n2), 
        .A2(n_majority7_module_30_n6), .ZN(
        n_majority7_module_30__or_module_3_res) );
  AND2_X1 u_majority7_module_30__and_module_4_U1 ( .A1(
        n_majority7_module_30__and_module_2_res), .A2(
        n_majority7_module_30__and_module_1_res), .ZN(
        n_majority7_module_30__and_module_4_res) );
  OR2_X1 u_majority7_module_30__or_module_4_U1 ( .A1(
        n_majority7_module_30__and_module_1_res), .A2(
        n_majority7_module_30__and_module_2_res), .ZN(
        n_majority7_module_30__or_module_4_res) );
  AND2_X1 u_majority7_module_30__and_module_5_U1 ( .A1(
        n_majority7_module_30__and_module_3_res), .A2(n_majority7_module_30_n4), .ZN(n_majority7_module_30__and_module_5_res) );
  OR2_X1 u_majority7_module_30__or_module_5_U1 ( .A1(n_majority7_module_30_n4), 
        .A2(n_majority7_module_30__and_module_3_res), .ZN(
        n_majority7_module_30__or_module_5_res) );
  AND2_X1 u_majority7_module_30__and_module_6_U1 ( .A1(
        n_majority7_module_30__or_module_1_res), .A2(
        n_majority7_module_30__or_module_2_res), .ZN(
        n_majority7_module_30__and_module_6_res) );
  OR2_X1 u_majority7_module_30__or_module_6_U1 ( .A1(
        n_majority7_module_30__or_module_2_res), .A2(
        n_majority7_module_30__or_module_1_res), .ZN(
        n_majority7_module_30__or_module_6_res) );
  OR2_X1 u_majority7_module_30__or_module_7_U1 ( .A1(
        n_majority7_module_30__and_module_4_res), .A2(
        n_majority7_module_30__and_module_5_res), .ZN(
        n_majority7_module_30__or_module_7_res) );
  AND2_X1 u_majority7_module_30__and_module_7_U1 ( .A1(
        n_majority7_module_30__or_module_3_res), .A2(
        n_majority7_module_30__or_module_4_res), .ZN(
        n_majority7_module_30__and_module_7_res) );
  OR2_X1 u_majority7_module_30__or_module_8_U1 ( .A1(
        n_majority7_module_30__or_module_4_res), .A2(
        n_majority7_module_30__or_module_3_res), .ZN(
        n_majority7_module_30__or_module_8_res) );
  AND2_X1 u_majority7_module_30__and_module_8_U1 ( .A1(
        n_majority7_module_30__or_module_5_res), .A2(
        n_majority7_module_30__and_module_6_res), .ZN(
        n_majority7_module_30__and_module_8_res) );
  OR2_X1 u_majority7_module_30__or_module_9_U1 ( .A1(
        n_majority7_module_30__and_module_6_res), .A2(
        n_majority7_module_30__or_module_5_res), .ZN(
        n_majority7_module_30__or_module_9_res) );
  OR2_X1 u_majority7_module_30__or_module_10_U1 ( .A1(
        n_majority7_module_30__or_module_7_res), .A2(
        n_majority7_module_30__and_module_7_res), .ZN(
        n_majority7_module_30__or_module_10_res) );
  AND2_X1 u_majority7_module_30__and_module_9_U1 ( .A1(
        n_majority7_module_30__or_module_6_res), .A2(
        n_majority7_module_30__or_module_9_res), .ZN(
        n_majority7_module_30__and_module_9_res) );
  OR2_X1 u_majority7_module_30__or_module_11_U1 ( .A1(
        n_majority7_module_30__or_module_10_res), .A2(
        n_majority7_module_30__and_module_8_res), .ZN(
        n_majority7_module_30__or_module_11_res) );
  AND2_X1 u_majority7_module_30__and_module_10_U1 ( .A1(
        n_majority7_module_30__or_module_8_res), .A2(
        n_majority7_module_30__and_module_9_res), .ZN(
        n_majority7_module_30__and_module_10_res) );
  AND2_X1 u_majority7_module_30__and_module_11_U1 ( .A1(
        n_majority7_module_30__and_module_10_res), .A2(
        n_majority7_module_30__or_module_11_res), .ZN(
        n_majority7_module_30_res) );
  DFF_X1 u_reg_module_31__cini_mul_v000_reg ( .D(n_majority7_module_30_res), 
        .CK(clock_1), .Q(n_reg_module_31_res), .QN() );
  BUF_X1 u_majority7_module_31_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_31_n7) );
  BUF_X1 u_majority7_module_31_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_31_n6) );
  BUF_X1 u_majority7_module_31_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_31_n5) );
  BUF_X1 u_majority7_module_31_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_31_n4) );
  BUF_X1 u_majority7_module_31_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_31_n3) );
  BUF_X1 u_majority7_module_31_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_31_n2) );
  BUF_X1 u_majority7_module_31_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_31_n1) );
  AND2_X1 u_majority7_module_31__and_module_1_U1 ( .A1(
        n_majority7_module_31_n1), .A2(n_majority7_module_31_n5), .ZN(
        n_majority7_module_31__and_module_1_res) );
  OR2_X1 u_majority7_module_31__or_module_1_U1 ( .A1(n_majority7_module_31_n5), 
        .A2(n_majority7_module_31_n1), .ZN(
        n_majority7_module_31__or_module_1_res) );
  AND2_X1 u_majority7_module_31__and_module_2_U1 ( .A1(
        n_majority7_module_31_n7), .A2(n_majority7_module_31_n3), .ZN(
        n_majority7_module_31__and_module_2_res) );
  OR2_X1 u_majority7_module_31__or_module_2_U1 ( .A1(n_majority7_module_31_n3), 
        .A2(n_majority7_module_31_n7), .ZN(
        n_majority7_module_31__or_module_2_res) );
  AND2_X1 u_majority7_module_31__and_module_3_U1 ( .A1(
        n_majority7_module_31_n6), .A2(n_majority7_module_31_n2), .ZN(
        n_majority7_module_31__and_module_3_res) );
  OR2_X1 u_majority7_module_31__or_module_3_U1 ( .A1(n_majority7_module_31_n2), 
        .A2(n_majority7_module_31_n6), .ZN(
        n_majority7_module_31__or_module_3_res) );
  AND2_X1 u_majority7_module_31__and_module_4_U1 ( .A1(
        n_majority7_module_31__and_module_2_res), .A2(
        n_majority7_module_31__and_module_1_res), .ZN(
        n_majority7_module_31__and_module_4_res) );
  OR2_X1 u_majority7_module_31__or_module_4_U1 ( .A1(
        n_majority7_module_31__and_module_1_res), .A2(
        n_majority7_module_31__and_module_2_res), .ZN(
        n_majority7_module_31__or_module_4_res) );
  AND2_X1 u_majority7_module_31__and_module_5_U1 ( .A1(
        n_majority7_module_31__and_module_3_res), .A2(n_majority7_module_31_n4), .ZN(n_majority7_module_31__and_module_5_res) );
  OR2_X1 u_majority7_module_31__or_module_5_U1 ( .A1(n_majority7_module_31_n4), 
        .A2(n_majority7_module_31__and_module_3_res), .ZN(
        n_majority7_module_31__or_module_5_res) );
  AND2_X1 u_majority7_module_31__and_module_6_U1 ( .A1(
        n_majority7_module_31__or_module_1_res), .A2(
        n_majority7_module_31__or_module_2_res), .ZN(
        n_majority7_module_31__and_module_6_res) );
  OR2_X1 u_majority7_module_31__or_module_6_U1 ( .A1(
        n_majority7_module_31__or_module_2_res), .A2(
        n_majority7_module_31__or_module_1_res), .ZN(
        n_majority7_module_31__or_module_6_res) );
  OR2_X1 u_majority7_module_31__or_module_7_U1 ( .A1(
        n_majority7_module_31__and_module_4_res), .A2(
        n_majority7_module_31__and_module_5_res), .ZN(
        n_majority7_module_31__or_module_7_res) );
  AND2_X1 u_majority7_module_31__and_module_7_U1 ( .A1(
        n_majority7_module_31__or_module_3_res), .A2(
        n_majority7_module_31__or_module_4_res), .ZN(
        n_majority7_module_31__and_module_7_res) );
  OR2_X1 u_majority7_module_31__or_module_8_U1 ( .A1(
        n_majority7_module_31__or_module_4_res), .A2(
        n_majority7_module_31__or_module_3_res), .ZN(
        n_majority7_module_31__or_module_8_res) );
  AND2_X1 u_majority7_module_31__and_module_8_U1 ( .A1(
        n_majority7_module_31__or_module_5_res), .A2(
        n_majority7_module_31__and_module_6_res), .ZN(
        n_majority7_module_31__and_module_8_res) );
  OR2_X1 u_majority7_module_31__or_module_9_U1 ( .A1(
        n_majority7_module_31__and_module_6_res), .A2(
        n_majority7_module_31__or_module_5_res), .ZN(
        n_majority7_module_31__or_module_9_res) );
  OR2_X1 u_majority7_module_31__or_module_10_U1 ( .A1(
        n_majority7_module_31__or_module_7_res), .A2(
        n_majority7_module_31__and_module_7_res), .ZN(
        n_majority7_module_31__or_module_10_res) );
  AND2_X1 u_majority7_module_31__and_module_9_U1 ( .A1(
        n_majority7_module_31__or_module_6_res), .A2(
        n_majority7_module_31__or_module_9_res), .ZN(
        n_majority7_module_31__and_module_9_res) );
  OR2_X1 u_majority7_module_31__or_module_11_U1 ( .A1(
        n_majority7_module_31__or_module_10_res), .A2(
        n_majority7_module_31__and_module_8_res), .ZN(
        n_majority7_module_31__or_module_11_res) );
  AND2_X1 u_majority7_module_31__and_module_10_U1 ( .A1(
        n_majority7_module_31__or_module_8_res), .A2(
        n_majority7_module_31__and_module_9_res), .ZN(
        n_majority7_module_31__and_module_10_res) );
  AND2_X1 u_majority7_module_31__and_module_11_U1 ( .A1(
        n_majority7_module_31__and_module_10_res), .A2(
        n_majority7_module_31__or_module_11_res), .ZN(
        n_majority7_module_31_res) );
  DFF_X1 u_reg_module_32__cini_mul_v000_reg ( .D(n_majority7_module_31_res), 
        .CK(clock_1), .Q(n_reg_module_32_res), .QN() );
  BUF_X1 u_majority7_module_32_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_32_n7) );
  BUF_X1 u_majority7_module_32_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_32_n6) );
  BUF_X1 u_majority7_module_32_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_32_n5) );
  BUF_X1 u_majority7_module_32_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_32_n4) );
  BUF_X1 u_majority7_module_32_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_32_n3) );
  BUF_X1 u_majority7_module_32_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_32_n2) );
  BUF_X1 u_majority7_module_32_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_32_n1) );
  AND2_X1 u_majority7_module_32__and_module_1_U1 ( .A1(
        n_majority7_module_32_n5), .A2(n_majority7_module_32_n4), .ZN(
        n_majority7_module_32__and_module_1_res) );
  OR2_X1 u_majority7_module_32__or_module_1_U1 ( .A1(n_majority7_module_32_n4), 
        .A2(n_majority7_module_32_n5), .ZN(
        n_majority7_module_32__or_module_1_res) );
  AND2_X1 u_majority7_module_32__and_module_2_U1 ( .A1(
        n_majority7_module_32_n7), .A2(n_majority7_module_32_n2), .ZN(
        n_majority7_module_32__and_module_2_res) );
  OR2_X1 u_majority7_module_32__or_module_2_U1 ( .A1(n_majority7_module_32_n2), 
        .A2(n_majority7_module_32_n7), .ZN(
        n_majority7_module_32__or_module_2_res) );
  AND2_X1 u_majority7_module_32__and_module_3_U1 ( .A1(
        n_majority7_module_32_n6), .A2(n_majority7_module_32_n1), .ZN(
        n_majority7_module_32__and_module_3_res) );
  OR2_X1 u_majority7_module_32__or_module_3_U1 ( .A1(n_majority7_module_32_n1), 
        .A2(n_majority7_module_32_n6), .ZN(
        n_majority7_module_32__or_module_3_res) );
  AND2_X1 u_majority7_module_32__and_module_4_U1 ( .A1(
        n_majority7_module_32__and_module_2_res), .A2(
        n_majority7_module_32__and_module_1_res), .ZN(
        n_majority7_module_32__and_module_4_res) );
  OR2_X1 u_majority7_module_32__or_module_4_U1 ( .A1(
        n_majority7_module_32__and_module_1_res), .A2(
        n_majority7_module_32__and_module_2_res), .ZN(
        n_majority7_module_32__or_module_4_res) );
  AND2_X1 u_majority7_module_32__and_module_5_U1 ( .A1(
        n_majority7_module_32__and_module_3_res), .A2(n_majority7_module_32_n3), .ZN(n_majority7_module_32__and_module_5_res) );
  OR2_X1 u_majority7_module_32__or_module_5_U1 ( .A1(n_majority7_module_32_n3), 
        .A2(n_majority7_module_32__and_module_3_res), .ZN(
        n_majority7_module_32__or_module_5_res) );
  AND2_X1 u_majority7_module_32__and_module_6_U1 ( .A1(
        n_majority7_module_32__or_module_1_res), .A2(
        n_majority7_module_32__or_module_2_res), .ZN(
        n_majority7_module_32__and_module_6_res) );
  OR2_X1 u_majority7_module_32__or_module_6_U1 ( .A1(
        n_majority7_module_32__or_module_2_res), .A2(
        n_majority7_module_32__or_module_1_res), .ZN(
        n_majority7_module_32__or_module_6_res) );
  OR2_X1 u_majority7_module_32__or_module_7_U1 ( .A1(
        n_majority7_module_32__and_module_4_res), .A2(
        n_majority7_module_32__and_module_5_res), .ZN(
        n_majority7_module_32__or_module_7_res) );
  AND2_X1 u_majority7_module_32__and_module_7_U1 ( .A1(
        n_majority7_module_32__or_module_3_res), .A2(
        n_majority7_module_32__or_module_4_res), .ZN(
        n_majority7_module_32__and_module_7_res) );
  OR2_X1 u_majority7_module_32__or_module_8_U1 ( .A1(
        n_majority7_module_32__or_module_4_res), .A2(
        n_majority7_module_32__or_module_3_res), .ZN(
        n_majority7_module_32__or_module_8_res) );
  AND2_X1 u_majority7_module_32__and_module_8_U1 ( .A1(
        n_majority7_module_32__or_module_5_res), .A2(
        n_majority7_module_32__and_module_6_res), .ZN(
        n_majority7_module_32__and_module_8_res) );
  OR2_X1 u_majority7_module_32__or_module_9_U1 ( .A1(
        n_majority7_module_32__and_module_6_res), .A2(
        n_majority7_module_32__or_module_5_res), .ZN(
        n_majority7_module_32__or_module_9_res) );
  OR2_X1 u_majority7_module_32__or_module_10_U1 ( .A1(
        n_majority7_module_32__or_module_7_res), .A2(
        n_majority7_module_32__and_module_7_res), .ZN(
        n_majority7_module_32__or_module_10_res) );
  AND2_X1 u_majority7_module_32__and_module_9_U1 ( .A1(
        n_majority7_module_32__or_module_6_res), .A2(
        n_majority7_module_32__or_module_9_res), .ZN(
        n_majority7_module_32__and_module_9_res) );
  OR2_X1 u_majority7_module_32__or_module_11_U1 ( .A1(
        n_majority7_module_32__or_module_10_res), .A2(
        n_majority7_module_32__and_module_8_res), .ZN(
        n_majority7_module_32__or_module_11_res) );
  AND2_X1 u_majority7_module_32__and_module_10_U1 ( .A1(
        n_majority7_module_32__or_module_8_res), .A2(
        n_majority7_module_32__and_module_9_res), .ZN(
        n_majority7_module_32__and_module_10_res) );
  AND2_X1 u_majority7_module_32__and_module_11_U1 ( .A1(
        n_majority7_module_32__and_module_10_res), .A2(
        n_majority7_module_32__or_module_11_res), .ZN(
        n_majority7_module_32_res) );
  DFF_X1 u_reg_module_33__cini_mul_v000_reg ( .D(n_majority7_module_32_res), 
        .CK(clock_2), .Q(n_reg_module_33_res), .QN() );
  BUF_X1 u_majority7_module_33_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_33_n7) );
  BUF_X1 u_majority7_module_33_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_33_n6) );
  BUF_X1 u_majority7_module_33_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_33_n5) );
  BUF_X1 u_majority7_module_33_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_33_n4) );
  BUF_X1 u_majority7_module_33_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_33_n3) );
  BUF_X1 u_majority7_module_33_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_33_n2) );
  BUF_X1 u_majority7_module_33_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_33_n1) );
  AND2_X1 u_majority7_module_33__and_module_1_U1 ( .A1(
        n_majority7_module_33_n5), .A2(n_majority7_module_33_n4), .ZN(
        n_majority7_module_33__and_module_1_res) );
  OR2_X1 u_majority7_module_33__or_module_1_U1 ( .A1(n_majority7_module_33_n4), 
        .A2(n_majority7_module_33_n5), .ZN(
        n_majority7_module_33__or_module_1_res) );
  AND2_X1 u_majority7_module_33__and_module_2_U1 ( .A1(
        n_majority7_module_33_n7), .A2(n_majority7_module_33_n2), .ZN(
        n_majority7_module_33__and_module_2_res) );
  OR2_X1 u_majority7_module_33__or_module_2_U1 ( .A1(n_majority7_module_33_n2), 
        .A2(n_majority7_module_33_n7), .ZN(
        n_majority7_module_33__or_module_2_res) );
  AND2_X1 u_majority7_module_33__and_module_3_U1 ( .A1(
        n_majority7_module_33_n6), .A2(n_majority7_module_33_n1), .ZN(
        n_majority7_module_33__and_module_3_res) );
  OR2_X1 u_majority7_module_33__or_module_3_U1 ( .A1(n_majority7_module_33_n1), 
        .A2(n_majority7_module_33_n6), .ZN(
        n_majority7_module_33__or_module_3_res) );
  AND2_X1 u_majority7_module_33__and_module_4_U1 ( .A1(
        n_majority7_module_33__and_module_2_res), .A2(
        n_majority7_module_33__and_module_1_res), .ZN(
        n_majority7_module_33__and_module_4_res) );
  OR2_X1 u_majority7_module_33__or_module_4_U1 ( .A1(
        n_majority7_module_33__and_module_1_res), .A2(
        n_majority7_module_33__and_module_2_res), .ZN(
        n_majority7_module_33__or_module_4_res) );
  AND2_X1 u_majority7_module_33__and_module_5_U1 ( .A1(
        n_majority7_module_33__and_module_3_res), .A2(n_majority7_module_33_n3), .ZN(n_majority7_module_33__and_module_5_res) );
  OR2_X1 u_majority7_module_33__or_module_5_U1 ( .A1(n_majority7_module_33_n3), 
        .A2(n_majority7_module_33__and_module_3_res), .ZN(
        n_majority7_module_33__or_module_5_res) );
  AND2_X1 u_majority7_module_33__and_module_6_U1 ( .A1(
        n_majority7_module_33__or_module_1_res), .A2(
        n_majority7_module_33__or_module_2_res), .ZN(
        n_majority7_module_33__and_module_6_res) );
  OR2_X1 u_majority7_module_33__or_module_6_U1 ( .A1(
        n_majority7_module_33__or_module_2_res), .A2(
        n_majority7_module_33__or_module_1_res), .ZN(
        n_majority7_module_33__or_module_6_res) );
  OR2_X1 u_majority7_module_33__or_module_7_U1 ( .A1(
        n_majority7_module_33__and_module_4_res), .A2(
        n_majority7_module_33__and_module_5_res), .ZN(
        n_majority7_module_33__or_module_7_res) );
  AND2_X1 u_majority7_module_33__and_module_7_U1 ( .A1(
        n_majority7_module_33__or_module_3_res), .A2(
        n_majority7_module_33__or_module_4_res), .ZN(
        n_majority7_module_33__and_module_7_res) );
  OR2_X1 u_majority7_module_33__or_module_8_U1 ( .A1(
        n_majority7_module_33__or_module_4_res), .A2(
        n_majority7_module_33__or_module_3_res), .ZN(
        n_majority7_module_33__or_module_8_res) );
  AND2_X1 u_majority7_module_33__and_module_8_U1 ( .A1(
        n_majority7_module_33__or_module_5_res), .A2(
        n_majority7_module_33__and_module_6_res), .ZN(
        n_majority7_module_33__and_module_8_res) );
  OR2_X1 u_majority7_module_33__or_module_9_U1 ( .A1(
        n_majority7_module_33__and_module_6_res), .A2(
        n_majority7_module_33__or_module_5_res), .ZN(
        n_majority7_module_33__or_module_9_res) );
  OR2_X1 u_majority7_module_33__or_module_10_U1 ( .A1(
        n_majority7_module_33__or_module_7_res), .A2(
        n_majority7_module_33__and_module_7_res), .ZN(
        n_majority7_module_33__or_module_10_res) );
  AND2_X1 u_majority7_module_33__and_module_9_U1 ( .A1(
        n_majority7_module_33__or_module_6_res), .A2(
        n_majority7_module_33__or_module_9_res), .ZN(
        n_majority7_module_33__and_module_9_res) );
  OR2_X1 u_majority7_module_33__or_module_11_U1 ( .A1(
        n_majority7_module_33__or_module_10_res), .A2(
        n_majority7_module_33__and_module_8_res), .ZN(
        n_majority7_module_33__or_module_11_res) );
  AND2_X1 u_majority7_module_33__and_module_10_U1 ( .A1(
        n_majority7_module_33__or_module_8_res), .A2(
        n_majority7_module_33__and_module_9_res), .ZN(
        n_majority7_module_33__and_module_10_res) );
  AND2_X1 u_majority7_module_33__and_module_11_U1 ( .A1(
        n_majority7_module_33__and_module_10_res), .A2(
        n_majority7_module_33__or_module_11_res), .ZN(
        n_majority7_module_33_res) );
  DFF_X1 u_reg_module_34__cini_mul_v000_reg ( .D(n_majority7_module_33_res), 
        .CK(clock_2), .Q(n_reg_module_34_res), .QN() );
  BUF_X1 u_majority7_module_34_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_34_n7) );
  BUF_X1 u_majority7_module_34_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_34_n6) );
  BUF_X1 u_majority7_module_34_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_34_n5) );
  BUF_X1 u_majority7_module_34_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_34_n4) );
  BUF_X1 u_majority7_module_34_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_34_n3) );
  BUF_X1 u_majority7_module_34_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_34_n2) );
  BUF_X1 u_majority7_module_34_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_34_n1) );
  AND2_X1 u_majority7_module_34__and_module_1_U1 ( .A1(
        n_majority7_module_34_n5), .A2(n_majority7_module_34_n4), .ZN(
        n_majority7_module_34__and_module_1_res) );
  OR2_X1 u_majority7_module_34__or_module_1_U1 ( .A1(n_majority7_module_34_n4), 
        .A2(n_majority7_module_34_n5), .ZN(
        n_majority7_module_34__or_module_1_res) );
  AND2_X1 u_majority7_module_34__and_module_2_U1 ( .A1(
        n_majority7_module_34_n7), .A2(n_majority7_module_34_n2), .ZN(
        n_majority7_module_34__and_module_2_res) );
  OR2_X1 u_majority7_module_34__or_module_2_U1 ( .A1(n_majority7_module_34_n2), 
        .A2(n_majority7_module_34_n7), .ZN(
        n_majority7_module_34__or_module_2_res) );
  AND2_X1 u_majority7_module_34__and_module_3_U1 ( .A1(
        n_majority7_module_34_n6), .A2(n_majority7_module_34_n1), .ZN(
        n_majority7_module_34__and_module_3_res) );
  OR2_X1 u_majority7_module_34__or_module_3_U1 ( .A1(n_majority7_module_34_n1), 
        .A2(n_majority7_module_34_n6), .ZN(
        n_majority7_module_34__or_module_3_res) );
  AND2_X1 u_majority7_module_34__and_module_4_U1 ( .A1(
        n_majority7_module_34__and_module_2_res), .A2(
        n_majority7_module_34__and_module_1_res), .ZN(
        n_majority7_module_34__and_module_4_res) );
  OR2_X1 u_majority7_module_34__or_module_4_U1 ( .A1(
        n_majority7_module_34__and_module_1_res), .A2(
        n_majority7_module_34__and_module_2_res), .ZN(
        n_majority7_module_34__or_module_4_res) );
  AND2_X1 u_majority7_module_34__and_module_5_U1 ( .A1(
        n_majority7_module_34__and_module_3_res), .A2(n_majority7_module_34_n3), .ZN(n_majority7_module_34__and_module_5_res) );
  OR2_X1 u_majority7_module_34__or_module_5_U1 ( .A1(n_majority7_module_34_n3), 
        .A2(n_majority7_module_34__and_module_3_res), .ZN(
        n_majority7_module_34__or_module_5_res) );
  AND2_X1 u_majority7_module_34__and_module_6_U1 ( .A1(
        n_majority7_module_34__or_module_1_res), .A2(
        n_majority7_module_34__or_module_2_res), .ZN(
        n_majority7_module_34__and_module_6_res) );
  OR2_X1 u_majority7_module_34__or_module_6_U1 ( .A1(
        n_majority7_module_34__or_module_2_res), .A2(
        n_majority7_module_34__or_module_1_res), .ZN(
        n_majority7_module_34__or_module_6_res) );
  OR2_X1 u_majority7_module_34__or_module_7_U1 ( .A1(
        n_majority7_module_34__and_module_4_res), .A2(
        n_majority7_module_34__and_module_5_res), .ZN(
        n_majority7_module_34__or_module_7_res) );
  AND2_X1 u_majority7_module_34__and_module_7_U1 ( .A1(
        n_majority7_module_34__or_module_3_res), .A2(
        n_majority7_module_34__or_module_4_res), .ZN(
        n_majority7_module_34__and_module_7_res) );
  OR2_X1 u_majority7_module_34__or_module_8_U1 ( .A1(
        n_majority7_module_34__or_module_4_res), .A2(
        n_majority7_module_34__or_module_3_res), .ZN(
        n_majority7_module_34__or_module_8_res) );
  AND2_X1 u_majority7_module_34__and_module_8_U1 ( .A1(
        n_majority7_module_34__or_module_5_res), .A2(
        n_majority7_module_34__and_module_6_res), .ZN(
        n_majority7_module_34__and_module_8_res) );
  OR2_X1 u_majority7_module_34__or_module_9_U1 ( .A1(
        n_majority7_module_34__and_module_6_res), .A2(
        n_majority7_module_34__or_module_5_res), .ZN(
        n_majority7_module_34__or_module_9_res) );
  OR2_X1 u_majority7_module_34__or_module_10_U1 ( .A1(
        n_majority7_module_34__or_module_7_res), .A2(
        n_majority7_module_34__and_module_7_res), .ZN(
        n_majority7_module_34__or_module_10_res) );
  AND2_X1 u_majority7_module_34__and_module_9_U1 ( .A1(
        n_majority7_module_34__or_module_6_res), .A2(
        n_majority7_module_34__or_module_9_res), .ZN(
        n_majority7_module_34__and_module_9_res) );
  OR2_X1 u_majority7_module_34__or_module_11_U1 ( .A1(
        n_majority7_module_34__or_module_10_res), .A2(
        n_majority7_module_34__and_module_8_res), .ZN(
        n_majority7_module_34__or_module_11_res) );
  AND2_X1 u_majority7_module_34__and_module_10_U1 ( .A1(
        n_majority7_module_34__or_module_8_res), .A2(
        n_majority7_module_34__and_module_9_res), .ZN(
        n_majority7_module_34__and_module_10_res) );
  AND2_X1 u_majority7_module_34__and_module_11_U1 ( .A1(
        n_majority7_module_34__and_module_10_res), .A2(
        n_majority7_module_34__or_module_11_res), .ZN(
        n_majority7_module_34_res) );
  DFF_X1 u_reg_module_35__cini_mul_v000_reg ( .D(n_majority7_module_34_res), 
        .CK(clock_2), .Q(n_reg_module_35_res), .QN() );
  BUF_X1 u_majority7_module_35_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_35_n7) );
  BUF_X1 u_majority7_module_35_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_35_n6) );
  BUF_X1 u_majority7_module_35_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_35_n5) );
  BUF_X1 u_majority7_module_35_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_35_n4) );
  BUF_X1 u_majority7_module_35_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_35_n3) );
  BUF_X1 u_majority7_module_35_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_35_n2) );
  BUF_X1 u_majority7_module_35_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_35_n1) );
  AND2_X1 u_majority7_module_35__and_module_1_U1 ( .A1(
        n_majority7_module_35_n5), .A2(n_majority7_module_35_n4), .ZN(
        n_majority7_module_35__and_module_1_res) );
  OR2_X1 u_majority7_module_35__or_module_1_U1 ( .A1(n_majority7_module_35_n4), 
        .A2(n_majority7_module_35_n5), .ZN(
        n_majority7_module_35__or_module_1_res) );
  AND2_X1 u_majority7_module_35__and_module_2_U1 ( .A1(
        n_majority7_module_35_n7), .A2(n_majority7_module_35_n2), .ZN(
        n_majority7_module_35__and_module_2_res) );
  OR2_X1 u_majority7_module_35__or_module_2_U1 ( .A1(n_majority7_module_35_n2), 
        .A2(n_majority7_module_35_n7), .ZN(
        n_majority7_module_35__or_module_2_res) );
  AND2_X1 u_majority7_module_35__and_module_3_U1 ( .A1(
        n_majority7_module_35_n6), .A2(n_majority7_module_35_n1), .ZN(
        n_majority7_module_35__and_module_3_res) );
  OR2_X1 u_majority7_module_35__or_module_3_U1 ( .A1(n_majority7_module_35_n1), 
        .A2(n_majority7_module_35_n6), .ZN(
        n_majority7_module_35__or_module_3_res) );
  AND2_X1 u_majority7_module_35__and_module_4_U1 ( .A1(
        n_majority7_module_35__and_module_2_res), .A2(
        n_majority7_module_35__and_module_1_res), .ZN(
        n_majority7_module_35__and_module_4_res) );
  OR2_X1 u_majority7_module_35__or_module_4_U1 ( .A1(
        n_majority7_module_35__and_module_1_res), .A2(
        n_majority7_module_35__and_module_2_res), .ZN(
        n_majority7_module_35__or_module_4_res) );
  AND2_X1 u_majority7_module_35__and_module_5_U1 ( .A1(
        n_majority7_module_35__and_module_3_res), .A2(n_majority7_module_35_n3), .ZN(n_majority7_module_35__and_module_5_res) );
  OR2_X1 u_majority7_module_35__or_module_5_U1 ( .A1(n_majority7_module_35_n3), 
        .A2(n_majority7_module_35__and_module_3_res), .ZN(
        n_majority7_module_35__or_module_5_res) );
  AND2_X1 u_majority7_module_35__and_module_6_U1 ( .A1(
        n_majority7_module_35__or_module_1_res), .A2(
        n_majority7_module_35__or_module_2_res), .ZN(
        n_majority7_module_35__and_module_6_res) );
  OR2_X1 u_majority7_module_35__or_module_6_U1 ( .A1(
        n_majority7_module_35__or_module_2_res), .A2(
        n_majority7_module_35__or_module_1_res), .ZN(
        n_majority7_module_35__or_module_6_res) );
  OR2_X1 u_majority7_module_35__or_module_7_U1 ( .A1(
        n_majority7_module_35__and_module_4_res), .A2(
        n_majority7_module_35__and_module_5_res), .ZN(
        n_majority7_module_35__or_module_7_res) );
  AND2_X1 u_majority7_module_35__and_module_7_U1 ( .A1(
        n_majority7_module_35__or_module_3_res), .A2(
        n_majority7_module_35__or_module_4_res), .ZN(
        n_majority7_module_35__and_module_7_res) );
  OR2_X1 u_majority7_module_35__or_module_8_U1 ( .A1(
        n_majority7_module_35__or_module_4_res), .A2(
        n_majority7_module_35__or_module_3_res), .ZN(
        n_majority7_module_35__or_module_8_res) );
  AND2_X1 u_majority7_module_35__and_module_8_U1 ( .A1(
        n_majority7_module_35__or_module_5_res), .A2(
        n_majority7_module_35__and_module_6_res), .ZN(
        n_majority7_module_35__and_module_8_res) );
  OR2_X1 u_majority7_module_35__or_module_9_U1 ( .A1(
        n_majority7_module_35__and_module_6_res), .A2(
        n_majority7_module_35__or_module_5_res), .ZN(
        n_majority7_module_35__or_module_9_res) );
  OR2_X1 u_majority7_module_35__or_module_10_U1 ( .A1(
        n_majority7_module_35__or_module_7_res), .A2(
        n_majority7_module_35__and_module_7_res), .ZN(
        n_majority7_module_35__or_module_10_res) );
  AND2_X1 u_majority7_module_35__and_module_9_U1 ( .A1(
        n_majority7_module_35__or_module_6_res), .A2(
        n_majority7_module_35__or_module_9_res), .ZN(
        n_majority7_module_35__and_module_9_res) );
  OR2_X1 u_majority7_module_35__or_module_11_U1 ( .A1(
        n_majority7_module_35__or_module_10_res), .A2(
        n_majority7_module_35__and_module_8_res), .ZN(
        n_majority7_module_35__or_module_11_res) );
  AND2_X1 u_majority7_module_35__and_module_10_U1 ( .A1(
        n_majority7_module_35__or_module_8_res), .A2(
        n_majority7_module_35__and_module_9_res), .ZN(
        n_majority7_module_35__and_module_10_res) );
  AND2_X1 u_majority7_module_35__and_module_11_U1 ( .A1(
        n_majority7_module_35__and_module_10_res), .A2(
        n_majority7_module_35__or_module_11_res), .ZN(
        n_majority7_module_35_res) );
  DFF_X1 u_reg_module_36__cini_mul_v000_reg ( .D(n_majority7_module_35_res), 
        .CK(clock_2), .Q(n_reg_module_36_res), .QN() );
  BUF_X1 u_majority7_module_36_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_36_n7) );
  BUF_X1 u_majority7_module_36_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_36_n6) );
  BUF_X1 u_majority7_module_36_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_36_n5) );
  BUF_X1 u_majority7_module_36_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_36_n4) );
  BUF_X1 u_majority7_module_36_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_36_n3) );
  BUF_X1 u_majority7_module_36_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_36_n2) );
  BUF_X1 u_majority7_module_36_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_36_n1) );
  AND2_X1 u_majority7_module_36__and_module_1_U1 ( .A1(
        n_majority7_module_36_n5), .A2(n_majority7_module_36_n4), .ZN(
        n_majority7_module_36__and_module_1_res) );
  OR2_X1 u_majority7_module_36__or_module_1_U1 ( .A1(n_majority7_module_36_n4), 
        .A2(n_majority7_module_36_n5), .ZN(
        n_majority7_module_36__or_module_1_res) );
  AND2_X1 u_majority7_module_36__and_module_2_U1 ( .A1(
        n_majority7_module_36_n7), .A2(n_majority7_module_36_n2), .ZN(
        n_majority7_module_36__and_module_2_res) );
  OR2_X1 u_majority7_module_36__or_module_2_U1 ( .A1(n_majority7_module_36_n2), 
        .A2(n_majority7_module_36_n7), .ZN(
        n_majority7_module_36__or_module_2_res) );
  AND2_X1 u_majority7_module_36__and_module_3_U1 ( .A1(
        n_majority7_module_36_n6), .A2(n_majority7_module_36_n1), .ZN(
        n_majority7_module_36__and_module_3_res) );
  OR2_X1 u_majority7_module_36__or_module_3_U1 ( .A1(n_majority7_module_36_n1), 
        .A2(n_majority7_module_36_n6), .ZN(
        n_majority7_module_36__or_module_3_res) );
  AND2_X1 u_majority7_module_36__and_module_4_U1 ( .A1(
        n_majority7_module_36__and_module_2_res), .A2(
        n_majority7_module_36__and_module_1_res), .ZN(
        n_majority7_module_36__and_module_4_res) );
  OR2_X1 u_majority7_module_36__or_module_4_U1 ( .A1(
        n_majority7_module_36__and_module_1_res), .A2(
        n_majority7_module_36__and_module_2_res), .ZN(
        n_majority7_module_36__or_module_4_res) );
  AND2_X1 u_majority7_module_36__and_module_5_U1 ( .A1(
        n_majority7_module_36__and_module_3_res), .A2(n_majority7_module_36_n3), .ZN(n_majority7_module_36__and_module_5_res) );
  OR2_X1 u_majority7_module_36__or_module_5_U1 ( .A1(n_majority7_module_36_n3), 
        .A2(n_majority7_module_36__and_module_3_res), .ZN(
        n_majority7_module_36__or_module_5_res) );
  AND2_X1 u_majority7_module_36__and_module_6_U1 ( .A1(
        n_majority7_module_36__or_module_1_res), .A2(
        n_majority7_module_36__or_module_2_res), .ZN(
        n_majority7_module_36__and_module_6_res) );
  OR2_X1 u_majority7_module_36__or_module_6_U1 ( .A1(
        n_majority7_module_36__or_module_2_res), .A2(
        n_majority7_module_36__or_module_1_res), .ZN(
        n_majority7_module_36__or_module_6_res) );
  OR2_X1 u_majority7_module_36__or_module_7_U1 ( .A1(
        n_majority7_module_36__and_module_4_res), .A2(
        n_majority7_module_36__and_module_5_res), .ZN(
        n_majority7_module_36__or_module_7_res) );
  AND2_X1 u_majority7_module_36__and_module_7_U1 ( .A1(
        n_majority7_module_36__or_module_3_res), .A2(
        n_majority7_module_36__or_module_4_res), .ZN(
        n_majority7_module_36__and_module_7_res) );
  OR2_X1 u_majority7_module_36__or_module_8_U1 ( .A1(
        n_majority7_module_36__or_module_4_res), .A2(
        n_majority7_module_36__or_module_3_res), .ZN(
        n_majority7_module_36__or_module_8_res) );
  AND2_X1 u_majority7_module_36__and_module_8_U1 ( .A1(
        n_majority7_module_36__or_module_5_res), .A2(
        n_majority7_module_36__and_module_6_res), .ZN(
        n_majority7_module_36__and_module_8_res) );
  OR2_X1 u_majority7_module_36__or_module_9_U1 ( .A1(
        n_majority7_module_36__and_module_6_res), .A2(
        n_majority7_module_36__or_module_5_res), .ZN(
        n_majority7_module_36__or_module_9_res) );
  OR2_X1 u_majority7_module_36__or_module_10_U1 ( .A1(
        n_majority7_module_36__or_module_7_res), .A2(
        n_majority7_module_36__and_module_7_res), .ZN(
        n_majority7_module_36__or_module_10_res) );
  AND2_X1 u_majority7_module_36__and_module_9_U1 ( .A1(
        n_majority7_module_36__or_module_6_res), .A2(
        n_majority7_module_36__or_module_9_res), .ZN(
        n_majority7_module_36__and_module_9_res) );
  OR2_X1 u_majority7_module_36__or_module_11_U1 ( .A1(
        n_majority7_module_36__or_module_10_res), .A2(
        n_majority7_module_36__and_module_8_res), .ZN(
        n_majority7_module_36__or_module_11_res) );
  AND2_X1 u_majority7_module_36__and_module_10_U1 ( .A1(
        n_majority7_module_36__or_module_8_res), .A2(
        n_majority7_module_36__and_module_9_res), .ZN(
        n_majority7_module_36__and_module_10_res) );
  AND2_X1 u_majority7_module_36__and_module_11_U1 ( .A1(
        n_majority7_module_36__and_module_10_res), .A2(
        n_majority7_module_36__or_module_11_res), .ZN(
        n_majority7_module_36_res) );
  DFF_X1 u_reg_module_37__cini_mul_v000_reg ( .D(n_majority7_module_36_res), 
        .CK(clock_2), .Q(n_reg_module_37_res), .QN() );
  BUF_X1 u_majority7_module_37_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_37_n7) );
  BUF_X1 u_majority7_module_37_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_37_n6) );
  BUF_X1 u_majority7_module_37_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_37_n5) );
  BUF_X1 u_majority7_module_37_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_37_n4) );
  BUF_X1 u_majority7_module_37_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_37_n3) );
  BUF_X1 u_majority7_module_37_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_37_n2) );
  BUF_X1 u_majority7_module_37_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_37_n1) );
  AND2_X1 u_majority7_module_37__and_module_1_U1 ( .A1(
        n_majority7_module_37_n5), .A2(n_majority7_module_37_n4), .ZN(
        n_majority7_module_37__and_module_1_res) );
  OR2_X1 u_majority7_module_37__or_module_1_U1 ( .A1(n_majority7_module_37_n4), 
        .A2(n_majority7_module_37_n5), .ZN(
        n_majority7_module_37__or_module_1_res) );
  AND2_X1 u_majority7_module_37__and_module_2_U1 ( .A1(
        n_majority7_module_37_n7), .A2(n_majority7_module_37_n2), .ZN(
        n_majority7_module_37__and_module_2_res) );
  OR2_X1 u_majority7_module_37__or_module_2_U1 ( .A1(n_majority7_module_37_n2), 
        .A2(n_majority7_module_37_n7), .ZN(
        n_majority7_module_37__or_module_2_res) );
  AND2_X1 u_majority7_module_37__and_module_3_U1 ( .A1(
        n_majority7_module_37_n6), .A2(n_majority7_module_37_n1), .ZN(
        n_majority7_module_37__and_module_3_res) );
  OR2_X1 u_majority7_module_37__or_module_3_U1 ( .A1(n_majority7_module_37_n1), 
        .A2(n_majority7_module_37_n6), .ZN(
        n_majority7_module_37__or_module_3_res) );
  AND2_X1 u_majority7_module_37__and_module_4_U1 ( .A1(
        n_majority7_module_37__and_module_2_res), .A2(
        n_majority7_module_37__and_module_1_res), .ZN(
        n_majority7_module_37__and_module_4_res) );
  OR2_X1 u_majority7_module_37__or_module_4_U1 ( .A1(
        n_majority7_module_37__and_module_1_res), .A2(
        n_majority7_module_37__and_module_2_res), .ZN(
        n_majority7_module_37__or_module_4_res) );
  AND2_X1 u_majority7_module_37__and_module_5_U1 ( .A1(
        n_majority7_module_37__and_module_3_res), .A2(n_majority7_module_37_n3), .ZN(n_majority7_module_37__and_module_5_res) );
  OR2_X1 u_majority7_module_37__or_module_5_U1 ( .A1(n_majority7_module_37_n3), 
        .A2(n_majority7_module_37__and_module_3_res), .ZN(
        n_majority7_module_37__or_module_5_res) );
  AND2_X1 u_majority7_module_37__and_module_6_U1 ( .A1(
        n_majority7_module_37__or_module_1_res), .A2(
        n_majority7_module_37__or_module_2_res), .ZN(
        n_majority7_module_37__and_module_6_res) );
  OR2_X1 u_majority7_module_37__or_module_6_U1 ( .A1(
        n_majority7_module_37__or_module_2_res), .A2(
        n_majority7_module_37__or_module_1_res), .ZN(
        n_majority7_module_37__or_module_6_res) );
  OR2_X1 u_majority7_module_37__or_module_7_U1 ( .A1(
        n_majority7_module_37__and_module_4_res), .A2(
        n_majority7_module_37__and_module_5_res), .ZN(
        n_majority7_module_37__or_module_7_res) );
  AND2_X1 u_majority7_module_37__and_module_7_U1 ( .A1(
        n_majority7_module_37__or_module_3_res), .A2(
        n_majority7_module_37__or_module_4_res), .ZN(
        n_majority7_module_37__and_module_7_res) );
  OR2_X1 u_majority7_module_37__or_module_8_U1 ( .A1(
        n_majority7_module_37__or_module_4_res), .A2(
        n_majority7_module_37__or_module_3_res), .ZN(
        n_majority7_module_37__or_module_8_res) );
  AND2_X1 u_majority7_module_37__and_module_8_U1 ( .A1(
        n_majority7_module_37__or_module_5_res), .A2(
        n_majority7_module_37__and_module_6_res), .ZN(
        n_majority7_module_37__and_module_8_res) );
  OR2_X1 u_majority7_module_37__or_module_9_U1 ( .A1(
        n_majority7_module_37__and_module_6_res), .A2(
        n_majority7_module_37__or_module_5_res), .ZN(
        n_majority7_module_37__or_module_9_res) );
  OR2_X1 u_majority7_module_37__or_module_10_U1 ( .A1(
        n_majority7_module_37__or_module_7_res), .A2(
        n_majority7_module_37__and_module_7_res), .ZN(
        n_majority7_module_37__or_module_10_res) );
  AND2_X1 u_majority7_module_37__and_module_9_U1 ( .A1(
        n_majority7_module_37__or_module_6_res), .A2(
        n_majority7_module_37__or_module_9_res), .ZN(
        n_majority7_module_37__and_module_9_res) );
  OR2_X1 u_majority7_module_37__or_module_11_U1 ( .A1(
        n_majority7_module_37__or_module_10_res), .A2(
        n_majority7_module_37__and_module_8_res), .ZN(
        n_majority7_module_37__or_module_11_res) );
  AND2_X1 u_majority7_module_37__and_module_10_U1 ( .A1(
        n_majority7_module_37__or_module_8_res), .A2(
        n_majority7_module_37__and_module_9_res), .ZN(
        n_majority7_module_37__and_module_10_res) );
  AND2_X1 u_majority7_module_37__and_module_11_U1 ( .A1(
        n_majority7_module_37__and_module_10_res), .A2(
        n_majority7_module_37__or_module_11_res), .ZN(
        n_majority7_module_37_res) );
  DFF_X1 u_reg_module_38__cini_mul_v000_reg ( .D(n_majority7_module_37_res), 
        .CK(clock_2), .Q(n_reg_module_38_res), .QN() );
  BUF_X1 u_majority7_module_38_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_38_n7) );
  BUF_X1 u_majority7_module_38_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_38_n6) );
  BUF_X1 u_majority7_module_38_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_38_n5) );
  BUF_X1 u_majority7_module_38_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_38_n4) );
  BUF_X1 u_majority7_module_38_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_38_n3) );
  BUF_X1 u_majority7_module_38_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_38_n2) );
  BUF_X1 u_majority7_module_38_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_38_n1) );
  AND2_X1 u_majority7_module_38__and_module_1_U1 ( .A1(
        n_majority7_module_38_n5), .A2(n_majority7_module_38_n4), .ZN(
        n_majority7_module_38__and_module_1_res) );
  OR2_X1 u_majority7_module_38__or_module_1_U1 ( .A1(n_majority7_module_38_n4), 
        .A2(n_majority7_module_38_n5), .ZN(
        n_majority7_module_38__or_module_1_res) );
  AND2_X1 u_majority7_module_38__and_module_2_U1 ( .A1(
        n_majority7_module_38_n7), .A2(n_majority7_module_38_n2), .ZN(
        n_majority7_module_38__and_module_2_res) );
  OR2_X1 u_majority7_module_38__or_module_2_U1 ( .A1(n_majority7_module_38_n2), 
        .A2(n_majority7_module_38_n7), .ZN(
        n_majority7_module_38__or_module_2_res) );
  AND2_X1 u_majority7_module_38__and_module_3_U1 ( .A1(
        n_majority7_module_38_n6), .A2(n_majority7_module_38_n1), .ZN(
        n_majority7_module_38__and_module_3_res) );
  OR2_X1 u_majority7_module_38__or_module_3_U1 ( .A1(n_majority7_module_38_n1), 
        .A2(n_majority7_module_38_n6), .ZN(
        n_majority7_module_38__or_module_3_res) );
  AND2_X1 u_majority7_module_38__and_module_4_U1 ( .A1(
        n_majority7_module_38__and_module_2_res), .A2(
        n_majority7_module_38__and_module_1_res), .ZN(
        n_majority7_module_38__and_module_4_res) );
  OR2_X1 u_majority7_module_38__or_module_4_U1 ( .A1(
        n_majority7_module_38__and_module_1_res), .A2(
        n_majority7_module_38__and_module_2_res), .ZN(
        n_majority7_module_38__or_module_4_res) );
  AND2_X1 u_majority7_module_38__and_module_5_U1 ( .A1(
        n_majority7_module_38__and_module_3_res), .A2(n_majority7_module_38_n3), .ZN(n_majority7_module_38__and_module_5_res) );
  OR2_X1 u_majority7_module_38__or_module_5_U1 ( .A1(n_majority7_module_38_n3), 
        .A2(n_majority7_module_38__and_module_3_res), .ZN(
        n_majority7_module_38__or_module_5_res) );
  AND2_X1 u_majority7_module_38__and_module_6_U1 ( .A1(
        n_majority7_module_38__or_module_1_res), .A2(
        n_majority7_module_38__or_module_2_res), .ZN(
        n_majority7_module_38__and_module_6_res) );
  OR2_X1 u_majority7_module_38__or_module_6_U1 ( .A1(
        n_majority7_module_38__or_module_2_res), .A2(
        n_majority7_module_38__or_module_1_res), .ZN(
        n_majority7_module_38__or_module_6_res) );
  OR2_X1 u_majority7_module_38__or_module_7_U1 ( .A1(
        n_majority7_module_38__and_module_4_res), .A2(
        n_majority7_module_38__and_module_5_res), .ZN(
        n_majority7_module_38__or_module_7_res) );
  AND2_X1 u_majority7_module_38__and_module_7_U1 ( .A1(
        n_majority7_module_38__or_module_3_res), .A2(
        n_majority7_module_38__or_module_4_res), .ZN(
        n_majority7_module_38__and_module_7_res) );
  OR2_X1 u_majority7_module_38__or_module_8_U1 ( .A1(
        n_majority7_module_38__or_module_4_res), .A2(
        n_majority7_module_38__or_module_3_res), .ZN(
        n_majority7_module_38__or_module_8_res) );
  AND2_X1 u_majority7_module_38__and_module_8_U1 ( .A1(
        n_majority7_module_38__or_module_5_res), .A2(
        n_majority7_module_38__and_module_6_res), .ZN(
        n_majority7_module_38__and_module_8_res) );
  OR2_X1 u_majority7_module_38__or_module_9_U1 ( .A1(
        n_majority7_module_38__and_module_6_res), .A2(
        n_majority7_module_38__or_module_5_res), .ZN(
        n_majority7_module_38__or_module_9_res) );
  OR2_X1 u_majority7_module_38__or_module_10_U1 ( .A1(
        n_majority7_module_38__or_module_7_res), .A2(
        n_majority7_module_38__and_module_7_res), .ZN(
        n_majority7_module_38__or_module_10_res) );
  AND2_X1 u_majority7_module_38__and_module_9_U1 ( .A1(
        n_majority7_module_38__or_module_6_res), .A2(
        n_majority7_module_38__or_module_9_res), .ZN(
        n_majority7_module_38__and_module_9_res) );
  OR2_X1 u_majority7_module_38__or_module_11_U1 ( .A1(
        n_majority7_module_38__or_module_10_res), .A2(
        n_majority7_module_38__and_module_8_res), .ZN(
        n_majority7_module_38__or_module_11_res) );
  AND2_X1 u_majority7_module_38__and_module_10_U1 ( .A1(
        n_majority7_module_38__or_module_8_res), .A2(
        n_majority7_module_38__and_module_9_res), .ZN(
        n_majority7_module_38__and_module_10_res) );
  AND2_X1 u_majority7_module_38__and_module_11_U1 ( .A1(
        n_majority7_module_38__and_module_10_res), .A2(
        n_majority7_module_38__or_module_11_res), .ZN(
        n_majority7_module_38_res) );
  DFF_X1 u_reg_module_39__cini_mul_v000_reg ( .D(n_majority7_module_38_res), 
        .CK(clock_2), .Q(n_reg_module_39_res), .QN() );
  BUF_X1 u_majority7_module_39_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_39_n7) );
  BUF_X1 u_majority7_module_39_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_39_n6) );
  BUF_X1 u_majority7_module_39_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_39_n5) );
  BUF_X1 u_majority7_module_39_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_39_n4) );
  BUF_X1 u_majority7_module_39_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_39_n3) );
  BUF_X1 u_majority7_module_39_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_39_n2) );
  BUF_X1 u_majority7_module_39_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_39_n1) );
  AND2_X1 u_majority7_module_39__and_module_1_U1 ( .A1(
        n_majority7_module_39_n5), .A2(n_majority7_module_39_n4), .ZN(
        n_majority7_module_39__and_module_1_res) );
  OR2_X1 u_majority7_module_39__or_module_1_U1 ( .A1(n_majority7_module_39_n4), 
        .A2(n_majority7_module_39_n5), .ZN(
        n_majority7_module_39__or_module_1_res) );
  AND2_X1 u_majority7_module_39__and_module_2_U1 ( .A1(
        n_majority7_module_39_n7), .A2(n_majority7_module_39_n2), .ZN(
        n_majority7_module_39__and_module_2_res) );
  OR2_X1 u_majority7_module_39__or_module_2_U1 ( .A1(n_majority7_module_39_n2), 
        .A2(n_majority7_module_39_n7), .ZN(
        n_majority7_module_39__or_module_2_res) );
  AND2_X1 u_majority7_module_39__and_module_3_U1 ( .A1(
        n_majority7_module_39_n6), .A2(n_majority7_module_39_n1), .ZN(
        n_majority7_module_39__and_module_3_res) );
  OR2_X1 u_majority7_module_39__or_module_3_U1 ( .A1(n_majority7_module_39_n1), 
        .A2(n_majority7_module_39_n6), .ZN(
        n_majority7_module_39__or_module_3_res) );
  AND2_X1 u_majority7_module_39__and_module_4_U1 ( .A1(
        n_majority7_module_39__and_module_2_res), .A2(
        n_majority7_module_39__and_module_1_res), .ZN(
        n_majority7_module_39__and_module_4_res) );
  OR2_X1 u_majority7_module_39__or_module_4_U1 ( .A1(
        n_majority7_module_39__and_module_1_res), .A2(
        n_majority7_module_39__and_module_2_res), .ZN(
        n_majority7_module_39__or_module_4_res) );
  AND2_X1 u_majority7_module_39__and_module_5_U1 ( .A1(
        n_majority7_module_39__and_module_3_res), .A2(n_majority7_module_39_n3), .ZN(n_majority7_module_39__and_module_5_res) );
  OR2_X1 u_majority7_module_39__or_module_5_U1 ( .A1(n_majority7_module_39_n3), 
        .A2(n_majority7_module_39__and_module_3_res), .ZN(
        n_majority7_module_39__or_module_5_res) );
  AND2_X1 u_majority7_module_39__and_module_6_U1 ( .A1(
        n_majority7_module_39__or_module_1_res), .A2(
        n_majority7_module_39__or_module_2_res), .ZN(
        n_majority7_module_39__and_module_6_res) );
  OR2_X1 u_majority7_module_39__or_module_6_U1 ( .A1(
        n_majority7_module_39__or_module_2_res), .A2(
        n_majority7_module_39__or_module_1_res), .ZN(
        n_majority7_module_39__or_module_6_res) );
  OR2_X1 u_majority7_module_39__or_module_7_U1 ( .A1(
        n_majority7_module_39__and_module_4_res), .A2(
        n_majority7_module_39__and_module_5_res), .ZN(
        n_majority7_module_39__or_module_7_res) );
  AND2_X1 u_majority7_module_39__and_module_7_U1 ( .A1(
        n_majority7_module_39__or_module_3_res), .A2(
        n_majority7_module_39__or_module_4_res), .ZN(
        n_majority7_module_39__and_module_7_res) );
  OR2_X1 u_majority7_module_39__or_module_8_U1 ( .A1(
        n_majority7_module_39__or_module_4_res), .A2(
        n_majority7_module_39__or_module_3_res), .ZN(
        n_majority7_module_39__or_module_8_res) );
  AND2_X1 u_majority7_module_39__and_module_8_U1 ( .A1(
        n_majority7_module_39__or_module_5_res), .A2(
        n_majority7_module_39__and_module_6_res), .ZN(
        n_majority7_module_39__and_module_8_res) );
  OR2_X1 u_majority7_module_39__or_module_9_U1 ( .A1(
        n_majority7_module_39__and_module_6_res), .A2(
        n_majority7_module_39__or_module_5_res), .ZN(
        n_majority7_module_39__or_module_9_res) );
  OR2_X1 u_majority7_module_39__or_module_10_U1 ( .A1(
        n_majority7_module_39__or_module_7_res), .A2(
        n_majority7_module_39__and_module_7_res), .ZN(
        n_majority7_module_39__or_module_10_res) );
  AND2_X1 u_majority7_module_39__and_module_9_U1 ( .A1(
        n_majority7_module_39__or_module_6_res), .A2(
        n_majority7_module_39__or_module_9_res), .ZN(
        n_majority7_module_39__and_module_9_res) );
  OR2_X1 u_majority7_module_39__or_module_11_U1 ( .A1(
        n_majority7_module_39__or_module_10_res), .A2(
        n_majority7_module_39__and_module_8_res), .ZN(
        n_majority7_module_39__or_module_11_res) );
  AND2_X1 u_majority7_module_39__and_module_10_U1 ( .A1(
        n_majority7_module_39__or_module_8_res), .A2(
        n_majority7_module_39__and_module_9_res), .ZN(
        n_majority7_module_39__and_module_10_res) );
  AND2_X1 u_majority7_module_39__and_module_11_U1 ( .A1(
        n_majority7_module_39__and_module_10_res), .A2(
        n_majority7_module_39__or_module_11_res), .ZN(
        n_majority7_module_39_res) );
  DFF_X1 u_reg_module_40__cini_mul_v000_reg ( .D(n_majority7_module_39_res), 
        .CK(clock_2), .Q(n_reg_module_40_res), .QN() );
  BUF_X1 u_majority7_module_40_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_40_n7) );
  BUF_X1 u_majority7_module_40_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_40_n6) );
  BUF_X1 u_majority7_module_40_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_40_n5) );
  BUF_X1 u_majority7_module_40_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_40_n4) );
  BUF_X1 u_majority7_module_40_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_40_n3) );
  BUF_X1 u_majority7_module_40_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_40_n2) );
  BUF_X1 u_majority7_module_40_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_40_n1) );
  AND2_X1 u_majority7_module_40__and_module_1_U1 ( .A1(
        n_majority7_module_40_n5), .A2(n_majority7_module_40_n4), .ZN(
        n_majority7_module_40__and_module_1_res) );
  OR2_X1 u_majority7_module_40__or_module_1_U1 ( .A1(n_majority7_module_40_n4), 
        .A2(n_majority7_module_40_n5), .ZN(
        n_majority7_module_40__or_module_1_res) );
  AND2_X1 u_majority7_module_40__and_module_2_U1 ( .A1(
        n_majority7_module_40_n7), .A2(n_majority7_module_40_n2), .ZN(
        n_majority7_module_40__and_module_2_res) );
  OR2_X1 u_majority7_module_40__or_module_2_U1 ( .A1(n_majority7_module_40_n2), 
        .A2(n_majority7_module_40_n7), .ZN(
        n_majority7_module_40__or_module_2_res) );
  AND2_X1 u_majority7_module_40__and_module_3_U1 ( .A1(
        n_majority7_module_40_n6), .A2(n_majority7_module_40_n1), .ZN(
        n_majority7_module_40__and_module_3_res) );
  OR2_X1 u_majority7_module_40__or_module_3_U1 ( .A1(n_majority7_module_40_n1), 
        .A2(n_majority7_module_40_n6), .ZN(
        n_majority7_module_40__or_module_3_res) );
  AND2_X1 u_majority7_module_40__and_module_4_U1 ( .A1(
        n_majority7_module_40__and_module_2_res), .A2(
        n_majority7_module_40__and_module_1_res), .ZN(
        n_majority7_module_40__and_module_4_res) );
  OR2_X1 u_majority7_module_40__or_module_4_U1 ( .A1(
        n_majority7_module_40__and_module_1_res), .A2(
        n_majority7_module_40__and_module_2_res), .ZN(
        n_majority7_module_40__or_module_4_res) );
  AND2_X1 u_majority7_module_40__and_module_5_U1 ( .A1(
        n_majority7_module_40__and_module_3_res), .A2(n_majority7_module_40_n3), .ZN(n_majority7_module_40__and_module_5_res) );
  OR2_X1 u_majority7_module_40__or_module_5_U1 ( .A1(n_majority7_module_40_n3), 
        .A2(n_majority7_module_40__and_module_3_res), .ZN(
        n_majority7_module_40__or_module_5_res) );
  AND2_X1 u_majority7_module_40__and_module_6_U1 ( .A1(
        n_majority7_module_40__or_module_1_res), .A2(
        n_majority7_module_40__or_module_2_res), .ZN(
        n_majority7_module_40__and_module_6_res) );
  OR2_X1 u_majority7_module_40__or_module_6_U1 ( .A1(
        n_majority7_module_40__or_module_2_res), .A2(
        n_majority7_module_40__or_module_1_res), .ZN(
        n_majority7_module_40__or_module_6_res) );
  OR2_X1 u_majority7_module_40__or_module_7_U1 ( .A1(
        n_majority7_module_40__and_module_4_res), .A2(
        n_majority7_module_40__and_module_5_res), .ZN(
        n_majority7_module_40__or_module_7_res) );
  AND2_X1 u_majority7_module_40__and_module_7_U1 ( .A1(
        n_majority7_module_40__or_module_3_res), .A2(
        n_majority7_module_40__or_module_4_res), .ZN(
        n_majority7_module_40__and_module_7_res) );
  OR2_X1 u_majority7_module_40__or_module_8_U1 ( .A1(
        n_majority7_module_40__or_module_4_res), .A2(
        n_majority7_module_40__or_module_3_res), .ZN(
        n_majority7_module_40__or_module_8_res) );
  AND2_X1 u_majority7_module_40__and_module_8_U1 ( .A1(
        n_majority7_module_40__or_module_5_res), .A2(
        n_majority7_module_40__and_module_6_res), .ZN(
        n_majority7_module_40__and_module_8_res) );
  OR2_X1 u_majority7_module_40__or_module_9_U1 ( .A1(
        n_majority7_module_40__and_module_6_res), .A2(
        n_majority7_module_40__or_module_5_res), .ZN(
        n_majority7_module_40__or_module_9_res) );
  OR2_X1 u_majority7_module_40__or_module_10_U1 ( .A1(
        n_majority7_module_40__or_module_7_res), .A2(
        n_majority7_module_40__and_module_7_res), .ZN(
        n_majority7_module_40__or_module_10_res) );
  AND2_X1 u_majority7_module_40__and_module_9_U1 ( .A1(
        n_majority7_module_40__or_module_6_res), .A2(
        n_majority7_module_40__or_module_9_res), .ZN(
        n_majority7_module_40__and_module_9_res) );
  OR2_X1 u_majority7_module_40__or_module_11_U1 ( .A1(
        n_majority7_module_40__or_module_10_res), .A2(
        n_majority7_module_40__and_module_8_res), .ZN(
        n_majority7_module_40__or_module_11_res) );
  AND2_X1 u_majority7_module_40__and_module_10_U1 ( .A1(
        n_majority7_module_40__or_module_8_res), .A2(
        n_majority7_module_40__and_module_9_res), .ZN(
        n_majority7_module_40__and_module_10_res) );
  AND2_X1 u_majority7_module_40__and_module_11_U1 ( .A1(
        n_majority7_module_40__and_module_10_res), .A2(
        n_majority7_module_40__or_module_11_res), .ZN(
        n_majority7_module_40_res) );
  DFF_X1 u_reg_module_41__cini_mul_v000_reg ( .D(n_majority7_module_40_res), 
        .CK(clock_2), .Q(n_reg_module_41_res), .QN() );
  BUF_X1 u_majority7_module_41_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_41_n7) );
  BUF_X1 u_majority7_module_41_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_41_n6) );
  BUF_X1 u_majority7_module_41_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_41_n5) );
  BUF_X1 u_majority7_module_41_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_41_n4) );
  BUF_X1 u_majority7_module_41_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_41_n3) );
  BUF_X1 u_majority7_module_41_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_41_n2) );
  BUF_X1 u_majority7_module_41_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_41_n1) );
  AND2_X1 u_majority7_module_41__and_module_1_U1 ( .A1(
        n_majority7_module_41_n5), .A2(n_majority7_module_41_n4), .ZN(
        n_majority7_module_41__and_module_1_res) );
  OR2_X1 u_majority7_module_41__or_module_1_U1 ( .A1(n_majority7_module_41_n4), 
        .A2(n_majority7_module_41_n5), .ZN(
        n_majority7_module_41__or_module_1_res) );
  AND2_X1 u_majority7_module_41__and_module_2_U1 ( .A1(
        n_majority7_module_41_n7), .A2(n_majority7_module_41_n2), .ZN(
        n_majority7_module_41__and_module_2_res) );
  OR2_X1 u_majority7_module_41__or_module_2_U1 ( .A1(n_majority7_module_41_n2), 
        .A2(n_majority7_module_41_n7), .ZN(
        n_majority7_module_41__or_module_2_res) );
  AND2_X1 u_majority7_module_41__and_module_3_U1 ( .A1(
        n_majority7_module_41_n6), .A2(n_majority7_module_41_n1), .ZN(
        n_majority7_module_41__and_module_3_res) );
  OR2_X1 u_majority7_module_41__or_module_3_U1 ( .A1(n_majority7_module_41_n1), 
        .A2(n_majority7_module_41_n6), .ZN(
        n_majority7_module_41__or_module_3_res) );
  AND2_X1 u_majority7_module_41__and_module_4_U1 ( .A1(
        n_majority7_module_41__and_module_2_res), .A2(
        n_majority7_module_41__and_module_1_res), .ZN(
        n_majority7_module_41__and_module_4_res) );
  OR2_X1 u_majority7_module_41__or_module_4_U1 ( .A1(
        n_majority7_module_41__and_module_1_res), .A2(
        n_majority7_module_41__and_module_2_res), .ZN(
        n_majority7_module_41__or_module_4_res) );
  AND2_X1 u_majority7_module_41__and_module_5_U1 ( .A1(
        n_majority7_module_41__and_module_3_res), .A2(n_majority7_module_41_n3), .ZN(n_majority7_module_41__and_module_5_res) );
  OR2_X1 u_majority7_module_41__or_module_5_U1 ( .A1(n_majority7_module_41_n3), 
        .A2(n_majority7_module_41__and_module_3_res), .ZN(
        n_majority7_module_41__or_module_5_res) );
  AND2_X1 u_majority7_module_41__and_module_6_U1 ( .A1(
        n_majority7_module_41__or_module_1_res), .A2(
        n_majority7_module_41__or_module_2_res), .ZN(
        n_majority7_module_41__and_module_6_res) );
  OR2_X1 u_majority7_module_41__or_module_6_U1 ( .A1(
        n_majority7_module_41__or_module_2_res), .A2(
        n_majority7_module_41__or_module_1_res), .ZN(
        n_majority7_module_41__or_module_6_res) );
  OR2_X1 u_majority7_module_41__or_module_7_U1 ( .A1(
        n_majority7_module_41__and_module_4_res), .A2(
        n_majority7_module_41__and_module_5_res), .ZN(
        n_majority7_module_41__or_module_7_res) );
  AND2_X1 u_majority7_module_41__and_module_7_U1 ( .A1(
        n_majority7_module_41__or_module_3_res), .A2(
        n_majority7_module_41__or_module_4_res), .ZN(
        n_majority7_module_41__and_module_7_res) );
  OR2_X1 u_majority7_module_41__or_module_8_U1 ( .A1(
        n_majority7_module_41__or_module_4_res), .A2(
        n_majority7_module_41__or_module_3_res), .ZN(
        n_majority7_module_41__or_module_8_res) );
  AND2_X1 u_majority7_module_41__and_module_8_U1 ( .A1(
        n_majority7_module_41__or_module_5_res), .A2(
        n_majority7_module_41__and_module_6_res), .ZN(
        n_majority7_module_41__and_module_8_res) );
  OR2_X1 u_majority7_module_41__or_module_9_U1 ( .A1(
        n_majority7_module_41__and_module_6_res), .A2(
        n_majority7_module_41__or_module_5_res), .ZN(
        n_majority7_module_41__or_module_9_res) );
  OR2_X1 u_majority7_module_41__or_module_10_U1 ( .A1(
        n_majority7_module_41__or_module_7_res), .A2(
        n_majority7_module_41__and_module_7_res), .ZN(
        n_majority7_module_41__or_module_10_res) );
  AND2_X1 u_majority7_module_41__and_module_9_U1 ( .A1(
        n_majority7_module_41__or_module_6_res), .A2(
        n_majority7_module_41__or_module_9_res), .ZN(
        n_majority7_module_41__and_module_9_res) );
  OR2_X1 u_majority7_module_41__or_module_11_U1 ( .A1(
        n_majority7_module_41__or_module_10_res), .A2(
        n_majority7_module_41__and_module_8_res), .ZN(
        n_majority7_module_41__or_module_11_res) );
  AND2_X1 u_majority7_module_41__and_module_10_U1 ( .A1(
        n_majority7_module_41__or_module_8_res), .A2(
        n_majority7_module_41__and_module_9_res), .ZN(
        n_majority7_module_41__and_module_10_res) );
  AND2_X1 u_majority7_module_41__and_module_11_U1 ( .A1(
        n_majority7_module_41__and_module_10_res), .A2(
        n_majority7_module_41__or_module_11_res), .ZN(
        n_majority7_module_41_res) );
  DFF_X1 u_reg_module_42__cini_mul_v000_reg ( .D(n_majority7_module_41_res), 
        .CK(clock_2), .Q(n_reg_module_42_res), .QN() );
  BUF_X1 u_majority7_module_42_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_42_n7) );
  BUF_X1 u_majority7_module_42_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_42_n6) );
  BUF_X1 u_majority7_module_42_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_42_n5) );
  BUF_X1 u_majority7_module_42_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_42_n4) );
  BUF_X1 u_majority7_module_42_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_42_n3) );
  BUF_X1 u_majority7_module_42_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_42_n2) );
  BUF_X1 u_majority7_module_42_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_42_n1) );
  AND2_X1 u_majority7_module_42__and_module_1_U1 ( .A1(
        n_majority7_module_42_n5), .A2(n_majority7_module_42_n4), .ZN(
        n_majority7_module_42__and_module_1_res) );
  OR2_X1 u_majority7_module_42__or_module_1_U1 ( .A1(n_majority7_module_42_n4), 
        .A2(n_majority7_module_42_n5), .ZN(
        n_majority7_module_42__or_module_1_res) );
  AND2_X1 u_majority7_module_42__and_module_2_U1 ( .A1(
        n_majority7_module_42_n7), .A2(n_majority7_module_42_n2), .ZN(
        n_majority7_module_42__and_module_2_res) );
  OR2_X1 u_majority7_module_42__or_module_2_U1 ( .A1(n_majority7_module_42_n2), 
        .A2(n_majority7_module_42_n7), .ZN(
        n_majority7_module_42__or_module_2_res) );
  AND2_X1 u_majority7_module_42__and_module_3_U1 ( .A1(
        n_majority7_module_42_n6), .A2(n_majority7_module_42_n1), .ZN(
        n_majority7_module_42__and_module_3_res) );
  OR2_X1 u_majority7_module_42__or_module_3_U1 ( .A1(n_majority7_module_42_n1), 
        .A2(n_majority7_module_42_n6), .ZN(
        n_majority7_module_42__or_module_3_res) );
  AND2_X1 u_majority7_module_42__and_module_4_U1 ( .A1(
        n_majority7_module_42__and_module_2_res), .A2(
        n_majority7_module_42__and_module_1_res), .ZN(
        n_majority7_module_42__and_module_4_res) );
  OR2_X1 u_majority7_module_42__or_module_4_U1 ( .A1(
        n_majority7_module_42__and_module_1_res), .A2(
        n_majority7_module_42__and_module_2_res), .ZN(
        n_majority7_module_42__or_module_4_res) );
  AND2_X1 u_majority7_module_42__and_module_5_U1 ( .A1(
        n_majority7_module_42__and_module_3_res), .A2(n_majority7_module_42_n3), .ZN(n_majority7_module_42__and_module_5_res) );
  OR2_X1 u_majority7_module_42__or_module_5_U1 ( .A1(n_majority7_module_42_n3), 
        .A2(n_majority7_module_42__and_module_3_res), .ZN(
        n_majority7_module_42__or_module_5_res) );
  AND2_X1 u_majority7_module_42__and_module_6_U1 ( .A1(
        n_majority7_module_42__or_module_1_res), .A2(
        n_majority7_module_42__or_module_2_res), .ZN(
        n_majority7_module_42__and_module_6_res) );
  OR2_X1 u_majority7_module_42__or_module_6_U1 ( .A1(
        n_majority7_module_42__or_module_2_res), .A2(
        n_majority7_module_42__or_module_1_res), .ZN(
        n_majority7_module_42__or_module_6_res) );
  OR2_X1 u_majority7_module_42__or_module_7_U1 ( .A1(
        n_majority7_module_42__and_module_4_res), .A2(
        n_majority7_module_42__and_module_5_res), .ZN(
        n_majority7_module_42__or_module_7_res) );
  AND2_X1 u_majority7_module_42__and_module_7_U1 ( .A1(
        n_majority7_module_42__or_module_3_res), .A2(
        n_majority7_module_42__or_module_4_res), .ZN(
        n_majority7_module_42__and_module_7_res) );
  OR2_X1 u_majority7_module_42__or_module_8_U1 ( .A1(
        n_majority7_module_42__or_module_4_res), .A2(
        n_majority7_module_42__or_module_3_res), .ZN(
        n_majority7_module_42__or_module_8_res) );
  AND2_X1 u_majority7_module_42__and_module_8_U1 ( .A1(
        n_majority7_module_42__or_module_5_res), .A2(
        n_majority7_module_42__and_module_6_res), .ZN(
        n_majority7_module_42__and_module_8_res) );
  OR2_X1 u_majority7_module_42__or_module_9_U1 ( .A1(
        n_majority7_module_42__and_module_6_res), .A2(
        n_majority7_module_42__or_module_5_res), .ZN(
        n_majority7_module_42__or_module_9_res) );
  OR2_X1 u_majority7_module_42__or_module_10_U1 ( .A1(
        n_majority7_module_42__or_module_7_res), .A2(
        n_majority7_module_42__and_module_7_res), .ZN(
        n_majority7_module_42__or_module_10_res) );
  AND2_X1 u_majority7_module_42__and_module_9_U1 ( .A1(
        n_majority7_module_42__or_module_6_res), .A2(
        n_majority7_module_42__or_module_9_res), .ZN(
        n_majority7_module_42__and_module_9_res) );
  OR2_X1 u_majority7_module_42__or_module_11_U1 ( .A1(
        n_majority7_module_42__or_module_10_res), .A2(
        n_majority7_module_42__and_module_8_res), .ZN(
        n_majority7_module_42__or_module_11_res) );
  AND2_X1 u_majority7_module_42__and_module_10_U1 ( .A1(
        n_majority7_module_42__or_module_8_res), .A2(
        n_majority7_module_42__and_module_9_res), .ZN(
        n_majority7_module_42__and_module_10_res) );
  AND2_X1 u_majority7_module_42__and_module_11_U1 ( .A1(
        n_majority7_module_42__and_module_10_res), .A2(
        n_majority7_module_42__or_module_11_res), .ZN(
        n_majority7_module_42_res) );
  DFF_X1 u_reg_module_43__cini_mul_v000_reg ( .D(n_majority7_module_42_res), 
        .CK(clock_2), .Q(n_reg_module_43_res), .QN() );
  BUF_X1 u_majority7_module_43_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_43_n7) );
  BUF_X1 u_majority7_module_43_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_43_n6) );
  BUF_X1 u_majority7_module_43_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_43_n5) );
  BUF_X1 u_majority7_module_43_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_43_n4) );
  BUF_X1 u_majority7_module_43_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_43_n3) );
  BUF_X1 u_majority7_module_43_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_43_n2) );
  BUF_X1 u_majority7_module_43_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_43_n1) );
  AND2_X1 u_majority7_module_43__and_module_1_U1 ( .A1(
        n_majority7_module_43_n5), .A2(n_majority7_module_43_n4), .ZN(
        n_majority7_module_43__and_module_1_res) );
  OR2_X1 u_majority7_module_43__or_module_1_U1 ( .A1(n_majority7_module_43_n4), 
        .A2(n_majority7_module_43_n5), .ZN(
        n_majority7_module_43__or_module_1_res) );
  AND2_X1 u_majority7_module_43__and_module_2_U1 ( .A1(
        n_majority7_module_43_n7), .A2(n_majority7_module_43_n2), .ZN(
        n_majority7_module_43__and_module_2_res) );
  OR2_X1 u_majority7_module_43__or_module_2_U1 ( .A1(n_majority7_module_43_n2), 
        .A2(n_majority7_module_43_n7), .ZN(
        n_majority7_module_43__or_module_2_res) );
  AND2_X1 u_majority7_module_43__and_module_3_U1 ( .A1(
        n_majority7_module_43_n6), .A2(n_majority7_module_43_n1), .ZN(
        n_majority7_module_43__and_module_3_res) );
  OR2_X1 u_majority7_module_43__or_module_3_U1 ( .A1(n_majority7_module_43_n1), 
        .A2(n_majority7_module_43_n6), .ZN(
        n_majority7_module_43__or_module_3_res) );
  AND2_X1 u_majority7_module_43__and_module_4_U1 ( .A1(
        n_majority7_module_43__and_module_2_res), .A2(
        n_majority7_module_43__and_module_1_res), .ZN(
        n_majority7_module_43__and_module_4_res) );
  OR2_X1 u_majority7_module_43__or_module_4_U1 ( .A1(
        n_majority7_module_43__and_module_1_res), .A2(
        n_majority7_module_43__and_module_2_res), .ZN(
        n_majority7_module_43__or_module_4_res) );
  AND2_X1 u_majority7_module_43__and_module_5_U1 ( .A1(
        n_majority7_module_43__and_module_3_res), .A2(n_majority7_module_43_n3), .ZN(n_majority7_module_43__and_module_5_res) );
  OR2_X1 u_majority7_module_43__or_module_5_U1 ( .A1(n_majority7_module_43_n3), 
        .A2(n_majority7_module_43__and_module_3_res), .ZN(
        n_majority7_module_43__or_module_5_res) );
  AND2_X1 u_majority7_module_43__and_module_6_U1 ( .A1(
        n_majority7_module_43__or_module_1_res), .A2(
        n_majority7_module_43__or_module_2_res), .ZN(
        n_majority7_module_43__and_module_6_res) );
  OR2_X1 u_majority7_module_43__or_module_6_U1 ( .A1(
        n_majority7_module_43__or_module_2_res), .A2(
        n_majority7_module_43__or_module_1_res), .ZN(
        n_majority7_module_43__or_module_6_res) );
  OR2_X1 u_majority7_module_43__or_module_7_U1 ( .A1(
        n_majority7_module_43__and_module_4_res), .A2(
        n_majority7_module_43__and_module_5_res), .ZN(
        n_majority7_module_43__or_module_7_res) );
  AND2_X1 u_majority7_module_43__and_module_7_U1 ( .A1(
        n_majority7_module_43__or_module_3_res), .A2(
        n_majority7_module_43__or_module_4_res), .ZN(
        n_majority7_module_43__and_module_7_res) );
  OR2_X1 u_majority7_module_43__or_module_8_U1 ( .A1(
        n_majority7_module_43__or_module_4_res), .A2(
        n_majority7_module_43__or_module_3_res), .ZN(
        n_majority7_module_43__or_module_8_res) );
  AND2_X1 u_majority7_module_43__and_module_8_U1 ( .A1(
        n_majority7_module_43__or_module_5_res), .A2(
        n_majority7_module_43__and_module_6_res), .ZN(
        n_majority7_module_43__and_module_8_res) );
  OR2_X1 u_majority7_module_43__or_module_9_U1 ( .A1(
        n_majority7_module_43__and_module_6_res), .A2(
        n_majority7_module_43__or_module_5_res), .ZN(
        n_majority7_module_43__or_module_9_res) );
  OR2_X1 u_majority7_module_43__or_module_10_U1 ( .A1(
        n_majority7_module_43__or_module_7_res), .A2(
        n_majority7_module_43__and_module_7_res), .ZN(
        n_majority7_module_43__or_module_10_res) );
  AND2_X1 u_majority7_module_43__and_module_9_U1 ( .A1(
        n_majority7_module_43__or_module_6_res), .A2(
        n_majority7_module_43__or_module_9_res), .ZN(
        n_majority7_module_43__and_module_9_res) );
  OR2_X1 u_majority7_module_43__or_module_11_U1 ( .A1(
        n_majority7_module_43__or_module_10_res), .A2(
        n_majority7_module_43__and_module_8_res), .ZN(
        n_majority7_module_43__or_module_11_res) );
  AND2_X1 u_majority7_module_43__and_module_10_U1 ( .A1(
        n_majority7_module_43__or_module_8_res), .A2(
        n_majority7_module_43__and_module_9_res), .ZN(
        n_majority7_module_43__and_module_10_res) );
  AND2_X1 u_majority7_module_43__and_module_11_U1 ( .A1(
        n_majority7_module_43__and_module_10_res), .A2(
        n_majority7_module_43__or_module_11_res), .ZN(
        n_majority7_module_43_res) );
  DFF_X1 u_reg_module_44__cini_mul_v000_reg ( .D(n_majority7_module_43_res), 
        .CK(clock_2), .Q(n_reg_module_44_res), .QN() );
  BUF_X1 u_majority7_module_44_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_44_n7) );
  BUF_X1 u_majority7_module_44_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_44_n6) );
  BUF_X1 u_majority7_module_44_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_44_n5) );
  BUF_X1 u_majority7_module_44_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_44_n4) );
  BUF_X1 u_majority7_module_44_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_44_n3) );
  BUF_X1 u_majority7_module_44_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_44_n2) );
  BUF_X1 u_majority7_module_44_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_44_n1) );
  AND2_X1 u_majority7_module_44__and_module_1_U1 ( .A1(
        n_majority7_module_44_n1), .A2(n_majority7_module_44_n5), .ZN(
        n_majority7_module_44__and_module_1_res) );
  OR2_X1 u_majority7_module_44__or_module_1_U1 ( .A1(n_majority7_module_44_n5), 
        .A2(n_majority7_module_44_n1), .ZN(
        n_majority7_module_44__or_module_1_res) );
  AND2_X1 u_majority7_module_44__and_module_2_U1 ( .A1(
        n_majority7_module_44_n7), .A2(n_majority7_module_44_n3), .ZN(
        n_majority7_module_44__and_module_2_res) );
  OR2_X1 u_majority7_module_44__or_module_2_U1 ( .A1(n_majority7_module_44_n3), 
        .A2(n_majority7_module_44_n7), .ZN(
        n_majority7_module_44__or_module_2_res) );
  AND2_X1 u_majority7_module_44__and_module_3_U1 ( .A1(
        n_majority7_module_44_n6), .A2(n_majority7_module_44_n2), .ZN(
        n_majority7_module_44__and_module_3_res) );
  OR2_X1 u_majority7_module_44__or_module_3_U1 ( .A1(n_majority7_module_44_n2), 
        .A2(n_majority7_module_44_n6), .ZN(
        n_majority7_module_44__or_module_3_res) );
  AND2_X1 u_majority7_module_44__and_module_4_U1 ( .A1(
        n_majority7_module_44__and_module_2_res), .A2(
        n_majority7_module_44__and_module_1_res), .ZN(
        n_majority7_module_44__and_module_4_res) );
  OR2_X1 u_majority7_module_44__or_module_4_U1 ( .A1(
        n_majority7_module_44__and_module_1_res), .A2(
        n_majority7_module_44__and_module_2_res), .ZN(
        n_majority7_module_44__or_module_4_res) );
  AND2_X1 u_majority7_module_44__and_module_5_U1 ( .A1(
        n_majority7_module_44__and_module_3_res), .A2(n_majority7_module_44_n4), .ZN(n_majority7_module_44__and_module_5_res) );
  OR2_X1 u_majority7_module_44__or_module_5_U1 ( .A1(n_majority7_module_44_n4), 
        .A2(n_majority7_module_44__and_module_3_res), .ZN(
        n_majority7_module_44__or_module_5_res) );
  AND2_X1 u_majority7_module_44__and_module_6_U1 ( .A1(
        n_majority7_module_44__or_module_1_res), .A2(
        n_majority7_module_44__or_module_2_res), .ZN(
        n_majority7_module_44__and_module_6_res) );
  OR2_X1 u_majority7_module_44__or_module_6_U1 ( .A1(
        n_majority7_module_44__or_module_2_res), .A2(
        n_majority7_module_44__or_module_1_res), .ZN(
        n_majority7_module_44__or_module_6_res) );
  OR2_X1 u_majority7_module_44__or_module_7_U1 ( .A1(
        n_majority7_module_44__and_module_4_res), .A2(
        n_majority7_module_44__and_module_5_res), .ZN(
        n_majority7_module_44__or_module_7_res) );
  AND2_X1 u_majority7_module_44__and_module_7_U1 ( .A1(
        n_majority7_module_44__or_module_3_res), .A2(
        n_majority7_module_44__or_module_4_res), .ZN(
        n_majority7_module_44__and_module_7_res) );
  OR2_X1 u_majority7_module_44__or_module_8_U1 ( .A1(
        n_majority7_module_44__or_module_4_res), .A2(
        n_majority7_module_44__or_module_3_res), .ZN(
        n_majority7_module_44__or_module_8_res) );
  AND2_X1 u_majority7_module_44__and_module_8_U1 ( .A1(
        n_majority7_module_44__or_module_5_res), .A2(
        n_majority7_module_44__and_module_6_res), .ZN(
        n_majority7_module_44__and_module_8_res) );
  OR2_X1 u_majority7_module_44__or_module_9_U1 ( .A1(
        n_majority7_module_44__and_module_6_res), .A2(
        n_majority7_module_44__or_module_5_res), .ZN(
        n_majority7_module_44__or_module_9_res) );
  OR2_X1 u_majority7_module_44__or_module_10_U1 ( .A1(
        n_majority7_module_44__or_module_7_res), .A2(
        n_majority7_module_44__and_module_7_res), .ZN(
        n_majority7_module_44__or_module_10_res) );
  AND2_X1 u_majority7_module_44__and_module_9_U1 ( .A1(
        n_majority7_module_44__or_module_6_res), .A2(
        n_majority7_module_44__or_module_9_res), .ZN(
        n_majority7_module_44__and_module_9_res) );
  OR2_X1 u_majority7_module_44__or_module_11_U1 ( .A1(
        n_majority7_module_44__or_module_10_res), .A2(
        n_majority7_module_44__and_module_8_res), .ZN(
        n_majority7_module_44__or_module_11_res) );
  AND2_X1 u_majority7_module_44__and_module_10_U1 ( .A1(
        n_majority7_module_44__or_module_8_res), .A2(
        n_majority7_module_44__and_module_9_res), .ZN(
        n_majority7_module_44__and_module_10_res) );
  AND2_X1 u_majority7_module_44__and_module_11_U1 ( .A1(
        n_majority7_module_44__and_module_10_res), .A2(
        n_majority7_module_44__or_module_11_res), .ZN(
        n_majority7_module_44_res) );
  DFF_X1 u_reg_module_45__cini_mul_v000_reg ( .D(n_majority7_module_44_res), 
        .CK(clock_2), .Q(n_reg_module_45_res), .QN() );
  BUF_X1 u_majority7_module_45_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_45_n7) );
  BUF_X1 u_majority7_module_45_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_45_n6) );
  BUF_X1 u_majority7_module_45_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_45_n5) );
  BUF_X1 u_majority7_module_45_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_45_n4) );
  BUF_X1 u_majority7_module_45_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_45_n3) );
  BUF_X1 u_majority7_module_45_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_45_n2) );
  BUF_X1 u_majority7_module_45_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_45_n1) );
  AND2_X1 u_majority7_module_45__and_module_1_U1 ( .A1(
        n_majority7_module_45_n1), .A2(n_majority7_module_45_n5), .ZN(
        n_majority7_module_45__and_module_1_res) );
  OR2_X1 u_majority7_module_45__or_module_1_U1 ( .A1(n_majority7_module_45_n5), 
        .A2(n_majority7_module_45_n1), .ZN(
        n_majority7_module_45__or_module_1_res) );
  AND2_X1 u_majority7_module_45__and_module_2_U1 ( .A1(
        n_majority7_module_45_n7), .A2(n_majority7_module_45_n3), .ZN(
        n_majority7_module_45__and_module_2_res) );
  OR2_X1 u_majority7_module_45__or_module_2_U1 ( .A1(n_majority7_module_45_n3), 
        .A2(n_majority7_module_45_n7), .ZN(
        n_majority7_module_45__or_module_2_res) );
  AND2_X1 u_majority7_module_45__and_module_3_U1 ( .A1(
        n_majority7_module_45_n6), .A2(n_majority7_module_45_n2), .ZN(
        n_majority7_module_45__and_module_3_res) );
  OR2_X1 u_majority7_module_45__or_module_3_U1 ( .A1(n_majority7_module_45_n2), 
        .A2(n_majority7_module_45_n6), .ZN(
        n_majority7_module_45__or_module_3_res) );
  AND2_X1 u_majority7_module_45__and_module_4_U1 ( .A1(
        n_majority7_module_45__and_module_2_res), .A2(
        n_majority7_module_45__and_module_1_res), .ZN(
        n_majority7_module_45__and_module_4_res) );
  OR2_X1 u_majority7_module_45__or_module_4_U1 ( .A1(
        n_majority7_module_45__and_module_1_res), .A2(
        n_majority7_module_45__and_module_2_res), .ZN(
        n_majority7_module_45__or_module_4_res) );
  AND2_X1 u_majority7_module_45__and_module_5_U1 ( .A1(
        n_majority7_module_45__and_module_3_res), .A2(n_majority7_module_45_n4), .ZN(n_majority7_module_45__and_module_5_res) );
  OR2_X1 u_majority7_module_45__or_module_5_U1 ( .A1(n_majority7_module_45_n4), 
        .A2(n_majority7_module_45__and_module_3_res), .ZN(
        n_majority7_module_45__or_module_5_res) );
  AND2_X1 u_majority7_module_45__and_module_6_U1 ( .A1(
        n_majority7_module_45__or_module_1_res), .A2(
        n_majority7_module_45__or_module_2_res), .ZN(
        n_majority7_module_45__and_module_6_res) );
  OR2_X1 u_majority7_module_45__or_module_6_U1 ( .A1(
        n_majority7_module_45__or_module_2_res), .A2(
        n_majority7_module_45__or_module_1_res), .ZN(
        n_majority7_module_45__or_module_6_res) );
  OR2_X1 u_majority7_module_45__or_module_7_U1 ( .A1(
        n_majority7_module_45__and_module_4_res), .A2(
        n_majority7_module_45__and_module_5_res), .ZN(
        n_majority7_module_45__or_module_7_res) );
  AND2_X1 u_majority7_module_45__and_module_7_U1 ( .A1(
        n_majority7_module_45__or_module_3_res), .A2(
        n_majority7_module_45__or_module_4_res), .ZN(
        n_majority7_module_45__and_module_7_res) );
  OR2_X1 u_majority7_module_45__or_module_8_U1 ( .A1(
        n_majority7_module_45__or_module_4_res), .A2(
        n_majority7_module_45__or_module_3_res), .ZN(
        n_majority7_module_45__or_module_8_res) );
  AND2_X1 u_majority7_module_45__and_module_8_U1 ( .A1(
        n_majority7_module_45__or_module_5_res), .A2(
        n_majority7_module_45__and_module_6_res), .ZN(
        n_majority7_module_45__and_module_8_res) );
  OR2_X1 u_majority7_module_45__or_module_9_U1 ( .A1(
        n_majority7_module_45__and_module_6_res), .A2(
        n_majority7_module_45__or_module_5_res), .ZN(
        n_majority7_module_45__or_module_9_res) );
  OR2_X1 u_majority7_module_45__or_module_10_U1 ( .A1(
        n_majority7_module_45__or_module_7_res), .A2(
        n_majority7_module_45__and_module_7_res), .ZN(
        n_majority7_module_45__or_module_10_res) );
  AND2_X1 u_majority7_module_45__and_module_9_U1 ( .A1(
        n_majority7_module_45__or_module_6_res), .A2(
        n_majority7_module_45__or_module_9_res), .ZN(
        n_majority7_module_45__and_module_9_res) );
  OR2_X1 u_majority7_module_45__or_module_11_U1 ( .A1(
        n_majority7_module_45__or_module_10_res), .A2(
        n_majority7_module_45__and_module_8_res), .ZN(
        n_majority7_module_45__or_module_11_res) );
  AND2_X1 u_majority7_module_45__and_module_10_U1 ( .A1(
        n_majority7_module_45__or_module_8_res), .A2(
        n_majority7_module_45__and_module_9_res), .ZN(
        n_majority7_module_45__and_module_10_res) );
  AND2_X1 u_majority7_module_45__and_module_11_U1 ( .A1(
        n_majority7_module_45__and_module_10_res), .A2(
        n_majority7_module_45__or_module_11_res), .ZN(
        n_majority7_module_45_res) );
  DFF_X1 u_reg_module_46__cini_mul_v000_reg ( .D(n_majority7_module_45_res), 
        .CK(clock_2), .Q(n_reg_module_46_res), .QN() );
  BUF_X1 u_majority7_module_46_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_46_n7) );
  BUF_X1 u_majority7_module_46_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_46_n6) );
  BUF_X1 u_majority7_module_46_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_46_n5) );
  BUF_X1 u_majority7_module_46_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_46_n4) );
  BUF_X1 u_majority7_module_46_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_46_n3) );
  BUF_X1 u_majority7_module_46_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_46_n2) );
  BUF_X1 u_majority7_module_46_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_46_n1) );
  AND2_X1 u_majority7_module_46__and_module_1_U1 ( .A1(
        n_majority7_module_46_n1), .A2(n_majority7_module_46_n5), .ZN(
        n_majority7_module_46__and_module_1_res) );
  OR2_X1 u_majority7_module_46__or_module_1_U1 ( .A1(n_majority7_module_46_n5), 
        .A2(n_majority7_module_46_n1), .ZN(
        n_majority7_module_46__or_module_1_res) );
  AND2_X1 u_majority7_module_46__and_module_2_U1 ( .A1(
        n_majority7_module_46_n7), .A2(n_majority7_module_46_n3), .ZN(
        n_majority7_module_46__and_module_2_res) );
  OR2_X1 u_majority7_module_46__or_module_2_U1 ( .A1(n_majority7_module_46_n3), 
        .A2(n_majority7_module_46_n7), .ZN(
        n_majority7_module_46__or_module_2_res) );
  AND2_X1 u_majority7_module_46__and_module_3_U1 ( .A1(
        n_majority7_module_46_n6), .A2(n_majority7_module_46_n2), .ZN(
        n_majority7_module_46__and_module_3_res) );
  OR2_X1 u_majority7_module_46__or_module_3_U1 ( .A1(n_majority7_module_46_n2), 
        .A2(n_majority7_module_46_n6), .ZN(
        n_majority7_module_46__or_module_3_res) );
  AND2_X1 u_majority7_module_46__and_module_4_U1 ( .A1(
        n_majority7_module_46__and_module_2_res), .A2(
        n_majority7_module_46__and_module_1_res), .ZN(
        n_majority7_module_46__and_module_4_res) );
  OR2_X1 u_majority7_module_46__or_module_4_U1 ( .A1(
        n_majority7_module_46__and_module_1_res), .A2(
        n_majority7_module_46__and_module_2_res), .ZN(
        n_majority7_module_46__or_module_4_res) );
  AND2_X1 u_majority7_module_46__and_module_5_U1 ( .A1(
        n_majority7_module_46__and_module_3_res), .A2(n_majority7_module_46_n4), .ZN(n_majority7_module_46__and_module_5_res) );
  OR2_X1 u_majority7_module_46__or_module_5_U1 ( .A1(n_majority7_module_46_n4), 
        .A2(n_majority7_module_46__and_module_3_res), .ZN(
        n_majority7_module_46__or_module_5_res) );
  AND2_X1 u_majority7_module_46__and_module_6_U1 ( .A1(
        n_majority7_module_46__or_module_1_res), .A2(
        n_majority7_module_46__or_module_2_res), .ZN(
        n_majority7_module_46__and_module_6_res) );
  OR2_X1 u_majority7_module_46__or_module_6_U1 ( .A1(
        n_majority7_module_46__or_module_2_res), .A2(
        n_majority7_module_46__or_module_1_res), .ZN(
        n_majority7_module_46__or_module_6_res) );
  OR2_X1 u_majority7_module_46__or_module_7_U1 ( .A1(
        n_majority7_module_46__and_module_4_res), .A2(
        n_majority7_module_46__and_module_5_res), .ZN(
        n_majority7_module_46__or_module_7_res) );
  AND2_X1 u_majority7_module_46__and_module_7_U1 ( .A1(
        n_majority7_module_46__or_module_3_res), .A2(
        n_majority7_module_46__or_module_4_res), .ZN(
        n_majority7_module_46__and_module_7_res) );
  OR2_X1 u_majority7_module_46__or_module_8_U1 ( .A1(
        n_majority7_module_46__or_module_4_res), .A2(
        n_majority7_module_46__or_module_3_res), .ZN(
        n_majority7_module_46__or_module_8_res) );
  AND2_X1 u_majority7_module_46__and_module_8_U1 ( .A1(
        n_majority7_module_46__or_module_5_res), .A2(
        n_majority7_module_46__and_module_6_res), .ZN(
        n_majority7_module_46__and_module_8_res) );
  OR2_X1 u_majority7_module_46__or_module_9_U1 ( .A1(
        n_majority7_module_46__and_module_6_res), .A2(
        n_majority7_module_46__or_module_5_res), .ZN(
        n_majority7_module_46__or_module_9_res) );
  OR2_X1 u_majority7_module_46__or_module_10_U1 ( .A1(
        n_majority7_module_46__or_module_7_res), .A2(
        n_majority7_module_46__and_module_7_res), .ZN(
        n_majority7_module_46__or_module_10_res) );
  AND2_X1 u_majority7_module_46__and_module_9_U1 ( .A1(
        n_majority7_module_46__or_module_6_res), .A2(
        n_majority7_module_46__or_module_9_res), .ZN(
        n_majority7_module_46__and_module_9_res) );
  OR2_X1 u_majority7_module_46__or_module_11_U1 ( .A1(
        n_majority7_module_46__or_module_10_res), .A2(
        n_majority7_module_46__and_module_8_res), .ZN(
        n_majority7_module_46__or_module_11_res) );
  AND2_X1 u_majority7_module_46__and_module_10_U1 ( .A1(
        n_majority7_module_46__or_module_8_res), .A2(
        n_majority7_module_46__and_module_9_res), .ZN(
        n_majority7_module_46__and_module_10_res) );
  AND2_X1 u_majority7_module_46__and_module_11_U1 ( .A1(
        n_majority7_module_46__and_module_10_res), .A2(
        n_majority7_module_46__or_module_11_res), .ZN(
        n_majority7_module_46_res) );
  DFF_X1 u_reg_module_47__cini_mul_v000_reg ( .D(n_majority7_module_46_res), 
        .CK(clock_2), .Q(n_reg_module_47_res), .QN() );
  BUF_X1 u_majority7_module_47_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_47_n7) );
  BUF_X1 u_majority7_module_47_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_47_n6) );
  BUF_X1 u_majority7_module_47_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_47_n5) );
  BUF_X1 u_majority7_module_47_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_47_n4) );
  BUF_X1 u_majority7_module_47_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_47_n3) );
  BUF_X1 u_majority7_module_47_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_47_n2) );
  BUF_X1 u_majority7_module_47_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_47_n1) );
  AND2_X1 u_majority7_module_47__and_module_1_U1 ( .A1(
        n_majority7_module_47_n1), .A2(n_majority7_module_47_n5), .ZN(
        n_majority7_module_47__and_module_1_res) );
  OR2_X1 u_majority7_module_47__or_module_1_U1 ( .A1(n_majority7_module_47_n5), 
        .A2(n_majority7_module_47_n1), .ZN(
        n_majority7_module_47__or_module_1_res) );
  AND2_X1 u_majority7_module_47__and_module_2_U1 ( .A1(
        n_majority7_module_47_n7), .A2(n_majority7_module_47_n3), .ZN(
        n_majority7_module_47__and_module_2_res) );
  OR2_X1 u_majority7_module_47__or_module_2_U1 ( .A1(n_majority7_module_47_n3), 
        .A2(n_majority7_module_47_n7), .ZN(
        n_majority7_module_47__or_module_2_res) );
  AND2_X1 u_majority7_module_47__and_module_3_U1 ( .A1(
        n_majority7_module_47_n6), .A2(n_majority7_module_47_n2), .ZN(
        n_majority7_module_47__and_module_3_res) );
  OR2_X1 u_majority7_module_47__or_module_3_U1 ( .A1(n_majority7_module_47_n2), 
        .A2(n_majority7_module_47_n6), .ZN(
        n_majority7_module_47__or_module_3_res) );
  AND2_X1 u_majority7_module_47__and_module_4_U1 ( .A1(
        n_majority7_module_47__and_module_2_res), .A2(
        n_majority7_module_47__and_module_1_res), .ZN(
        n_majority7_module_47__and_module_4_res) );
  OR2_X1 u_majority7_module_47__or_module_4_U1 ( .A1(
        n_majority7_module_47__and_module_1_res), .A2(
        n_majority7_module_47__and_module_2_res), .ZN(
        n_majority7_module_47__or_module_4_res) );
  AND2_X1 u_majority7_module_47__and_module_5_U1 ( .A1(
        n_majority7_module_47__and_module_3_res), .A2(n_majority7_module_47_n4), .ZN(n_majority7_module_47__and_module_5_res) );
  OR2_X1 u_majority7_module_47__or_module_5_U1 ( .A1(n_majority7_module_47_n4), 
        .A2(n_majority7_module_47__and_module_3_res), .ZN(
        n_majority7_module_47__or_module_5_res) );
  AND2_X1 u_majority7_module_47__and_module_6_U1 ( .A1(
        n_majority7_module_47__or_module_1_res), .A2(
        n_majority7_module_47__or_module_2_res), .ZN(
        n_majority7_module_47__and_module_6_res) );
  OR2_X1 u_majority7_module_47__or_module_6_U1 ( .A1(
        n_majority7_module_47__or_module_2_res), .A2(
        n_majority7_module_47__or_module_1_res), .ZN(
        n_majority7_module_47__or_module_6_res) );
  OR2_X1 u_majority7_module_47__or_module_7_U1 ( .A1(
        n_majority7_module_47__and_module_4_res), .A2(
        n_majority7_module_47__and_module_5_res), .ZN(
        n_majority7_module_47__or_module_7_res) );
  AND2_X1 u_majority7_module_47__and_module_7_U1 ( .A1(
        n_majority7_module_47__or_module_3_res), .A2(
        n_majority7_module_47__or_module_4_res), .ZN(
        n_majority7_module_47__and_module_7_res) );
  OR2_X1 u_majority7_module_47__or_module_8_U1 ( .A1(
        n_majority7_module_47__or_module_4_res), .A2(
        n_majority7_module_47__or_module_3_res), .ZN(
        n_majority7_module_47__or_module_8_res) );
  AND2_X1 u_majority7_module_47__and_module_8_U1 ( .A1(
        n_majority7_module_47__or_module_5_res), .A2(
        n_majority7_module_47__and_module_6_res), .ZN(
        n_majority7_module_47__and_module_8_res) );
  OR2_X1 u_majority7_module_47__or_module_9_U1 ( .A1(
        n_majority7_module_47__and_module_6_res), .A2(
        n_majority7_module_47__or_module_5_res), .ZN(
        n_majority7_module_47__or_module_9_res) );
  OR2_X1 u_majority7_module_47__or_module_10_U1 ( .A1(
        n_majority7_module_47__or_module_7_res), .A2(
        n_majority7_module_47__and_module_7_res), .ZN(
        n_majority7_module_47__or_module_10_res) );
  AND2_X1 u_majority7_module_47__and_module_9_U1 ( .A1(
        n_majority7_module_47__or_module_6_res), .A2(
        n_majority7_module_47__or_module_9_res), .ZN(
        n_majority7_module_47__and_module_9_res) );
  OR2_X1 u_majority7_module_47__or_module_11_U1 ( .A1(
        n_majority7_module_47__or_module_10_res), .A2(
        n_majority7_module_47__and_module_8_res), .ZN(
        n_majority7_module_47__or_module_11_res) );
  AND2_X1 u_majority7_module_47__and_module_10_U1 ( .A1(
        n_majority7_module_47__or_module_8_res), .A2(
        n_majority7_module_47__and_module_9_res), .ZN(
        n_majority7_module_47__and_module_10_res) );
  AND2_X1 u_majority7_module_47__and_module_11_U1 ( .A1(
        n_majority7_module_47__and_module_10_res), .A2(
        n_majority7_module_47__or_module_11_res), .ZN(
        n_majority7_module_47_res) );
  DFF_X1 u_reg_module_48__cini_mul_v000_reg ( .D(n_majority7_module_47_res), 
        .CK(clock_2), .Q(n_reg_module_48_res), .QN() );
  BUF_X1 u_majority7_module_48_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_48_n7) );
  BUF_X1 u_majority7_module_48_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_48_n6) );
  BUF_X1 u_majority7_module_48_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_48_n5) );
  BUF_X1 u_majority7_module_48_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_48_n4) );
  BUF_X1 u_majority7_module_48_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_48_n3) );
  BUF_X1 u_majority7_module_48_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_48_n2) );
  BUF_X1 u_majority7_module_48_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_48_n1) );
  AND2_X1 u_majority7_module_48__and_module_1_U1 ( .A1(
        n_majority7_module_48_n5), .A2(n_majority7_module_48_n4), .ZN(
        n_majority7_module_48__and_module_1_res) );
  OR2_X1 u_majority7_module_48__or_module_1_U1 ( .A1(n_majority7_module_48_n4), 
        .A2(n_majority7_module_48_n5), .ZN(
        n_majority7_module_48__or_module_1_res) );
  AND2_X1 u_majority7_module_48__and_module_2_U1 ( .A1(
        n_majority7_module_48_n7), .A2(n_majority7_module_48_n2), .ZN(
        n_majority7_module_48__and_module_2_res) );
  OR2_X1 u_majority7_module_48__or_module_2_U1 ( .A1(n_majority7_module_48_n2), 
        .A2(n_majority7_module_48_n7), .ZN(
        n_majority7_module_48__or_module_2_res) );
  AND2_X1 u_majority7_module_48__and_module_3_U1 ( .A1(
        n_majority7_module_48_n6), .A2(n_majority7_module_48_n1), .ZN(
        n_majority7_module_48__and_module_3_res) );
  OR2_X1 u_majority7_module_48__or_module_3_U1 ( .A1(n_majority7_module_48_n1), 
        .A2(n_majority7_module_48_n6), .ZN(
        n_majority7_module_48__or_module_3_res) );
  AND2_X1 u_majority7_module_48__and_module_4_U1 ( .A1(
        n_majority7_module_48__and_module_2_res), .A2(
        n_majority7_module_48__and_module_1_res), .ZN(
        n_majority7_module_48__and_module_4_res) );
  OR2_X1 u_majority7_module_48__or_module_4_U1 ( .A1(
        n_majority7_module_48__and_module_1_res), .A2(
        n_majority7_module_48__and_module_2_res), .ZN(
        n_majority7_module_48__or_module_4_res) );
  AND2_X1 u_majority7_module_48__and_module_5_U1 ( .A1(
        n_majority7_module_48__and_module_3_res), .A2(n_majority7_module_48_n3), .ZN(n_majority7_module_48__and_module_5_res) );
  OR2_X1 u_majority7_module_48__or_module_5_U1 ( .A1(n_majority7_module_48_n3), 
        .A2(n_majority7_module_48__and_module_3_res), .ZN(
        n_majority7_module_48__or_module_5_res) );
  AND2_X1 u_majority7_module_48__and_module_6_U1 ( .A1(
        n_majority7_module_48__or_module_1_res), .A2(
        n_majority7_module_48__or_module_2_res), .ZN(
        n_majority7_module_48__and_module_6_res) );
  OR2_X1 u_majority7_module_48__or_module_6_U1 ( .A1(
        n_majority7_module_48__or_module_2_res), .A2(
        n_majority7_module_48__or_module_1_res), .ZN(
        n_majority7_module_48__or_module_6_res) );
  OR2_X1 u_majority7_module_48__or_module_7_U1 ( .A1(
        n_majority7_module_48__and_module_4_res), .A2(
        n_majority7_module_48__and_module_5_res), .ZN(
        n_majority7_module_48__or_module_7_res) );
  AND2_X1 u_majority7_module_48__and_module_7_U1 ( .A1(
        n_majority7_module_48__or_module_3_res), .A2(
        n_majority7_module_48__or_module_4_res), .ZN(
        n_majority7_module_48__and_module_7_res) );
  OR2_X1 u_majority7_module_48__or_module_8_U1 ( .A1(
        n_majority7_module_48__or_module_4_res), .A2(
        n_majority7_module_48__or_module_3_res), .ZN(
        n_majority7_module_48__or_module_8_res) );
  AND2_X1 u_majority7_module_48__and_module_8_U1 ( .A1(
        n_majority7_module_48__or_module_5_res), .A2(
        n_majority7_module_48__and_module_6_res), .ZN(
        n_majority7_module_48__and_module_8_res) );
  OR2_X1 u_majority7_module_48__or_module_9_U1 ( .A1(
        n_majority7_module_48__and_module_6_res), .A2(
        n_majority7_module_48__or_module_5_res), .ZN(
        n_majority7_module_48__or_module_9_res) );
  OR2_X1 u_majority7_module_48__or_module_10_U1 ( .A1(
        n_majority7_module_48__or_module_7_res), .A2(
        n_majority7_module_48__and_module_7_res), .ZN(
        n_majority7_module_48__or_module_10_res) );
  AND2_X1 u_majority7_module_48__and_module_9_U1 ( .A1(
        n_majority7_module_48__or_module_6_res), .A2(
        n_majority7_module_48__or_module_9_res), .ZN(
        n_majority7_module_48__and_module_9_res) );
  OR2_X1 u_majority7_module_48__or_module_11_U1 ( .A1(
        n_majority7_module_48__or_module_10_res), .A2(
        n_majority7_module_48__and_module_8_res), .ZN(
        n_majority7_module_48__or_module_11_res) );
  AND2_X1 u_majority7_module_48__and_module_10_U1 ( .A1(
        n_majority7_module_48__or_module_8_res), .A2(
        n_majority7_module_48__and_module_9_res), .ZN(
        n_majority7_module_48__and_module_10_res) );
  AND2_X1 u_majority7_module_48__and_module_11_U1 ( .A1(
        n_majority7_module_48__and_module_10_res), .A2(
        n_majority7_module_48__or_module_11_res), .ZN(
        n_majority7_module_48_res) );
  DFF_X1 u_reg_module_49__cini_mul_v000_reg ( .D(n_majority7_module_48_res), 
        .CK(clock_3), .Q(n_reg_module_49_res), .QN() );
  BUF_X1 u_majority7_module_49_U7 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_49_n7) );
  BUF_X1 u_majority7_module_49_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_49_n6) );
  BUF_X1 u_majority7_module_49_U5 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_49_n5) );
  BUF_X1 u_majority7_module_49_U4 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_49_n4) );
  BUF_X1 u_majority7_module_49_U3 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_49_n3) );
  BUF_X1 u_majority7_module_49_U2 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_49_n2) );
  BUF_X1 u_majority7_module_49_U1 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_49_n1) );
  AND2_X1 u_majority7_module_49__and_module_1_U1 ( .A1(
        n_majority7_module_49_n5), .A2(n_majority7_module_49_n4), .ZN(
        n_majority7_module_49__and_module_1_res) );
  OR2_X1 u_majority7_module_49__or_module_1_U1 ( .A1(n_majority7_module_49_n4), 
        .A2(n_majority7_module_49_n5), .ZN(
        n_majority7_module_49__or_module_1_res) );
  AND2_X1 u_majority7_module_49__and_module_2_U1 ( .A1(
        n_majority7_module_49_n7), .A2(n_majority7_module_49_n2), .ZN(
        n_majority7_module_49__and_module_2_res) );
  OR2_X1 u_majority7_module_49__or_module_2_U1 ( .A1(n_majority7_module_49_n2), 
        .A2(n_majority7_module_49_n7), .ZN(
        n_majority7_module_49__or_module_2_res) );
  AND2_X1 u_majority7_module_49__and_module_3_U1 ( .A1(
        n_majority7_module_49_n6), .A2(n_majority7_module_49_n1), .ZN(
        n_majority7_module_49__and_module_3_res) );
  OR2_X1 u_majority7_module_49__or_module_3_U1 ( .A1(n_majority7_module_49_n1), 
        .A2(n_majority7_module_49_n6), .ZN(
        n_majority7_module_49__or_module_3_res) );
  AND2_X1 u_majority7_module_49__and_module_4_U1 ( .A1(
        n_majority7_module_49__and_module_2_res), .A2(
        n_majority7_module_49__and_module_1_res), .ZN(
        n_majority7_module_49__and_module_4_res) );
  OR2_X1 u_majority7_module_49__or_module_4_U1 ( .A1(
        n_majority7_module_49__and_module_1_res), .A2(
        n_majority7_module_49__and_module_2_res), .ZN(
        n_majority7_module_49__or_module_4_res) );
  AND2_X1 u_majority7_module_49__and_module_5_U1 ( .A1(
        n_majority7_module_49__and_module_3_res), .A2(n_majority7_module_49_n3), .ZN(n_majority7_module_49__and_module_5_res) );
  OR2_X1 u_majority7_module_49__or_module_5_U1 ( .A1(n_majority7_module_49_n3), 
        .A2(n_majority7_module_49__and_module_3_res), .ZN(
        n_majority7_module_49__or_module_5_res) );
  AND2_X1 u_majority7_module_49__and_module_6_U1 ( .A1(
        n_majority7_module_49__or_module_1_res), .A2(
        n_majority7_module_49__or_module_2_res), .ZN(
        n_majority7_module_49__and_module_6_res) );
  OR2_X1 u_majority7_module_49__or_module_6_U1 ( .A1(
        n_majority7_module_49__or_module_2_res), .A2(
        n_majority7_module_49__or_module_1_res), .ZN(
        n_majority7_module_49__or_module_6_res) );
  OR2_X1 u_majority7_module_49__or_module_7_U1 ( .A1(
        n_majority7_module_49__and_module_4_res), .A2(
        n_majority7_module_49__and_module_5_res), .ZN(
        n_majority7_module_49__or_module_7_res) );
  AND2_X1 u_majority7_module_49__and_module_7_U1 ( .A1(
        n_majority7_module_49__or_module_3_res), .A2(
        n_majority7_module_49__or_module_4_res), .ZN(
        n_majority7_module_49__and_module_7_res) );
  OR2_X1 u_majority7_module_49__or_module_8_U1 ( .A1(
        n_majority7_module_49__or_module_4_res), .A2(
        n_majority7_module_49__or_module_3_res), .ZN(
        n_majority7_module_49__or_module_8_res) );
  AND2_X1 u_majority7_module_49__and_module_8_U1 ( .A1(
        n_majority7_module_49__or_module_5_res), .A2(
        n_majority7_module_49__and_module_6_res), .ZN(
        n_majority7_module_49__and_module_8_res) );
  OR2_X1 u_majority7_module_49__or_module_9_U1 ( .A1(
        n_majority7_module_49__and_module_6_res), .A2(
        n_majority7_module_49__or_module_5_res), .ZN(
        n_majority7_module_49__or_module_9_res) );
  OR2_X1 u_majority7_module_49__or_module_10_U1 ( .A1(
        n_majority7_module_49__or_module_7_res), .A2(
        n_majority7_module_49__and_module_7_res), .ZN(
        n_majority7_module_49__or_module_10_res) );
  AND2_X1 u_majority7_module_49__and_module_9_U1 ( .A1(
        n_majority7_module_49__or_module_6_res), .A2(
        n_majority7_module_49__or_module_9_res), .ZN(
        n_majority7_module_49__and_module_9_res) );
  OR2_X1 u_majority7_module_49__or_module_11_U1 ( .A1(
        n_majority7_module_49__or_module_10_res), .A2(
        n_majority7_module_49__and_module_8_res), .ZN(
        n_majority7_module_49__or_module_11_res) );
  AND2_X1 u_majority7_module_49__and_module_10_U1 ( .A1(
        n_majority7_module_49__or_module_8_res), .A2(
        n_majority7_module_49__and_module_9_res), .ZN(
        n_majority7_module_49__and_module_10_res) );
  AND2_X1 u_majority7_module_49__and_module_11_U1 ( .A1(
        n_majority7_module_49__and_module_10_res), .A2(
        n_majority7_module_49__or_module_11_res), .ZN(
        n_majority7_module_49_res) );
  DFF_X1 u_reg_module_50__cini_mul_v000_reg ( .D(n_majority7_module_49_res), 
        .CK(clock_3), .Q(n_reg_module_50_res), .QN() );
  BUF_X1 u_majority7_module_50_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_50_n7) );
  BUF_X1 u_majority7_module_50_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_50_n6) );
  BUF_X1 u_majority7_module_50_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_50_n5) );
  BUF_X1 u_majority7_module_50_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_50_n4) );
  BUF_X1 u_majority7_module_50_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_50_n3) );
  BUF_X1 u_majority7_module_50_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_50_n2) );
  BUF_X1 u_majority7_module_50_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_50_n1) );
  AND2_X1 u_majority7_module_50__and_module_1_U1 ( .A1(
        n_majority7_module_50_n7), .A2(n_majority7_module_50_n1), .ZN(
        n_majority7_module_50__and_module_1_res) );
  OR2_X1 u_majority7_module_50__or_module_1_U1 ( .A1(n_majority7_module_50_n1), 
        .A2(n_majority7_module_50_n7), .ZN(
        n_majority7_module_50__or_module_1_res) );
  AND2_X1 u_majority7_module_50__and_module_2_U1 ( .A1(
        n_majority7_module_50_n5), .A2(n_majority7_module_50_n3), .ZN(
        n_majority7_module_50__and_module_2_res) );
  OR2_X1 u_majority7_module_50__or_module_2_U1 ( .A1(n_majority7_module_50_n3), 
        .A2(n_majority7_module_50_n5), .ZN(
        n_majority7_module_50__or_module_2_res) );
  AND2_X1 u_majority7_module_50__and_module_3_U1 ( .A1(
        n_majority7_module_50_n6), .A2(n_majority7_module_50_n4), .ZN(
        n_majority7_module_50__and_module_3_res) );
  OR2_X1 u_majority7_module_50__or_module_3_U1 ( .A1(n_majority7_module_50_n4), 
        .A2(n_majority7_module_50_n6), .ZN(
        n_majority7_module_50__or_module_3_res) );
  AND2_X1 u_majority7_module_50__and_module_4_U1 ( .A1(
        n_majority7_module_50__and_module_2_res), .A2(
        n_majority7_module_50__and_module_1_res), .ZN(
        n_majority7_module_50__and_module_4_res) );
  OR2_X1 u_majority7_module_50__or_module_4_U1 ( .A1(
        n_majority7_module_50__and_module_1_res), .A2(
        n_majority7_module_50__and_module_2_res), .ZN(
        n_majority7_module_50__or_module_4_res) );
  AND2_X1 u_majority7_module_50__and_module_5_U1 ( .A1(
        n_majority7_module_50__and_module_3_res), .A2(n_majority7_module_50_n2), .ZN(n_majority7_module_50__and_module_5_res) );
  OR2_X1 u_majority7_module_50__or_module_5_U1 ( .A1(n_majority7_module_50_n2), 
        .A2(n_majority7_module_50__and_module_3_res), .ZN(
        n_majority7_module_50__or_module_5_res) );
  AND2_X1 u_majority7_module_50__and_module_6_U1 ( .A1(
        n_majority7_module_50__or_module_1_res), .A2(
        n_majority7_module_50__or_module_2_res), .ZN(
        n_majority7_module_50__and_module_6_res) );
  OR2_X1 u_majority7_module_50__or_module_6_U1 ( .A1(
        n_majority7_module_50__or_module_2_res), .A2(
        n_majority7_module_50__or_module_1_res), .ZN(
        n_majority7_module_50__or_module_6_res) );
  OR2_X1 u_majority7_module_50__or_module_7_U1 ( .A1(
        n_majority7_module_50__and_module_4_res), .A2(
        n_majority7_module_50__and_module_5_res), .ZN(
        n_majority7_module_50__or_module_7_res) );
  AND2_X1 u_majority7_module_50__and_module_7_U1 ( .A1(
        n_majority7_module_50__or_module_3_res), .A2(
        n_majority7_module_50__or_module_4_res), .ZN(
        n_majority7_module_50__and_module_7_res) );
  OR2_X1 u_majority7_module_50__or_module_8_U1 ( .A1(
        n_majority7_module_50__or_module_4_res), .A2(
        n_majority7_module_50__or_module_3_res), .ZN(
        n_majority7_module_50__or_module_8_res) );
  AND2_X1 u_majority7_module_50__and_module_8_U1 ( .A1(
        n_majority7_module_50__or_module_5_res), .A2(
        n_majority7_module_50__and_module_6_res), .ZN(
        n_majority7_module_50__and_module_8_res) );
  OR2_X1 u_majority7_module_50__or_module_9_U1 ( .A1(
        n_majority7_module_50__and_module_6_res), .A2(
        n_majority7_module_50__or_module_5_res), .ZN(
        n_majority7_module_50__or_module_9_res) );
  OR2_X1 u_majority7_module_50__or_module_10_U1 ( .A1(
        n_majority7_module_50__or_module_7_res), .A2(
        n_majority7_module_50__and_module_7_res), .ZN(
        n_majority7_module_50__or_module_10_res) );
  AND2_X1 u_majority7_module_50__and_module_9_U1 ( .A1(
        n_majority7_module_50__or_module_6_res), .A2(
        n_majority7_module_50__or_module_9_res), .ZN(
        n_majority7_module_50__and_module_9_res) );
  OR2_X1 u_majority7_module_50__or_module_11_U1 ( .A1(
        n_majority7_module_50__or_module_10_res), .A2(
        n_majority7_module_50__and_module_8_res), .ZN(
        n_majority7_module_50__or_module_11_res) );
  AND2_X1 u_majority7_module_50__and_module_10_U1 ( .A1(
        n_majority7_module_50__or_module_8_res), .A2(
        n_majority7_module_50__and_module_9_res), .ZN(
        n_majority7_module_50__and_module_10_res) );
  AND2_X1 u_majority7_module_50__and_module_11_U1 ( .A1(
        n_majority7_module_50__and_module_10_res), .A2(
        n_majority7_module_50__or_module_11_res), .ZN(
        n_majority7_module_50_res) );
  DFF_X1 u_reg_module_51__cini_mul_v000_reg ( .D(n_majority7_module_50_res), 
        .CK(clock_3), .Q(n_reg_module_51_res), .QN() );
  BUF_X1 u_majority7_module_51_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_51_n7) );
  BUF_X1 u_majority7_module_51_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_51_n6) );
  BUF_X1 u_majority7_module_51_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_51_n5) );
  BUF_X1 u_majority7_module_51_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_51_n4) );
  BUF_X1 u_majority7_module_51_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_51_n3) );
  BUF_X1 u_majority7_module_51_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_51_n2) );
  BUF_X1 u_majority7_module_51_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_51_n1) );
  AND2_X1 u_majority7_module_51__and_module_1_U1 ( .A1(
        n_majority7_module_51_n7), .A2(n_majority7_module_51_n1), .ZN(
        n_majority7_module_51__and_module_1_res) );
  OR2_X1 u_majority7_module_51__or_module_1_U1 ( .A1(n_majority7_module_51_n1), 
        .A2(n_majority7_module_51_n7), .ZN(
        n_majority7_module_51__or_module_1_res) );
  AND2_X1 u_majority7_module_51__and_module_2_U1 ( .A1(
        n_majority7_module_51_n5), .A2(n_majority7_module_51_n3), .ZN(
        n_majority7_module_51__and_module_2_res) );
  OR2_X1 u_majority7_module_51__or_module_2_U1 ( .A1(n_majority7_module_51_n3), 
        .A2(n_majority7_module_51_n5), .ZN(
        n_majority7_module_51__or_module_2_res) );
  AND2_X1 u_majority7_module_51__and_module_3_U1 ( .A1(
        n_majority7_module_51_n6), .A2(n_majority7_module_51_n4), .ZN(
        n_majority7_module_51__and_module_3_res) );
  OR2_X1 u_majority7_module_51__or_module_3_U1 ( .A1(n_majority7_module_51_n4), 
        .A2(n_majority7_module_51_n6), .ZN(
        n_majority7_module_51__or_module_3_res) );
  AND2_X1 u_majority7_module_51__and_module_4_U1 ( .A1(
        n_majority7_module_51__and_module_2_res), .A2(
        n_majority7_module_51__and_module_1_res), .ZN(
        n_majority7_module_51__and_module_4_res) );
  OR2_X1 u_majority7_module_51__or_module_4_U1 ( .A1(
        n_majority7_module_51__and_module_1_res), .A2(
        n_majority7_module_51__and_module_2_res), .ZN(
        n_majority7_module_51__or_module_4_res) );
  AND2_X1 u_majority7_module_51__and_module_5_U1 ( .A1(
        n_majority7_module_51__and_module_3_res), .A2(n_majority7_module_51_n2), .ZN(n_majority7_module_51__and_module_5_res) );
  OR2_X1 u_majority7_module_51__or_module_5_U1 ( .A1(n_majority7_module_51_n2), 
        .A2(n_majority7_module_51__and_module_3_res), .ZN(
        n_majority7_module_51__or_module_5_res) );
  AND2_X1 u_majority7_module_51__and_module_6_U1 ( .A1(
        n_majority7_module_51__or_module_1_res), .A2(
        n_majority7_module_51__or_module_2_res), .ZN(
        n_majority7_module_51__and_module_6_res) );
  OR2_X1 u_majority7_module_51__or_module_6_U1 ( .A1(
        n_majority7_module_51__or_module_2_res), .A2(
        n_majority7_module_51__or_module_1_res), .ZN(
        n_majority7_module_51__or_module_6_res) );
  OR2_X1 u_majority7_module_51__or_module_7_U1 ( .A1(
        n_majority7_module_51__and_module_4_res), .A2(
        n_majority7_module_51__and_module_5_res), .ZN(
        n_majority7_module_51__or_module_7_res) );
  AND2_X1 u_majority7_module_51__and_module_7_U1 ( .A1(
        n_majority7_module_51__or_module_3_res), .A2(
        n_majority7_module_51__or_module_4_res), .ZN(
        n_majority7_module_51__and_module_7_res) );
  OR2_X1 u_majority7_module_51__or_module_8_U1 ( .A1(
        n_majority7_module_51__or_module_4_res), .A2(
        n_majority7_module_51__or_module_3_res), .ZN(
        n_majority7_module_51__or_module_8_res) );
  AND2_X1 u_majority7_module_51__and_module_8_U1 ( .A1(
        n_majority7_module_51__or_module_5_res), .A2(
        n_majority7_module_51__and_module_6_res), .ZN(
        n_majority7_module_51__and_module_8_res) );
  OR2_X1 u_majority7_module_51__or_module_9_U1 ( .A1(
        n_majority7_module_51__and_module_6_res), .A2(
        n_majority7_module_51__or_module_5_res), .ZN(
        n_majority7_module_51__or_module_9_res) );
  OR2_X1 u_majority7_module_51__or_module_10_U1 ( .A1(
        n_majority7_module_51__or_module_7_res), .A2(
        n_majority7_module_51__and_module_7_res), .ZN(
        n_majority7_module_51__or_module_10_res) );
  AND2_X1 u_majority7_module_51__and_module_9_U1 ( .A1(
        n_majority7_module_51__or_module_6_res), .A2(
        n_majority7_module_51__or_module_9_res), .ZN(
        n_majority7_module_51__and_module_9_res) );
  OR2_X1 u_majority7_module_51__or_module_11_U1 ( .A1(
        n_majority7_module_51__or_module_10_res), .A2(
        n_majority7_module_51__and_module_8_res), .ZN(
        n_majority7_module_51__or_module_11_res) );
  AND2_X1 u_majority7_module_51__and_module_10_U1 ( .A1(
        n_majority7_module_51__or_module_8_res), .A2(
        n_majority7_module_51__and_module_9_res), .ZN(
        n_majority7_module_51__and_module_10_res) );
  AND2_X1 u_majority7_module_51__and_module_11_U1 ( .A1(
        n_majority7_module_51__and_module_10_res), .A2(
        n_majority7_module_51__or_module_11_res), .ZN(
        n_majority7_module_51_res) );
  DFF_X1 u_reg_module_52__cini_mul_v000_reg ( .D(n_majority7_module_51_res), 
        .CK(clock_3), .Q(n_reg_module_52_res), .QN() );
  BUF_X1 u_majority7_module_52_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_52_n7) );
  BUF_X1 u_majority7_module_52_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_52_n6) );
  BUF_X1 u_majority7_module_52_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_52_n5) );
  BUF_X1 u_majority7_module_52_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_52_n4) );
  BUF_X1 u_majority7_module_52_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_52_n3) );
  BUF_X1 u_majority7_module_52_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_52_n2) );
  BUF_X1 u_majority7_module_52_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_52_n1) );
  AND2_X1 u_majority7_module_52__and_module_1_U1 ( .A1(
        n_majority7_module_52_n5), .A2(n_majority7_module_52_n4), .ZN(
        n_majority7_module_52__and_module_1_res) );
  OR2_X1 u_majority7_module_52__or_module_1_U1 ( .A1(n_majority7_module_52_n4), 
        .A2(n_majority7_module_52_n5), .ZN(
        n_majority7_module_52__or_module_1_res) );
  AND2_X1 u_majority7_module_52__and_module_2_U1 ( .A1(
        n_majority7_module_52_n7), .A2(n_majority7_module_52_n2), .ZN(
        n_majority7_module_52__and_module_2_res) );
  OR2_X1 u_majority7_module_52__or_module_2_U1 ( .A1(n_majority7_module_52_n2), 
        .A2(n_majority7_module_52_n7), .ZN(
        n_majority7_module_52__or_module_2_res) );
  AND2_X1 u_majority7_module_52__and_module_3_U1 ( .A1(
        n_majority7_module_52_n6), .A2(n_majority7_module_52_n1), .ZN(
        n_majority7_module_52__and_module_3_res) );
  OR2_X1 u_majority7_module_52__or_module_3_U1 ( .A1(n_majority7_module_52_n1), 
        .A2(n_majority7_module_52_n6), .ZN(
        n_majority7_module_52__or_module_3_res) );
  AND2_X1 u_majority7_module_52__and_module_4_U1 ( .A1(
        n_majority7_module_52__and_module_2_res), .A2(
        n_majority7_module_52__and_module_1_res), .ZN(
        n_majority7_module_52__and_module_4_res) );
  OR2_X1 u_majority7_module_52__or_module_4_U1 ( .A1(
        n_majority7_module_52__and_module_1_res), .A2(
        n_majority7_module_52__and_module_2_res), .ZN(
        n_majority7_module_52__or_module_4_res) );
  AND2_X1 u_majority7_module_52__and_module_5_U1 ( .A1(
        n_majority7_module_52__and_module_3_res), .A2(n_majority7_module_52_n3), .ZN(n_majority7_module_52__and_module_5_res) );
  OR2_X1 u_majority7_module_52__or_module_5_U1 ( .A1(n_majority7_module_52_n3), 
        .A2(n_majority7_module_52__and_module_3_res), .ZN(
        n_majority7_module_52__or_module_5_res) );
  AND2_X1 u_majority7_module_52__and_module_6_U1 ( .A1(
        n_majority7_module_52__or_module_1_res), .A2(
        n_majority7_module_52__or_module_2_res), .ZN(
        n_majority7_module_52__and_module_6_res) );
  OR2_X1 u_majority7_module_52__or_module_6_U1 ( .A1(
        n_majority7_module_52__or_module_2_res), .A2(
        n_majority7_module_52__or_module_1_res), .ZN(
        n_majority7_module_52__or_module_6_res) );
  OR2_X1 u_majority7_module_52__or_module_7_U1 ( .A1(
        n_majority7_module_52__and_module_4_res), .A2(
        n_majority7_module_52__and_module_5_res), .ZN(
        n_majority7_module_52__or_module_7_res) );
  AND2_X1 u_majority7_module_52__and_module_7_U1 ( .A1(
        n_majority7_module_52__or_module_3_res), .A2(
        n_majority7_module_52__or_module_4_res), .ZN(
        n_majority7_module_52__and_module_7_res) );
  OR2_X1 u_majority7_module_52__or_module_8_U1 ( .A1(
        n_majority7_module_52__or_module_4_res), .A2(
        n_majority7_module_52__or_module_3_res), .ZN(
        n_majority7_module_52__or_module_8_res) );
  AND2_X1 u_majority7_module_52__and_module_8_U1 ( .A1(
        n_majority7_module_52__or_module_5_res), .A2(
        n_majority7_module_52__and_module_6_res), .ZN(
        n_majority7_module_52__and_module_8_res) );
  OR2_X1 u_majority7_module_52__or_module_9_U1 ( .A1(
        n_majority7_module_52__and_module_6_res), .A2(
        n_majority7_module_52__or_module_5_res), .ZN(
        n_majority7_module_52__or_module_9_res) );
  OR2_X1 u_majority7_module_52__or_module_10_U1 ( .A1(
        n_majority7_module_52__or_module_7_res), .A2(
        n_majority7_module_52__and_module_7_res), .ZN(
        n_majority7_module_52__or_module_10_res) );
  AND2_X1 u_majority7_module_52__and_module_9_U1 ( .A1(
        n_majority7_module_52__or_module_6_res), .A2(
        n_majority7_module_52__or_module_9_res), .ZN(
        n_majority7_module_52__and_module_9_res) );
  OR2_X1 u_majority7_module_52__or_module_11_U1 ( .A1(
        n_majority7_module_52__or_module_10_res), .A2(
        n_majority7_module_52__and_module_8_res), .ZN(
        n_majority7_module_52__or_module_11_res) );
  AND2_X1 u_majority7_module_52__and_module_10_U1 ( .A1(
        n_majority7_module_52__or_module_8_res), .A2(
        n_majority7_module_52__and_module_9_res), .ZN(
        n_majority7_module_52__and_module_10_res) );
  AND2_X1 u_majority7_module_52__and_module_11_U1 ( .A1(
        n_majority7_module_52__and_module_10_res), .A2(
        n_majority7_module_52__or_module_11_res), .ZN(
        n_majority7_module_52_res) );
  DFF_X1 u_reg_module_53__cini_mul_v000_reg ( .D(n_majority7_module_52_res), 
        .CK(clock_3), .Q(n_reg_module_53_res), .QN() );
  BUF_X1 u_majority7_module_53_U7 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_53_n7) );
  BUF_X1 u_majority7_module_53_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_53_n6) );
  BUF_X1 u_majority7_module_53_U5 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_53_n5) );
  BUF_X1 u_majority7_module_53_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_53_n4) );
  BUF_X1 u_majority7_module_53_U3 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_53_n3) );
  BUF_X1 u_majority7_module_53_U2 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_53_n2) );
  BUF_X1 u_majority7_module_53_U1 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_53_n1) );
  AND2_X1 u_majority7_module_53__and_module_1_U1 ( .A1(
        n_majority7_module_53_n5), .A2(n_majority7_module_53_n4), .ZN(
        n_majority7_module_53__and_module_1_res) );
  OR2_X1 u_majority7_module_53__or_module_1_U1 ( .A1(n_majority7_module_53_n4), 
        .A2(n_majority7_module_53_n5), .ZN(
        n_majority7_module_53__or_module_1_res) );
  AND2_X1 u_majority7_module_53__and_module_2_U1 ( .A1(
        n_majority7_module_53_n7), .A2(n_majority7_module_53_n2), .ZN(
        n_majority7_module_53__and_module_2_res) );
  OR2_X1 u_majority7_module_53__or_module_2_U1 ( .A1(n_majority7_module_53_n2), 
        .A2(n_majority7_module_53_n7), .ZN(
        n_majority7_module_53__or_module_2_res) );
  AND2_X1 u_majority7_module_53__and_module_3_U1 ( .A1(
        n_majority7_module_53_n6), .A2(n_majority7_module_53_n1), .ZN(
        n_majority7_module_53__and_module_3_res) );
  OR2_X1 u_majority7_module_53__or_module_3_U1 ( .A1(n_majority7_module_53_n1), 
        .A2(n_majority7_module_53_n6), .ZN(
        n_majority7_module_53__or_module_3_res) );
  AND2_X1 u_majority7_module_53__and_module_4_U1 ( .A1(
        n_majority7_module_53__and_module_2_res), .A2(
        n_majority7_module_53__and_module_1_res), .ZN(
        n_majority7_module_53__and_module_4_res) );
  OR2_X1 u_majority7_module_53__or_module_4_U1 ( .A1(
        n_majority7_module_53__and_module_1_res), .A2(
        n_majority7_module_53__and_module_2_res), .ZN(
        n_majority7_module_53__or_module_4_res) );
  AND2_X1 u_majority7_module_53__and_module_5_U1 ( .A1(
        n_majority7_module_53__and_module_3_res), .A2(n_majority7_module_53_n3), .ZN(n_majority7_module_53__and_module_5_res) );
  OR2_X1 u_majority7_module_53__or_module_5_U1 ( .A1(n_majority7_module_53_n3), 
        .A2(n_majority7_module_53__and_module_3_res), .ZN(
        n_majority7_module_53__or_module_5_res) );
  AND2_X1 u_majority7_module_53__and_module_6_U1 ( .A1(
        n_majority7_module_53__or_module_1_res), .A2(
        n_majority7_module_53__or_module_2_res), .ZN(
        n_majority7_module_53__and_module_6_res) );
  OR2_X1 u_majority7_module_53__or_module_6_U1 ( .A1(
        n_majority7_module_53__or_module_2_res), .A2(
        n_majority7_module_53__or_module_1_res), .ZN(
        n_majority7_module_53__or_module_6_res) );
  OR2_X1 u_majority7_module_53__or_module_7_U1 ( .A1(
        n_majority7_module_53__and_module_4_res), .A2(
        n_majority7_module_53__and_module_5_res), .ZN(
        n_majority7_module_53__or_module_7_res) );
  AND2_X1 u_majority7_module_53__and_module_7_U1 ( .A1(
        n_majority7_module_53__or_module_3_res), .A2(
        n_majority7_module_53__or_module_4_res), .ZN(
        n_majority7_module_53__and_module_7_res) );
  OR2_X1 u_majority7_module_53__or_module_8_U1 ( .A1(
        n_majority7_module_53__or_module_4_res), .A2(
        n_majority7_module_53__or_module_3_res), .ZN(
        n_majority7_module_53__or_module_8_res) );
  AND2_X1 u_majority7_module_53__and_module_8_U1 ( .A1(
        n_majority7_module_53__or_module_5_res), .A2(
        n_majority7_module_53__and_module_6_res), .ZN(
        n_majority7_module_53__and_module_8_res) );
  OR2_X1 u_majority7_module_53__or_module_9_U1 ( .A1(
        n_majority7_module_53__and_module_6_res), .A2(
        n_majority7_module_53__or_module_5_res), .ZN(
        n_majority7_module_53__or_module_9_res) );
  OR2_X1 u_majority7_module_53__or_module_10_U1 ( .A1(
        n_majority7_module_53__or_module_7_res), .A2(
        n_majority7_module_53__and_module_7_res), .ZN(
        n_majority7_module_53__or_module_10_res) );
  AND2_X1 u_majority7_module_53__and_module_9_U1 ( .A1(
        n_majority7_module_53__or_module_6_res), .A2(
        n_majority7_module_53__or_module_9_res), .ZN(
        n_majority7_module_53__and_module_9_res) );
  OR2_X1 u_majority7_module_53__or_module_11_U1 ( .A1(
        n_majority7_module_53__or_module_10_res), .A2(
        n_majority7_module_53__and_module_8_res), .ZN(
        n_majority7_module_53__or_module_11_res) );
  AND2_X1 u_majority7_module_53__and_module_10_U1 ( .A1(
        n_majority7_module_53__or_module_8_res), .A2(
        n_majority7_module_53__and_module_9_res), .ZN(
        n_majority7_module_53__and_module_10_res) );
  AND2_X1 u_majority7_module_53__and_module_11_U1 ( .A1(
        n_majority7_module_53__and_module_10_res), .A2(
        n_majority7_module_53__or_module_11_res), .ZN(
        n_majority7_module_53_res) );
  DFF_X1 u_reg_module_54__cini_mul_v000_reg ( .D(n_majority7_module_53_res), 
        .CK(clock_3), .Q(n_reg_module_54_res), .QN() );
  BUF_X1 u_majority7_module_54_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_54_n7) );
  BUF_X1 u_majority7_module_54_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_54_n6) );
  BUF_X1 u_majority7_module_54_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_54_n5) );
  BUF_X1 u_majority7_module_54_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_54_n4) );
  BUF_X1 u_majority7_module_54_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_54_n3) );
  BUF_X1 u_majority7_module_54_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_54_n2) );
  BUF_X1 u_majority7_module_54_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_54_n1) );
  AND2_X1 u_majority7_module_54__and_module_1_U1 ( .A1(
        n_majority7_module_54_n7), .A2(n_majority7_module_54_n1), .ZN(
        n_majority7_module_54__and_module_1_res) );
  OR2_X1 u_majority7_module_54__or_module_1_U1 ( .A1(n_majority7_module_54_n1), 
        .A2(n_majority7_module_54_n7), .ZN(
        n_majority7_module_54__or_module_1_res) );
  AND2_X1 u_majority7_module_54__and_module_2_U1 ( .A1(
        n_majority7_module_54_n5), .A2(n_majority7_module_54_n3), .ZN(
        n_majority7_module_54__and_module_2_res) );
  OR2_X1 u_majority7_module_54__or_module_2_U1 ( .A1(n_majority7_module_54_n3), 
        .A2(n_majority7_module_54_n5), .ZN(
        n_majority7_module_54__or_module_2_res) );
  AND2_X1 u_majority7_module_54__and_module_3_U1 ( .A1(
        n_majority7_module_54_n6), .A2(n_majority7_module_54_n4), .ZN(
        n_majority7_module_54__and_module_3_res) );
  OR2_X1 u_majority7_module_54__or_module_3_U1 ( .A1(n_majority7_module_54_n4), 
        .A2(n_majority7_module_54_n6), .ZN(
        n_majority7_module_54__or_module_3_res) );
  AND2_X1 u_majority7_module_54__and_module_4_U1 ( .A1(
        n_majority7_module_54__and_module_2_res), .A2(
        n_majority7_module_54__and_module_1_res), .ZN(
        n_majority7_module_54__and_module_4_res) );
  OR2_X1 u_majority7_module_54__or_module_4_U1 ( .A1(
        n_majority7_module_54__and_module_1_res), .A2(
        n_majority7_module_54__and_module_2_res), .ZN(
        n_majority7_module_54__or_module_4_res) );
  AND2_X1 u_majority7_module_54__and_module_5_U1 ( .A1(
        n_majority7_module_54__and_module_3_res), .A2(n_majority7_module_54_n2), .ZN(n_majority7_module_54__and_module_5_res) );
  OR2_X1 u_majority7_module_54__or_module_5_U1 ( .A1(n_majority7_module_54_n2), 
        .A2(n_majority7_module_54__and_module_3_res), .ZN(
        n_majority7_module_54__or_module_5_res) );
  AND2_X1 u_majority7_module_54__and_module_6_U1 ( .A1(
        n_majority7_module_54__or_module_1_res), .A2(
        n_majority7_module_54__or_module_2_res), .ZN(
        n_majority7_module_54__and_module_6_res) );
  OR2_X1 u_majority7_module_54__or_module_6_U1 ( .A1(
        n_majority7_module_54__or_module_2_res), .A2(
        n_majority7_module_54__or_module_1_res), .ZN(
        n_majority7_module_54__or_module_6_res) );
  OR2_X1 u_majority7_module_54__or_module_7_U1 ( .A1(
        n_majority7_module_54__and_module_4_res), .A2(
        n_majority7_module_54__and_module_5_res), .ZN(
        n_majority7_module_54__or_module_7_res) );
  AND2_X1 u_majority7_module_54__and_module_7_U1 ( .A1(
        n_majority7_module_54__or_module_3_res), .A2(
        n_majority7_module_54__or_module_4_res), .ZN(
        n_majority7_module_54__and_module_7_res) );
  OR2_X1 u_majority7_module_54__or_module_8_U1 ( .A1(
        n_majority7_module_54__or_module_4_res), .A2(
        n_majority7_module_54__or_module_3_res), .ZN(
        n_majority7_module_54__or_module_8_res) );
  AND2_X1 u_majority7_module_54__and_module_8_U1 ( .A1(
        n_majority7_module_54__or_module_5_res), .A2(
        n_majority7_module_54__and_module_6_res), .ZN(
        n_majority7_module_54__and_module_8_res) );
  OR2_X1 u_majority7_module_54__or_module_9_U1 ( .A1(
        n_majority7_module_54__and_module_6_res), .A2(
        n_majority7_module_54__or_module_5_res), .ZN(
        n_majority7_module_54__or_module_9_res) );
  OR2_X1 u_majority7_module_54__or_module_10_U1 ( .A1(
        n_majority7_module_54__or_module_7_res), .A2(
        n_majority7_module_54__and_module_7_res), .ZN(
        n_majority7_module_54__or_module_10_res) );
  AND2_X1 u_majority7_module_54__and_module_9_U1 ( .A1(
        n_majority7_module_54__or_module_6_res), .A2(
        n_majority7_module_54__or_module_9_res), .ZN(
        n_majority7_module_54__and_module_9_res) );
  OR2_X1 u_majority7_module_54__or_module_11_U1 ( .A1(
        n_majority7_module_54__or_module_10_res), .A2(
        n_majority7_module_54__and_module_8_res), .ZN(
        n_majority7_module_54__or_module_11_res) );
  AND2_X1 u_majority7_module_54__and_module_10_U1 ( .A1(
        n_majority7_module_54__or_module_8_res), .A2(
        n_majority7_module_54__and_module_9_res), .ZN(
        n_majority7_module_54__and_module_10_res) );
  AND2_X1 u_majority7_module_54__and_module_11_U1 ( .A1(
        n_majority7_module_54__and_module_10_res), .A2(
        n_majority7_module_54__or_module_11_res), .ZN(
        n_majority7_module_54_res) );
  DFF_X1 u_reg_module_55__cini_mul_v000_reg ( .D(n_majority7_module_54_res), 
        .CK(clock_3), .Q(n_reg_module_55_res), .QN() );
  BUF_X1 u_majority7_module_55_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_55_n7) );
  BUF_X1 u_majority7_module_55_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_55_n6) );
  BUF_X1 u_majority7_module_55_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_55_n5) );
  BUF_X1 u_majority7_module_55_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_55_n4) );
  BUF_X1 u_majority7_module_55_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_55_n3) );
  BUF_X1 u_majority7_module_55_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_55_n2) );
  BUF_X1 u_majority7_module_55_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_55_n1) );
  AND2_X1 u_majority7_module_55__and_module_1_U1 ( .A1(
        n_majority7_module_55_n7), .A2(n_majority7_module_55_n1), .ZN(
        n_majority7_module_55__and_module_1_res) );
  OR2_X1 u_majority7_module_55__or_module_1_U1 ( .A1(n_majority7_module_55_n1), 
        .A2(n_majority7_module_55_n7), .ZN(
        n_majority7_module_55__or_module_1_res) );
  AND2_X1 u_majority7_module_55__and_module_2_U1 ( .A1(
        n_majority7_module_55_n5), .A2(n_majority7_module_55_n3), .ZN(
        n_majority7_module_55__and_module_2_res) );
  OR2_X1 u_majority7_module_55__or_module_2_U1 ( .A1(n_majority7_module_55_n3), 
        .A2(n_majority7_module_55_n5), .ZN(
        n_majority7_module_55__or_module_2_res) );
  AND2_X1 u_majority7_module_55__and_module_3_U1 ( .A1(
        n_majority7_module_55_n6), .A2(n_majority7_module_55_n4), .ZN(
        n_majority7_module_55__and_module_3_res) );
  OR2_X1 u_majority7_module_55__or_module_3_U1 ( .A1(n_majority7_module_55_n4), 
        .A2(n_majority7_module_55_n6), .ZN(
        n_majority7_module_55__or_module_3_res) );
  AND2_X1 u_majority7_module_55__and_module_4_U1 ( .A1(
        n_majority7_module_55__and_module_2_res), .A2(
        n_majority7_module_55__and_module_1_res), .ZN(
        n_majority7_module_55__and_module_4_res) );
  OR2_X1 u_majority7_module_55__or_module_4_U1 ( .A1(
        n_majority7_module_55__and_module_1_res), .A2(
        n_majority7_module_55__and_module_2_res), .ZN(
        n_majority7_module_55__or_module_4_res) );
  AND2_X1 u_majority7_module_55__and_module_5_U1 ( .A1(
        n_majority7_module_55__and_module_3_res), .A2(n_majority7_module_55_n2), .ZN(n_majority7_module_55__and_module_5_res) );
  OR2_X1 u_majority7_module_55__or_module_5_U1 ( .A1(n_majority7_module_55_n2), 
        .A2(n_majority7_module_55__and_module_3_res), .ZN(
        n_majority7_module_55__or_module_5_res) );
  AND2_X1 u_majority7_module_55__and_module_6_U1 ( .A1(
        n_majority7_module_55__or_module_1_res), .A2(
        n_majority7_module_55__or_module_2_res), .ZN(
        n_majority7_module_55__and_module_6_res) );
  OR2_X1 u_majority7_module_55__or_module_6_U1 ( .A1(
        n_majority7_module_55__or_module_2_res), .A2(
        n_majority7_module_55__or_module_1_res), .ZN(
        n_majority7_module_55__or_module_6_res) );
  OR2_X1 u_majority7_module_55__or_module_7_U1 ( .A1(
        n_majority7_module_55__and_module_4_res), .A2(
        n_majority7_module_55__and_module_5_res), .ZN(
        n_majority7_module_55__or_module_7_res) );
  AND2_X1 u_majority7_module_55__and_module_7_U1 ( .A1(
        n_majority7_module_55__or_module_3_res), .A2(
        n_majority7_module_55__or_module_4_res), .ZN(
        n_majority7_module_55__and_module_7_res) );
  OR2_X1 u_majority7_module_55__or_module_8_U1 ( .A1(
        n_majority7_module_55__or_module_4_res), .A2(
        n_majority7_module_55__or_module_3_res), .ZN(
        n_majority7_module_55__or_module_8_res) );
  AND2_X1 u_majority7_module_55__and_module_8_U1 ( .A1(
        n_majority7_module_55__or_module_5_res), .A2(
        n_majority7_module_55__and_module_6_res), .ZN(
        n_majority7_module_55__and_module_8_res) );
  OR2_X1 u_majority7_module_55__or_module_9_U1 ( .A1(
        n_majority7_module_55__and_module_6_res), .A2(
        n_majority7_module_55__or_module_5_res), .ZN(
        n_majority7_module_55__or_module_9_res) );
  OR2_X1 u_majority7_module_55__or_module_10_U1 ( .A1(
        n_majority7_module_55__or_module_7_res), .A2(
        n_majority7_module_55__and_module_7_res), .ZN(
        n_majority7_module_55__or_module_10_res) );
  AND2_X1 u_majority7_module_55__and_module_9_U1 ( .A1(
        n_majority7_module_55__or_module_6_res), .A2(
        n_majority7_module_55__or_module_9_res), .ZN(
        n_majority7_module_55__and_module_9_res) );
  OR2_X1 u_majority7_module_55__or_module_11_U1 ( .A1(
        n_majority7_module_55__or_module_10_res), .A2(
        n_majority7_module_55__and_module_8_res), .ZN(
        n_majority7_module_55__or_module_11_res) );
  AND2_X1 u_majority7_module_55__and_module_10_U1 ( .A1(
        n_majority7_module_55__or_module_8_res), .A2(
        n_majority7_module_55__and_module_9_res), .ZN(
        n_majority7_module_55__and_module_10_res) );
  AND2_X1 u_majority7_module_55__and_module_11_U1 ( .A1(
        n_majority7_module_55__and_module_10_res), .A2(
        n_majority7_module_55__or_module_11_res), .ZN(
        n_majority7_module_55_res) );
  DFF_X1 u_reg_module_56__cini_mul_v000_reg ( .D(n_majority7_module_55_res), 
        .CK(clock_3), .Q(n_reg_module_56_res), .QN() );
  BUF_X1 u_majority7_module_56_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_56_n7) );
  BUF_X1 u_majority7_module_56_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_56_n6) );
  BUF_X1 u_majority7_module_56_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_56_n5) );
  BUF_X1 u_majority7_module_56_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_56_n4) );
  BUF_X1 u_majority7_module_56_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_56_n3) );
  BUF_X1 u_majority7_module_56_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_56_n2) );
  BUF_X1 u_majority7_module_56_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_56_n1) );
  AND2_X1 u_majority7_module_56__and_module_1_U1 ( .A1(
        n_majority7_module_56_n5), .A2(n_majority7_module_56_n4), .ZN(
        n_majority7_module_56__and_module_1_res) );
  OR2_X1 u_majority7_module_56__or_module_1_U1 ( .A1(n_majority7_module_56_n4), 
        .A2(n_majority7_module_56_n5), .ZN(
        n_majority7_module_56__or_module_1_res) );
  AND2_X1 u_majority7_module_56__and_module_2_U1 ( .A1(
        n_majority7_module_56_n7), .A2(n_majority7_module_56_n2), .ZN(
        n_majority7_module_56__and_module_2_res) );
  OR2_X1 u_majority7_module_56__or_module_2_U1 ( .A1(n_majority7_module_56_n2), 
        .A2(n_majority7_module_56_n7), .ZN(
        n_majority7_module_56__or_module_2_res) );
  AND2_X1 u_majority7_module_56__and_module_3_U1 ( .A1(
        n_majority7_module_56_n6), .A2(n_majority7_module_56_n1), .ZN(
        n_majority7_module_56__and_module_3_res) );
  OR2_X1 u_majority7_module_56__or_module_3_U1 ( .A1(n_majority7_module_56_n1), 
        .A2(n_majority7_module_56_n6), .ZN(
        n_majority7_module_56__or_module_3_res) );
  AND2_X1 u_majority7_module_56__and_module_4_U1 ( .A1(
        n_majority7_module_56__and_module_2_res), .A2(
        n_majority7_module_56__and_module_1_res), .ZN(
        n_majority7_module_56__and_module_4_res) );
  OR2_X1 u_majority7_module_56__or_module_4_U1 ( .A1(
        n_majority7_module_56__and_module_1_res), .A2(
        n_majority7_module_56__and_module_2_res), .ZN(
        n_majority7_module_56__or_module_4_res) );
  AND2_X1 u_majority7_module_56__and_module_5_U1 ( .A1(
        n_majority7_module_56__and_module_3_res), .A2(n_majority7_module_56_n3), .ZN(n_majority7_module_56__and_module_5_res) );
  OR2_X1 u_majority7_module_56__or_module_5_U1 ( .A1(n_majority7_module_56_n3), 
        .A2(n_majority7_module_56__and_module_3_res), .ZN(
        n_majority7_module_56__or_module_5_res) );
  AND2_X1 u_majority7_module_56__and_module_6_U1 ( .A1(
        n_majority7_module_56__or_module_1_res), .A2(
        n_majority7_module_56__or_module_2_res), .ZN(
        n_majority7_module_56__and_module_6_res) );
  OR2_X1 u_majority7_module_56__or_module_6_U1 ( .A1(
        n_majority7_module_56__or_module_2_res), .A2(
        n_majority7_module_56__or_module_1_res), .ZN(
        n_majority7_module_56__or_module_6_res) );
  OR2_X1 u_majority7_module_56__or_module_7_U1 ( .A1(
        n_majority7_module_56__and_module_4_res), .A2(
        n_majority7_module_56__and_module_5_res), .ZN(
        n_majority7_module_56__or_module_7_res) );
  AND2_X1 u_majority7_module_56__and_module_7_U1 ( .A1(
        n_majority7_module_56__or_module_3_res), .A2(
        n_majority7_module_56__or_module_4_res), .ZN(
        n_majority7_module_56__and_module_7_res) );
  OR2_X1 u_majority7_module_56__or_module_8_U1 ( .A1(
        n_majority7_module_56__or_module_4_res), .A2(
        n_majority7_module_56__or_module_3_res), .ZN(
        n_majority7_module_56__or_module_8_res) );
  AND2_X1 u_majority7_module_56__and_module_8_U1 ( .A1(
        n_majority7_module_56__or_module_5_res), .A2(
        n_majority7_module_56__and_module_6_res), .ZN(
        n_majority7_module_56__and_module_8_res) );
  OR2_X1 u_majority7_module_56__or_module_9_U1 ( .A1(
        n_majority7_module_56__and_module_6_res), .A2(
        n_majority7_module_56__or_module_5_res), .ZN(
        n_majority7_module_56__or_module_9_res) );
  OR2_X1 u_majority7_module_56__or_module_10_U1 ( .A1(
        n_majority7_module_56__or_module_7_res), .A2(
        n_majority7_module_56__and_module_7_res), .ZN(
        n_majority7_module_56__or_module_10_res) );
  AND2_X1 u_majority7_module_56__and_module_9_U1 ( .A1(
        n_majority7_module_56__or_module_6_res), .A2(
        n_majority7_module_56__or_module_9_res), .ZN(
        n_majority7_module_56__and_module_9_res) );
  OR2_X1 u_majority7_module_56__or_module_11_U1 ( .A1(
        n_majority7_module_56__or_module_10_res), .A2(
        n_majority7_module_56__and_module_8_res), .ZN(
        n_majority7_module_56__or_module_11_res) );
  AND2_X1 u_majority7_module_56__and_module_10_U1 ( .A1(
        n_majority7_module_56__or_module_8_res), .A2(
        n_majority7_module_56__and_module_9_res), .ZN(
        n_majority7_module_56__and_module_10_res) );
  AND2_X1 u_majority7_module_56__and_module_11_U1 ( .A1(
        n_majority7_module_56__and_module_10_res), .A2(
        n_majority7_module_56__or_module_11_res), .ZN(
        n_majority7_module_56_res) );
  DFF_X1 u_reg_module_57__cini_mul_v000_reg ( .D(n_majority7_module_56_res), 
        .CK(clock_3), .Q(n_reg_module_57_res), .QN() );
  BUF_X1 u_majority7_module_57_U7 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_57_n7) );
  BUF_X1 u_majority7_module_57_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_57_n6) );
  BUF_X1 u_majority7_module_57_U5 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_57_n5) );
  BUF_X1 u_majority7_module_57_U4 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_57_n4) );
  BUF_X1 u_majority7_module_57_U3 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_57_n3) );
  BUF_X1 u_majority7_module_57_U2 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_57_n2) );
  BUF_X1 u_majority7_module_57_U1 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_57_n1) );
  AND2_X1 u_majority7_module_57__and_module_1_U1 ( .A1(
        n_majority7_module_57_n5), .A2(n_majority7_module_57_n4), .ZN(
        n_majority7_module_57__and_module_1_res) );
  OR2_X1 u_majority7_module_57__or_module_1_U1 ( .A1(n_majority7_module_57_n4), 
        .A2(n_majority7_module_57_n5), .ZN(
        n_majority7_module_57__or_module_1_res) );
  AND2_X1 u_majority7_module_57__and_module_2_U1 ( .A1(
        n_majority7_module_57_n7), .A2(n_majority7_module_57_n2), .ZN(
        n_majority7_module_57__and_module_2_res) );
  OR2_X1 u_majority7_module_57__or_module_2_U1 ( .A1(n_majority7_module_57_n2), 
        .A2(n_majority7_module_57_n7), .ZN(
        n_majority7_module_57__or_module_2_res) );
  AND2_X1 u_majority7_module_57__and_module_3_U1 ( .A1(
        n_majority7_module_57_n6), .A2(n_majority7_module_57_n1), .ZN(
        n_majority7_module_57__and_module_3_res) );
  OR2_X1 u_majority7_module_57__or_module_3_U1 ( .A1(n_majority7_module_57_n1), 
        .A2(n_majority7_module_57_n6), .ZN(
        n_majority7_module_57__or_module_3_res) );
  AND2_X1 u_majority7_module_57__and_module_4_U1 ( .A1(
        n_majority7_module_57__and_module_2_res), .A2(
        n_majority7_module_57__and_module_1_res), .ZN(
        n_majority7_module_57__and_module_4_res) );
  OR2_X1 u_majority7_module_57__or_module_4_U1 ( .A1(
        n_majority7_module_57__and_module_1_res), .A2(
        n_majority7_module_57__and_module_2_res), .ZN(
        n_majority7_module_57__or_module_4_res) );
  AND2_X1 u_majority7_module_57__and_module_5_U1 ( .A1(
        n_majority7_module_57__and_module_3_res), .A2(n_majority7_module_57_n3), .ZN(n_majority7_module_57__and_module_5_res) );
  OR2_X1 u_majority7_module_57__or_module_5_U1 ( .A1(n_majority7_module_57_n3), 
        .A2(n_majority7_module_57__and_module_3_res), .ZN(
        n_majority7_module_57__or_module_5_res) );
  AND2_X1 u_majority7_module_57__and_module_6_U1 ( .A1(
        n_majority7_module_57__or_module_1_res), .A2(
        n_majority7_module_57__or_module_2_res), .ZN(
        n_majority7_module_57__and_module_6_res) );
  OR2_X1 u_majority7_module_57__or_module_6_U1 ( .A1(
        n_majority7_module_57__or_module_2_res), .A2(
        n_majority7_module_57__or_module_1_res), .ZN(
        n_majority7_module_57__or_module_6_res) );
  OR2_X1 u_majority7_module_57__or_module_7_U1 ( .A1(
        n_majority7_module_57__and_module_4_res), .A2(
        n_majority7_module_57__and_module_5_res), .ZN(
        n_majority7_module_57__or_module_7_res) );
  AND2_X1 u_majority7_module_57__and_module_7_U1 ( .A1(
        n_majority7_module_57__or_module_3_res), .A2(
        n_majority7_module_57__or_module_4_res), .ZN(
        n_majority7_module_57__and_module_7_res) );
  OR2_X1 u_majority7_module_57__or_module_8_U1 ( .A1(
        n_majority7_module_57__or_module_4_res), .A2(
        n_majority7_module_57__or_module_3_res), .ZN(
        n_majority7_module_57__or_module_8_res) );
  AND2_X1 u_majority7_module_57__and_module_8_U1 ( .A1(
        n_majority7_module_57__or_module_5_res), .A2(
        n_majority7_module_57__and_module_6_res), .ZN(
        n_majority7_module_57__and_module_8_res) );
  OR2_X1 u_majority7_module_57__or_module_9_U1 ( .A1(
        n_majority7_module_57__and_module_6_res), .A2(
        n_majority7_module_57__or_module_5_res), .ZN(
        n_majority7_module_57__or_module_9_res) );
  OR2_X1 u_majority7_module_57__or_module_10_U1 ( .A1(
        n_majority7_module_57__or_module_7_res), .A2(
        n_majority7_module_57__and_module_7_res), .ZN(
        n_majority7_module_57__or_module_10_res) );
  AND2_X1 u_majority7_module_57__and_module_9_U1 ( .A1(
        n_majority7_module_57__or_module_6_res), .A2(
        n_majority7_module_57__or_module_9_res), .ZN(
        n_majority7_module_57__and_module_9_res) );
  OR2_X1 u_majority7_module_57__or_module_11_U1 ( .A1(
        n_majority7_module_57__or_module_10_res), .A2(
        n_majority7_module_57__and_module_8_res), .ZN(
        n_majority7_module_57__or_module_11_res) );
  AND2_X1 u_majority7_module_57__and_module_10_U1 ( .A1(
        n_majority7_module_57__or_module_8_res), .A2(
        n_majority7_module_57__and_module_9_res), .ZN(
        n_majority7_module_57__and_module_10_res) );
  AND2_X1 u_majority7_module_57__and_module_11_U1 ( .A1(
        n_majority7_module_57__and_module_10_res), .A2(
        n_majority7_module_57__or_module_11_res), .ZN(
        n_majority7_module_57_res) );
  DFF_X1 u_reg_module_58__cini_mul_v000_reg ( .D(n_majority7_module_57_res), 
        .CK(clock_3), .Q(n_reg_module_58_res), .QN() );
  BUF_X1 u_majority7_module_58_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_58_n7) );
  BUF_X1 u_majority7_module_58_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_58_n6) );
  BUF_X1 u_majority7_module_58_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_58_n5) );
  BUF_X1 u_majority7_module_58_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_58_n4) );
  BUF_X1 u_majority7_module_58_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_58_n3) );
  BUF_X1 u_majority7_module_58_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_58_n2) );
  BUF_X1 u_majority7_module_58_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_58_n1) );
  AND2_X1 u_majority7_module_58__and_module_1_U1 ( .A1(
        n_majority7_module_58_n7), .A2(n_majority7_module_58_n1), .ZN(
        n_majority7_module_58__and_module_1_res) );
  OR2_X1 u_majority7_module_58__or_module_1_U1 ( .A1(n_majority7_module_58_n1), 
        .A2(n_majority7_module_58_n7), .ZN(
        n_majority7_module_58__or_module_1_res) );
  AND2_X1 u_majority7_module_58__and_module_2_U1 ( .A1(
        n_majority7_module_58_n5), .A2(n_majority7_module_58_n3), .ZN(
        n_majority7_module_58__and_module_2_res) );
  OR2_X1 u_majority7_module_58__or_module_2_U1 ( .A1(n_majority7_module_58_n3), 
        .A2(n_majority7_module_58_n5), .ZN(
        n_majority7_module_58__or_module_2_res) );
  AND2_X1 u_majority7_module_58__and_module_3_U1 ( .A1(
        n_majority7_module_58_n6), .A2(n_majority7_module_58_n4), .ZN(
        n_majority7_module_58__and_module_3_res) );
  OR2_X1 u_majority7_module_58__or_module_3_U1 ( .A1(n_majority7_module_58_n4), 
        .A2(n_majority7_module_58_n6), .ZN(
        n_majority7_module_58__or_module_3_res) );
  AND2_X1 u_majority7_module_58__and_module_4_U1 ( .A1(
        n_majority7_module_58__and_module_2_res), .A2(
        n_majority7_module_58__and_module_1_res), .ZN(
        n_majority7_module_58__and_module_4_res) );
  OR2_X1 u_majority7_module_58__or_module_4_U1 ( .A1(
        n_majority7_module_58__and_module_1_res), .A2(
        n_majority7_module_58__and_module_2_res), .ZN(
        n_majority7_module_58__or_module_4_res) );
  AND2_X1 u_majority7_module_58__and_module_5_U1 ( .A1(
        n_majority7_module_58__and_module_3_res), .A2(n_majority7_module_58_n2), .ZN(n_majority7_module_58__and_module_5_res) );
  OR2_X1 u_majority7_module_58__or_module_5_U1 ( .A1(n_majority7_module_58_n2), 
        .A2(n_majority7_module_58__and_module_3_res), .ZN(
        n_majority7_module_58__or_module_5_res) );
  AND2_X1 u_majority7_module_58__and_module_6_U1 ( .A1(
        n_majority7_module_58__or_module_1_res), .A2(
        n_majority7_module_58__or_module_2_res), .ZN(
        n_majority7_module_58__and_module_6_res) );
  OR2_X1 u_majority7_module_58__or_module_6_U1 ( .A1(
        n_majority7_module_58__or_module_2_res), .A2(
        n_majority7_module_58__or_module_1_res), .ZN(
        n_majority7_module_58__or_module_6_res) );
  OR2_X1 u_majority7_module_58__or_module_7_U1 ( .A1(
        n_majority7_module_58__and_module_4_res), .A2(
        n_majority7_module_58__and_module_5_res), .ZN(
        n_majority7_module_58__or_module_7_res) );
  AND2_X1 u_majority7_module_58__and_module_7_U1 ( .A1(
        n_majority7_module_58__or_module_3_res), .A2(
        n_majority7_module_58__or_module_4_res), .ZN(
        n_majority7_module_58__and_module_7_res) );
  OR2_X1 u_majority7_module_58__or_module_8_U1 ( .A1(
        n_majority7_module_58__or_module_4_res), .A2(
        n_majority7_module_58__or_module_3_res), .ZN(
        n_majority7_module_58__or_module_8_res) );
  AND2_X1 u_majority7_module_58__and_module_8_U1 ( .A1(
        n_majority7_module_58__or_module_5_res), .A2(
        n_majority7_module_58__and_module_6_res), .ZN(
        n_majority7_module_58__and_module_8_res) );
  OR2_X1 u_majority7_module_58__or_module_9_U1 ( .A1(
        n_majority7_module_58__and_module_6_res), .A2(
        n_majority7_module_58__or_module_5_res), .ZN(
        n_majority7_module_58__or_module_9_res) );
  OR2_X1 u_majority7_module_58__or_module_10_U1 ( .A1(
        n_majority7_module_58__or_module_7_res), .A2(
        n_majority7_module_58__and_module_7_res), .ZN(
        n_majority7_module_58__or_module_10_res) );
  AND2_X1 u_majority7_module_58__and_module_9_U1 ( .A1(
        n_majority7_module_58__or_module_6_res), .A2(
        n_majority7_module_58__or_module_9_res), .ZN(
        n_majority7_module_58__and_module_9_res) );
  OR2_X1 u_majority7_module_58__or_module_11_U1 ( .A1(
        n_majority7_module_58__or_module_10_res), .A2(
        n_majority7_module_58__and_module_8_res), .ZN(
        n_majority7_module_58__or_module_11_res) );
  AND2_X1 u_majority7_module_58__and_module_10_U1 ( .A1(
        n_majority7_module_58__or_module_8_res), .A2(
        n_majority7_module_58__and_module_9_res), .ZN(
        n_majority7_module_58__and_module_10_res) );
  AND2_X1 u_majority7_module_58__and_module_11_U1 ( .A1(
        n_majority7_module_58__and_module_10_res), .A2(
        n_majority7_module_58__or_module_11_res), .ZN(
        n_majority7_module_58_res) );
  DFF_X1 u_reg_module_59__cini_mul_v000_reg ( .D(n_majority7_module_58_res), 
        .CK(clock_3), .Q(n_reg_module_59_res), .QN() );
  BUF_X1 u_majority7_module_59_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_59_n7) );
  BUF_X1 u_majority7_module_59_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_59_n6) );
  BUF_X1 u_majority7_module_59_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_59_n5) );
  BUF_X1 u_majority7_module_59_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_59_n4) );
  BUF_X1 u_majority7_module_59_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_59_n3) );
  BUF_X1 u_majority7_module_59_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_59_n2) );
  BUF_X1 u_majority7_module_59_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_59_n1) );
  AND2_X1 u_majority7_module_59__and_module_1_U1 ( .A1(
        n_majority7_module_59_n7), .A2(n_majority7_module_59_n1), .ZN(
        n_majority7_module_59__and_module_1_res) );
  OR2_X1 u_majority7_module_59__or_module_1_U1 ( .A1(n_majority7_module_59_n1), 
        .A2(n_majority7_module_59_n7), .ZN(
        n_majority7_module_59__or_module_1_res) );
  AND2_X1 u_majority7_module_59__and_module_2_U1 ( .A1(
        n_majority7_module_59_n5), .A2(n_majority7_module_59_n3), .ZN(
        n_majority7_module_59__and_module_2_res) );
  OR2_X1 u_majority7_module_59__or_module_2_U1 ( .A1(n_majority7_module_59_n3), 
        .A2(n_majority7_module_59_n5), .ZN(
        n_majority7_module_59__or_module_2_res) );
  AND2_X1 u_majority7_module_59__and_module_3_U1 ( .A1(
        n_majority7_module_59_n6), .A2(n_majority7_module_59_n4), .ZN(
        n_majority7_module_59__and_module_3_res) );
  OR2_X1 u_majority7_module_59__or_module_3_U1 ( .A1(n_majority7_module_59_n4), 
        .A2(n_majority7_module_59_n6), .ZN(
        n_majority7_module_59__or_module_3_res) );
  AND2_X1 u_majority7_module_59__and_module_4_U1 ( .A1(
        n_majority7_module_59__and_module_2_res), .A2(
        n_majority7_module_59__and_module_1_res), .ZN(
        n_majority7_module_59__and_module_4_res) );
  OR2_X1 u_majority7_module_59__or_module_4_U1 ( .A1(
        n_majority7_module_59__and_module_1_res), .A2(
        n_majority7_module_59__and_module_2_res), .ZN(
        n_majority7_module_59__or_module_4_res) );
  AND2_X1 u_majority7_module_59__and_module_5_U1 ( .A1(
        n_majority7_module_59__and_module_3_res), .A2(n_majority7_module_59_n2), .ZN(n_majority7_module_59__and_module_5_res) );
  OR2_X1 u_majority7_module_59__or_module_5_U1 ( .A1(n_majority7_module_59_n2), 
        .A2(n_majority7_module_59__and_module_3_res), .ZN(
        n_majority7_module_59__or_module_5_res) );
  AND2_X1 u_majority7_module_59__and_module_6_U1 ( .A1(
        n_majority7_module_59__or_module_1_res), .A2(
        n_majority7_module_59__or_module_2_res), .ZN(
        n_majority7_module_59__and_module_6_res) );
  OR2_X1 u_majority7_module_59__or_module_6_U1 ( .A1(
        n_majority7_module_59__or_module_2_res), .A2(
        n_majority7_module_59__or_module_1_res), .ZN(
        n_majority7_module_59__or_module_6_res) );
  OR2_X1 u_majority7_module_59__or_module_7_U1 ( .A1(
        n_majority7_module_59__and_module_4_res), .A2(
        n_majority7_module_59__and_module_5_res), .ZN(
        n_majority7_module_59__or_module_7_res) );
  AND2_X1 u_majority7_module_59__and_module_7_U1 ( .A1(
        n_majority7_module_59__or_module_3_res), .A2(
        n_majority7_module_59__or_module_4_res), .ZN(
        n_majority7_module_59__and_module_7_res) );
  OR2_X1 u_majority7_module_59__or_module_8_U1 ( .A1(
        n_majority7_module_59__or_module_4_res), .A2(
        n_majority7_module_59__or_module_3_res), .ZN(
        n_majority7_module_59__or_module_8_res) );
  AND2_X1 u_majority7_module_59__and_module_8_U1 ( .A1(
        n_majority7_module_59__or_module_5_res), .A2(
        n_majority7_module_59__and_module_6_res), .ZN(
        n_majority7_module_59__and_module_8_res) );
  OR2_X1 u_majority7_module_59__or_module_9_U1 ( .A1(
        n_majority7_module_59__and_module_6_res), .A2(
        n_majority7_module_59__or_module_5_res), .ZN(
        n_majority7_module_59__or_module_9_res) );
  OR2_X1 u_majority7_module_59__or_module_10_U1 ( .A1(
        n_majority7_module_59__or_module_7_res), .A2(
        n_majority7_module_59__and_module_7_res), .ZN(
        n_majority7_module_59__or_module_10_res) );
  AND2_X1 u_majority7_module_59__and_module_9_U1 ( .A1(
        n_majority7_module_59__or_module_6_res), .A2(
        n_majority7_module_59__or_module_9_res), .ZN(
        n_majority7_module_59__and_module_9_res) );
  OR2_X1 u_majority7_module_59__or_module_11_U1 ( .A1(
        n_majority7_module_59__or_module_10_res), .A2(
        n_majority7_module_59__and_module_8_res), .ZN(
        n_majority7_module_59__or_module_11_res) );
  AND2_X1 u_majority7_module_59__and_module_10_U1 ( .A1(
        n_majority7_module_59__or_module_8_res), .A2(
        n_majority7_module_59__and_module_9_res), .ZN(
        n_majority7_module_59__and_module_10_res) );
  AND2_X1 u_majority7_module_59__and_module_11_U1 ( .A1(
        n_majority7_module_59__and_module_10_res), .A2(
        n_majority7_module_59__or_module_11_res), .ZN(
        n_majority7_module_59_res) );
  DFF_X1 u_reg_module_60__cini_mul_v000_reg ( .D(n_majority7_module_59_res), 
        .CK(clock_3), .Q(n_reg_module_60_res), .QN() );
  BUF_X1 u_majority7_module_60_U7 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_60_n7) );
  BUF_X1 u_majority7_module_60_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_60_n6) );
  BUF_X1 u_majority7_module_60_U5 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_60_n5) );
  BUF_X1 u_majority7_module_60_U4 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_60_n4) );
  BUF_X1 u_majority7_module_60_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_60_n3) );
  BUF_X1 u_majority7_module_60_U2 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_60_n2) );
  BUF_X1 u_majority7_module_60_U1 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_60_n1) );
  AND2_X1 u_majority7_module_60__and_module_1_U1 ( .A1(
        n_majority7_module_60_n1), .A2(n_majority7_module_60_n5), .ZN(
        n_majority7_module_60__and_module_1_res) );
  OR2_X1 u_majority7_module_60__or_module_1_U1 ( .A1(n_majority7_module_60_n5), 
        .A2(n_majority7_module_60_n1), .ZN(
        n_majority7_module_60__or_module_1_res) );
  AND2_X1 u_majority7_module_60__and_module_2_U1 ( .A1(
        n_majority7_module_60_n7), .A2(n_majority7_module_60_n3), .ZN(
        n_majority7_module_60__and_module_2_res) );
  OR2_X1 u_majority7_module_60__or_module_2_U1 ( .A1(n_majority7_module_60_n3), 
        .A2(n_majority7_module_60_n7), .ZN(
        n_majority7_module_60__or_module_2_res) );
  AND2_X1 u_majority7_module_60__and_module_3_U1 ( .A1(
        n_majority7_module_60_n6), .A2(n_majority7_module_60_n2), .ZN(
        n_majority7_module_60__and_module_3_res) );
  OR2_X1 u_majority7_module_60__or_module_3_U1 ( .A1(n_majority7_module_60_n2), 
        .A2(n_majority7_module_60_n6), .ZN(
        n_majority7_module_60__or_module_3_res) );
  AND2_X1 u_majority7_module_60__and_module_4_U1 ( .A1(
        n_majority7_module_60__and_module_2_res), .A2(
        n_majority7_module_60__and_module_1_res), .ZN(
        n_majority7_module_60__and_module_4_res) );
  OR2_X1 u_majority7_module_60__or_module_4_U1 ( .A1(
        n_majority7_module_60__and_module_1_res), .A2(
        n_majority7_module_60__and_module_2_res), .ZN(
        n_majority7_module_60__or_module_4_res) );
  AND2_X1 u_majority7_module_60__and_module_5_U1 ( .A1(
        n_majority7_module_60__and_module_3_res), .A2(n_majority7_module_60_n4), .ZN(n_majority7_module_60__and_module_5_res) );
  OR2_X1 u_majority7_module_60__or_module_5_U1 ( .A1(n_majority7_module_60_n4), 
        .A2(n_majority7_module_60__and_module_3_res), .ZN(
        n_majority7_module_60__or_module_5_res) );
  AND2_X1 u_majority7_module_60__and_module_6_U1 ( .A1(
        n_majority7_module_60__or_module_1_res), .A2(
        n_majority7_module_60__or_module_2_res), .ZN(
        n_majority7_module_60__and_module_6_res) );
  OR2_X1 u_majority7_module_60__or_module_6_U1 ( .A1(
        n_majority7_module_60__or_module_2_res), .A2(
        n_majority7_module_60__or_module_1_res), .ZN(
        n_majority7_module_60__or_module_6_res) );
  OR2_X1 u_majority7_module_60__or_module_7_U1 ( .A1(
        n_majority7_module_60__and_module_4_res), .A2(
        n_majority7_module_60__and_module_5_res), .ZN(
        n_majority7_module_60__or_module_7_res) );
  AND2_X1 u_majority7_module_60__and_module_7_U1 ( .A1(
        n_majority7_module_60__or_module_3_res), .A2(
        n_majority7_module_60__or_module_4_res), .ZN(
        n_majority7_module_60__and_module_7_res) );
  OR2_X1 u_majority7_module_60__or_module_8_U1 ( .A1(
        n_majority7_module_60__or_module_4_res), .A2(
        n_majority7_module_60__or_module_3_res), .ZN(
        n_majority7_module_60__or_module_8_res) );
  AND2_X1 u_majority7_module_60__and_module_8_U1 ( .A1(
        n_majority7_module_60__or_module_5_res), .A2(
        n_majority7_module_60__and_module_6_res), .ZN(
        n_majority7_module_60__and_module_8_res) );
  OR2_X1 u_majority7_module_60__or_module_9_U1 ( .A1(
        n_majority7_module_60__and_module_6_res), .A2(
        n_majority7_module_60__or_module_5_res), .ZN(
        n_majority7_module_60__or_module_9_res) );
  OR2_X1 u_majority7_module_60__or_module_10_U1 ( .A1(
        n_majority7_module_60__or_module_7_res), .A2(
        n_majority7_module_60__and_module_7_res), .ZN(
        n_majority7_module_60__or_module_10_res) );
  AND2_X1 u_majority7_module_60__and_module_9_U1 ( .A1(
        n_majority7_module_60__or_module_6_res), .A2(
        n_majority7_module_60__or_module_9_res), .ZN(
        n_majority7_module_60__and_module_9_res) );
  OR2_X1 u_majority7_module_60__or_module_11_U1 ( .A1(
        n_majority7_module_60__or_module_10_res), .A2(
        n_majority7_module_60__and_module_8_res), .ZN(
        n_majority7_module_60__or_module_11_res) );
  AND2_X1 u_majority7_module_60__and_module_10_U1 ( .A1(
        n_majority7_module_60__or_module_8_res), .A2(
        n_majority7_module_60__and_module_9_res), .ZN(
        n_majority7_module_60__and_module_10_res) );
  AND2_X1 u_majority7_module_60__and_module_11_U1 ( .A1(
        n_majority7_module_60__and_module_10_res), .A2(
        n_majority7_module_60__or_module_11_res), .ZN(
        n_majority7_module_60_res) );
  DFF_X1 u_reg_module_61__cini_mul_v000_reg ( .D(n_majority7_module_60_res), 
        .CK(clock_3), .Q(n_reg_module_61_res), .QN() );
  BUF_X1 u_majority7_module_61_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_61_n7) );
  BUF_X1 u_majority7_module_61_U6 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_61_n6) );
  BUF_X1 u_majority7_module_61_U5 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_61_n5) );
  BUF_X1 u_majority7_module_61_U4 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_61_n4) );
  BUF_X1 u_majority7_module_61_U3 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_61_n3) );
  BUF_X1 u_majority7_module_61_U2 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_61_n2) );
  BUF_X1 u_majority7_module_61_U1 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_61_n1) );
  AND2_X1 u_majority7_module_61__and_module_1_U1 ( .A1(
        n_majority7_module_61_n7), .A2(n_majority7_module_61_n4), .ZN(
        n_majority7_module_61__and_module_1_res) );
  OR2_X1 u_majority7_module_61__or_module_1_U1 ( .A1(n_majority7_module_61_n4), 
        .A2(n_majority7_module_61_n7), .ZN(
        n_majority7_module_61__or_module_1_res) );
  AND2_X1 u_majority7_module_61__and_module_2_U1 ( .A1(
        n_majority7_module_61_n6), .A2(n_majority7_module_61_n2), .ZN(
        n_majority7_module_61__and_module_2_res) );
  OR2_X1 u_majority7_module_61__or_module_2_U1 ( .A1(n_majority7_module_61_n2), 
        .A2(n_majority7_module_61_n6), .ZN(
        n_majority7_module_61__or_module_2_res) );
  AND2_X1 u_majority7_module_61__and_module_3_U1 ( .A1(
        n_majority7_module_61_n5), .A2(n_majority7_module_61_n1), .ZN(
        n_majority7_module_61__and_module_3_res) );
  OR2_X1 u_majority7_module_61__or_module_3_U1 ( .A1(n_majority7_module_61_n1), 
        .A2(n_majority7_module_61_n5), .ZN(
        n_majority7_module_61__or_module_3_res) );
  AND2_X1 u_majority7_module_61__and_module_4_U1 ( .A1(
        n_majority7_module_61__and_module_2_res), .A2(
        n_majority7_module_61__and_module_1_res), .ZN(
        n_majority7_module_61__and_module_4_res) );
  OR2_X1 u_majority7_module_61__or_module_4_U1 ( .A1(
        n_majority7_module_61__and_module_1_res), .A2(
        n_majority7_module_61__and_module_2_res), .ZN(
        n_majority7_module_61__or_module_4_res) );
  AND2_X1 u_majority7_module_61__and_module_5_U1 ( .A1(
        n_majority7_module_61__and_module_3_res), .A2(n_majority7_module_61_n3), .ZN(n_majority7_module_61__and_module_5_res) );
  OR2_X1 u_majority7_module_61__or_module_5_U1 ( .A1(n_majority7_module_61_n3), 
        .A2(n_majority7_module_61__and_module_3_res), .ZN(
        n_majority7_module_61__or_module_5_res) );
  AND2_X1 u_majority7_module_61__and_module_6_U1 ( .A1(
        n_majority7_module_61__or_module_1_res), .A2(
        n_majority7_module_61__or_module_2_res), .ZN(
        n_majority7_module_61__and_module_6_res) );
  OR2_X1 u_majority7_module_61__or_module_6_U1 ( .A1(
        n_majority7_module_61__or_module_2_res), .A2(
        n_majority7_module_61__or_module_1_res), .ZN(
        n_majority7_module_61__or_module_6_res) );
  OR2_X1 u_majority7_module_61__or_module_7_U1 ( .A1(
        n_majority7_module_61__and_module_4_res), .A2(
        n_majority7_module_61__and_module_5_res), .ZN(
        n_majority7_module_61__or_module_7_res) );
  AND2_X1 u_majority7_module_61__and_module_7_U1 ( .A1(
        n_majority7_module_61__or_module_3_res), .A2(
        n_majority7_module_61__or_module_4_res), .ZN(
        n_majority7_module_61__and_module_7_res) );
  OR2_X1 u_majority7_module_61__or_module_8_U1 ( .A1(
        n_majority7_module_61__or_module_4_res), .A2(
        n_majority7_module_61__or_module_3_res), .ZN(
        n_majority7_module_61__or_module_8_res) );
  AND2_X1 u_majority7_module_61__and_module_8_U1 ( .A1(
        n_majority7_module_61__or_module_5_res), .A2(
        n_majority7_module_61__and_module_6_res), .ZN(
        n_majority7_module_61__and_module_8_res) );
  OR2_X1 u_majority7_module_61__or_module_9_U1 ( .A1(
        n_majority7_module_61__and_module_6_res), .A2(
        n_majority7_module_61__or_module_5_res), .ZN(
        n_majority7_module_61__or_module_9_res) );
  OR2_X1 u_majority7_module_61__or_module_10_U1 ( .A1(
        n_majority7_module_61__or_module_7_res), .A2(
        n_majority7_module_61__and_module_7_res), .ZN(
        n_majority7_module_61__or_module_10_res) );
  AND2_X1 u_majority7_module_61__and_module_9_U1 ( .A1(
        n_majority7_module_61__or_module_6_res), .A2(
        n_majority7_module_61__or_module_9_res), .ZN(
        n_majority7_module_61__and_module_9_res) );
  OR2_X1 u_majority7_module_61__or_module_11_U1 ( .A1(
        n_majority7_module_61__or_module_10_res), .A2(
        n_majority7_module_61__and_module_8_res), .ZN(
        n_majority7_module_61__or_module_11_res) );
  AND2_X1 u_majority7_module_61__and_module_10_U1 ( .A1(
        n_majority7_module_61__or_module_8_res), .A2(
        n_majority7_module_61__and_module_9_res), .ZN(
        n_majority7_module_61__and_module_10_res) );
  AND2_X1 u_majority7_module_61__and_module_11_U1 ( .A1(
        n_majority7_module_61__and_module_10_res), .A2(
        n_majority7_module_61__or_module_11_res), .ZN(
        n_majority7_module_61_res) );
  DFF_X1 u_reg_module_62__cini_mul_v000_reg ( .D(n_majority7_module_61_res), 
        .CK(clock_3), .Q(n_reg_module_62_res), .QN() );
  BUF_X1 u_majority7_module_62_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_62_n7) );
  BUF_X1 u_majority7_module_62_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_62_n6) );
  BUF_X1 u_majority7_module_62_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_62_n5) );
  BUF_X1 u_majority7_module_62_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_62_n4) );
  BUF_X1 u_majority7_module_62_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_62_n3) );
  BUF_X1 u_majority7_module_62_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_62_n2) );
  BUF_X1 u_majority7_module_62_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_62_n1) );
  AND2_X1 u_majority7_module_62__and_module_1_U1 ( .A1(
        n_majority7_module_62_n7), .A2(n_majority7_module_62_n1), .ZN(
        n_majority7_module_62__and_module_1_res) );
  OR2_X1 u_majority7_module_62__or_module_1_U1 ( .A1(n_majority7_module_62_n1), 
        .A2(n_majority7_module_62_n7), .ZN(
        n_majority7_module_62__or_module_1_res) );
  AND2_X1 u_majority7_module_62__and_module_2_U1 ( .A1(
        n_majority7_module_62_n5), .A2(n_majority7_module_62_n3), .ZN(
        n_majority7_module_62__and_module_2_res) );
  OR2_X1 u_majority7_module_62__or_module_2_U1 ( .A1(n_majority7_module_62_n3), 
        .A2(n_majority7_module_62_n5), .ZN(
        n_majority7_module_62__or_module_2_res) );
  AND2_X1 u_majority7_module_62__and_module_3_U1 ( .A1(
        n_majority7_module_62_n6), .A2(n_majority7_module_62_n4), .ZN(
        n_majority7_module_62__and_module_3_res) );
  OR2_X1 u_majority7_module_62__or_module_3_U1 ( .A1(n_majority7_module_62_n4), 
        .A2(n_majority7_module_62_n6), .ZN(
        n_majority7_module_62__or_module_3_res) );
  AND2_X1 u_majority7_module_62__and_module_4_U1 ( .A1(
        n_majority7_module_62__and_module_2_res), .A2(
        n_majority7_module_62__and_module_1_res), .ZN(
        n_majority7_module_62__and_module_4_res) );
  OR2_X1 u_majority7_module_62__or_module_4_U1 ( .A1(
        n_majority7_module_62__and_module_1_res), .A2(
        n_majority7_module_62__and_module_2_res), .ZN(
        n_majority7_module_62__or_module_4_res) );
  AND2_X1 u_majority7_module_62__and_module_5_U1 ( .A1(
        n_majority7_module_62__and_module_3_res), .A2(n_majority7_module_62_n2), .ZN(n_majority7_module_62__and_module_5_res) );
  OR2_X1 u_majority7_module_62__or_module_5_U1 ( .A1(n_majority7_module_62_n2), 
        .A2(n_majority7_module_62__and_module_3_res), .ZN(
        n_majority7_module_62__or_module_5_res) );
  AND2_X1 u_majority7_module_62__and_module_6_U1 ( .A1(
        n_majority7_module_62__or_module_1_res), .A2(
        n_majority7_module_62__or_module_2_res), .ZN(
        n_majority7_module_62__and_module_6_res) );
  OR2_X1 u_majority7_module_62__or_module_6_U1 ( .A1(
        n_majority7_module_62__or_module_2_res), .A2(
        n_majority7_module_62__or_module_1_res), .ZN(
        n_majority7_module_62__or_module_6_res) );
  OR2_X1 u_majority7_module_62__or_module_7_U1 ( .A1(
        n_majority7_module_62__and_module_4_res), .A2(
        n_majority7_module_62__and_module_5_res), .ZN(
        n_majority7_module_62__or_module_7_res) );
  AND2_X1 u_majority7_module_62__and_module_7_U1 ( .A1(
        n_majority7_module_62__or_module_3_res), .A2(
        n_majority7_module_62__or_module_4_res), .ZN(
        n_majority7_module_62__and_module_7_res) );
  OR2_X1 u_majority7_module_62__or_module_8_U1 ( .A1(
        n_majority7_module_62__or_module_4_res), .A2(
        n_majority7_module_62__or_module_3_res), .ZN(
        n_majority7_module_62__or_module_8_res) );
  AND2_X1 u_majority7_module_62__and_module_8_U1 ( .A1(
        n_majority7_module_62__or_module_5_res), .A2(
        n_majority7_module_62__and_module_6_res), .ZN(
        n_majority7_module_62__and_module_8_res) );
  OR2_X1 u_majority7_module_62__or_module_9_U1 ( .A1(
        n_majority7_module_62__and_module_6_res), .A2(
        n_majority7_module_62__or_module_5_res), .ZN(
        n_majority7_module_62__or_module_9_res) );
  OR2_X1 u_majority7_module_62__or_module_10_U1 ( .A1(
        n_majority7_module_62__or_module_7_res), .A2(
        n_majority7_module_62__and_module_7_res), .ZN(
        n_majority7_module_62__or_module_10_res) );
  AND2_X1 u_majority7_module_62__and_module_9_U1 ( .A1(
        n_majority7_module_62__or_module_6_res), .A2(
        n_majority7_module_62__or_module_9_res), .ZN(
        n_majority7_module_62__and_module_9_res) );
  OR2_X1 u_majority7_module_62__or_module_11_U1 ( .A1(
        n_majority7_module_62__or_module_10_res), .A2(
        n_majority7_module_62__and_module_8_res), .ZN(
        n_majority7_module_62__or_module_11_res) );
  AND2_X1 u_majority7_module_62__and_module_10_U1 ( .A1(
        n_majority7_module_62__or_module_8_res), .A2(
        n_majority7_module_62__and_module_9_res), .ZN(
        n_majority7_module_62__and_module_10_res) );
  AND2_X1 u_majority7_module_62__and_module_11_U1 ( .A1(
        n_majority7_module_62__and_module_10_res), .A2(
        n_majority7_module_62__or_module_11_res), .ZN(
        n_majority7_module_62_res) );
  DFF_X1 u_reg_module_63__cini_mul_v000_reg ( .D(n_majority7_module_62_res), 
        .CK(clock_3), .Q(n_reg_module_63_res), .QN() );
  BUF_X1 u_majority7_module_63_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_63_n7) );
  BUF_X1 u_majority7_module_63_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_63_n6) );
  BUF_X1 u_majority7_module_63_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_63_n5) );
  BUF_X1 u_majority7_module_63_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_63_n4) );
  BUF_X1 u_majority7_module_63_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_63_n3) );
  BUF_X1 u_majority7_module_63_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_63_n2) );
  BUF_X1 u_majority7_module_63_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_63_n1) );
  AND2_X1 u_majority7_module_63__and_module_1_U1 ( .A1(
        n_majority7_module_63_n7), .A2(n_majority7_module_63_n1), .ZN(
        n_majority7_module_63__and_module_1_res) );
  OR2_X1 u_majority7_module_63__or_module_1_U1 ( .A1(n_majority7_module_63_n1), 
        .A2(n_majority7_module_63_n7), .ZN(
        n_majority7_module_63__or_module_1_res) );
  AND2_X1 u_majority7_module_63__and_module_2_U1 ( .A1(
        n_majority7_module_63_n5), .A2(n_majority7_module_63_n3), .ZN(
        n_majority7_module_63__and_module_2_res) );
  OR2_X1 u_majority7_module_63__or_module_2_U1 ( .A1(n_majority7_module_63_n3), 
        .A2(n_majority7_module_63_n5), .ZN(
        n_majority7_module_63__or_module_2_res) );
  AND2_X1 u_majority7_module_63__and_module_3_U1 ( .A1(
        n_majority7_module_63_n6), .A2(n_majority7_module_63_n4), .ZN(
        n_majority7_module_63__and_module_3_res) );
  OR2_X1 u_majority7_module_63__or_module_3_U1 ( .A1(n_majority7_module_63_n4), 
        .A2(n_majority7_module_63_n6), .ZN(
        n_majority7_module_63__or_module_3_res) );
  AND2_X1 u_majority7_module_63__and_module_4_U1 ( .A1(
        n_majority7_module_63__and_module_2_res), .A2(
        n_majority7_module_63__and_module_1_res), .ZN(
        n_majority7_module_63__and_module_4_res) );
  OR2_X1 u_majority7_module_63__or_module_4_U1 ( .A1(
        n_majority7_module_63__and_module_1_res), .A2(
        n_majority7_module_63__and_module_2_res), .ZN(
        n_majority7_module_63__or_module_4_res) );
  AND2_X1 u_majority7_module_63__and_module_5_U1 ( .A1(
        n_majority7_module_63__and_module_3_res), .A2(n_majority7_module_63_n2), .ZN(n_majority7_module_63__and_module_5_res) );
  OR2_X1 u_majority7_module_63__or_module_5_U1 ( .A1(n_majority7_module_63_n2), 
        .A2(n_majority7_module_63__and_module_3_res), .ZN(
        n_majority7_module_63__or_module_5_res) );
  AND2_X1 u_majority7_module_63__and_module_6_U1 ( .A1(
        n_majority7_module_63__or_module_1_res), .A2(
        n_majority7_module_63__or_module_2_res), .ZN(
        n_majority7_module_63__and_module_6_res) );
  OR2_X1 u_majority7_module_63__or_module_6_U1 ( .A1(
        n_majority7_module_63__or_module_2_res), .A2(
        n_majority7_module_63__or_module_1_res), .ZN(
        n_majority7_module_63__or_module_6_res) );
  OR2_X1 u_majority7_module_63__or_module_7_U1 ( .A1(
        n_majority7_module_63__and_module_4_res), .A2(
        n_majority7_module_63__and_module_5_res), .ZN(
        n_majority7_module_63__or_module_7_res) );
  AND2_X1 u_majority7_module_63__and_module_7_U1 ( .A1(
        n_majority7_module_63__or_module_3_res), .A2(
        n_majority7_module_63__or_module_4_res), .ZN(
        n_majority7_module_63__and_module_7_res) );
  OR2_X1 u_majority7_module_63__or_module_8_U1 ( .A1(
        n_majority7_module_63__or_module_4_res), .A2(
        n_majority7_module_63__or_module_3_res), .ZN(
        n_majority7_module_63__or_module_8_res) );
  AND2_X1 u_majority7_module_63__and_module_8_U1 ( .A1(
        n_majority7_module_63__or_module_5_res), .A2(
        n_majority7_module_63__and_module_6_res), .ZN(
        n_majority7_module_63__and_module_8_res) );
  OR2_X1 u_majority7_module_63__or_module_9_U1 ( .A1(
        n_majority7_module_63__and_module_6_res), .A2(
        n_majority7_module_63__or_module_5_res), .ZN(
        n_majority7_module_63__or_module_9_res) );
  OR2_X1 u_majority7_module_63__or_module_10_U1 ( .A1(
        n_majority7_module_63__or_module_7_res), .A2(
        n_majority7_module_63__and_module_7_res), .ZN(
        n_majority7_module_63__or_module_10_res) );
  AND2_X1 u_majority7_module_63__and_module_9_U1 ( .A1(
        n_majority7_module_63__or_module_6_res), .A2(
        n_majority7_module_63__or_module_9_res), .ZN(
        n_majority7_module_63__and_module_9_res) );
  OR2_X1 u_majority7_module_63__or_module_11_U1 ( .A1(
        n_majority7_module_63__or_module_10_res), .A2(
        n_majority7_module_63__and_module_8_res), .ZN(
        n_majority7_module_63__or_module_11_res) );
  AND2_X1 u_majority7_module_63__and_module_10_U1 ( .A1(
        n_majority7_module_63__or_module_8_res), .A2(
        n_majority7_module_63__and_module_9_res), .ZN(
        n_majority7_module_63__and_module_10_res) );
  AND2_X1 u_majority7_module_63__and_module_11_U1 ( .A1(
        n_majority7_module_63__and_module_10_res), .A2(
        n_majority7_module_63__or_module_11_res), .ZN(
        n_majority7_module_63_res) );
  DFF_X1 u_reg_module_64__cini_mul_v000_reg ( .D(n_majority7_module_63_res), 
        .CK(clock_3), .Q(n_reg_module_64_res), .QN() );
  BUF_X1 u_majority7_module_64_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_64_n7) );
  BUF_X1 u_majority7_module_64_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_64_n6) );
  BUF_X1 u_majority7_module_64_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_64_n5) );
  BUF_X1 u_majority7_module_64_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_64_n4) );
  BUF_X1 u_majority7_module_64_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_64_n3) );
  BUF_X1 u_majority7_module_64_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_64_n2) );
  BUF_X1 u_majority7_module_64_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_64_n1) );
  AND2_X1 u_majority7_module_64__and_module_1_U1 ( .A1(
        n_majority7_module_64_n7), .A2(n_majority7_module_64_n1), .ZN(
        n_majority7_module_64__and_module_1_res) );
  OR2_X1 u_majority7_module_64__or_module_1_U1 ( .A1(n_majority7_module_64_n1), 
        .A2(n_majority7_module_64_n7), .ZN(
        n_majority7_module_64__or_module_1_res) );
  AND2_X1 u_majority7_module_64__and_module_2_U1 ( .A1(
        n_majority7_module_64_n5), .A2(n_majority7_module_64_n3), .ZN(
        n_majority7_module_64__and_module_2_res) );
  OR2_X1 u_majority7_module_64__or_module_2_U1 ( .A1(n_majority7_module_64_n3), 
        .A2(n_majority7_module_64_n5), .ZN(
        n_majority7_module_64__or_module_2_res) );
  AND2_X1 u_majority7_module_64__and_module_3_U1 ( .A1(
        n_majority7_module_64_n6), .A2(n_majority7_module_64_n4), .ZN(
        n_majority7_module_64__and_module_3_res) );
  OR2_X1 u_majority7_module_64__or_module_3_U1 ( .A1(n_majority7_module_64_n4), 
        .A2(n_majority7_module_64_n6), .ZN(
        n_majority7_module_64__or_module_3_res) );
  AND2_X1 u_majority7_module_64__and_module_4_U1 ( .A1(
        n_majority7_module_64__and_module_2_res), .A2(
        n_majority7_module_64__and_module_1_res), .ZN(
        n_majority7_module_64__and_module_4_res) );
  OR2_X1 u_majority7_module_64__or_module_4_U1 ( .A1(
        n_majority7_module_64__and_module_1_res), .A2(
        n_majority7_module_64__and_module_2_res), .ZN(
        n_majority7_module_64__or_module_4_res) );
  AND2_X1 u_majority7_module_64__and_module_5_U1 ( .A1(
        n_majority7_module_64__and_module_3_res), .A2(n_majority7_module_64_n2), .ZN(n_majority7_module_64__and_module_5_res) );
  OR2_X1 u_majority7_module_64__or_module_5_U1 ( .A1(n_majority7_module_64_n2), 
        .A2(n_majority7_module_64__and_module_3_res), .ZN(
        n_majority7_module_64__or_module_5_res) );
  AND2_X1 u_majority7_module_64__and_module_6_U1 ( .A1(
        n_majority7_module_64__or_module_1_res), .A2(
        n_majority7_module_64__or_module_2_res), .ZN(
        n_majority7_module_64__and_module_6_res) );
  OR2_X1 u_majority7_module_64__or_module_6_U1 ( .A1(
        n_majority7_module_64__or_module_2_res), .A2(
        n_majority7_module_64__or_module_1_res), .ZN(
        n_majority7_module_64__or_module_6_res) );
  OR2_X1 u_majority7_module_64__or_module_7_U1 ( .A1(
        n_majority7_module_64__and_module_4_res), .A2(
        n_majority7_module_64__and_module_5_res), .ZN(
        n_majority7_module_64__or_module_7_res) );
  AND2_X1 u_majority7_module_64__and_module_7_U1 ( .A1(
        n_majority7_module_64__or_module_3_res), .A2(
        n_majority7_module_64__or_module_4_res), .ZN(
        n_majority7_module_64__and_module_7_res) );
  OR2_X1 u_majority7_module_64__or_module_8_U1 ( .A1(
        n_majority7_module_64__or_module_4_res), .A2(
        n_majority7_module_64__or_module_3_res), .ZN(
        n_majority7_module_64__or_module_8_res) );
  AND2_X1 u_majority7_module_64__and_module_8_U1 ( .A1(
        n_majority7_module_64__or_module_5_res), .A2(
        n_majority7_module_64__and_module_6_res), .ZN(
        n_majority7_module_64__and_module_8_res) );
  OR2_X1 u_majority7_module_64__or_module_9_U1 ( .A1(
        n_majority7_module_64__and_module_6_res), .A2(
        n_majority7_module_64__or_module_5_res), .ZN(
        n_majority7_module_64__or_module_9_res) );
  OR2_X1 u_majority7_module_64__or_module_10_U1 ( .A1(
        n_majority7_module_64__or_module_7_res), .A2(
        n_majority7_module_64__and_module_7_res), .ZN(
        n_majority7_module_64__or_module_10_res) );
  AND2_X1 u_majority7_module_64__and_module_9_U1 ( .A1(
        n_majority7_module_64__or_module_6_res), .A2(
        n_majority7_module_64__or_module_9_res), .ZN(
        n_majority7_module_64__and_module_9_res) );
  OR2_X1 u_majority7_module_64__or_module_11_U1 ( .A1(
        n_majority7_module_64__or_module_10_res), .A2(
        n_majority7_module_64__and_module_8_res), .ZN(
        n_majority7_module_64__or_module_11_res) );
  AND2_X1 u_majority7_module_64__and_module_10_U1 ( .A1(
        n_majority7_module_64__or_module_8_res), .A2(
        n_majority7_module_64__and_module_9_res), .ZN(
        n_majority7_module_64__and_module_10_res) );
  AND2_X1 u_majority7_module_64__and_module_11_U1 ( .A1(
        n_majority7_module_64__and_module_10_res), .A2(
        n_majority7_module_64__or_module_11_res), .ZN(
        n_majority7_module_64_res) );
  DFF_X1 u_reg_module_65__cini_mul_v000_reg ( .D(n_majority7_module_64_res), 
        .CK(clock_4), .Q(n_reg_module_65_res), .QN() );
  BUF_X1 u_majority7_module_65_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_65_n7) );
  BUF_X1 u_majority7_module_65_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_65_n6) );
  BUF_X1 u_majority7_module_65_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_65_n5) );
  BUF_X1 u_majority7_module_65_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_65_n4) );
  BUF_X1 u_majority7_module_65_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_65_n3) );
  BUF_X1 u_majority7_module_65_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_65_n2) );
  BUF_X1 u_majority7_module_65_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_65_n1) );
  AND2_X1 u_majority7_module_65__and_module_1_U1 ( .A1(
        n_majority7_module_65_n7), .A2(n_majority7_module_65_n1), .ZN(
        n_majority7_module_65__and_module_1_res) );
  OR2_X1 u_majority7_module_65__or_module_1_U1 ( .A1(n_majority7_module_65_n1), 
        .A2(n_majority7_module_65_n7), .ZN(
        n_majority7_module_65__or_module_1_res) );
  AND2_X1 u_majority7_module_65__and_module_2_U1 ( .A1(
        n_majority7_module_65_n5), .A2(n_majority7_module_65_n3), .ZN(
        n_majority7_module_65__and_module_2_res) );
  OR2_X1 u_majority7_module_65__or_module_2_U1 ( .A1(n_majority7_module_65_n3), 
        .A2(n_majority7_module_65_n5), .ZN(
        n_majority7_module_65__or_module_2_res) );
  AND2_X1 u_majority7_module_65__and_module_3_U1 ( .A1(
        n_majority7_module_65_n6), .A2(n_majority7_module_65_n4), .ZN(
        n_majority7_module_65__and_module_3_res) );
  OR2_X1 u_majority7_module_65__or_module_3_U1 ( .A1(n_majority7_module_65_n4), 
        .A2(n_majority7_module_65_n6), .ZN(
        n_majority7_module_65__or_module_3_res) );
  AND2_X1 u_majority7_module_65__and_module_4_U1 ( .A1(
        n_majority7_module_65__and_module_2_res), .A2(
        n_majority7_module_65__and_module_1_res), .ZN(
        n_majority7_module_65__and_module_4_res) );
  OR2_X1 u_majority7_module_65__or_module_4_U1 ( .A1(
        n_majority7_module_65__and_module_1_res), .A2(
        n_majority7_module_65__and_module_2_res), .ZN(
        n_majority7_module_65__or_module_4_res) );
  AND2_X1 u_majority7_module_65__and_module_5_U1 ( .A1(
        n_majority7_module_65__and_module_3_res), .A2(n_majority7_module_65_n2), .ZN(n_majority7_module_65__and_module_5_res) );
  OR2_X1 u_majority7_module_65__or_module_5_U1 ( .A1(n_majority7_module_65_n2), 
        .A2(n_majority7_module_65__and_module_3_res), .ZN(
        n_majority7_module_65__or_module_5_res) );
  AND2_X1 u_majority7_module_65__and_module_6_U1 ( .A1(
        n_majority7_module_65__or_module_1_res), .A2(
        n_majority7_module_65__or_module_2_res), .ZN(
        n_majority7_module_65__and_module_6_res) );
  OR2_X1 u_majority7_module_65__or_module_6_U1 ( .A1(
        n_majority7_module_65__or_module_2_res), .A2(
        n_majority7_module_65__or_module_1_res), .ZN(
        n_majority7_module_65__or_module_6_res) );
  OR2_X1 u_majority7_module_65__or_module_7_U1 ( .A1(
        n_majority7_module_65__and_module_4_res), .A2(
        n_majority7_module_65__and_module_5_res), .ZN(
        n_majority7_module_65__or_module_7_res) );
  AND2_X1 u_majority7_module_65__and_module_7_U1 ( .A1(
        n_majority7_module_65__or_module_3_res), .A2(
        n_majority7_module_65__or_module_4_res), .ZN(
        n_majority7_module_65__and_module_7_res) );
  OR2_X1 u_majority7_module_65__or_module_8_U1 ( .A1(
        n_majority7_module_65__or_module_4_res), .A2(
        n_majority7_module_65__or_module_3_res), .ZN(
        n_majority7_module_65__or_module_8_res) );
  AND2_X1 u_majority7_module_65__and_module_8_U1 ( .A1(
        n_majority7_module_65__or_module_5_res), .A2(
        n_majority7_module_65__and_module_6_res), .ZN(
        n_majority7_module_65__and_module_8_res) );
  OR2_X1 u_majority7_module_65__or_module_9_U1 ( .A1(
        n_majority7_module_65__and_module_6_res), .A2(
        n_majority7_module_65__or_module_5_res), .ZN(
        n_majority7_module_65__or_module_9_res) );
  OR2_X1 u_majority7_module_65__or_module_10_U1 ( .A1(
        n_majority7_module_65__or_module_7_res), .A2(
        n_majority7_module_65__and_module_7_res), .ZN(
        n_majority7_module_65__or_module_10_res) );
  AND2_X1 u_majority7_module_65__and_module_9_U1 ( .A1(
        n_majority7_module_65__or_module_6_res), .A2(
        n_majority7_module_65__or_module_9_res), .ZN(
        n_majority7_module_65__and_module_9_res) );
  OR2_X1 u_majority7_module_65__or_module_11_U1 ( .A1(
        n_majority7_module_65__or_module_10_res), .A2(
        n_majority7_module_65__and_module_8_res), .ZN(
        n_majority7_module_65__or_module_11_res) );
  AND2_X1 u_majority7_module_65__and_module_10_U1 ( .A1(
        n_majority7_module_65__or_module_8_res), .A2(
        n_majority7_module_65__and_module_9_res), .ZN(
        n_majority7_module_65__and_module_10_res) );
  AND2_X1 u_majority7_module_65__and_module_11_U1 ( .A1(
        n_majority7_module_65__and_module_10_res), .A2(
        n_majority7_module_65__or_module_11_res), .ZN(
        n_majority7_module_65_res) );
  DFF_X1 u_reg_module_66__cini_mul_v000_reg ( .D(n_majority7_module_65_res), 
        .CK(clock_4), .Q(n_reg_module_66_res), .QN() );
  BUF_X1 u_majority7_module_66_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_66_n7) );
  BUF_X1 u_majority7_module_66_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_66_n6) );
  BUF_X1 u_majority7_module_66_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_66_n5) );
  BUF_X1 u_majority7_module_66_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_66_n4) );
  BUF_X1 u_majority7_module_66_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_66_n3) );
  BUF_X1 u_majority7_module_66_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_66_n2) );
  BUF_X1 u_majority7_module_66_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_66_n1) );
  AND2_X1 u_majority7_module_66__and_module_1_U1 ( .A1(
        n_majority7_module_66_n7), .A2(n_majority7_module_66_n1), .ZN(
        n_majority7_module_66__and_module_1_res) );
  OR2_X1 u_majority7_module_66__or_module_1_U1 ( .A1(n_majority7_module_66_n1), 
        .A2(n_majority7_module_66_n7), .ZN(
        n_majority7_module_66__or_module_1_res) );
  AND2_X1 u_majority7_module_66__and_module_2_U1 ( .A1(
        n_majority7_module_66_n5), .A2(n_majority7_module_66_n3), .ZN(
        n_majority7_module_66__and_module_2_res) );
  OR2_X1 u_majority7_module_66__or_module_2_U1 ( .A1(n_majority7_module_66_n3), 
        .A2(n_majority7_module_66_n5), .ZN(
        n_majority7_module_66__or_module_2_res) );
  AND2_X1 u_majority7_module_66__and_module_3_U1 ( .A1(
        n_majority7_module_66_n6), .A2(n_majority7_module_66_n4), .ZN(
        n_majority7_module_66__and_module_3_res) );
  OR2_X1 u_majority7_module_66__or_module_3_U1 ( .A1(n_majority7_module_66_n4), 
        .A2(n_majority7_module_66_n6), .ZN(
        n_majority7_module_66__or_module_3_res) );
  AND2_X1 u_majority7_module_66__and_module_4_U1 ( .A1(
        n_majority7_module_66__and_module_2_res), .A2(
        n_majority7_module_66__and_module_1_res), .ZN(
        n_majority7_module_66__and_module_4_res) );
  OR2_X1 u_majority7_module_66__or_module_4_U1 ( .A1(
        n_majority7_module_66__and_module_1_res), .A2(
        n_majority7_module_66__and_module_2_res), .ZN(
        n_majority7_module_66__or_module_4_res) );
  AND2_X1 u_majority7_module_66__and_module_5_U1 ( .A1(
        n_majority7_module_66__and_module_3_res), .A2(n_majority7_module_66_n2), .ZN(n_majority7_module_66__and_module_5_res) );
  OR2_X1 u_majority7_module_66__or_module_5_U1 ( .A1(n_majority7_module_66_n2), 
        .A2(n_majority7_module_66__and_module_3_res), .ZN(
        n_majority7_module_66__or_module_5_res) );
  AND2_X1 u_majority7_module_66__and_module_6_U1 ( .A1(
        n_majority7_module_66__or_module_1_res), .A2(
        n_majority7_module_66__or_module_2_res), .ZN(
        n_majority7_module_66__and_module_6_res) );
  OR2_X1 u_majority7_module_66__or_module_6_U1 ( .A1(
        n_majority7_module_66__or_module_2_res), .A2(
        n_majority7_module_66__or_module_1_res), .ZN(
        n_majority7_module_66__or_module_6_res) );
  OR2_X1 u_majority7_module_66__or_module_7_U1 ( .A1(
        n_majority7_module_66__and_module_4_res), .A2(
        n_majority7_module_66__and_module_5_res), .ZN(
        n_majority7_module_66__or_module_7_res) );
  AND2_X1 u_majority7_module_66__and_module_7_U1 ( .A1(
        n_majority7_module_66__or_module_3_res), .A2(
        n_majority7_module_66__or_module_4_res), .ZN(
        n_majority7_module_66__and_module_7_res) );
  OR2_X1 u_majority7_module_66__or_module_8_U1 ( .A1(
        n_majority7_module_66__or_module_4_res), .A2(
        n_majority7_module_66__or_module_3_res), .ZN(
        n_majority7_module_66__or_module_8_res) );
  AND2_X1 u_majority7_module_66__and_module_8_U1 ( .A1(
        n_majority7_module_66__or_module_5_res), .A2(
        n_majority7_module_66__and_module_6_res), .ZN(
        n_majority7_module_66__and_module_8_res) );
  OR2_X1 u_majority7_module_66__or_module_9_U1 ( .A1(
        n_majority7_module_66__and_module_6_res), .A2(
        n_majority7_module_66__or_module_5_res), .ZN(
        n_majority7_module_66__or_module_9_res) );
  OR2_X1 u_majority7_module_66__or_module_10_U1 ( .A1(
        n_majority7_module_66__or_module_7_res), .A2(
        n_majority7_module_66__and_module_7_res), .ZN(
        n_majority7_module_66__or_module_10_res) );
  AND2_X1 u_majority7_module_66__and_module_9_U1 ( .A1(
        n_majority7_module_66__or_module_6_res), .A2(
        n_majority7_module_66__or_module_9_res), .ZN(
        n_majority7_module_66__and_module_9_res) );
  OR2_X1 u_majority7_module_66__or_module_11_U1 ( .A1(
        n_majority7_module_66__or_module_10_res), .A2(
        n_majority7_module_66__and_module_8_res), .ZN(
        n_majority7_module_66__or_module_11_res) );
  AND2_X1 u_majority7_module_66__and_module_10_U1 ( .A1(
        n_majority7_module_66__or_module_8_res), .A2(
        n_majority7_module_66__and_module_9_res), .ZN(
        n_majority7_module_66__and_module_10_res) );
  AND2_X1 u_majority7_module_66__and_module_11_U1 ( .A1(
        n_majority7_module_66__and_module_10_res), .A2(
        n_majority7_module_66__or_module_11_res), .ZN(
        n_majority7_module_66_res) );
  DFF_X1 u_reg_module_67__cini_mul_v000_reg ( .D(n_majority7_module_66_res), 
        .CK(clock_4), .Q(n_reg_module_67_res), .QN() );
  BUF_X1 u_majority7_module_67_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_67_n7) );
  BUF_X1 u_majority7_module_67_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_67_n6) );
  BUF_X1 u_majority7_module_67_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_67_n5) );
  BUF_X1 u_majority7_module_67_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_67_n4) );
  BUF_X1 u_majority7_module_67_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_67_n3) );
  BUF_X1 u_majority7_module_67_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_67_n2) );
  BUF_X1 u_majority7_module_67_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_67_n1) );
  AND2_X1 u_majority7_module_67__and_module_1_U1 ( .A1(
        n_majority7_module_67_n7), .A2(n_majority7_module_67_n1), .ZN(
        n_majority7_module_67__and_module_1_res) );
  OR2_X1 u_majority7_module_67__or_module_1_U1 ( .A1(n_majority7_module_67_n1), 
        .A2(n_majority7_module_67_n7), .ZN(
        n_majority7_module_67__or_module_1_res) );
  AND2_X1 u_majority7_module_67__and_module_2_U1 ( .A1(
        n_majority7_module_67_n5), .A2(n_majority7_module_67_n3), .ZN(
        n_majority7_module_67__and_module_2_res) );
  OR2_X1 u_majority7_module_67__or_module_2_U1 ( .A1(n_majority7_module_67_n3), 
        .A2(n_majority7_module_67_n5), .ZN(
        n_majority7_module_67__or_module_2_res) );
  AND2_X1 u_majority7_module_67__and_module_3_U1 ( .A1(
        n_majority7_module_67_n6), .A2(n_majority7_module_67_n4), .ZN(
        n_majority7_module_67__and_module_3_res) );
  OR2_X1 u_majority7_module_67__or_module_3_U1 ( .A1(n_majority7_module_67_n4), 
        .A2(n_majority7_module_67_n6), .ZN(
        n_majority7_module_67__or_module_3_res) );
  AND2_X1 u_majority7_module_67__and_module_4_U1 ( .A1(
        n_majority7_module_67__and_module_2_res), .A2(
        n_majority7_module_67__and_module_1_res), .ZN(
        n_majority7_module_67__and_module_4_res) );
  OR2_X1 u_majority7_module_67__or_module_4_U1 ( .A1(
        n_majority7_module_67__and_module_1_res), .A2(
        n_majority7_module_67__and_module_2_res), .ZN(
        n_majority7_module_67__or_module_4_res) );
  AND2_X1 u_majority7_module_67__and_module_5_U1 ( .A1(
        n_majority7_module_67__and_module_3_res), .A2(n_majority7_module_67_n2), .ZN(n_majority7_module_67__and_module_5_res) );
  OR2_X1 u_majority7_module_67__or_module_5_U1 ( .A1(n_majority7_module_67_n2), 
        .A2(n_majority7_module_67__and_module_3_res), .ZN(
        n_majority7_module_67__or_module_5_res) );
  AND2_X1 u_majority7_module_67__and_module_6_U1 ( .A1(
        n_majority7_module_67__or_module_1_res), .A2(
        n_majority7_module_67__or_module_2_res), .ZN(
        n_majority7_module_67__and_module_6_res) );
  OR2_X1 u_majority7_module_67__or_module_6_U1 ( .A1(
        n_majority7_module_67__or_module_2_res), .A2(
        n_majority7_module_67__or_module_1_res), .ZN(
        n_majority7_module_67__or_module_6_res) );
  OR2_X1 u_majority7_module_67__or_module_7_U1 ( .A1(
        n_majority7_module_67__and_module_4_res), .A2(
        n_majority7_module_67__and_module_5_res), .ZN(
        n_majority7_module_67__or_module_7_res) );
  AND2_X1 u_majority7_module_67__and_module_7_U1 ( .A1(
        n_majority7_module_67__or_module_3_res), .A2(
        n_majority7_module_67__or_module_4_res), .ZN(
        n_majority7_module_67__and_module_7_res) );
  OR2_X1 u_majority7_module_67__or_module_8_U1 ( .A1(
        n_majority7_module_67__or_module_4_res), .A2(
        n_majority7_module_67__or_module_3_res), .ZN(
        n_majority7_module_67__or_module_8_res) );
  AND2_X1 u_majority7_module_67__and_module_8_U1 ( .A1(
        n_majority7_module_67__or_module_5_res), .A2(
        n_majority7_module_67__and_module_6_res), .ZN(
        n_majority7_module_67__and_module_8_res) );
  OR2_X1 u_majority7_module_67__or_module_9_U1 ( .A1(
        n_majority7_module_67__and_module_6_res), .A2(
        n_majority7_module_67__or_module_5_res), .ZN(
        n_majority7_module_67__or_module_9_res) );
  OR2_X1 u_majority7_module_67__or_module_10_U1 ( .A1(
        n_majority7_module_67__or_module_7_res), .A2(
        n_majority7_module_67__and_module_7_res), .ZN(
        n_majority7_module_67__or_module_10_res) );
  AND2_X1 u_majority7_module_67__and_module_9_U1 ( .A1(
        n_majority7_module_67__or_module_6_res), .A2(
        n_majority7_module_67__or_module_9_res), .ZN(
        n_majority7_module_67__and_module_9_res) );
  OR2_X1 u_majority7_module_67__or_module_11_U1 ( .A1(
        n_majority7_module_67__or_module_10_res), .A2(
        n_majority7_module_67__and_module_8_res), .ZN(
        n_majority7_module_67__or_module_11_res) );
  AND2_X1 u_majority7_module_67__and_module_10_U1 ( .A1(
        n_majority7_module_67__or_module_8_res), .A2(
        n_majority7_module_67__and_module_9_res), .ZN(
        n_majority7_module_67__and_module_10_res) );
  AND2_X1 u_majority7_module_67__and_module_11_U1 ( .A1(
        n_majority7_module_67__and_module_10_res), .A2(
        n_majority7_module_67__or_module_11_res), .ZN(
        n_majority7_module_67_res) );
  DFF_X1 u_reg_module_68__cini_mul_v000_reg ( .D(n_majority7_module_67_res), 
        .CK(clock_4), .Q(n_reg_module_68_res), .QN() );
  BUF_X1 u_majority7_module_68_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_68_n7) );
  BUF_X1 u_majority7_module_68_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_68_n6) );
  BUF_X1 u_majority7_module_68_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_68_n5) );
  BUF_X1 u_majority7_module_68_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_68_n4) );
  BUF_X1 u_majority7_module_68_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_68_n3) );
  BUF_X1 u_majority7_module_68_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_68_n2) );
  BUF_X1 u_majority7_module_68_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_68_n1) );
  AND2_X1 u_majority7_module_68__and_module_1_U1 ( .A1(
        n_majority7_module_68_n7), .A2(n_majority7_module_68_n1), .ZN(
        n_majority7_module_68__and_module_1_res) );
  OR2_X1 u_majority7_module_68__or_module_1_U1 ( .A1(n_majority7_module_68_n1), 
        .A2(n_majority7_module_68_n7), .ZN(
        n_majority7_module_68__or_module_1_res) );
  AND2_X1 u_majority7_module_68__and_module_2_U1 ( .A1(
        n_majority7_module_68_n5), .A2(n_majority7_module_68_n3), .ZN(
        n_majority7_module_68__and_module_2_res) );
  OR2_X1 u_majority7_module_68__or_module_2_U1 ( .A1(n_majority7_module_68_n3), 
        .A2(n_majority7_module_68_n5), .ZN(
        n_majority7_module_68__or_module_2_res) );
  AND2_X1 u_majority7_module_68__and_module_3_U1 ( .A1(
        n_majority7_module_68_n6), .A2(n_majority7_module_68_n4), .ZN(
        n_majority7_module_68__and_module_3_res) );
  OR2_X1 u_majority7_module_68__or_module_3_U1 ( .A1(n_majority7_module_68_n4), 
        .A2(n_majority7_module_68_n6), .ZN(
        n_majority7_module_68__or_module_3_res) );
  AND2_X1 u_majority7_module_68__and_module_4_U1 ( .A1(
        n_majority7_module_68__and_module_2_res), .A2(
        n_majority7_module_68__and_module_1_res), .ZN(
        n_majority7_module_68__and_module_4_res) );
  OR2_X1 u_majority7_module_68__or_module_4_U1 ( .A1(
        n_majority7_module_68__and_module_1_res), .A2(
        n_majority7_module_68__and_module_2_res), .ZN(
        n_majority7_module_68__or_module_4_res) );
  AND2_X1 u_majority7_module_68__and_module_5_U1 ( .A1(
        n_majority7_module_68__and_module_3_res), .A2(n_majority7_module_68_n2), .ZN(n_majority7_module_68__and_module_5_res) );
  OR2_X1 u_majority7_module_68__or_module_5_U1 ( .A1(n_majority7_module_68_n2), 
        .A2(n_majority7_module_68__and_module_3_res), .ZN(
        n_majority7_module_68__or_module_5_res) );
  AND2_X1 u_majority7_module_68__and_module_6_U1 ( .A1(
        n_majority7_module_68__or_module_1_res), .A2(
        n_majority7_module_68__or_module_2_res), .ZN(
        n_majority7_module_68__and_module_6_res) );
  OR2_X1 u_majority7_module_68__or_module_6_U1 ( .A1(
        n_majority7_module_68__or_module_2_res), .A2(
        n_majority7_module_68__or_module_1_res), .ZN(
        n_majority7_module_68__or_module_6_res) );
  OR2_X1 u_majority7_module_68__or_module_7_U1 ( .A1(
        n_majority7_module_68__and_module_4_res), .A2(
        n_majority7_module_68__and_module_5_res), .ZN(
        n_majority7_module_68__or_module_7_res) );
  AND2_X1 u_majority7_module_68__and_module_7_U1 ( .A1(
        n_majority7_module_68__or_module_3_res), .A2(
        n_majority7_module_68__or_module_4_res), .ZN(
        n_majority7_module_68__and_module_7_res) );
  OR2_X1 u_majority7_module_68__or_module_8_U1 ( .A1(
        n_majority7_module_68__or_module_4_res), .A2(
        n_majority7_module_68__or_module_3_res), .ZN(
        n_majority7_module_68__or_module_8_res) );
  AND2_X1 u_majority7_module_68__and_module_8_U1 ( .A1(
        n_majority7_module_68__or_module_5_res), .A2(
        n_majority7_module_68__and_module_6_res), .ZN(
        n_majority7_module_68__and_module_8_res) );
  OR2_X1 u_majority7_module_68__or_module_9_U1 ( .A1(
        n_majority7_module_68__and_module_6_res), .A2(
        n_majority7_module_68__or_module_5_res), .ZN(
        n_majority7_module_68__or_module_9_res) );
  OR2_X1 u_majority7_module_68__or_module_10_U1 ( .A1(
        n_majority7_module_68__or_module_7_res), .A2(
        n_majority7_module_68__and_module_7_res), .ZN(
        n_majority7_module_68__or_module_10_res) );
  AND2_X1 u_majority7_module_68__and_module_9_U1 ( .A1(
        n_majority7_module_68__or_module_6_res), .A2(
        n_majority7_module_68__or_module_9_res), .ZN(
        n_majority7_module_68__and_module_9_res) );
  OR2_X1 u_majority7_module_68__or_module_11_U1 ( .A1(
        n_majority7_module_68__or_module_10_res), .A2(
        n_majority7_module_68__and_module_8_res), .ZN(
        n_majority7_module_68__or_module_11_res) );
  AND2_X1 u_majority7_module_68__and_module_10_U1 ( .A1(
        n_majority7_module_68__or_module_8_res), .A2(
        n_majority7_module_68__and_module_9_res), .ZN(
        n_majority7_module_68__and_module_10_res) );
  AND2_X1 u_majority7_module_68__and_module_11_U1 ( .A1(
        n_majority7_module_68__and_module_10_res), .A2(
        n_majority7_module_68__or_module_11_res), .ZN(
        n_majority7_module_68_res) );
  DFF_X1 u_reg_module_69__cini_mul_v000_reg ( .D(n_majority7_module_68_res), 
        .CK(clock_4), .Q(n_reg_module_69_res), .QN() );
  BUF_X1 u_majority7_module_69_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_69_n7) );
  BUF_X1 u_majority7_module_69_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_69_n6) );
  BUF_X1 u_majority7_module_69_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_69_n5) );
  BUF_X1 u_majority7_module_69_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_69_n4) );
  BUF_X1 u_majority7_module_69_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_69_n3) );
  BUF_X1 u_majority7_module_69_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_69_n2) );
  BUF_X1 u_majority7_module_69_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_69_n1) );
  AND2_X1 u_majority7_module_69__and_module_1_U1 ( .A1(
        n_majority7_module_69_n7), .A2(n_majority7_module_69_n1), .ZN(
        n_majority7_module_69__and_module_1_res) );
  OR2_X1 u_majority7_module_69__or_module_1_U1 ( .A1(n_majority7_module_69_n1), 
        .A2(n_majority7_module_69_n7), .ZN(
        n_majority7_module_69__or_module_1_res) );
  AND2_X1 u_majority7_module_69__and_module_2_U1 ( .A1(
        n_majority7_module_69_n5), .A2(n_majority7_module_69_n3), .ZN(
        n_majority7_module_69__and_module_2_res) );
  OR2_X1 u_majority7_module_69__or_module_2_U1 ( .A1(n_majority7_module_69_n3), 
        .A2(n_majority7_module_69_n5), .ZN(
        n_majority7_module_69__or_module_2_res) );
  AND2_X1 u_majority7_module_69__and_module_3_U1 ( .A1(
        n_majority7_module_69_n6), .A2(n_majority7_module_69_n4), .ZN(
        n_majority7_module_69__and_module_3_res) );
  OR2_X1 u_majority7_module_69__or_module_3_U1 ( .A1(n_majority7_module_69_n4), 
        .A2(n_majority7_module_69_n6), .ZN(
        n_majority7_module_69__or_module_3_res) );
  AND2_X1 u_majority7_module_69__and_module_4_U1 ( .A1(
        n_majority7_module_69__and_module_2_res), .A2(
        n_majority7_module_69__and_module_1_res), .ZN(
        n_majority7_module_69__and_module_4_res) );
  OR2_X1 u_majority7_module_69__or_module_4_U1 ( .A1(
        n_majority7_module_69__and_module_1_res), .A2(
        n_majority7_module_69__and_module_2_res), .ZN(
        n_majority7_module_69__or_module_4_res) );
  AND2_X1 u_majority7_module_69__and_module_5_U1 ( .A1(
        n_majority7_module_69__and_module_3_res), .A2(n_majority7_module_69_n2), .ZN(n_majority7_module_69__and_module_5_res) );
  OR2_X1 u_majority7_module_69__or_module_5_U1 ( .A1(n_majority7_module_69_n2), 
        .A2(n_majority7_module_69__and_module_3_res), .ZN(
        n_majority7_module_69__or_module_5_res) );
  AND2_X1 u_majority7_module_69__and_module_6_U1 ( .A1(
        n_majority7_module_69__or_module_1_res), .A2(
        n_majority7_module_69__or_module_2_res), .ZN(
        n_majority7_module_69__and_module_6_res) );
  OR2_X1 u_majority7_module_69__or_module_6_U1 ( .A1(
        n_majority7_module_69__or_module_2_res), .A2(
        n_majority7_module_69__or_module_1_res), .ZN(
        n_majority7_module_69__or_module_6_res) );
  OR2_X1 u_majority7_module_69__or_module_7_U1 ( .A1(
        n_majority7_module_69__and_module_4_res), .A2(
        n_majority7_module_69__and_module_5_res), .ZN(
        n_majority7_module_69__or_module_7_res) );
  AND2_X1 u_majority7_module_69__and_module_7_U1 ( .A1(
        n_majority7_module_69__or_module_3_res), .A2(
        n_majority7_module_69__or_module_4_res), .ZN(
        n_majority7_module_69__and_module_7_res) );
  OR2_X1 u_majority7_module_69__or_module_8_U1 ( .A1(
        n_majority7_module_69__or_module_4_res), .A2(
        n_majority7_module_69__or_module_3_res), .ZN(
        n_majority7_module_69__or_module_8_res) );
  AND2_X1 u_majority7_module_69__and_module_8_U1 ( .A1(
        n_majority7_module_69__or_module_5_res), .A2(
        n_majority7_module_69__and_module_6_res), .ZN(
        n_majority7_module_69__and_module_8_res) );
  OR2_X1 u_majority7_module_69__or_module_9_U1 ( .A1(
        n_majority7_module_69__and_module_6_res), .A2(
        n_majority7_module_69__or_module_5_res), .ZN(
        n_majority7_module_69__or_module_9_res) );
  OR2_X1 u_majority7_module_69__or_module_10_U1 ( .A1(
        n_majority7_module_69__or_module_7_res), .A2(
        n_majority7_module_69__and_module_7_res), .ZN(
        n_majority7_module_69__or_module_10_res) );
  AND2_X1 u_majority7_module_69__and_module_9_U1 ( .A1(
        n_majority7_module_69__or_module_6_res), .A2(
        n_majority7_module_69__or_module_9_res), .ZN(
        n_majority7_module_69__and_module_9_res) );
  OR2_X1 u_majority7_module_69__or_module_11_U1 ( .A1(
        n_majority7_module_69__or_module_10_res), .A2(
        n_majority7_module_69__and_module_8_res), .ZN(
        n_majority7_module_69__or_module_11_res) );
  AND2_X1 u_majority7_module_69__and_module_10_U1 ( .A1(
        n_majority7_module_69__or_module_8_res), .A2(
        n_majority7_module_69__and_module_9_res), .ZN(
        n_majority7_module_69__and_module_10_res) );
  AND2_X1 u_majority7_module_69__and_module_11_U1 ( .A1(
        n_majority7_module_69__and_module_10_res), .A2(
        n_majority7_module_69__or_module_11_res), .ZN(
        n_majority7_module_69_res) );
  DFF_X1 u_reg_module_70__cini_mul_v000_reg ( .D(n_majority7_module_69_res), 
        .CK(clock_4), .Q(n_reg_module_70_res), .QN() );
  BUF_X1 u_majority7_module_70_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_70_n7) );
  BUF_X1 u_majority7_module_70_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_70_n6) );
  BUF_X1 u_majority7_module_70_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_70_n5) );
  BUF_X1 u_majority7_module_70_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_70_n4) );
  BUF_X1 u_majority7_module_70_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_70_n3) );
  BUF_X1 u_majority7_module_70_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_70_n2) );
  BUF_X1 u_majority7_module_70_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_70_n1) );
  AND2_X1 u_majority7_module_70__and_module_1_U1 ( .A1(
        n_majority7_module_70_n7), .A2(n_majority7_module_70_n1), .ZN(
        n_majority7_module_70__and_module_1_res) );
  OR2_X1 u_majority7_module_70__or_module_1_U1 ( .A1(n_majority7_module_70_n1), 
        .A2(n_majority7_module_70_n7), .ZN(
        n_majority7_module_70__or_module_1_res) );
  AND2_X1 u_majority7_module_70__and_module_2_U1 ( .A1(
        n_majority7_module_70_n5), .A2(n_majority7_module_70_n3), .ZN(
        n_majority7_module_70__and_module_2_res) );
  OR2_X1 u_majority7_module_70__or_module_2_U1 ( .A1(n_majority7_module_70_n3), 
        .A2(n_majority7_module_70_n5), .ZN(
        n_majority7_module_70__or_module_2_res) );
  AND2_X1 u_majority7_module_70__and_module_3_U1 ( .A1(
        n_majority7_module_70_n6), .A2(n_majority7_module_70_n4), .ZN(
        n_majority7_module_70__and_module_3_res) );
  OR2_X1 u_majority7_module_70__or_module_3_U1 ( .A1(n_majority7_module_70_n4), 
        .A2(n_majority7_module_70_n6), .ZN(
        n_majority7_module_70__or_module_3_res) );
  AND2_X1 u_majority7_module_70__and_module_4_U1 ( .A1(
        n_majority7_module_70__and_module_2_res), .A2(
        n_majority7_module_70__and_module_1_res), .ZN(
        n_majority7_module_70__and_module_4_res) );
  OR2_X1 u_majority7_module_70__or_module_4_U1 ( .A1(
        n_majority7_module_70__and_module_1_res), .A2(
        n_majority7_module_70__and_module_2_res), .ZN(
        n_majority7_module_70__or_module_4_res) );
  AND2_X1 u_majority7_module_70__and_module_5_U1 ( .A1(
        n_majority7_module_70__and_module_3_res), .A2(n_majority7_module_70_n2), .ZN(n_majority7_module_70__and_module_5_res) );
  OR2_X1 u_majority7_module_70__or_module_5_U1 ( .A1(n_majority7_module_70_n2), 
        .A2(n_majority7_module_70__and_module_3_res), .ZN(
        n_majority7_module_70__or_module_5_res) );
  AND2_X1 u_majority7_module_70__and_module_6_U1 ( .A1(
        n_majority7_module_70__or_module_1_res), .A2(
        n_majority7_module_70__or_module_2_res), .ZN(
        n_majority7_module_70__and_module_6_res) );
  OR2_X1 u_majority7_module_70__or_module_6_U1 ( .A1(
        n_majority7_module_70__or_module_2_res), .A2(
        n_majority7_module_70__or_module_1_res), .ZN(
        n_majority7_module_70__or_module_6_res) );
  OR2_X1 u_majority7_module_70__or_module_7_U1 ( .A1(
        n_majority7_module_70__and_module_4_res), .A2(
        n_majority7_module_70__and_module_5_res), .ZN(
        n_majority7_module_70__or_module_7_res) );
  AND2_X1 u_majority7_module_70__and_module_7_U1 ( .A1(
        n_majority7_module_70__or_module_3_res), .A2(
        n_majority7_module_70__or_module_4_res), .ZN(
        n_majority7_module_70__and_module_7_res) );
  OR2_X1 u_majority7_module_70__or_module_8_U1 ( .A1(
        n_majority7_module_70__or_module_4_res), .A2(
        n_majority7_module_70__or_module_3_res), .ZN(
        n_majority7_module_70__or_module_8_res) );
  AND2_X1 u_majority7_module_70__and_module_8_U1 ( .A1(
        n_majority7_module_70__or_module_5_res), .A2(
        n_majority7_module_70__and_module_6_res), .ZN(
        n_majority7_module_70__and_module_8_res) );
  OR2_X1 u_majority7_module_70__or_module_9_U1 ( .A1(
        n_majority7_module_70__and_module_6_res), .A2(
        n_majority7_module_70__or_module_5_res), .ZN(
        n_majority7_module_70__or_module_9_res) );
  OR2_X1 u_majority7_module_70__or_module_10_U1 ( .A1(
        n_majority7_module_70__or_module_7_res), .A2(
        n_majority7_module_70__and_module_7_res), .ZN(
        n_majority7_module_70__or_module_10_res) );
  AND2_X1 u_majority7_module_70__and_module_9_U1 ( .A1(
        n_majority7_module_70__or_module_6_res), .A2(
        n_majority7_module_70__or_module_9_res), .ZN(
        n_majority7_module_70__and_module_9_res) );
  OR2_X1 u_majority7_module_70__or_module_11_U1 ( .A1(
        n_majority7_module_70__or_module_10_res), .A2(
        n_majority7_module_70__and_module_8_res), .ZN(
        n_majority7_module_70__or_module_11_res) );
  AND2_X1 u_majority7_module_70__and_module_10_U1 ( .A1(
        n_majority7_module_70__or_module_8_res), .A2(
        n_majority7_module_70__and_module_9_res), .ZN(
        n_majority7_module_70__and_module_10_res) );
  AND2_X1 u_majority7_module_70__and_module_11_U1 ( .A1(
        n_majority7_module_70__and_module_10_res), .A2(
        n_majority7_module_70__or_module_11_res), .ZN(
        n_majority7_module_70_res) );
  DFF_X1 u_reg_module_71__cini_mul_v000_reg ( .D(n_majority7_module_70_res), 
        .CK(clock_4), .Q(n_reg_module_71_res), .QN() );
  BUF_X1 u_majority7_module_71_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_71_n7) );
  BUF_X1 u_majority7_module_71_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_71_n6) );
  BUF_X1 u_majority7_module_71_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_71_n5) );
  BUF_X1 u_majority7_module_71_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_71_n4) );
  BUF_X1 u_majority7_module_71_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_71_n3) );
  BUF_X1 u_majority7_module_71_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_71_n2) );
  BUF_X1 u_majority7_module_71_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_71_n1) );
  AND2_X1 u_majority7_module_71__and_module_1_U1 ( .A1(
        n_majority7_module_71_n7), .A2(n_majority7_module_71_n1), .ZN(
        n_majority7_module_71__and_module_1_res) );
  OR2_X1 u_majority7_module_71__or_module_1_U1 ( .A1(n_majority7_module_71_n1), 
        .A2(n_majority7_module_71_n7), .ZN(
        n_majority7_module_71__or_module_1_res) );
  AND2_X1 u_majority7_module_71__and_module_2_U1 ( .A1(
        n_majority7_module_71_n5), .A2(n_majority7_module_71_n3), .ZN(
        n_majority7_module_71__and_module_2_res) );
  OR2_X1 u_majority7_module_71__or_module_2_U1 ( .A1(n_majority7_module_71_n3), 
        .A2(n_majority7_module_71_n5), .ZN(
        n_majority7_module_71__or_module_2_res) );
  AND2_X1 u_majority7_module_71__and_module_3_U1 ( .A1(
        n_majority7_module_71_n6), .A2(n_majority7_module_71_n4), .ZN(
        n_majority7_module_71__and_module_3_res) );
  OR2_X1 u_majority7_module_71__or_module_3_U1 ( .A1(n_majority7_module_71_n4), 
        .A2(n_majority7_module_71_n6), .ZN(
        n_majority7_module_71__or_module_3_res) );
  AND2_X1 u_majority7_module_71__and_module_4_U1 ( .A1(
        n_majority7_module_71__and_module_2_res), .A2(
        n_majority7_module_71__and_module_1_res), .ZN(
        n_majority7_module_71__and_module_4_res) );
  OR2_X1 u_majority7_module_71__or_module_4_U1 ( .A1(
        n_majority7_module_71__and_module_1_res), .A2(
        n_majority7_module_71__and_module_2_res), .ZN(
        n_majority7_module_71__or_module_4_res) );
  AND2_X1 u_majority7_module_71__and_module_5_U1 ( .A1(
        n_majority7_module_71__and_module_3_res), .A2(n_majority7_module_71_n2), .ZN(n_majority7_module_71__and_module_5_res) );
  OR2_X1 u_majority7_module_71__or_module_5_U1 ( .A1(n_majority7_module_71_n2), 
        .A2(n_majority7_module_71__and_module_3_res), .ZN(
        n_majority7_module_71__or_module_5_res) );
  AND2_X1 u_majority7_module_71__and_module_6_U1 ( .A1(
        n_majority7_module_71__or_module_1_res), .A2(
        n_majority7_module_71__or_module_2_res), .ZN(
        n_majority7_module_71__and_module_6_res) );
  OR2_X1 u_majority7_module_71__or_module_6_U1 ( .A1(
        n_majority7_module_71__or_module_2_res), .A2(
        n_majority7_module_71__or_module_1_res), .ZN(
        n_majority7_module_71__or_module_6_res) );
  OR2_X1 u_majority7_module_71__or_module_7_U1 ( .A1(
        n_majority7_module_71__and_module_4_res), .A2(
        n_majority7_module_71__and_module_5_res), .ZN(
        n_majority7_module_71__or_module_7_res) );
  AND2_X1 u_majority7_module_71__and_module_7_U1 ( .A1(
        n_majority7_module_71__or_module_3_res), .A2(
        n_majority7_module_71__or_module_4_res), .ZN(
        n_majority7_module_71__and_module_7_res) );
  OR2_X1 u_majority7_module_71__or_module_8_U1 ( .A1(
        n_majority7_module_71__or_module_4_res), .A2(
        n_majority7_module_71__or_module_3_res), .ZN(
        n_majority7_module_71__or_module_8_res) );
  AND2_X1 u_majority7_module_71__and_module_8_U1 ( .A1(
        n_majority7_module_71__or_module_5_res), .A2(
        n_majority7_module_71__and_module_6_res), .ZN(
        n_majority7_module_71__and_module_8_res) );
  OR2_X1 u_majority7_module_71__or_module_9_U1 ( .A1(
        n_majority7_module_71__and_module_6_res), .A2(
        n_majority7_module_71__or_module_5_res), .ZN(
        n_majority7_module_71__or_module_9_res) );
  OR2_X1 u_majority7_module_71__or_module_10_U1 ( .A1(
        n_majority7_module_71__or_module_7_res), .A2(
        n_majority7_module_71__and_module_7_res), .ZN(
        n_majority7_module_71__or_module_10_res) );
  AND2_X1 u_majority7_module_71__and_module_9_U1 ( .A1(
        n_majority7_module_71__or_module_6_res), .A2(
        n_majority7_module_71__or_module_9_res), .ZN(
        n_majority7_module_71__and_module_9_res) );
  OR2_X1 u_majority7_module_71__or_module_11_U1 ( .A1(
        n_majority7_module_71__or_module_10_res), .A2(
        n_majority7_module_71__and_module_8_res), .ZN(
        n_majority7_module_71__or_module_11_res) );
  AND2_X1 u_majority7_module_71__and_module_10_U1 ( .A1(
        n_majority7_module_71__or_module_8_res), .A2(
        n_majority7_module_71__and_module_9_res), .ZN(
        n_majority7_module_71__and_module_10_res) );
  AND2_X1 u_majority7_module_71__and_module_11_U1 ( .A1(
        n_majority7_module_71__and_module_10_res), .A2(
        n_majority7_module_71__or_module_11_res), .ZN(
        n_majority7_module_71_res) );
  DFF_X1 u_reg_module_72__cini_mul_v000_reg ( .D(n_majority7_module_71_res), 
        .CK(clock_4), .Q(n_reg_module_72_res), .QN() );
  BUF_X1 u_majority7_module_72_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_72_n7) );
  BUF_X1 u_majority7_module_72_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_72_n6) );
  BUF_X1 u_majority7_module_72_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_72_n5) );
  BUF_X1 u_majority7_module_72_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_72_n4) );
  BUF_X1 u_majority7_module_72_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_72_n3) );
  BUF_X1 u_majority7_module_72_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_72_n2) );
  BUF_X1 u_majority7_module_72_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_72_n1) );
  AND2_X1 u_majority7_module_72__and_module_1_U1 ( .A1(
        n_majority7_module_72_n7), .A2(n_majority7_module_72_n1), .ZN(
        n_majority7_module_72__and_module_1_res) );
  OR2_X1 u_majority7_module_72__or_module_1_U1 ( .A1(n_majority7_module_72_n1), 
        .A2(n_majority7_module_72_n7), .ZN(
        n_majority7_module_72__or_module_1_res) );
  AND2_X1 u_majority7_module_72__and_module_2_U1 ( .A1(
        n_majority7_module_72_n5), .A2(n_majority7_module_72_n3), .ZN(
        n_majority7_module_72__and_module_2_res) );
  OR2_X1 u_majority7_module_72__or_module_2_U1 ( .A1(n_majority7_module_72_n3), 
        .A2(n_majority7_module_72_n5), .ZN(
        n_majority7_module_72__or_module_2_res) );
  AND2_X1 u_majority7_module_72__and_module_3_U1 ( .A1(
        n_majority7_module_72_n6), .A2(n_majority7_module_72_n4), .ZN(
        n_majority7_module_72__and_module_3_res) );
  OR2_X1 u_majority7_module_72__or_module_3_U1 ( .A1(n_majority7_module_72_n4), 
        .A2(n_majority7_module_72_n6), .ZN(
        n_majority7_module_72__or_module_3_res) );
  AND2_X1 u_majority7_module_72__and_module_4_U1 ( .A1(
        n_majority7_module_72__and_module_2_res), .A2(
        n_majority7_module_72__and_module_1_res), .ZN(
        n_majority7_module_72__and_module_4_res) );
  OR2_X1 u_majority7_module_72__or_module_4_U1 ( .A1(
        n_majority7_module_72__and_module_1_res), .A2(
        n_majority7_module_72__and_module_2_res), .ZN(
        n_majority7_module_72__or_module_4_res) );
  AND2_X1 u_majority7_module_72__and_module_5_U1 ( .A1(
        n_majority7_module_72__and_module_3_res), .A2(n_majority7_module_72_n2), .ZN(n_majority7_module_72__and_module_5_res) );
  OR2_X1 u_majority7_module_72__or_module_5_U1 ( .A1(n_majority7_module_72_n2), 
        .A2(n_majority7_module_72__and_module_3_res), .ZN(
        n_majority7_module_72__or_module_5_res) );
  AND2_X1 u_majority7_module_72__and_module_6_U1 ( .A1(
        n_majority7_module_72__or_module_1_res), .A2(
        n_majority7_module_72__or_module_2_res), .ZN(
        n_majority7_module_72__and_module_6_res) );
  OR2_X1 u_majority7_module_72__or_module_6_U1 ( .A1(
        n_majority7_module_72__or_module_2_res), .A2(
        n_majority7_module_72__or_module_1_res), .ZN(
        n_majority7_module_72__or_module_6_res) );
  OR2_X1 u_majority7_module_72__or_module_7_U1 ( .A1(
        n_majority7_module_72__and_module_4_res), .A2(
        n_majority7_module_72__and_module_5_res), .ZN(
        n_majority7_module_72__or_module_7_res) );
  AND2_X1 u_majority7_module_72__and_module_7_U1 ( .A1(
        n_majority7_module_72__or_module_3_res), .A2(
        n_majority7_module_72__or_module_4_res), .ZN(
        n_majority7_module_72__and_module_7_res) );
  OR2_X1 u_majority7_module_72__or_module_8_U1 ( .A1(
        n_majority7_module_72__or_module_4_res), .A2(
        n_majority7_module_72__or_module_3_res), .ZN(
        n_majority7_module_72__or_module_8_res) );
  AND2_X1 u_majority7_module_72__and_module_8_U1 ( .A1(
        n_majority7_module_72__or_module_5_res), .A2(
        n_majority7_module_72__and_module_6_res), .ZN(
        n_majority7_module_72__and_module_8_res) );
  OR2_X1 u_majority7_module_72__or_module_9_U1 ( .A1(
        n_majority7_module_72__and_module_6_res), .A2(
        n_majority7_module_72__or_module_5_res), .ZN(
        n_majority7_module_72__or_module_9_res) );
  OR2_X1 u_majority7_module_72__or_module_10_U1 ( .A1(
        n_majority7_module_72__or_module_7_res), .A2(
        n_majority7_module_72__and_module_7_res), .ZN(
        n_majority7_module_72__or_module_10_res) );
  AND2_X1 u_majority7_module_72__and_module_9_U1 ( .A1(
        n_majority7_module_72__or_module_6_res), .A2(
        n_majority7_module_72__or_module_9_res), .ZN(
        n_majority7_module_72__and_module_9_res) );
  OR2_X1 u_majority7_module_72__or_module_11_U1 ( .A1(
        n_majority7_module_72__or_module_10_res), .A2(
        n_majority7_module_72__and_module_8_res), .ZN(
        n_majority7_module_72__or_module_11_res) );
  AND2_X1 u_majority7_module_72__and_module_10_U1 ( .A1(
        n_majority7_module_72__or_module_8_res), .A2(
        n_majority7_module_72__and_module_9_res), .ZN(
        n_majority7_module_72__and_module_10_res) );
  AND2_X1 u_majority7_module_72__and_module_11_U1 ( .A1(
        n_majority7_module_72__and_module_10_res), .A2(
        n_majority7_module_72__or_module_11_res), .ZN(
        n_majority7_module_72_res) );
  DFF_X1 u_reg_module_73__cini_mul_v000_reg ( .D(n_majority7_module_72_res), 
        .CK(clock_4), .Q(n_reg_module_73_res), .QN() );
  BUF_X1 u_majority7_module_73_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_73_n7) );
  BUF_X1 u_majority7_module_73_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_73_n6) );
  BUF_X1 u_majority7_module_73_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_73_n5) );
  BUF_X1 u_majority7_module_73_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_73_n4) );
  BUF_X1 u_majority7_module_73_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_73_n3) );
  BUF_X1 u_majority7_module_73_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_73_n2) );
  BUF_X1 u_majority7_module_73_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_73_n1) );
  AND2_X1 u_majority7_module_73__and_module_1_U1 ( .A1(
        n_majority7_module_73_n7), .A2(n_majority7_module_73_n1), .ZN(
        n_majority7_module_73__and_module_1_res) );
  OR2_X1 u_majority7_module_73__or_module_1_U1 ( .A1(n_majority7_module_73_n1), 
        .A2(n_majority7_module_73_n7), .ZN(
        n_majority7_module_73__or_module_1_res) );
  AND2_X1 u_majority7_module_73__and_module_2_U1 ( .A1(
        n_majority7_module_73_n5), .A2(n_majority7_module_73_n3), .ZN(
        n_majority7_module_73__and_module_2_res) );
  OR2_X1 u_majority7_module_73__or_module_2_U1 ( .A1(n_majority7_module_73_n3), 
        .A2(n_majority7_module_73_n5), .ZN(
        n_majority7_module_73__or_module_2_res) );
  AND2_X1 u_majority7_module_73__and_module_3_U1 ( .A1(
        n_majority7_module_73_n6), .A2(n_majority7_module_73_n4), .ZN(
        n_majority7_module_73__and_module_3_res) );
  OR2_X1 u_majority7_module_73__or_module_3_U1 ( .A1(n_majority7_module_73_n4), 
        .A2(n_majority7_module_73_n6), .ZN(
        n_majority7_module_73__or_module_3_res) );
  AND2_X1 u_majority7_module_73__and_module_4_U1 ( .A1(
        n_majority7_module_73__and_module_2_res), .A2(
        n_majority7_module_73__and_module_1_res), .ZN(
        n_majority7_module_73__and_module_4_res) );
  OR2_X1 u_majority7_module_73__or_module_4_U1 ( .A1(
        n_majority7_module_73__and_module_1_res), .A2(
        n_majority7_module_73__and_module_2_res), .ZN(
        n_majority7_module_73__or_module_4_res) );
  AND2_X1 u_majority7_module_73__and_module_5_U1 ( .A1(
        n_majority7_module_73__and_module_3_res), .A2(n_majority7_module_73_n2), .ZN(n_majority7_module_73__and_module_5_res) );
  OR2_X1 u_majority7_module_73__or_module_5_U1 ( .A1(n_majority7_module_73_n2), 
        .A2(n_majority7_module_73__and_module_3_res), .ZN(
        n_majority7_module_73__or_module_5_res) );
  AND2_X1 u_majority7_module_73__and_module_6_U1 ( .A1(
        n_majority7_module_73__or_module_1_res), .A2(
        n_majority7_module_73__or_module_2_res), .ZN(
        n_majority7_module_73__and_module_6_res) );
  OR2_X1 u_majority7_module_73__or_module_6_U1 ( .A1(
        n_majority7_module_73__or_module_2_res), .A2(
        n_majority7_module_73__or_module_1_res), .ZN(
        n_majority7_module_73__or_module_6_res) );
  OR2_X1 u_majority7_module_73__or_module_7_U1 ( .A1(
        n_majority7_module_73__and_module_4_res), .A2(
        n_majority7_module_73__and_module_5_res), .ZN(
        n_majority7_module_73__or_module_7_res) );
  AND2_X1 u_majority7_module_73__and_module_7_U1 ( .A1(
        n_majority7_module_73__or_module_3_res), .A2(
        n_majority7_module_73__or_module_4_res), .ZN(
        n_majority7_module_73__and_module_7_res) );
  OR2_X1 u_majority7_module_73__or_module_8_U1 ( .A1(
        n_majority7_module_73__or_module_4_res), .A2(
        n_majority7_module_73__or_module_3_res), .ZN(
        n_majority7_module_73__or_module_8_res) );
  AND2_X1 u_majority7_module_73__and_module_8_U1 ( .A1(
        n_majority7_module_73__or_module_5_res), .A2(
        n_majority7_module_73__and_module_6_res), .ZN(
        n_majority7_module_73__and_module_8_res) );
  OR2_X1 u_majority7_module_73__or_module_9_U1 ( .A1(
        n_majority7_module_73__and_module_6_res), .A2(
        n_majority7_module_73__or_module_5_res), .ZN(
        n_majority7_module_73__or_module_9_res) );
  OR2_X1 u_majority7_module_73__or_module_10_U1 ( .A1(
        n_majority7_module_73__or_module_7_res), .A2(
        n_majority7_module_73__and_module_7_res), .ZN(
        n_majority7_module_73__or_module_10_res) );
  AND2_X1 u_majority7_module_73__and_module_9_U1 ( .A1(
        n_majority7_module_73__or_module_6_res), .A2(
        n_majority7_module_73__or_module_9_res), .ZN(
        n_majority7_module_73__and_module_9_res) );
  OR2_X1 u_majority7_module_73__or_module_11_U1 ( .A1(
        n_majority7_module_73__or_module_10_res), .A2(
        n_majority7_module_73__and_module_8_res), .ZN(
        n_majority7_module_73__or_module_11_res) );
  AND2_X1 u_majority7_module_73__and_module_10_U1 ( .A1(
        n_majority7_module_73__or_module_8_res), .A2(
        n_majority7_module_73__and_module_9_res), .ZN(
        n_majority7_module_73__and_module_10_res) );
  AND2_X1 u_majority7_module_73__and_module_11_U1 ( .A1(
        n_majority7_module_73__and_module_10_res), .A2(
        n_majority7_module_73__or_module_11_res), .ZN(
        n_majority7_module_73_res) );
  DFF_X1 u_reg_module_74__cini_mul_v000_reg ( .D(n_majority7_module_73_res), 
        .CK(clock_4), .Q(n_reg_module_74_res), .QN() );
  BUF_X1 u_majority7_module_74_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_74_n7) );
  BUF_X1 u_majority7_module_74_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_74_n6) );
  BUF_X1 u_majority7_module_74_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_74_n5) );
  BUF_X1 u_majority7_module_74_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_74_n4) );
  BUF_X1 u_majority7_module_74_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_74_n3) );
  BUF_X1 u_majority7_module_74_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_74_n2) );
  BUF_X1 u_majority7_module_74_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_74_n1) );
  AND2_X1 u_majority7_module_74__and_module_1_U1 ( .A1(
        n_majority7_module_74_n7), .A2(n_majority7_module_74_n1), .ZN(
        n_majority7_module_74__and_module_1_res) );
  OR2_X1 u_majority7_module_74__or_module_1_U1 ( .A1(n_majority7_module_74_n1), 
        .A2(n_majority7_module_74_n7), .ZN(
        n_majority7_module_74__or_module_1_res) );
  AND2_X1 u_majority7_module_74__and_module_2_U1 ( .A1(
        n_majority7_module_74_n5), .A2(n_majority7_module_74_n3), .ZN(
        n_majority7_module_74__and_module_2_res) );
  OR2_X1 u_majority7_module_74__or_module_2_U1 ( .A1(n_majority7_module_74_n3), 
        .A2(n_majority7_module_74_n5), .ZN(
        n_majority7_module_74__or_module_2_res) );
  AND2_X1 u_majority7_module_74__and_module_3_U1 ( .A1(
        n_majority7_module_74_n6), .A2(n_majority7_module_74_n4), .ZN(
        n_majority7_module_74__and_module_3_res) );
  OR2_X1 u_majority7_module_74__or_module_3_U1 ( .A1(n_majority7_module_74_n4), 
        .A2(n_majority7_module_74_n6), .ZN(
        n_majority7_module_74__or_module_3_res) );
  AND2_X1 u_majority7_module_74__and_module_4_U1 ( .A1(
        n_majority7_module_74__and_module_2_res), .A2(
        n_majority7_module_74__and_module_1_res), .ZN(
        n_majority7_module_74__and_module_4_res) );
  OR2_X1 u_majority7_module_74__or_module_4_U1 ( .A1(
        n_majority7_module_74__and_module_1_res), .A2(
        n_majority7_module_74__and_module_2_res), .ZN(
        n_majority7_module_74__or_module_4_res) );
  AND2_X1 u_majority7_module_74__and_module_5_U1 ( .A1(
        n_majority7_module_74__and_module_3_res), .A2(n_majority7_module_74_n2), .ZN(n_majority7_module_74__and_module_5_res) );
  OR2_X1 u_majority7_module_74__or_module_5_U1 ( .A1(n_majority7_module_74_n2), 
        .A2(n_majority7_module_74__and_module_3_res), .ZN(
        n_majority7_module_74__or_module_5_res) );
  AND2_X1 u_majority7_module_74__and_module_6_U1 ( .A1(
        n_majority7_module_74__or_module_1_res), .A2(
        n_majority7_module_74__or_module_2_res), .ZN(
        n_majority7_module_74__and_module_6_res) );
  OR2_X1 u_majority7_module_74__or_module_6_U1 ( .A1(
        n_majority7_module_74__or_module_2_res), .A2(
        n_majority7_module_74__or_module_1_res), .ZN(
        n_majority7_module_74__or_module_6_res) );
  OR2_X1 u_majority7_module_74__or_module_7_U1 ( .A1(
        n_majority7_module_74__and_module_4_res), .A2(
        n_majority7_module_74__and_module_5_res), .ZN(
        n_majority7_module_74__or_module_7_res) );
  AND2_X1 u_majority7_module_74__and_module_7_U1 ( .A1(
        n_majority7_module_74__or_module_3_res), .A2(
        n_majority7_module_74__or_module_4_res), .ZN(
        n_majority7_module_74__and_module_7_res) );
  OR2_X1 u_majority7_module_74__or_module_8_U1 ( .A1(
        n_majority7_module_74__or_module_4_res), .A2(
        n_majority7_module_74__or_module_3_res), .ZN(
        n_majority7_module_74__or_module_8_res) );
  AND2_X1 u_majority7_module_74__and_module_8_U1 ( .A1(
        n_majority7_module_74__or_module_5_res), .A2(
        n_majority7_module_74__and_module_6_res), .ZN(
        n_majority7_module_74__and_module_8_res) );
  OR2_X1 u_majority7_module_74__or_module_9_U1 ( .A1(
        n_majority7_module_74__and_module_6_res), .A2(
        n_majority7_module_74__or_module_5_res), .ZN(
        n_majority7_module_74__or_module_9_res) );
  OR2_X1 u_majority7_module_74__or_module_10_U1 ( .A1(
        n_majority7_module_74__or_module_7_res), .A2(
        n_majority7_module_74__and_module_7_res), .ZN(
        n_majority7_module_74__or_module_10_res) );
  AND2_X1 u_majority7_module_74__and_module_9_U1 ( .A1(
        n_majority7_module_74__or_module_6_res), .A2(
        n_majority7_module_74__or_module_9_res), .ZN(
        n_majority7_module_74__and_module_9_res) );
  OR2_X1 u_majority7_module_74__or_module_11_U1 ( .A1(
        n_majority7_module_74__or_module_10_res), .A2(
        n_majority7_module_74__and_module_8_res), .ZN(
        n_majority7_module_74__or_module_11_res) );
  AND2_X1 u_majority7_module_74__and_module_10_U1 ( .A1(
        n_majority7_module_74__or_module_8_res), .A2(
        n_majority7_module_74__and_module_9_res), .ZN(
        n_majority7_module_74__and_module_10_res) );
  AND2_X1 u_majority7_module_74__and_module_11_U1 ( .A1(
        n_majority7_module_74__and_module_10_res), .A2(
        n_majority7_module_74__or_module_11_res), .ZN(
        n_majority7_module_74_res) );
  DFF_X1 u_reg_module_75__cini_mul_v000_reg ( .D(n_majority7_module_74_res), 
        .CK(clock_4), .Q(n_reg_module_75_res), .QN() );
  BUF_X1 u_majority7_module_75_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_75_n7) );
  BUF_X1 u_majority7_module_75_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_75_n6) );
  BUF_X1 u_majority7_module_75_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_75_n5) );
  BUF_X1 u_majority7_module_75_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_75_n4) );
  BUF_X1 u_majority7_module_75_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_75_n3) );
  BUF_X1 u_majority7_module_75_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_75_n2) );
  BUF_X1 u_majority7_module_75_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_75_n1) );
  AND2_X1 u_majority7_module_75__and_module_1_U1 ( .A1(
        n_majority7_module_75_n7), .A2(n_majority7_module_75_n1), .ZN(
        n_majority7_module_75__and_module_1_res) );
  OR2_X1 u_majority7_module_75__or_module_1_U1 ( .A1(n_majority7_module_75_n1), 
        .A2(n_majority7_module_75_n7), .ZN(
        n_majority7_module_75__or_module_1_res) );
  AND2_X1 u_majority7_module_75__and_module_2_U1 ( .A1(
        n_majority7_module_75_n5), .A2(n_majority7_module_75_n3), .ZN(
        n_majority7_module_75__and_module_2_res) );
  OR2_X1 u_majority7_module_75__or_module_2_U1 ( .A1(n_majority7_module_75_n3), 
        .A2(n_majority7_module_75_n5), .ZN(
        n_majority7_module_75__or_module_2_res) );
  AND2_X1 u_majority7_module_75__and_module_3_U1 ( .A1(
        n_majority7_module_75_n6), .A2(n_majority7_module_75_n4), .ZN(
        n_majority7_module_75__and_module_3_res) );
  OR2_X1 u_majority7_module_75__or_module_3_U1 ( .A1(n_majority7_module_75_n4), 
        .A2(n_majority7_module_75_n6), .ZN(
        n_majority7_module_75__or_module_3_res) );
  AND2_X1 u_majority7_module_75__and_module_4_U1 ( .A1(
        n_majority7_module_75__and_module_2_res), .A2(
        n_majority7_module_75__and_module_1_res), .ZN(
        n_majority7_module_75__and_module_4_res) );
  OR2_X1 u_majority7_module_75__or_module_4_U1 ( .A1(
        n_majority7_module_75__and_module_1_res), .A2(
        n_majority7_module_75__and_module_2_res), .ZN(
        n_majority7_module_75__or_module_4_res) );
  AND2_X1 u_majority7_module_75__and_module_5_U1 ( .A1(
        n_majority7_module_75__and_module_3_res), .A2(n_majority7_module_75_n2), .ZN(n_majority7_module_75__and_module_5_res) );
  OR2_X1 u_majority7_module_75__or_module_5_U1 ( .A1(n_majority7_module_75_n2), 
        .A2(n_majority7_module_75__and_module_3_res), .ZN(
        n_majority7_module_75__or_module_5_res) );
  AND2_X1 u_majority7_module_75__and_module_6_U1 ( .A1(
        n_majority7_module_75__or_module_1_res), .A2(
        n_majority7_module_75__or_module_2_res), .ZN(
        n_majority7_module_75__and_module_6_res) );
  OR2_X1 u_majority7_module_75__or_module_6_U1 ( .A1(
        n_majority7_module_75__or_module_2_res), .A2(
        n_majority7_module_75__or_module_1_res), .ZN(
        n_majority7_module_75__or_module_6_res) );
  OR2_X1 u_majority7_module_75__or_module_7_U1 ( .A1(
        n_majority7_module_75__and_module_4_res), .A2(
        n_majority7_module_75__and_module_5_res), .ZN(
        n_majority7_module_75__or_module_7_res) );
  AND2_X1 u_majority7_module_75__and_module_7_U1 ( .A1(
        n_majority7_module_75__or_module_3_res), .A2(
        n_majority7_module_75__or_module_4_res), .ZN(
        n_majority7_module_75__and_module_7_res) );
  OR2_X1 u_majority7_module_75__or_module_8_U1 ( .A1(
        n_majority7_module_75__or_module_4_res), .A2(
        n_majority7_module_75__or_module_3_res), .ZN(
        n_majority7_module_75__or_module_8_res) );
  AND2_X1 u_majority7_module_75__and_module_8_U1 ( .A1(
        n_majority7_module_75__or_module_5_res), .A2(
        n_majority7_module_75__and_module_6_res), .ZN(
        n_majority7_module_75__and_module_8_res) );
  OR2_X1 u_majority7_module_75__or_module_9_U1 ( .A1(
        n_majority7_module_75__and_module_6_res), .A2(
        n_majority7_module_75__or_module_5_res), .ZN(
        n_majority7_module_75__or_module_9_res) );
  OR2_X1 u_majority7_module_75__or_module_10_U1 ( .A1(
        n_majority7_module_75__or_module_7_res), .A2(
        n_majority7_module_75__and_module_7_res), .ZN(
        n_majority7_module_75__or_module_10_res) );
  AND2_X1 u_majority7_module_75__and_module_9_U1 ( .A1(
        n_majority7_module_75__or_module_6_res), .A2(
        n_majority7_module_75__or_module_9_res), .ZN(
        n_majority7_module_75__and_module_9_res) );
  OR2_X1 u_majority7_module_75__or_module_11_U1 ( .A1(
        n_majority7_module_75__or_module_10_res), .A2(
        n_majority7_module_75__and_module_8_res), .ZN(
        n_majority7_module_75__or_module_11_res) );
  AND2_X1 u_majority7_module_75__and_module_10_U1 ( .A1(
        n_majority7_module_75__or_module_8_res), .A2(
        n_majority7_module_75__and_module_9_res), .ZN(
        n_majority7_module_75__and_module_10_res) );
  AND2_X1 u_majority7_module_75__and_module_11_U1 ( .A1(
        n_majority7_module_75__and_module_10_res), .A2(
        n_majority7_module_75__or_module_11_res), .ZN(
        n_majority7_module_75_res) );
  DFF_X1 u_reg_module_76__cini_mul_v000_reg ( .D(n_majority7_module_75_res), 
        .CK(clock_4), .Q(n_reg_module_76_res), .QN() );
  BUF_X1 u_majority7_module_76_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_76_n7) );
  BUF_X1 u_majority7_module_76_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_76_n6) );
  BUF_X1 u_majority7_module_76_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_76_n5) );
  BUF_X1 u_majority7_module_76_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_76_n4) );
  BUF_X1 u_majority7_module_76_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_76_n3) );
  BUF_X1 u_majority7_module_76_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_76_n2) );
  BUF_X1 u_majority7_module_76_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_76_n1) );
  AND2_X1 u_majority7_module_76__and_module_1_U1 ( .A1(
        n_majority7_module_76_n7), .A2(n_majority7_module_76_n1), .ZN(
        n_majority7_module_76__and_module_1_res) );
  OR2_X1 u_majority7_module_76__or_module_1_U1 ( .A1(n_majority7_module_76_n1), 
        .A2(n_majority7_module_76_n7), .ZN(
        n_majority7_module_76__or_module_1_res) );
  AND2_X1 u_majority7_module_76__and_module_2_U1 ( .A1(
        n_majority7_module_76_n5), .A2(n_majority7_module_76_n3), .ZN(
        n_majority7_module_76__and_module_2_res) );
  OR2_X1 u_majority7_module_76__or_module_2_U1 ( .A1(n_majority7_module_76_n3), 
        .A2(n_majority7_module_76_n5), .ZN(
        n_majority7_module_76__or_module_2_res) );
  AND2_X1 u_majority7_module_76__and_module_3_U1 ( .A1(
        n_majority7_module_76_n6), .A2(n_majority7_module_76_n4), .ZN(
        n_majority7_module_76__and_module_3_res) );
  OR2_X1 u_majority7_module_76__or_module_3_U1 ( .A1(n_majority7_module_76_n4), 
        .A2(n_majority7_module_76_n6), .ZN(
        n_majority7_module_76__or_module_3_res) );
  AND2_X1 u_majority7_module_76__and_module_4_U1 ( .A1(
        n_majority7_module_76__and_module_2_res), .A2(
        n_majority7_module_76__and_module_1_res), .ZN(
        n_majority7_module_76__and_module_4_res) );
  OR2_X1 u_majority7_module_76__or_module_4_U1 ( .A1(
        n_majority7_module_76__and_module_1_res), .A2(
        n_majority7_module_76__and_module_2_res), .ZN(
        n_majority7_module_76__or_module_4_res) );
  AND2_X1 u_majority7_module_76__and_module_5_U1 ( .A1(
        n_majority7_module_76__and_module_3_res), .A2(n_majority7_module_76_n2), .ZN(n_majority7_module_76__and_module_5_res) );
  OR2_X1 u_majority7_module_76__or_module_5_U1 ( .A1(n_majority7_module_76_n2), 
        .A2(n_majority7_module_76__and_module_3_res), .ZN(
        n_majority7_module_76__or_module_5_res) );
  AND2_X1 u_majority7_module_76__and_module_6_U1 ( .A1(
        n_majority7_module_76__or_module_1_res), .A2(
        n_majority7_module_76__or_module_2_res), .ZN(
        n_majority7_module_76__and_module_6_res) );
  OR2_X1 u_majority7_module_76__or_module_6_U1 ( .A1(
        n_majority7_module_76__or_module_2_res), .A2(
        n_majority7_module_76__or_module_1_res), .ZN(
        n_majority7_module_76__or_module_6_res) );
  OR2_X1 u_majority7_module_76__or_module_7_U1 ( .A1(
        n_majority7_module_76__and_module_4_res), .A2(
        n_majority7_module_76__and_module_5_res), .ZN(
        n_majority7_module_76__or_module_7_res) );
  AND2_X1 u_majority7_module_76__and_module_7_U1 ( .A1(
        n_majority7_module_76__or_module_3_res), .A2(
        n_majority7_module_76__or_module_4_res), .ZN(
        n_majority7_module_76__and_module_7_res) );
  OR2_X1 u_majority7_module_76__or_module_8_U1 ( .A1(
        n_majority7_module_76__or_module_4_res), .A2(
        n_majority7_module_76__or_module_3_res), .ZN(
        n_majority7_module_76__or_module_8_res) );
  AND2_X1 u_majority7_module_76__and_module_8_U1 ( .A1(
        n_majority7_module_76__or_module_5_res), .A2(
        n_majority7_module_76__and_module_6_res), .ZN(
        n_majority7_module_76__and_module_8_res) );
  OR2_X1 u_majority7_module_76__or_module_9_U1 ( .A1(
        n_majority7_module_76__and_module_6_res), .A2(
        n_majority7_module_76__or_module_5_res), .ZN(
        n_majority7_module_76__or_module_9_res) );
  OR2_X1 u_majority7_module_76__or_module_10_U1 ( .A1(
        n_majority7_module_76__or_module_7_res), .A2(
        n_majority7_module_76__and_module_7_res), .ZN(
        n_majority7_module_76__or_module_10_res) );
  AND2_X1 u_majority7_module_76__and_module_9_U1 ( .A1(
        n_majority7_module_76__or_module_6_res), .A2(
        n_majority7_module_76__or_module_9_res), .ZN(
        n_majority7_module_76__and_module_9_res) );
  OR2_X1 u_majority7_module_76__or_module_11_U1 ( .A1(
        n_majority7_module_76__or_module_10_res), .A2(
        n_majority7_module_76__and_module_8_res), .ZN(
        n_majority7_module_76__or_module_11_res) );
  AND2_X1 u_majority7_module_76__and_module_10_U1 ( .A1(
        n_majority7_module_76__or_module_8_res), .A2(
        n_majority7_module_76__and_module_9_res), .ZN(
        n_majority7_module_76__and_module_10_res) );
  AND2_X1 u_majority7_module_76__and_module_11_U1 ( .A1(
        n_majority7_module_76__and_module_10_res), .A2(
        n_majority7_module_76__or_module_11_res), .ZN(
        n_majority7_module_76_res) );
  DFF_X1 u_reg_module_77__cini_mul_v000_reg ( .D(n_majority7_module_76_res), 
        .CK(clock_4), .Q(n_reg_module_77_res), .QN() );
  BUF_X1 u_majority7_module_77_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_77_n7) );
  BUF_X1 u_majority7_module_77_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_77_n6) );
  BUF_X1 u_majority7_module_77_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_77_n5) );
  BUF_X1 u_majority7_module_77_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_77_n4) );
  BUF_X1 u_majority7_module_77_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_77_n3) );
  BUF_X1 u_majority7_module_77_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_77_n2) );
  BUF_X1 u_majority7_module_77_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_77_n1) );
  AND2_X1 u_majority7_module_77__and_module_1_U1 ( .A1(
        n_majority7_module_77_n7), .A2(n_majority7_module_77_n1), .ZN(
        n_majority7_module_77__and_module_1_res) );
  OR2_X1 u_majority7_module_77__or_module_1_U1 ( .A1(n_majority7_module_77_n1), 
        .A2(n_majority7_module_77_n7), .ZN(
        n_majority7_module_77__or_module_1_res) );
  AND2_X1 u_majority7_module_77__and_module_2_U1 ( .A1(
        n_majority7_module_77_n5), .A2(n_majority7_module_77_n3), .ZN(
        n_majority7_module_77__and_module_2_res) );
  OR2_X1 u_majority7_module_77__or_module_2_U1 ( .A1(n_majority7_module_77_n3), 
        .A2(n_majority7_module_77_n5), .ZN(
        n_majority7_module_77__or_module_2_res) );
  AND2_X1 u_majority7_module_77__and_module_3_U1 ( .A1(
        n_majority7_module_77_n6), .A2(n_majority7_module_77_n4), .ZN(
        n_majority7_module_77__and_module_3_res) );
  OR2_X1 u_majority7_module_77__or_module_3_U1 ( .A1(n_majority7_module_77_n4), 
        .A2(n_majority7_module_77_n6), .ZN(
        n_majority7_module_77__or_module_3_res) );
  AND2_X1 u_majority7_module_77__and_module_4_U1 ( .A1(
        n_majority7_module_77__and_module_2_res), .A2(
        n_majority7_module_77__and_module_1_res), .ZN(
        n_majority7_module_77__and_module_4_res) );
  OR2_X1 u_majority7_module_77__or_module_4_U1 ( .A1(
        n_majority7_module_77__and_module_1_res), .A2(
        n_majority7_module_77__and_module_2_res), .ZN(
        n_majority7_module_77__or_module_4_res) );
  AND2_X1 u_majority7_module_77__and_module_5_U1 ( .A1(
        n_majority7_module_77__and_module_3_res), .A2(n_majority7_module_77_n2), .ZN(n_majority7_module_77__and_module_5_res) );
  OR2_X1 u_majority7_module_77__or_module_5_U1 ( .A1(n_majority7_module_77_n2), 
        .A2(n_majority7_module_77__and_module_3_res), .ZN(
        n_majority7_module_77__or_module_5_res) );
  AND2_X1 u_majority7_module_77__and_module_6_U1 ( .A1(
        n_majority7_module_77__or_module_1_res), .A2(
        n_majority7_module_77__or_module_2_res), .ZN(
        n_majority7_module_77__and_module_6_res) );
  OR2_X1 u_majority7_module_77__or_module_6_U1 ( .A1(
        n_majority7_module_77__or_module_2_res), .A2(
        n_majority7_module_77__or_module_1_res), .ZN(
        n_majority7_module_77__or_module_6_res) );
  OR2_X1 u_majority7_module_77__or_module_7_U1 ( .A1(
        n_majority7_module_77__and_module_4_res), .A2(
        n_majority7_module_77__and_module_5_res), .ZN(
        n_majority7_module_77__or_module_7_res) );
  AND2_X1 u_majority7_module_77__and_module_7_U1 ( .A1(
        n_majority7_module_77__or_module_3_res), .A2(
        n_majority7_module_77__or_module_4_res), .ZN(
        n_majority7_module_77__and_module_7_res) );
  OR2_X1 u_majority7_module_77__or_module_8_U1 ( .A1(
        n_majority7_module_77__or_module_4_res), .A2(
        n_majority7_module_77__or_module_3_res), .ZN(
        n_majority7_module_77__or_module_8_res) );
  AND2_X1 u_majority7_module_77__and_module_8_U1 ( .A1(
        n_majority7_module_77__or_module_5_res), .A2(
        n_majority7_module_77__and_module_6_res), .ZN(
        n_majority7_module_77__and_module_8_res) );
  OR2_X1 u_majority7_module_77__or_module_9_U1 ( .A1(
        n_majority7_module_77__and_module_6_res), .A2(
        n_majority7_module_77__or_module_5_res), .ZN(
        n_majority7_module_77__or_module_9_res) );
  OR2_X1 u_majority7_module_77__or_module_10_U1 ( .A1(
        n_majority7_module_77__or_module_7_res), .A2(
        n_majority7_module_77__and_module_7_res), .ZN(
        n_majority7_module_77__or_module_10_res) );
  AND2_X1 u_majority7_module_77__and_module_9_U1 ( .A1(
        n_majority7_module_77__or_module_6_res), .A2(
        n_majority7_module_77__or_module_9_res), .ZN(
        n_majority7_module_77__and_module_9_res) );
  OR2_X1 u_majority7_module_77__or_module_11_U1 ( .A1(
        n_majority7_module_77__or_module_10_res), .A2(
        n_majority7_module_77__and_module_8_res), .ZN(
        n_majority7_module_77__or_module_11_res) );
  AND2_X1 u_majority7_module_77__and_module_10_U1 ( .A1(
        n_majority7_module_77__or_module_8_res), .A2(
        n_majority7_module_77__and_module_9_res), .ZN(
        n_majority7_module_77__and_module_10_res) );
  AND2_X1 u_majority7_module_77__and_module_11_U1 ( .A1(
        n_majority7_module_77__and_module_10_res), .A2(
        n_majority7_module_77__or_module_11_res), .ZN(
        n_majority7_module_77_res) );
  DFF_X1 u_reg_module_78__cini_mul_v000_reg ( .D(n_majority7_module_77_res), 
        .CK(clock_4), .Q(n_reg_module_78_res), .QN() );
  BUF_X1 u_majority7_module_78_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_78_n7) );
  BUF_X1 u_majority7_module_78_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_78_n6) );
  BUF_X1 u_majority7_module_78_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_78_n5) );
  BUF_X1 u_majority7_module_78_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_78_n4) );
  BUF_X1 u_majority7_module_78_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_78_n3) );
  BUF_X1 u_majority7_module_78_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_78_n2) );
  BUF_X1 u_majority7_module_78_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_78_n1) );
  AND2_X1 u_majority7_module_78__and_module_1_U1 ( .A1(
        n_majority7_module_78_n7), .A2(n_majority7_module_78_n1), .ZN(
        n_majority7_module_78__and_module_1_res) );
  OR2_X1 u_majority7_module_78__or_module_1_U1 ( .A1(n_majority7_module_78_n1), 
        .A2(n_majority7_module_78_n7), .ZN(
        n_majority7_module_78__or_module_1_res) );
  AND2_X1 u_majority7_module_78__and_module_2_U1 ( .A1(
        n_majority7_module_78_n5), .A2(n_majority7_module_78_n3), .ZN(
        n_majority7_module_78__and_module_2_res) );
  OR2_X1 u_majority7_module_78__or_module_2_U1 ( .A1(n_majority7_module_78_n3), 
        .A2(n_majority7_module_78_n5), .ZN(
        n_majority7_module_78__or_module_2_res) );
  AND2_X1 u_majority7_module_78__and_module_3_U1 ( .A1(
        n_majority7_module_78_n6), .A2(n_majority7_module_78_n4), .ZN(
        n_majority7_module_78__and_module_3_res) );
  OR2_X1 u_majority7_module_78__or_module_3_U1 ( .A1(n_majority7_module_78_n4), 
        .A2(n_majority7_module_78_n6), .ZN(
        n_majority7_module_78__or_module_3_res) );
  AND2_X1 u_majority7_module_78__and_module_4_U1 ( .A1(
        n_majority7_module_78__and_module_2_res), .A2(
        n_majority7_module_78__and_module_1_res), .ZN(
        n_majority7_module_78__and_module_4_res) );
  OR2_X1 u_majority7_module_78__or_module_4_U1 ( .A1(
        n_majority7_module_78__and_module_1_res), .A2(
        n_majority7_module_78__and_module_2_res), .ZN(
        n_majority7_module_78__or_module_4_res) );
  AND2_X1 u_majority7_module_78__and_module_5_U1 ( .A1(
        n_majority7_module_78__and_module_3_res), .A2(n_majority7_module_78_n2), .ZN(n_majority7_module_78__and_module_5_res) );
  OR2_X1 u_majority7_module_78__or_module_5_U1 ( .A1(n_majority7_module_78_n2), 
        .A2(n_majority7_module_78__and_module_3_res), .ZN(
        n_majority7_module_78__or_module_5_res) );
  AND2_X1 u_majority7_module_78__and_module_6_U1 ( .A1(
        n_majority7_module_78__or_module_1_res), .A2(
        n_majority7_module_78__or_module_2_res), .ZN(
        n_majority7_module_78__and_module_6_res) );
  OR2_X1 u_majority7_module_78__or_module_6_U1 ( .A1(
        n_majority7_module_78__or_module_2_res), .A2(
        n_majority7_module_78__or_module_1_res), .ZN(
        n_majority7_module_78__or_module_6_res) );
  OR2_X1 u_majority7_module_78__or_module_7_U1 ( .A1(
        n_majority7_module_78__and_module_4_res), .A2(
        n_majority7_module_78__and_module_5_res), .ZN(
        n_majority7_module_78__or_module_7_res) );
  AND2_X1 u_majority7_module_78__and_module_7_U1 ( .A1(
        n_majority7_module_78__or_module_3_res), .A2(
        n_majority7_module_78__or_module_4_res), .ZN(
        n_majority7_module_78__and_module_7_res) );
  OR2_X1 u_majority7_module_78__or_module_8_U1 ( .A1(
        n_majority7_module_78__or_module_4_res), .A2(
        n_majority7_module_78__or_module_3_res), .ZN(
        n_majority7_module_78__or_module_8_res) );
  AND2_X1 u_majority7_module_78__and_module_8_U1 ( .A1(
        n_majority7_module_78__or_module_5_res), .A2(
        n_majority7_module_78__and_module_6_res), .ZN(
        n_majority7_module_78__and_module_8_res) );
  OR2_X1 u_majority7_module_78__or_module_9_U1 ( .A1(
        n_majority7_module_78__and_module_6_res), .A2(
        n_majority7_module_78__or_module_5_res), .ZN(
        n_majority7_module_78__or_module_9_res) );
  OR2_X1 u_majority7_module_78__or_module_10_U1 ( .A1(
        n_majority7_module_78__or_module_7_res), .A2(
        n_majority7_module_78__and_module_7_res), .ZN(
        n_majority7_module_78__or_module_10_res) );
  AND2_X1 u_majority7_module_78__and_module_9_U1 ( .A1(
        n_majority7_module_78__or_module_6_res), .A2(
        n_majority7_module_78__or_module_9_res), .ZN(
        n_majority7_module_78__and_module_9_res) );
  OR2_X1 u_majority7_module_78__or_module_11_U1 ( .A1(
        n_majority7_module_78__or_module_10_res), .A2(
        n_majority7_module_78__and_module_8_res), .ZN(
        n_majority7_module_78__or_module_11_res) );
  AND2_X1 u_majority7_module_78__and_module_10_U1 ( .A1(
        n_majority7_module_78__or_module_8_res), .A2(
        n_majority7_module_78__and_module_9_res), .ZN(
        n_majority7_module_78__and_module_10_res) );
  AND2_X1 u_majority7_module_78__and_module_11_U1 ( .A1(
        n_majority7_module_78__and_module_10_res), .A2(
        n_majority7_module_78__or_module_11_res), .ZN(
        n_majority7_module_78_res) );
  DFF_X1 u_reg_module_79__cini_mul_v000_reg ( .D(n_majority7_module_78_res), 
        .CK(clock_4), .Q(n_reg_module_79_res), .QN() );
  BUF_X1 u_majority7_module_79_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_79_n7) );
  BUF_X1 u_majority7_module_79_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_79_n6) );
  BUF_X1 u_majority7_module_79_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_79_n5) );
  BUF_X1 u_majority7_module_79_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_79_n4) );
  BUF_X1 u_majority7_module_79_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_79_n3) );
  BUF_X1 u_majority7_module_79_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_79_n2) );
  BUF_X1 u_majority7_module_79_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_79_n1) );
  AND2_X1 u_majority7_module_79__and_module_1_U1 ( .A1(
        n_majority7_module_79_n7), .A2(n_majority7_module_79_n1), .ZN(
        n_majority7_module_79__and_module_1_res) );
  OR2_X1 u_majority7_module_79__or_module_1_U1 ( .A1(n_majority7_module_79_n1), 
        .A2(n_majority7_module_79_n7), .ZN(
        n_majority7_module_79__or_module_1_res) );
  AND2_X1 u_majority7_module_79__and_module_2_U1 ( .A1(
        n_majority7_module_79_n5), .A2(n_majority7_module_79_n3), .ZN(
        n_majority7_module_79__and_module_2_res) );
  OR2_X1 u_majority7_module_79__or_module_2_U1 ( .A1(n_majority7_module_79_n3), 
        .A2(n_majority7_module_79_n5), .ZN(
        n_majority7_module_79__or_module_2_res) );
  AND2_X1 u_majority7_module_79__and_module_3_U1 ( .A1(
        n_majority7_module_79_n6), .A2(n_majority7_module_79_n4), .ZN(
        n_majority7_module_79__and_module_3_res) );
  OR2_X1 u_majority7_module_79__or_module_3_U1 ( .A1(n_majority7_module_79_n4), 
        .A2(n_majority7_module_79_n6), .ZN(
        n_majority7_module_79__or_module_3_res) );
  AND2_X1 u_majority7_module_79__and_module_4_U1 ( .A1(
        n_majority7_module_79__and_module_2_res), .A2(
        n_majority7_module_79__and_module_1_res), .ZN(
        n_majority7_module_79__and_module_4_res) );
  OR2_X1 u_majority7_module_79__or_module_4_U1 ( .A1(
        n_majority7_module_79__and_module_1_res), .A2(
        n_majority7_module_79__and_module_2_res), .ZN(
        n_majority7_module_79__or_module_4_res) );
  AND2_X1 u_majority7_module_79__and_module_5_U1 ( .A1(
        n_majority7_module_79__and_module_3_res), .A2(n_majority7_module_79_n2), .ZN(n_majority7_module_79__and_module_5_res) );
  OR2_X1 u_majority7_module_79__or_module_5_U1 ( .A1(n_majority7_module_79_n2), 
        .A2(n_majority7_module_79__and_module_3_res), .ZN(
        n_majority7_module_79__or_module_5_res) );
  AND2_X1 u_majority7_module_79__and_module_6_U1 ( .A1(
        n_majority7_module_79__or_module_1_res), .A2(
        n_majority7_module_79__or_module_2_res), .ZN(
        n_majority7_module_79__and_module_6_res) );
  OR2_X1 u_majority7_module_79__or_module_6_U1 ( .A1(
        n_majority7_module_79__or_module_2_res), .A2(
        n_majority7_module_79__or_module_1_res), .ZN(
        n_majority7_module_79__or_module_6_res) );
  OR2_X1 u_majority7_module_79__or_module_7_U1 ( .A1(
        n_majority7_module_79__and_module_4_res), .A2(
        n_majority7_module_79__and_module_5_res), .ZN(
        n_majority7_module_79__or_module_7_res) );
  AND2_X1 u_majority7_module_79__and_module_7_U1 ( .A1(
        n_majority7_module_79__or_module_3_res), .A2(
        n_majority7_module_79__or_module_4_res), .ZN(
        n_majority7_module_79__and_module_7_res) );
  OR2_X1 u_majority7_module_79__or_module_8_U1 ( .A1(
        n_majority7_module_79__or_module_4_res), .A2(
        n_majority7_module_79__or_module_3_res), .ZN(
        n_majority7_module_79__or_module_8_res) );
  AND2_X1 u_majority7_module_79__and_module_8_U1 ( .A1(
        n_majority7_module_79__or_module_5_res), .A2(
        n_majority7_module_79__and_module_6_res), .ZN(
        n_majority7_module_79__and_module_8_res) );
  OR2_X1 u_majority7_module_79__or_module_9_U1 ( .A1(
        n_majority7_module_79__and_module_6_res), .A2(
        n_majority7_module_79__or_module_5_res), .ZN(
        n_majority7_module_79__or_module_9_res) );
  OR2_X1 u_majority7_module_79__or_module_10_U1 ( .A1(
        n_majority7_module_79__or_module_7_res), .A2(
        n_majority7_module_79__and_module_7_res), .ZN(
        n_majority7_module_79__or_module_10_res) );
  AND2_X1 u_majority7_module_79__and_module_9_U1 ( .A1(
        n_majority7_module_79__or_module_6_res), .A2(
        n_majority7_module_79__or_module_9_res), .ZN(
        n_majority7_module_79__and_module_9_res) );
  OR2_X1 u_majority7_module_79__or_module_11_U1 ( .A1(
        n_majority7_module_79__or_module_10_res), .A2(
        n_majority7_module_79__and_module_8_res), .ZN(
        n_majority7_module_79__or_module_11_res) );
  AND2_X1 u_majority7_module_79__and_module_10_U1 ( .A1(
        n_majority7_module_79__or_module_8_res), .A2(
        n_majority7_module_79__and_module_9_res), .ZN(
        n_majority7_module_79__and_module_10_res) );
  AND2_X1 u_majority7_module_79__and_module_11_U1 ( .A1(
        n_majority7_module_79__and_module_10_res), .A2(
        n_majority7_module_79__or_module_11_res), .ZN(
        n_majority7_module_79_res) );
  DFF_X1 u_reg_module_80__cini_mul_v000_reg ( .D(n_majority7_module_79_res), 
        .CK(clock_4), .Q(n_reg_module_80_res), .QN() );
  BUF_X1 u_majority7_module_80_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_80_n7) );
  BUF_X1 u_majority7_module_80_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_80_n6) );
  BUF_X1 u_majority7_module_80_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_80_n5) );
  BUF_X1 u_majority7_module_80_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_80_n4) );
  BUF_X1 u_majority7_module_80_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_80_n3) );
  BUF_X1 u_majority7_module_80_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_80_n2) );
  BUF_X1 u_majority7_module_80_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_80_n1) );
  AND2_X1 u_majority7_module_80__and_module_1_U1 ( .A1(
        n_majority7_module_80_n7), .A2(n_majority7_module_80_n1), .ZN(
        n_majority7_module_80__and_module_1_res) );
  OR2_X1 u_majority7_module_80__or_module_1_U1 ( .A1(n_majority7_module_80_n1), 
        .A2(n_majority7_module_80_n7), .ZN(
        n_majority7_module_80__or_module_1_res) );
  AND2_X1 u_majority7_module_80__and_module_2_U1 ( .A1(
        n_majority7_module_80_n5), .A2(n_majority7_module_80_n3), .ZN(
        n_majority7_module_80__and_module_2_res) );
  OR2_X1 u_majority7_module_80__or_module_2_U1 ( .A1(n_majority7_module_80_n3), 
        .A2(n_majority7_module_80_n5), .ZN(
        n_majority7_module_80__or_module_2_res) );
  AND2_X1 u_majority7_module_80__and_module_3_U1 ( .A1(
        n_majority7_module_80_n6), .A2(n_majority7_module_80_n4), .ZN(
        n_majority7_module_80__and_module_3_res) );
  OR2_X1 u_majority7_module_80__or_module_3_U1 ( .A1(n_majority7_module_80_n4), 
        .A2(n_majority7_module_80_n6), .ZN(
        n_majority7_module_80__or_module_3_res) );
  AND2_X1 u_majority7_module_80__and_module_4_U1 ( .A1(
        n_majority7_module_80__and_module_2_res), .A2(
        n_majority7_module_80__and_module_1_res), .ZN(
        n_majority7_module_80__and_module_4_res) );
  OR2_X1 u_majority7_module_80__or_module_4_U1 ( .A1(
        n_majority7_module_80__and_module_1_res), .A2(
        n_majority7_module_80__and_module_2_res), .ZN(
        n_majority7_module_80__or_module_4_res) );
  AND2_X1 u_majority7_module_80__and_module_5_U1 ( .A1(
        n_majority7_module_80__and_module_3_res), .A2(n_majority7_module_80_n2), .ZN(n_majority7_module_80__and_module_5_res) );
  OR2_X1 u_majority7_module_80__or_module_5_U1 ( .A1(n_majority7_module_80_n2), 
        .A2(n_majority7_module_80__and_module_3_res), .ZN(
        n_majority7_module_80__or_module_5_res) );
  AND2_X1 u_majority7_module_80__and_module_6_U1 ( .A1(
        n_majority7_module_80__or_module_1_res), .A2(
        n_majority7_module_80__or_module_2_res), .ZN(
        n_majority7_module_80__and_module_6_res) );
  OR2_X1 u_majority7_module_80__or_module_6_U1 ( .A1(
        n_majority7_module_80__or_module_2_res), .A2(
        n_majority7_module_80__or_module_1_res), .ZN(
        n_majority7_module_80__or_module_6_res) );
  OR2_X1 u_majority7_module_80__or_module_7_U1 ( .A1(
        n_majority7_module_80__and_module_4_res), .A2(
        n_majority7_module_80__and_module_5_res), .ZN(
        n_majority7_module_80__or_module_7_res) );
  AND2_X1 u_majority7_module_80__and_module_7_U1 ( .A1(
        n_majority7_module_80__or_module_3_res), .A2(
        n_majority7_module_80__or_module_4_res), .ZN(
        n_majority7_module_80__and_module_7_res) );
  OR2_X1 u_majority7_module_80__or_module_8_U1 ( .A1(
        n_majority7_module_80__or_module_4_res), .A2(
        n_majority7_module_80__or_module_3_res), .ZN(
        n_majority7_module_80__or_module_8_res) );
  AND2_X1 u_majority7_module_80__and_module_8_U1 ( .A1(
        n_majority7_module_80__or_module_5_res), .A2(
        n_majority7_module_80__and_module_6_res), .ZN(
        n_majority7_module_80__and_module_8_res) );
  OR2_X1 u_majority7_module_80__or_module_9_U1 ( .A1(
        n_majority7_module_80__and_module_6_res), .A2(
        n_majority7_module_80__or_module_5_res), .ZN(
        n_majority7_module_80__or_module_9_res) );
  OR2_X1 u_majority7_module_80__or_module_10_U1 ( .A1(
        n_majority7_module_80__or_module_7_res), .A2(
        n_majority7_module_80__and_module_7_res), .ZN(
        n_majority7_module_80__or_module_10_res) );
  AND2_X1 u_majority7_module_80__and_module_9_U1 ( .A1(
        n_majority7_module_80__or_module_6_res), .A2(
        n_majority7_module_80__or_module_9_res), .ZN(
        n_majority7_module_80__and_module_9_res) );
  OR2_X1 u_majority7_module_80__or_module_11_U1 ( .A1(
        n_majority7_module_80__or_module_10_res), .A2(
        n_majority7_module_80__and_module_8_res), .ZN(
        n_majority7_module_80__or_module_11_res) );
  AND2_X1 u_majority7_module_80__and_module_10_U1 ( .A1(
        n_majority7_module_80__or_module_8_res), .A2(
        n_majority7_module_80__and_module_9_res), .ZN(
        n_majority7_module_80__and_module_10_res) );
  AND2_X1 u_majority7_module_80__and_module_11_U1 ( .A1(
        n_majority7_module_80__and_module_10_res), .A2(
        n_majority7_module_80__or_module_11_res), .ZN(
        n_majority7_module_80_res) );
  DFF_X1 u_reg_module_81__cini_mul_v000_reg ( .D(n_majority7_module_80_res), 
        .CK(clock_5), .Q(n_reg_module_81_res), .QN() );
  BUF_X1 u_majority7_module_81_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_81_n7) );
  BUF_X1 u_majority7_module_81_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_81_n6) );
  BUF_X1 u_majority7_module_81_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_81_n5) );
  BUF_X1 u_majority7_module_81_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_81_n4) );
  BUF_X1 u_majority7_module_81_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_81_n3) );
  BUF_X1 u_majority7_module_81_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_81_n2) );
  BUF_X1 u_majority7_module_81_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_81_n1) );
  AND2_X1 u_majority7_module_81__and_module_1_U1 ( .A1(
        n_majority7_module_81_n7), .A2(n_majority7_module_81_n1), .ZN(
        n_majority7_module_81__and_module_1_res) );
  OR2_X1 u_majority7_module_81__or_module_1_U1 ( .A1(n_majority7_module_81_n1), 
        .A2(n_majority7_module_81_n7), .ZN(
        n_majority7_module_81__or_module_1_res) );
  AND2_X1 u_majority7_module_81__and_module_2_U1 ( .A1(
        n_majority7_module_81_n5), .A2(n_majority7_module_81_n3), .ZN(
        n_majority7_module_81__and_module_2_res) );
  OR2_X1 u_majority7_module_81__or_module_2_U1 ( .A1(n_majority7_module_81_n3), 
        .A2(n_majority7_module_81_n5), .ZN(
        n_majority7_module_81__or_module_2_res) );
  AND2_X1 u_majority7_module_81__and_module_3_U1 ( .A1(
        n_majority7_module_81_n6), .A2(n_majority7_module_81_n4), .ZN(
        n_majority7_module_81__and_module_3_res) );
  OR2_X1 u_majority7_module_81__or_module_3_U1 ( .A1(n_majority7_module_81_n4), 
        .A2(n_majority7_module_81_n6), .ZN(
        n_majority7_module_81__or_module_3_res) );
  AND2_X1 u_majority7_module_81__and_module_4_U1 ( .A1(
        n_majority7_module_81__and_module_2_res), .A2(
        n_majority7_module_81__and_module_1_res), .ZN(
        n_majority7_module_81__and_module_4_res) );
  OR2_X1 u_majority7_module_81__or_module_4_U1 ( .A1(
        n_majority7_module_81__and_module_1_res), .A2(
        n_majority7_module_81__and_module_2_res), .ZN(
        n_majority7_module_81__or_module_4_res) );
  AND2_X1 u_majority7_module_81__and_module_5_U1 ( .A1(
        n_majority7_module_81__and_module_3_res), .A2(n_majority7_module_81_n2), .ZN(n_majority7_module_81__and_module_5_res) );
  OR2_X1 u_majority7_module_81__or_module_5_U1 ( .A1(n_majority7_module_81_n2), 
        .A2(n_majority7_module_81__and_module_3_res), .ZN(
        n_majority7_module_81__or_module_5_res) );
  AND2_X1 u_majority7_module_81__and_module_6_U1 ( .A1(
        n_majority7_module_81__or_module_1_res), .A2(
        n_majority7_module_81__or_module_2_res), .ZN(
        n_majority7_module_81__and_module_6_res) );
  OR2_X1 u_majority7_module_81__or_module_6_U1 ( .A1(
        n_majority7_module_81__or_module_2_res), .A2(
        n_majority7_module_81__or_module_1_res), .ZN(
        n_majority7_module_81__or_module_6_res) );
  OR2_X1 u_majority7_module_81__or_module_7_U1 ( .A1(
        n_majority7_module_81__and_module_4_res), .A2(
        n_majority7_module_81__and_module_5_res), .ZN(
        n_majority7_module_81__or_module_7_res) );
  AND2_X1 u_majority7_module_81__and_module_7_U1 ( .A1(
        n_majority7_module_81__or_module_3_res), .A2(
        n_majority7_module_81__or_module_4_res), .ZN(
        n_majority7_module_81__and_module_7_res) );
  OR2_X1 u_majority7_module_81__or_module_8_U1 ( .A1(
        n_majority7_module_81__or_module_4_res), .A2(
        n_majority7_module_81__or_module_3_res), .ZN(
        n_majority7_module_81__or_module_8_res) );
  AND2_X1 u_majority7_module_81__and_module_8_U1 ( .A1(
        n_majority7_module_81__or_module_5_res), .A2(
        n_majority7_module_81__and_module_6_res), .ZN(
        n_majority7_module_81__and_module_8_res) );
  OR2_X1 u_majority7_module_81__or_module_9_U1 ( .A1(
        n_majority7_module_81__and_module_6_res), .A2(
        n_majority7_module_81__or_module_5_res), .ZN(
        n_majority7_module_81__or_module_9_res) );
  OR2_X1 u_majority7_module_81__or_module_10_U1 ( .A1(
        n_majority7_module_81__or_module_7_res), .A2(
        n_majority7_module_81__and_module_7_res), .ZN(
        n_majority7_module_81__or_module_10_res) );
  AND2_X1 u_majority7_module_81__and_module_9_U1 ( .A1(
        n_majority7_module_81__or_module_6_res), .A2(
        n_majority7_module_81__or_module_9_res), .ZN(
        n_majority7_module_81__and_module_9_res) );
  OR2_X1 u_majority7_module_81__or_module_11_U1 ( .A1(
        n_majority7_module_81__or_module_10_res), .A2(
        n_majority7_module_81__and_module_8_res), .ZN(
        n_majority7_module_81__or_module_11_res) );
  AND2_X1 u_majority7_module_81__and_module_10_U1 ( .A1(
        n_majority7_module_81__or_module_8_res), .A2(
        n_majority7_module_81__and_module_9_res), .ZN(
        n_majority7_module_81__and_module_10_res) );
  AND2_X1 u_majority7_module_81__and_module_11_U1 ( .A1(
        n_majority7_module_81__and_module_10_res), .A2(
        n_majority7_module_81__or_module_11_res), .ZN(
        n_majority7_module_81_res) );
  DFF_X1 u_reg_module_82__cini_mul_v000_reg ( .D(n_majority7_module_81_res), 
        .CK(clock_5), .Q(n_reg_module_82_res), .QN() );
  BUF_X1 u_majority7_module_82_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_82_n7) );
  BUF_X1 u_majority7_module_82_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_82_n6) );
  BUF_X1 u_majority7_module_82_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_82_n5) );
  BUF_X1 u_majority7_module_82_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_82_n4) );
  BUF_X1 u_majority7_module_82_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_82_n3) );
  BUF_X1 u_majority7_module_82_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_82_n2) );
  BUF_X1 u_majority7_module_82_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_82_n1) );
  AND2_X1 u_majority7_module_82__and_module_1_U1 ( .A1(
        n_majority7_module_82_n7), .A2(n_majority7_module_82_n1), .ZN(
        n_majority7_module_82__and_module_1_res) );
  OR2_X1 u_majority7_module_82__or_module_1_U1 ( .A1(n_majority7_module_82_n1), 
        .A2(n_majority7_module_82_n7), .ZN(
        n_majority7_module_82__or_module_1_res) );
  AND2_X1 u_majority7_module_82__and_module_2_U1 ( .A1(
        n_majority7_module_82_n5), .A2(n_majority7_module_82_n3), .ZN(
        n_majority7_module_82__and_module_2_res) );
  OR2_X1 u_majority7_module_82__or_module_2_U1 ( .A1(n_majority7_module_82_n3), 
        .A2(n_majority7_module_82_n5), .ZN(
        n_majority7_module_82__or_module_2_res) );
  AND2_X1 u_majority7_module_82__and_module_3_U1 ( .A1(
        n_majority7_module_82_n6), .A2(n_majority7_module_82_n4), .ZN(
        n_majority7_module_82__and_module_3_res) );
  OR2_X1 u_majority7_module_82__or_module_3_U1 ( .A1(n_majority7_module_82_n4), 
        .A2(n_majority7_module_82_n6), .ZN(
        n_majority7_module_82__or_module_3_res) );
  AND2_X1 u_majority7_module_82__and_module_4_U1 ( .A1(
        n_majority7_module_82__and_module_2_res), .A2(
        n_majority7_module_82__and_module_1_res), .ZN(
        n_majority7_module_82__and_module_4_res) );
  OR2_X1 u_majority7_module_82__or_module_4_U1 ( .A1(
        n_majority7_module_82__and_module_1_res), .A2(
        n_majority7_module_82__and_module_2_res), .ZN(
        n_majority7_module_82__or_module_4_res) );
  AND2_X1 u_majority7_module_82__and_module_5_U1 ( .A1(
        n_majority7_module_82__and_module_3_res), .A2(n_majority7_module_82_n2), .ZN(n_majority7_module_82__and_module_5_res) );
  OR2_X1 u_majority7_module_82__or_module_5_U1 ( .A1(n_majority7_module_82_n2), 
        .A2(n_majority7_module_82__and_module_3_res), .ZN(
        n_majority7_module_82__or_module_5_res) );
  AND2_X1 u_majority7_module_82__and_module_6_U1 ( .A1(
        n_majority7_module_82__or_module_1_res), .A2(
        n_majority7_module_82__or_module_2_res), .ZN(
        n_majority7_module_82__and_module_6_res) );
  OR2_X1 u_majority7_module_82__or_module_6_U1 ( .A1(
        n_majority7_module_82__or_module_2_res), .A2(
        n_majority7_module_82__or_module_1_res), .ZN(
        n_majority7_module_82__or_module_6_res) );
  OR2_X1 u_majority7_module_82__or_module_7_U1 ( .A1(
        n_majority7_module_82__and_module_4_res), .A2(
        n_majority7_module_82__and_module_5_res), .ZN(
        n_majority7_module_82__or_module_7_res) );
  AND2_X1 u_majority7_module_82__and_module_7_U1 ( .A1(
        n_majority7_module_82__or_module_3_res), .A2(
        n_majority7_module_82__or_module_4_res), .ZN(
        n_majority7_module_82__and_module_7_res) );
  OR2_X1 u_majority7_module_82__or_module_8_U1 ( .A1(
        n_majority7_module_82__or_module_4_res), .A2(
        n_majority7_module_82__or_module_3_res), .ZN(
        n_majority7_module_82__or_module_8_res) );
  AND2_X1 u_majority7_module_82__and_module_8_U1 ( .A1(
        n_majority7_module_82__or_module_5_res), .A2(
        n_majority7_module_82__and_module_6_res), .ZN(
        n_majority7_module_82__and_module_8_res) );
  OR2_X1 u_majority7_module_82__or_module_9_U1 ( .A1(
        n_majority7_module_82__and_module_6_res), .A2(
        n_majority7_module_82__or_module_5_res), .ZN(
        n_majority7_module_82__or_module_9_res) );
  OR2_X1 u_majority7_module_82__or_module_10_U1 ( .A1(
        n_majority7_module_82__or_module_7_res), .A2(
        n_majority7_module_82__and_module_7_res), .ZN(
        n_majority7_module_82__or_module_10_res) );
  AND2_X1 u_majority7_module_82__and_module_9_U1 ( .A1(
        n_majority7_module_82__or_module_6_res), .A2(
        n_majority7_module_82__or_module_9_res), .ZN(
        n_majority7_module_82__and_module_9_res) );
  OR2_X1 u_majority7_module_82__or_module_11_U1 ( .A1(
        n_majority7_module_82__or_module_10_res), .A2(
        n_majority7_module_82__and_module_8_res), .ZN(
        n_majority7_module_82__or_module_11_res) );
  AND2_X1 u_majority7_module_82__and_module_10_U1 ( .A1(
        n_majority7_module_82__or_module_8_res), .A2(
        n_majority7_module_82__and_module_9_res), .ZN(
        n_majority7_module_82__and_module_10_res) );
  AND2_X1 u_majority7_module_82__and_module_11_U1 ( .A1(
        n_majority7_module_82__and_module_10_res), .A2(
        n_majority7_module_82__or_module_11_res), .ZN(
        n_majority7_module_82_res) );
  DFF_X1 u_reg_module_83__cini_mul_v000_reg ( .D(n_majority7_module_82_res), 
        .CK(clock_5), .Q(n_reg_module_83_res), .QN() );
  BUF_X1 u_majority7_module_83_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_83_n7) );
  BUF_X1 u_majority7_module_83_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_83_n6) );
  BUF_X1 u_majority7_module_83_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_83_n5) );
  BUF_X1 u_majority7_module_83_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_83_n4) );
  BUF_X1 u_majority7_module_83_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_83_n3) );
  BUF_X1 u_majority7_module_83_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_83_n2) );
  BUF_X1 u_majority7_module_83_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_83_n1) );
  AND2_X1 u_majority7_module_83__and_module_1_U1 ( .A1(
        n_majority7_module_83_n7), .A2(n_majority7_module_83_n1), .ZN(
        n_majority7_module_83__and_module_1_res) );
  OR2_X1 u_majority7_module_83__or_module_1_U1 ( .A1(n_majority7_module_83_n1), 
        .A2(n_majority7_module_83_n7), .ZN(
        n_majority7_module_83__or_module_1_res) );
  AND2_X1 u_majority7_module_83__and_module_2_U1 ( .A1(
        n_majority7_module_83_n5), .A2(n_majority7_module_83_n3), .ZN(
        n_majority7_module_83__and_module_2_res) );
  OR2_X1 u_majority7_module_83__or_module_2_U1 ( .A1(n_majority7_module_83_n3), 
        .A2(n_majority7_module_83_n5), .ZN(
        n_majority7_module_83__or_module_2_res) );
  AND2_X1 u_majority7_module_83__and_module_3_U1 ( .A1(
        n_majority7_module_83_n6), .A2(n_majority7_module_83_n4), .ZN(
        n_majority7_module_83__and_module_3_res) );
  OR2_X1 u_majority7_module_83__or_module_3_U1 ( .A1(n_majority7_module_83_n4), 
        .A2(n_majority7_module_83_n6), .ZN(
        n_majority7_module_83__or_module_3_res) );
  AND2_X1 u_majority7_module_83__and_module_4_U1 ( .A1(
        n_majority7_module_83__and_module_2_res), .A2(
        n_majority7_module_83__and_module_1_res), .ZN(
        n_majority7_module_83__and_module_4_res) );
  OR2_X1 u_majority7_module_83__or_module_4_U1 ( .A1(
        n_majority7_module_83__and_module_1_res), .A2(
        n_majority7_module_83__and_module_2_res), .ZN(
        n_majority7_module_83__or_module_4_res) );
  AND2_X1 u_majority7_module_83__and_module_5_U1 ( .A1(
        n_majority7_module_83__and_module_3_res), .A2(n_majority7_module_83_n2), .ZN(n_majority7_module_83__and_module_5_res) );
  OR2_X1 u_majority7_module_83__or_module_5_U1 ( .A1(n_majority7_module_83_n2), 
        .A2(n_majority7_module_83__and_module_3_res), .ZN(
        n_majority7_module_83__or_module_5_res) );
  AND2_X1 u_majority7_module_83__and_module_6_U1 ( .A1(
        n_majority7_module_83__or_module_1_res), .A2(
        n_majority7_module_83__or_module_2_res), .ZN(
        n_majority7_module_83__and_module_6_res) );
  OR2_X1 u_majority7_module_83__or_module_6_U1 ( .A1(
        n_majority7_module_83__or_module_2_res), .A2(
        n_majority7_module_83__or_module_1_res), .ZN(
        n_majority7_module_83__or_module_6_res) );
  OR2_X1 u_majority7_module_83__or_module_7_U1 ( .A1(
        n_majority7_module_83__and_module_4_res), .A2(
        n_majority7_module_83__and_module_5_res), .ZN(
        n_majority7_module_83__or_module_7_res) );
  AND2_X1 u_majority7_module_83__and_module_7_U1 ( .A1(
        n_majority7_module_83__or_module_3_res), .A2(
        n_majority7_module_83__or_module_4_res), .ZN(
        n_majority7_module_83__and_module_7_res) );
  OR2_X1 u_majority7_module_83__or_module_8_U1 ( .A1(
        n_majority7_module_83__or_module_4_res), .A2(
        n_majority7_module_83__or_module_3_res), .ZN(
        n_majority7_module_83__or_module_8_res) );
  AND2_X1 u_majority7_module_83__and_module_8_U1 ( .A1(
        n_majority7_module_83__or_module_5_res), .A2(
        n_majority7_module_83__and_module_6_res), .ZN(
        n_majority7_module_83__and_module_8_res) );
  OR2_X1 u_majority7_module_83__or_module_9_U1 ( .A1(
        n_majority7_module_83__and_module_6_res), .A2(
        n_majority7_module_83__or_module_5_res), .ZN(
        n_majority7_module_83__or_module_9_res) );
  OR2_X1 u_majority7_module_83__or_module_10_U1 ( .A1(
        n_majority7_module_83__or_module_7_res), .A2(
        n_majority7_module_83__and_module_7_res), .ZN(
        n_majority7_module_83__or_module_10_res) );
  AND2_X1 u_majority7_module_83__and_module_9_U1 ( .A1(
        n_majority7_module_83__or_module_6_res), .A2(
        n_majority7_module_83__or_module_9_res), .ZN(
        n_majority7_module_83__and_module_9_res) );
  OR2_X1 u_majority7_module_83__or_module_11_U1 ( .A1(
        n_majority7_module_83__or_module_10_res), .A2(
        n_majority7_module_83__and_module_8_res), .ZN(
        n_majority7_module_83__or_module_11_res) );
  AND2_X1 u_majority7_module_83__and_module_10_U1 ( .A1(
        n_majority7_module_83__or_module_8_res), .A2(
        n_majority7_module_83__and_module_9_res), .ZN(
        n_majority7_module_83__and_module_10_res) );
  AND2_X1 u_majority7_module_83__and_module_11_U1 ( .A1(
        n_majority7_module_83__and_module_10_res), .A2(
        n_majority7_module_83__or_module_11_res), .ZN(
        n_majority7_module_83_res) );
  DFF_X1 u_reg_module_84__cini_mul_v000_reg ( .D(n_majority7_module_83_res), 
        .CK(clock_5), .Q(n_reg_module_84_res), .QN() );
  BUF_X1 u_majority7_module_84_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_84_n7) );
  BUF_X1 u_majority7_module_84_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_84_n6) );
  BUF_X1 u_majority7_module_84_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_84_n5) );
  BUF_X1 u_majority7_module_84_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_84_n4) );
  BUF_X1 u_majority7_module_84_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_84_n3) );
  BUF_X1 u_majority7_module_84_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_84_n2) );
  BUF_X1 u_majority7_module_84_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_84_n1) );
  AND2_X1 u_majority7_module_84__and_module_1_U1 ( .A1(
        n_majority7_module_84_n7), .A2(n_majority7_module_84_n1), .ZN(
        n_majority7_module_84__and_module_1_res) );
  OR2_X1 u_majority7_module_84__or_module_1_U1 ( .A1(n_majority7_module_84_n1), 
        .A2(n_majority7_module_84_n7), .ZN(
        n_majority7_module_84__or_module_1_res) );
  AND2_X1 u_majority7_module_84__and_module_2_U1 ( .A1(
        n_majority7_module_84_n5), .A2(n_majority7_module_84_n3), .ZN(
        n_majority7_module_84__and_module_2_res) );
  OR2_X1 u_majority7_module_84__or_module_2_U1 ( .A1(n_majority7_module_84_n3), 
        .A2(n_majority7_module_84_n5), .ZN(
        n_majority7_module_84__or_module_2_res) );
  AND2_X1 u_majority7_module_84__and_module_3_U1 ( .A1(
        n_majority7_module_84_n6), .A2(n_majority7_module_84_n4), .ZN(
        n_majority7_module_84__and_module_3_res) );
  OR2_X1 u_majority7_module_84__or_module_3_U1 ( .A1(n_majority7_module_84_n4), 
        .A2(n_majority7_module_84_n6), .ZN(
        n_majority7_module_84__or_module_3_res) );
  AND2_X1 u_majority7_module_84__and_module_4_U1 ( .A1(
        n_majority7_module_84__and_module_2_res), .A2(
        n_majority7_module_84__and_module_1_res), .ZN(
        n_majority7_module_84__and_module_4_res) );
  OR2_X1 u_majority7_module_84__or_module_4_U1 ( .A1(
        n_majority7_module_84__and_module_1_res), .A2(
        n_majority7_module_84__and_module_2_res), .ZN(
        n_majority7_module_84__or_module_4_res) );
  AND2_X1 u_majority7_module_84__and_module_5_U1 ( .A1(
        n_majority7_module_84__and_module_3_res), .A2(n_majority7_module_84_n2), .ZN(n_majority7_module_84__and_module_5_res) );
  OR2_X1 u_majority7_module_84__or_module_5_U1 ( .A1(n_majority7_module_84_n2), 
        .A2(n_majority7_module_84__and_module_3_res), .ZN(
        n_majority7_module_84__or_module_5_res) );
  AND2_X1 u_majority7_module_84__and_module_6_U1 ( .A1(
        n_majority7_module_84__or_module_1_res), .A2(
        n_majority7_module_84__or_module_2_res), .ZN(
        n_majority7_module_84__and_module_6_res) );
  OR2_X1 u_majority7_module_84__or_module_6_U1 ( .A1(
        n_majority7_module_84__or_module_2_res), .A2(
        n_majority7_module_84__or_module_1_res), .ZN(
        n_majority7_module_84__or_module_6_res) );
  OR2_X1 u_majority7_module_84__or_module_7_U1 ( .A1(
        n_majority7_module_84__and_module_4_res), .A2(
        n_majority7_module_84__and_module_5_res), .ZN(
        n_majority7_module_84__or_module_7_res) );
  AND2_X1 u_majority7_module_84__and_module_7_U1 ( .A1(
        n_majority7_module_84__or_module_3_res), .A2(
        n_majority7_module_84__or_module_4_res), .ZN(
        n_majority7_module_84__and_module_7_res) );
  OR2_X1 u_majority7_module_84__or_module_8_U1 ( .A1(
        n_majority7_module_84__or_module_4_res), .A2(
        n_majority7_module_84__or_module_3_res), .ZN(
        n_majority7_module_84__or_module_8_res) );
  AND2_X1 u_majority7_module_84__and_module_8_U1 ( .A1(
        n_majority7_module_84__or_module_5_res), .A2(
        n_majority7_module_84__and_module_6_res), .ZN(
        n_majority7_module_84__and_module_8_res) );
  OR2_X1 u_majority7_module_84__or_module_9_U1 ( .A1(
        n_majority7_module_84__and_module_6_res), .A2(
        n_majority7_module_84__or_module_5_res), .ZN(
        n_majority7_module_84__or_module_9_res) );
  OR2_X1 u_majority7_module_84__or_module_10_U1 ( .A1(
        n_majority7_module_84__or_module_7_res), .A2(
        n_majority7_module_84__and_module_7_res), .ZN(
        n_majority7_module_84__or_module_10_res) );
  AND2_X1 u_majority7_module_84__and_module_9_U1 ( .A1(
        n_majority7_module_84__or_module_6_res), .A2(
        n_majority7_module_84__or_module_9_res), .ZN(
        n_majority7_module_84__and_module_9_res) );
  OR2_X1 u_majority7_module_84__or_module_11_U1 ( .A1(
        n_majority7_module_84__or_module_10_res), .A2(
        n_majority7_module_84__and_module_8_res), .ZN(
        n_majority7_module_84__or_module_11_res) );
  AND2_X1 u_majority7_module_84__and_module_10_U1 ( .A1(
        n_majority7_module_84__or_module_8_res), .A2(
        n_majority7_module_84__and_module_9_res), .ZN(
        n_majority7_module_84__and_module_10_res) );
  AND2_X1 u_majority7_module_84__and_module_11_U1 ( .A1(
        n_majority7_module_84__and_module_10_res), .A2(
        n_majority7_module_84__or_module_11_res), .ZN(
        n_majority7_module_84_res) );
  DFF_X1 u_reg_module_85__cini_mul_v000_reg ( .D(n_majority7_module_84_res), 
        .CK(clock_5), .Q(n_reg_module_85_res), .QN() );
  BUF_X1 u_majority7_module_85_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_85_n7) );
  BUF_X1 u_majority7_module_85_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_85_n6) );
  BUF_X1 u_majority7_module_85_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_85_n5) );
  BUF_X1 u_majority7_module_85_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_85_n4) );
  BUF_X1 u_majority7_module_85_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_85_n3) );
  BUF_X1 u_majority7_module_85_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_85_n2) );
  BUF_X1 u_majority7_module_85_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_85_n1) );
  AND2_X1 u_majority7_module_85__and_module_1_U1 ( .A1(
        n_majority7_module_85_n7), .A2(n_majority7_module_85_n1), .ZN(
        n_majority7_module_85__and_module_1_res) );
  OR2_X1 u_majority7_module_85__or_module_1_U1 ( .A1(n_majority7_module_85_n1), 
        .A2(n_majority7_module_85_n7), .ZN(
        n_majority7_module_85__or_module_1_res) );
  AND2_X1 u_majority7_module_85__and_module_2_U1 ( .A1(
        n_majority7_module_85_n5), .A2(n_majority7_module_85_n3), .ZN(
        n_majority7_module_85__and_module_2_res) );
  OR2_X1 u_majority7_module_85__or_module_2_U1 ( .A1(n_majority7_module_85_n3), 
        .A2(n_majority7_module_85_n5), .ZN(
        n_majority7_module_85__or_module_2_res) );
  AND2_X1 u_majority7_module_85__and_module_3_U1 ( .A1(
        n_majority7_module_85_n6), .A2(n_majority7_module_85_n4), .ZN(
        n_majority7_module_85__and_module_3_res) );
  OR2_X1 u_majority7_module_85__or_module_3_U1 ( .A1(n_majority7_module_85_n4), 
        .A2(n_majority7_module_85_n6), .ZN(
        n_majority7_module_85__or_module_3_res) );
  AND2_X1 u_majority7_module_85__and_module_4_U1 ( .A1(
        n_majority7_module_85__and_module_2_res), .A2(
        n_majority7_module_85__and_module_1_res), .ZN(
        n_majority7_module_85__and_module_4_res) );
  OR2_X1 u_majority7_module_85__or_module_4_U1 ( .A1(
        n_majority7_module_85__and_module_1_res), .A2(
        n_majority7_module_85__and_module_2_res), .ZN(
        n_majority7_module_85__or_module_4_res) );
  AND2_X1 u_majority7_module_85__and_module_5_U1 ( .A1(
        n_majority7_module_85__and_module_3_res), .A2(n_majority7_module_85_n2), .ZN(n_majority7_module_85__and_module_5_res) );
  OR2_X1 u_majority7_module_85__or_module_5_U1 ( .A1(n_majority7_module_85_n2), 
        .A2(n_majority7_module_85__and_module_3_res), .ZN(
        n_majority7_module_85__or_module_5_res) );
  AND2_X1 u_majority7_module_85__and_module_6_U1 ( .A1(
        n_majority7_module_85__or_module_1_res), .A2(
        n_majority7_module_85__or_module_2_res), .ZN(
        n_majority7_module_85__and_module_6_res) );
  OR2_X1 u_majority7_module_85__or_module_6_U1 ( .A1(
        n_majority7_module_85__or_module_2_res), .A2(
        n_majority7_module_85__or_module_1_res), .ZN(
        n_majority7_module_85__or_module_6_res) );
  OR2_X1 u_majority7_module_85__or_module_7_U1 ( .A1(
        n_majority7_module_85__and_module_4_res), .A2(
        n_majority7_module_85__and_module_5_res), .ZN(
        n_majority7_module_85__or_module_7_res) );
  AND2_X1 u_majority7_module_85__and_module_7_U1 ( .A1(
        n_majority7_module_85__or_module_3_res), .A2(
        n_majority7_module_85__or_module_4_res), .ZN(
        n_majority7_module_85__and_module_7_res) );
  OR2_X1 u_majority7_module_85__or_module_8_U1 ( .A1(
        n_majority7_module_85__or_module_4_res), .A2(
        n_majority7_module_85__or_module_3_res), .ZN(
        n_majority7_module_85__or_module_8_res) );
  AND2_X1 u_majority7_module_85__and_module_8_U1 ( .A1(
        n_majority7_module_85__or_module_5_res), .A2(
        n_majority7_module_85__and_module_6_res), .ZN(
        n_majority7_module_85__and_module_8_res) );
  OR2_X1 u_majority7_module_85__or_module_9_U1 ( .A1(
        n_majority7_module_85__and_module_6_res), .A2(
        n_majority7_module_85__or_module_5_res), .ZN(
        n_majority7_module_85__or_module_9_res) );
  OR2_X1 u_majority7_module_85__or_module_10_U1 ( .A1(
        n_majority7_module_85__or_module_7_res), .A2(
        n_majority7_module_85__and_module_7_res), .ZN(
        n_majority7_module_85__or_module_10_res) );
  AND2_X1 u_majority7_module_85__and_module_9_U1 ( .A1(
        n_majority7_module_85__or_module_6_res), .A2(
        n_majority7_module_85__or_module_9_res), .ZN(
        n_majority7_module_85__and_module_9_res) );
  OR2_X1 u_majority7_module_85__or_module_11_U1 ( .A1(
        n_majority7_module_85__or_module_10_res), .A2(
        n_majority7_module_85__and_module_8_res), .ZN(
        n_majority7_module_85__or_module_11_res) );
  AND2_X1 u_majority7_module_85__and_module_10_U1 ( .A1(
        n_majority7_module_85__or_module_8_res), .A2(
        n_majority7_module_85__and_module_9_res), .ZN(
        n_majority7_module_85__and_module_10_res) );
  AND2_X1 u_majority7_module_85__and_module_11_U1 ( .A1(
        n_majority7_module_85__and_module_10_res), .A2(
        n_majority7_module_85__or_module_11_res), .ZN(
        n_majority7_module_85_res) );
  DFF_X1 u_reg_module_86__cini_mul_v000_reg ( .D(n_majority7_module_85_res), 
        .CK(clock_5), .Q(n_reg_module_86_res), .QN() );
  BUF_X1 u_majority7_module_86_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_86_n7) );
  BUF_X1 u_majority7_module_86_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_86_n6) );
  BUF_X1 u_majority7_module_86_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_86_n5) );
  BUF_X1 u_majority7_module_86_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_86_n4) );
  BUF_X1 u_majority7_module_86_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_86_n3) );
  BUF_X1 u_majority7_module_86_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_86_n2) );
  BUF_X1 u_majority7_module_86_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_86_n1) );
  AND2_X1 u_majority7_module_86__and_module_1_U1 ( .A1(
        n_majority7_module_86_n7), .A2(n_majority7_module_86_n1), .ZN(
        n_majority7_module_86__and_module_1_res) );
  OR2_X1 u_majority7_module_86__or_module_1_U1 ( .A1(n_majority7_module_86_n1), 
        .A2(n_majority7_module_86_n7), .ZN(
        n_majority7_module_86__or_module_1_res) );
  AND2_X1 u_majority7_module_86__and_module_2_U1 ( .A1(
        n_majority7_module_86_n5), .A2(n_majority7_module_86_n3), .ZN(
        n_majority7_module_86__and_module_2_res) );
  OR2_X1 u_majority7_module_86__or_module_2_U1 ( .A1(n_majority7_module_86_n3), 
        .A2(n_majority7_module_86_n5), .ZN(
        n_majority7_module_86__or_module_2_res) );
  AND2_X1 u_majority7_module_86__and_module_3_U1 ( .A1(
        n_majority7_module_86_n6), .A2(n_majority7_module_86_n4), .ZN(
        n_majority7_module_86__and_module_3_res) );
  OR2_X1 u_majority7_module_86__or_module_3_U1 ( .A1(n_majority7_module_86_n4), 
        .A2(n_majority7_module_86_n6), .ZN(
        n_majority7_module_86__or_module_3_res) );
  AND2_X1 u_majority7_module_86__and_module_4_U1 ( .A1(
        n_majority7_module_86__and_module_2_res), .A2(
        n_majority7_module_86__and_module_1_res), .ZN(
        n_majority7_module_86__and_module_4_res) );
  OR2_X1 u_majority7_module_86__or_module_4_U1 ( .A1(
        n_majority7_module_86__and_module_1_res), .A2(
        n_majority7_module_86__and_module_2_res), .ZN(
        n_majority7_module_86__or_module_4_res) );
  AND2_X1 u_majority7_module_86__and_module_5_U1 ( .A1(
        n_majority7_module_86__and_module_3_res), .A2(n_majority7_module_86_n2), .ZN(n_majority7_module_86__and_module_5_res) );
  OR2_X1 u_majority7_module_86__or_module_5_U1 ( .A1(n_majority7_module_86_n2), 
        .A2(n_majority7_module_86__and_module_3_res), .ZN(
        n_majority7_module_86__or_module_5_res) );
  AND2_X1 u_majority7_module_86__and_module_6_U1 ( .A1(
        n_majority7_module_86__or_module_1_res), .A2(
        n_majority7_module_86__or_module_2_res), .ZN(
        n_majority7_module_86__and_module_6_res) );
  OR2_X1 u_majority7_module_86__or_module_6_U1 ( .A1(
        n_majority7_module_86__or_module_2_res), .A2(
        n_majority7_module_86__or_module_1_res), .ZN(
        n_majority7_module_86__or_module_6_res) );
  OR2_X1 u_majority7_module_86__or_module_7_U1 ( .A1(
        n_majority7_module_86__and_module_4_res), .A2(
        n_majority7_module_86__and_module_5_res), .ZN(
        n_majority7_module_86__or_module_7_res) );
  AND2_X1 u_majority7_module_86__and_module_7_U1 ( .A1(
        n_majority7_module_86__or_module_3_res), .A2(
        n_majority7_module_86__or_module_4_res), .ZN(
        n_majority7_module_86__and_module_7_res) );
  OR2_X1 u_majority7_module_86__or_module_8_U1 ( .A1(
        n_majority7_module_86__or_module_4_res), .A2(
        n_majority7_module_86__or_module_3_res), .ZN(
        n_majority7_module_86__or_module_8_res) );
  AND2_X1 u_majority7_module_86__and_module_8_U1 ( .A1(
        n_majority7_module_86__or_module_5_res), .A2(
        n_majority7_module_86__and_module_6_res), .ZN(
        n_majority7_module_86__and_module_8_res) );
  OR2_X1 u_majority7_module_86__or_module_9_U1 ( .A1(
        n_majority7_module_86__and_module_6_res), .A2(
        n_majority7_module_86__or_module_5_res), .ZN(
        n_majority7_module_86__or_module_9_res) );
  OR2_X1 u_majority7_module_86__or_module_10_U1 ( .A1(
        n_majority7_module_86__or_module_7_res), .A2(
        n_majority7_module_86__and_module_7_res), .ZN(
        n_majority7_module_86__or_module_10_res) );
  AND2_X1 u_majority7_module_86__and_module_9_U1 ( .A1(
        n_majority7_module_86__or_module_6_res), .A2(
        n_majority7_module_86__or_module_9_res), .ZN(
        n_majority7_module_86__and_module_9_res) );
  OR2_X1 u_majority7_module_86__or_module_11_U1 ( .A1(
        n_majority7_module_86__or_module_10_res), .A2(
        n_majority7_module_86__and_module_8_res), .ZN(
        n_majority7_module_86__or_module_11_res) );
  AND2_X1 u_majority7_module_86__and_module_10_U1 ( .A1(
        n_majority7_module_86__or_module_8_res), .A2(
        n_majority7_module_86__and_module_9_res), .ZN(
        n_majority7_module_86__and_module_10_res) );
  AND2_X1 u_majority7_module_86__and_module_11_U1 ( .A1(
        n_majority7_module_86__and_module_10_res), .A2(
        n_majority7_module_86__or_module_11_res), .ZN(
        n_majority7_module_86_res) );
  DFF_X1 u_reg_module_87__cini_mul_v000_reg ( .D(n_majority7_module_86_res), 
        .CK(clock_5), .Q(n_reg_module_87_res), .QN() );
  BUF_X1 u_majority7_module_87_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_87_n7) );
  BUF_X1 u_majority7_module_87_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_87_n6) );
  BUF_X1 u_majority7_module_87_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_87_n5) );
  BUF_X1 u_majority7_module_87_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_87_n4) );
  BUF_X1 u_majority7_module_87_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_87_n3) );
  BUF_X1 u_majority7_module_87_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_87_n2) );
  BUF_X1 u_majority7_module_87_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_87_n1) );
  AND2_X1 u_majority7_module_87__and_module_1_U1 ( .A1(
        n_majority7_module_87_n7), .A2(n_majority7_module_87_n1), .ZN(
        n_majority7_module_87__and_module_1_res) );
  OR2_X1 u_majority7_module_87__or_module_1_U1 ( .A1(n_majority7_module_87_n1), 
        .A2(n_majority7_module_87_n7), .ZN(
        n_majority7_module_87__or_module_1_res) );
  AND2_X1 u_majority7_module_87__and_module_2_U1 ( .A1(
        n_majority7_module_87_n5), .A2(n_majority7_module_87_n3), .ZN(
        n_majority7_module_87__and_module_2_res) );
  OR2_X1 u_majority7_module_87__or_module_2_U1 ( .A1(n_majority7_module_87_n3), 
        .A2(n_majority7_module_87_n5), .ZN(
        n_majority7_module_87__or_module_2_res) );
  AND2_X1 u_majority7_module_87__and_module_3_U1 ( .A1(
        n_majority7_module_87_n6), .A2(n_majority7_module_87_n4), .ZN(
        n_majority7_module_87__and_module_3_res) );
  OR2_X1 u_majority7_module_87__or_module_3_U1 ( .A1(n_majority7_module_87_n4), 
        .A2(n_majority7_module_87_n6), .ZN(
        n_majority7_module_87__or_module_3_res) );
  AND2_X1 u_majority7_module_87__and_module_4_U1 ( .A1(
        n_majority7_module_87__and_module_2_res), .A2(
        n_majority7_module_87__and_module_1_res), .ZN(
        n_majority7_module_87__and_module_4_res) );
  OR2_X1 u_majority7_module_87__or_module_4_U1 ( .A1(
        n_majority7_module_87__and_module_1_res), .A2(
        n_majority7_module_87__and_module_2_res), .ZN(
        n_majority7_module_87__or_module_4_res) );
  AND2_X1 u_majority7_module_87__and_module_5_U1 ( .A1(
        n_majority7_module_87__and_module_3_res), .A2(n_majority7_module_87_n2), .ZN(n_majority7_module_87__and_module_5_res) );
  OR2_X1 u_majority7_module_87__or_module_5_U1 ( .A1(n_majority7_module_87_n2), 
        .A2(n_majority7_module_87__and_module_3_res), .ZN(
        n_majority7_module_87__or_module_5_res) );
  AND2_X1 u_majority7_module_87__and_module_6_U1 ( .A1(
        n_majority7_module_87__or_module_1_res), .A2(
        n_majority7_module_87__or_module_2_res), .ZN(
        n_majority7_module_87__and_module_6_res) );
  OR2_X1 u_majority7_module_87__or_module_6_U1 ( .A1(
        n_majority7_module_87__or_module_2_res), .A2(
        n_majority7_module_87__or_module_1_res), .ZN(
        n_majority7_module_87__or_module_6_res) );
  OR2_X1 u_majority7_module_87__or_module_7_U1 ( .A1(
        n_majority7_module_87__and_module_4_res), .A2(
        n_majority7_module_87__and_module_5_res), .ZN(
        n_majority7_module_87__or_module_7_res) );
  AND2_X1 u_majority7_module_87__and_module_7_U1 ( .A1(
        n_majority7_module_87__or_module_3_res), .A2(
        n_majority7_module_87__or_module_4_res), .ZN(
        n_majority7_module_87__and_module_7_res) );
  OR2_X1 u_majority7_module_87__or_module_8_U1 ( .A1(
        n_majority7_module_87__or_module_4_res), .A2(
        n_majority7_module_87__or_module_3_res), .ZN(
        n_majority7_module_87__or_module_8_res) );
  AND2_X1 u_majority7_module_87__and_module_8_U1 ( .A1(
        n_majority7_module_87__or_module_5_res), .A2(
        n_majority7_module_87__and_module_6_res), .ZN(
        n_majority7_module_87__and_module_8_res) );
  OR2_X1 u_majority7_module_87__or_module_9_U1 ( .A1(
        n_majority7_module_87__and_module_6_res), .A2(
        n_majority7_module_87__or_module_5_res), .ZN(
        n_majority7_module_87__or_module_9_res) );
  OR2_X1 u_majority7_module_87__or_module_10_U1 ( .A1(
        n_majority7_module_87__or_module_7_res), .A2(
        n_majority7_module_87__and_module_7_res), .ZN(
        n_majority7_module_87__or_module_10_res) );
  AND2_X1 u_majority7_module_87__and_module_9_U1 ( .A1(
        n_majority7_module_87__or_module_6_res), .A2(
        n_majority7_module_87__or_module_9_res), .ZN(
        n_majority7_module_87__and_module_9_res) );
  OR2_X1 u_majority7_module_87__or_module_11_U1 ( .A1(
        n_majority7_module_87__or_module_10_res), .A2(
        n_majority7_module_87__and_module_8_res), .ZN(
        n_majority7_module_87__or_module_11_res) );
  AND2_X1 u_majority7_module_87__and_module_10_U1 ( .A1(
        n_majority7_module_87__or_module_8_res), .A2(
        n_majority7_module_87__and_module_9_res), .ZN(
        n_majority7_module_87__and_module_10_res) );
  AND2_X1 u_majority7_module_87__and_module_11_U1 ( .A1(
        n_majority7_module_87__and_module_10_res), .A2(
        n_majority7_module_87__or_module_11_res), .ZN(
        n_majority7_module_87_res) );
  DFF_X1 u_reg_module_88__cini_mul_v000_reg ( .D(n_majority7_module_87_res), 
        .CK(clock_5), .Q(n_reg_module_88_res), .QN() );
  BUF_X1 u_majority7_module_88_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_88_n7) );
  BUF_X1 u_majority7_module_88_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_88_n6) );
  BUF_X1 u_majority7_module_88_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_88_n5) );
  BUF_X1 u_majority7_module_88_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_88_n4) );
  BUF_X1 u_majority7_module_88_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_88_n3) );
  BUF_X1 u_majority7_module_88_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_88_n2) );
  BUF_X1 u_majority7_module_88_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_88_n1) );
  AND2_X1 u_majority7_module_88__and_module_1_U1 ( .A1(
        n_majority7_module_88_n7), .A2(n_majority7_module_88_n1), .ZN(
        n_majority7_module_88__and_module_1_res) );
  OR2_X1 u_majority7_module_88__or_module_1_U1 ( .A1(n_majority7_module_88_n1), 
        .A2(n_majority7_module_88_n7), .ZN(
        n_majority7_module_88__or_module_1_res) );
  AND2_X1 u_majority7_module_88__and_module_2_U1 ( .A1(
        n_majority7_module_88_n5), .A2(n_majority7_module_88_n3), .ZN(
        n_majority7_module_88__and_module_2_res) );
  OR2_X1 u_majority7_module_88__or_module_2_U1 ( .A1(n_majority7_module_88_n3), 
        .A2(n_majority7_module_88_n5), .ZN(
        n_majority7_module_88__or_module_2_res) );
  AND2_X1 u_majority7_module_88__and_module_3_U1 ( .A1(
        n_majority7_module_88_n6), .A2(n_majority7_module_88_n4), .ZN(
        n_majority7_module_88__and_module_3_res) );
  OR2_X1 u_majority7_module_88__or_module_3_U1 ( .A1(n_majority7_module_88_n4), 
        .A2(n_majority7_module_88_n6), .ZN(
        n_majority7_module_88__or_module_3_res) );
  AND2_X1 u_majority7_module_88__and_module_4_U1 ( .A1(
        n_majority7_module_88__and_module_2_res), .A2(
        n_majority7_module_88__and_module_1_res), .ZN(
        n_majority7_module_88__and_module_4_res) );
  OR2_X1 u_majority7_module_88__or_module_4_U1 ( .A1(
        n_majority7_module_88__and_module_1_res), .A2(
        n_majority7_module_88__and_module_2_res), .ZN(
        n_majority7_module_88__or_module_4_res) );
  AND2_X1 u_majority7_module_88__and_module_5_U1 ( .A1(
        n_majority7_module_88__and_module_3_res), .A2(n_majority7_module_88_n2), .ZN(n_majority7_module_88__and_module_5_res) );
  OR2_X1 u_majority7_module_88__or_module_5_U1 ( .A1(n_majority7_module_88_n2), 
        .A2(n_majority7_module_88__and_module_3_res), .ZN(
        n_majority7_module_88__or_module_5_res) );
  AND2_X1 u_majority7_module_88__and_module_6_U1 ( .A1(
        n_majority7_module_88__or_module_1_res), .A2(
        n_majority7_module_88__or_module_2_res), .ZN(
        n_majority7_module_88__and_module_6_res) );
  OR2_X1 u_majority7_module_88__or_module_6_U1 ( .A1(
        n_majority7_module_88__or_module_2_res), .A2(
        n_majority7_module_88__or_module_1_res), .ZN(
        n_majority7_module_88__or_module_6_res) );
  OR2_X1 u_majority7_module_88__or_module_7_U1 ( .A1(
        n_majority7_module_88__and_module_4_res), .A2(
        n_majority7_module_88__and_module_5_res), .ZN(
        n_majority7_module_88__or_module_7_res) );
  AND2_X1 u_majority7_module_88__and_module_7_U1 ( .A1(
        n_majority7_module_88__or_module_3_res), .A2(
        n_majority7_module_88__or_module_4_res), .ZN(
        n_majority7_module_88__and_module_7_res) );
  OR2_X1 u_majority7_module_88__or_module_8_U1 ( .A1(
        n_majority7_module_88__or_module_4_res), .A2(
        n_majority7_module_88__or_module_3_res), .ZN(
        n_majority7_module_88__or_module_8_res) );
  AND2_X1 u_majority7_module_88__and_module_8_U1 ( .A1(
        n_majority7_module_88__or_module_5_res), .A2(
        n_majority7_module_88__and_module_6_res), .ZN(
        n_majority7_module_88__and_module_8_res) );
  OR2_X1 u_majority7_module_88__or_module_9_U1 ( .A1(
        n_majority7_module_88__and_module_6_res), .A2(
        n_majority7_module_88__or_module_5_res), .ZN(
        n_majority7_module_88__or_module_9_res) );
  OR2_X1 u_majority7_module_88__or_module_10_U1 ( .A1(
        n_majority7_module_88__or_module_7_res), .A2(
        n_majority7_module_88__and_module_7_res), .ZN(
        n_majority7_module_88__or_module_10_res) );
  AND2_X1 u_majority7_module_88__and_module_9_U1 ( .A1(
        n_majority7_module_88__or_module_6_res), .A2(
        n_majority7_module_88__or_module_9_res), .ZN(
        n_majority7_module_88__and_module_9_res) );
  OR2_X1 u_majority7_module_88__or_module_11_U1 ( .A1(
        n_majority7_module_88__or_module_10_res), .A2(
        n_majority7_module_88__and_module_8_res), .ZN(
        n_majority7_module_88__or_module_11_res) );
  AND2_X1 u_majority7_module_88__and_module_10_U1 ( .A1(
        n_majority7_module_88__or_module_8_res), .A2(
        n_majority7_module_88__and_module_9_res), .ZN(
        n_majority7_module_88__and_module_10_res) );
  AND2_X1 u_majority7_module_88__and_module_11_U1 ( .A1(
        n_majority7_module_88__and_module_10_res), .A2(
        n_majority7_module_88__or_module_11_res), .ZN(
        n_majority7_module_88_res) );
  DFF_X1 u_reg_module_89__cini_mul_v000_reg ( .D(n_majority7_module_88_res), 
        .CK(clock_5), .Q(n_reg_module_89_res), .QN() );
  BUF_X1 u_majority7_module_89_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_89_n7) );
  BUF_X1 u_majority7_module_89_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_89_n6) );
  BUF_X1 u_majority7_module_89_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_89_n5) );
  BUF_X1 u_majority7_module_89_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_89_n4) );
  BUF_X1 u_majority7_module_89_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_89_n3) );
  BUF_X1 u_majority7_module_89_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_89_n2) );
  BUF_X1 u_majority7_module_89_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_89_n1) );
  AND2_X1 u_majority7_module_89__and_module_1_U1 ( .A1(
        n_majority7_module_89_n7), .A2(n_majority7_module_89_n1), .ZN(
        n_majority7_module_89__and_module_1_res) );
  OR2_X1 u_majority7_module_89__or_module_1_U1 ( .A1(n_majority7_module_89_n1), 
        .A2(n_majority7_module_89_n7), .ZN(
        n_majority7_module_89__or_module_1_res) );
  AND2_X1 u_majority7_module_89__and_module_2_U1 ( .A1(
        n_majority7_module_89_n5), .A2(n_majority7_module_89_n3), .ZN(
        n_majority7_module_89__and_module_2_res) );
  OR2_X1 u_majority7_module_89__or_module_2_U1 ( .A1(n_majority7_module_89_n3), 
        .A2(n_majority7_module_89_n5), .ZN(
        n_majority7_module_89__or_module_2_res) );
  AND2_X1 u_majority7_module_89__and_module_3_U1 ( .A1(
        n_majority7_module_89_n6), .A2(n_majority7_module_89_n4), .ZN(
        n_majority7_module_89__and_module_3_res) );
  OR2_X1 u_majority7_module_89__or_module_3_U1 ( .A1(n_majority7_module_89_n4), 
        .A2(n_majority7_module_89_n6), .ZN(
        n_majority7_module_89__or_module_3_res) );
  AND2_X1 u_majority7_module_89__and_module_4_U1 ( .A1(
        n_majority7_module_89__and_module_2_res), .A2(
        n_majority7_module_89__and_module_1_res), .ZN(
        n_majority7_module_89__and_module_4_res) );
  OR2_X1 u_majority7_module_89__or_module_4_U1 ( .A1(
        n_majority7_module_89__and_module_1_res), .A2(
        n_majority7_module_89__and_module_2_res), .ZN(
        n_majority7_module_89__or_module_4_res) );
  AND2_X1 u_majority7_module_89__and_module_5_U1 ( .A1(
        n_majority7_module_89__and_module_3_res), .A2(n_majority7_module_89_n2), .ZN(n_majority7_module_89__and_module_5_res) );
  OR2_X1 u_majority7_module_89__or_module_5_U1 ( .A1(n_majority7_module_89_n2), 
        .A2(n_majority7_module_89__and_module_3_res), .ZN(
        n_majority7_module_89__or_module_5_res) );
  AND2_X1 u_majority7_module_89__and_module_6_U1 ( .A1(
        n_majority7_module_89__or_module_1_res), .A2(
        n_majority7_module_89__or_module_2_res), .ZN(
        n_majority7_module_89__and_module_6_res) );
  OR2_X1 u_majority7_module_89__or_module_6_U1 ( .A1(
        n_majority7_module_89__or_module_2_res), .A2(
        n_majority7_module_89__or_module_1_res), .ZN(
        n_majority7_module_89__or_module_6_res) );
  OR2_X1 u_majority7_module_89__or_module_7_U1 ( .A1(
        n_majority7_module_89__and_module_4_res), .A2(
        n_majority7_module_89__and_module_5_res), .ZN(
        n_majority7_module_89__or_module_7_res) );
  AND2_X1 u_majority7_module_89__and_module_7_U1 ( .A1(
        n_majority7_module_89__or_module_3_res), .A2(
        n_majority7_module_89__or_module_4_res), .ZN(
        n_majority7_module_89__and_module_7_res) );
  OR2_X1 u_majority7_module_89__or_module_8_U1 ( .A1(
        n_majority7_module_89__or_module_4_res), .A2(
        n_majority7_module_89__or_module_3_res), .ZN(
        n_majority7_module_89__or_module_8_res) );
  AND2_X1 u_majority7_module_89__and_module_8_U1 ( .A1(
        n_majority7_module_89__or_module_5_res), .A2(
        n_majority7_module_89__and_module_6_res), .ZN(
        n_majority7_module_89__and_module_8_res) );
  OR2_X1 u_majority7_module_89__or_module_9_U1 ( .A1(
        n_majority7_module_89__and_module_6_res), .A2(
        n_majority7_module_89__or_module_5_res), .ZN(
        n_majority7_module_89__or_module_9_res) );
  OR2_X1 u_majority7_module_89__or_module_10_U1 ( .A1(
        n_majority7_module_89__or_module_7_res), .A2(
        n_majority7_module_89__and_module_7_res), .ZN(
        n_majority7_module_89__or_module_10_res) );
  AND2_X1 u_majority7_module_89__and_module_9_U1 ( .A1(
        n_majority7_module_89__or_module_6_res), .A2(
        n_majority7_module_89__or_module_9_res), .ZN(
        n_majority7_module_89__and_module_9_res) );
  OR2_X1 u_majority7_module_89__or_module_11_U1 ( .A1(
        n_majority7_module_89__or_module_10_res), .A2(
        n_majority7_module_89__and_module_8_res), .ZN(
        n_majority7_module_89__or_module_11_res) );
  AND2_X1 u_majority7_module_89__and_module_10_U1 ( .A1(
        n_majority7_module_89__or_module_8_res), .A2(
        n_majority7_module_89__and_module_9_res), .ZN(
        n_majority7_module_89__and_module_10_res) );
  AND2_X1 u_majority7_module_89__and_module_11_U1 ( .A1(
        n_majority7_module_89__and_module_10_res), .A2(
        n_majority7_module_89__or_module_11_res), .ZN(
        n_majority7_module_89_res) );
  DFF_X1 u_reg_module_90__cini_mul_v000_reg ( .D(n_majority7_module_89_res), 
        .CK(clock_5), .Q(n_reg_module_90_res), .QN() );
  BUF_X1 u_majority7_module_90_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_90_n7) );
  BUF_X1 u_majority7_module_90_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_90_n6) );
  BUF_X1 u_majority7_module_90_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_90_n5) );
  BUF_X1 u_majority7_module_90_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_90_n4) );
  BUF_X1 u_majority7_module_90_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_90_n3) );
  BUF_X1 u_majority7_module_90_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_90_n2) );
  BUF_X1 u_majority7_module_90_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_90_n1) );
  AND2_X1 u_majority7_module_90__and_module_1_U1 ( .A1(
        n_majority7_module_90_n7), .A2(n_majority7_module_90_n1), .ZN(
        n_majority7_module_90__and_module_1_res) );
  OR2_X1 u_majority7_module_90__or_module_1_U1 ( .A1(n_majority7_module_90_n1), 
        .A2(n_majority7_module_90_n7), .ZN(
        n_majority7_module_90__or_module_1_res) );
  AND2_X1 u_majority7_module_90__and_module_2_U1 ( .A1(
        n_majority7_module_90_n5), .A2(n_majority7_module_90_n3), .ZN(
        n_majority7_module_90__and_module_2_res) );
  OR2_X1 u_majority7_module_90__or_module_2_U1 ( .A1(n_majority7_module_90_n3), 
        .A2(n_majority7_module_90_n5), .ZN(
        n_majority7_module_90__or_module_2_res) );
  AND2_X1 u_majority7_module_90__and_module_3_U1 ( .A1(
        n_majority7_module_90_n6), .A2(n_majority7_module_90_n4), .ZN(
        n_majority7_module_90__and_module_3_res) );
  OR2_X1 u_majority7_module_90__or_module_3_U1 ( .A1(n_majority7_module_90_n4), 
        .A2(n_majority7_module_90_n6), .ZN(
        n_majority7_module_90__or_module_3_res) );
  AND2_X1 u_majority7_module_90__and_module_4_U1 ( .A1(
        n_majority7_module_90__and_module_2_res), .A2(
        n_majority7_module_90__and_module_1_res), .ZN(
        n_majority7_module_90__and_module_4_res) );
  OR2_X1 u_majority7_module_90__or_module_4_U1 ( .A1(
        n_majority7_module_90__and_module_1_res), .A2(
        n_majority7_module_90__and_module_2_res), .ZN(
        n_majority7_module_90__or_module_4_res) );
  AND2_X1 u_majority7_module_90__and_module_5_U1 ( .A1(
        n_majority7_module_90__and_module_3_res), .A2(n_majority7_module_90_n2), .ZN(n_majority7_module_90__and_module_5_res) );
  OR2_X1 u_majority7_module_90__or_module_5_U1 ( .A1(n_majority7_module_90_n2), 
        .A2(n_majority7_module_90__and_module_3_res), .ZN(
        n_majority7_module_90__or_module_5_res) );
  AND2_X1 u_majority7_module_90__and_module_6_U1 ( .A1(
        n_majority7_module_90__or_module_1_res), .A2(
        n_majority7_module_90__or_module_2_res), .ZN(
        n_majority7_module_90__and_module_6_res) );
  OR2_X1 u_majority7_module_90__or_module_6_U1 ( .A1(
        n_majority7_module_90__or_module_2_res), .A2(
        n_majority7_module_90__or_module_1_res), .ZN(
        n_majority7_module_90__or_module_6_res) );
  OR2_X1 u_majority7_module_90__or_module_7_U1 ( .A1(
        n_majority7_module_90__and_module_4_res), .A2(
        n_majority7_module_90__and_module_5_res), .ZN(
        n_majority7_module_90__or_module_7_res) );
  AND2_X1 u_majority7_module_90__and_module_7_U1 ( .A1(
        n_majority7_module_90__or_module_3_res), .A2(
        n_majority7_module_90__or_module_4_res), .ZN(
        n_majority7_module_90__and_module_7_res) );
  OR2_X1 u_majority7_module_90__or_module_8_U1 ( .A1(
        n_majority7_module_90__or_module_4_res), .A2(
        n_majority7_module_90__or_module_3_res), .ZN(
        n_majority7_module_90__or_module_8_res) );
  AND2_X1 u_majority7_module_90__and_module_8_U1 ( .A1(
        n_majority7_module_90__or_module_5_res), .A2(
        n_majority7_module_90__and_module_6_res), .ZN(
        n_majority7_module_90__and_module_8_res) );
  OR2_X1 u_majority7_module_90__or_module_9_U1 ( .A1(
        n_majority7_module_90__and_module_6_res), .A2(
        n_majority7_module_90__or_module_5_res), .ZN(
        n_majority7_module_90__or_module_9_res) );
  OR2_X1 u_majority7_module_90__or_module_10_U1 ( .A1(
        n_majority7_module_90__or_module_7_res), .A2(
        n_majority7_module_90__and_module_7_res), .ZN(
        n_majority7_module_90__or_module_10_res) );
  AND2_X1 u_majority7_module_90__and_module_9_U1 ( .A1(
        n_majority7_module_90__or_module_6_res), .A2(
        n_majority7_module_90__or_module_9_res), .ZN(
        n_majority7_module_90__and_module_9_res) );
  OR2_X1 u_majority7_module_90__or_module_11_U1 ( .A1(
        n_majority7_module_90__or_module_10_res), .A2(
        n_majority7_module_90__and_module_8_res), .ZN(
        n_majority7_module_90__or_module_11_res) );
  AND2_X1 u_majority7_module_90__and_module_10_U1 ( .A1(
        n_majority7_module_90__or_module_8_res), .A2(
        n_majority7_module_90__and_module_9_res), .ZN(
        n_majority7_module_90__and_module_10_res) );
  AND2_X1 u_majority7_module_90__and_module_11_U1 ( .A1(
        n_majority7_module_90__and_module_10_res), .A2(
        n_majority7_module_90__or_module_11_res), .ZN(
        n_majority7_module_90_res) );
  DFF_X1 u_reg_module_91__cini_mul_v000_reg ( .D(n_majority7_module_90_res), 
        .CK(clock_5), .Q(n_reg_module_91_res), .QN() );
  BUF_X1 u_majority7_module_91_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_91_n7) );
  BUF_X1 u_majority7_module_91_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_91_n6) );
  BUF_X1 u_majority7_module_91_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_91_n5) );
  BUF_X1 u_majority7_module_91_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_91_n4) );
  BUF_X1 u_majority7_module_91_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_91_n3) );
  BUF_X1 u_majority7_module_91_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_91_n2) );
  BUF_X1 u_majority7_module_91_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_91_n1) );
  AND2_X1 u_majority7_module_91__and_module_1_U1 ( .A1(
        n_majority7_module_91_n7), .A2(n_majority7_module_91_n1), .ZN(
        n_majority7_module_91__and_module_1_res) );
  OR2_X1 u_majority7_module_91__or_module_1_U1 ( .A1(n_majority7_module_91_n1), 
        .A2(n_majority7_module_91_n7), .ZN(
        n_majority7_module_91__or_module_1_res) );
  AND2_X1 u_majority7_module_91__and_module_2_U1 ( .A1(
        n_majority7_module_91_n5), .A2(n_majority7_module_91_n3), .ZN(
        n_majority7_module_91__and_module_2_res) );
  OR2_X1 u_majority7_module_91__or_module_2_U1 ( .A1(n_majority7_module_91_n3), 
        .A2(n_majority7_module_91_n5), .ZN(
        n_majority7_module_91__or_module_2_res) );
  AND2_X1 u_majority7_module_91__and_module_3_U1 ( .A1(
        n_majority7_module_91_n6), .A2(n_majority7_module_91_n4), .ZN(
        n_majority7_module_91__and_module_3_res) );
  OR2_X1 u_majority7_module_91__or_module_3_U1 ( .A1(n_majority7_module_91_n4), 
        .A2(n_majority7_module_91_n6), .ZN(
        n_majority7_module_91__or_module_3_res) );
  AND2_X1 u_majority7_module_91__and_module_4_U1 ( .A1(
        n_majority7_module_91__and_module_2_res), .A2(
        n_majority7_module_91__and_module_1_res), .ZN(
        n_majority7_module_91__and_module_4_res) );
  OR2_X1 u_majority7_module_91__or_module_4_U1 ( .A1(
        n_majority7_module_91__and_module_1_res), .A2(
        n_majority7_module_91__and_module_2_res), .ZN(
        n_majority7_module_91__or_module_4_res) );
  AND2_X1 u_majority7_module_91__and_module_5_U1 ( .A1(
        n_majority7_module_91__and_module_3_res), .A2(n_majority7_module_91_n2), .ZN(n_majority7_module_91__and_module_5_res) );
  OR2_X1 u_majority7_module_91__or_module_5_U1 ( .A1(n_majority7_module_91_n2), 
        .A2(n_majority7_module_91__and_module_3_res), .ZN(
        n_majority7_module_91__or_module_5_res) );
  AND2_X1 u_majority7_module_91__and_module_6_U1 ( .A1(
        n_majority7_module_91__or_module_1_res), .A2(
        n_majority7_module_91__or_module_2_res), .ZN(
        n_majority7_module_91__and_module_6_res) );
  OR2_X1 u_majority7_module_91__or_module_6_U1 ( .A1(
        n_majority7_module_91__or_module_2_res), .A2(
        n_majority7_module_91__or_module_1_res), .ZN(
        n_majority7_module_91__or_module_6_res) );
  OR2_X1 u_majority7_module_91__or_module_7_U1 ( .A1(
        n_majority7_module_91__and_module_4_res), .A2(
        n_majority7_module_91__and_module_5_res), .ZN(
        n_majority7_module_91__or_module_7_res) );
  AND2_X1 u_majority7_module_91__and_module_7_U1 ( .A1(
        n_majority7_module_91__or_module_3_res), .A2(
        n_majority7_module_91__or_module_4_res), .ZN(
        n_majority7_module_91__and_module_7_res) );
  OR2_X1 u_majority7_module_91__or_module_8_U1 ( .A1(
        n_majority7_module_91__or_module_4_res), .A2(
        n_majority7_module_91__or_module_3_res), .ZN(
        n_majority7_module_91__or_module_8_res) );
  AND2_X1 u_majority7_module_91__and_module_8_U1 ( .A1(
        n_majority7_module_91__or_module_5_res), .A2(
        n_majority7_module_91__and_module_6_res), .ZN(
        n_majority7_module_91__and_module_8_res) );
  OR2_X1 u_majority7_module_91__or_module_9_U1 ( .A1(
        n_majority7_module_91__and_module_6_res), .A2(
        n_majority7_module_91__or_module_5_res), .ZN(
        n_majority7_module_91__or_module_9_res) );
  OR2_X1 u_majority7_module_91__or_module_10_U1 ( .A1(
        n_majority7_module_91__or_module_7_res), .A2(
        n_majority7_module_91__and_module_7_res), .ZN(
        n_majority7_module_91__or_module_10_res) );
  AND2_X1 u_majority7_module_91__and_module_9_U1 ( .A1(
        n_majority7_module_91__or_module_6_res), .A2(
        n_majority7_module_91__or_module_9_res), .ZN(
        n_majority7_module_91__and_module_9_res) );
  OR2_X1 u_majority7_module_91__or_module_11_U1 ( .A1(
        n_majority7_module_91__or_module_10_res), .A2(
        n_majority7_module_91__and_module_8_res), .ZN(
        n_majority7_module_91__or_module_11_res) );
  AND2_X1 u_majority7_module_91__and_module_10_U1 ( .A1(
        n_majority7_module_91__or_module_8_res), .A2(
        n_majority7_module_91__and_module_9_res), .ZN(
        n_majority7_module_91__and_module_10_res) );
  AND2_X1 u_majority7_module_91__and_module_11_U1 ( .A1(
        n_majority7_module_91__and_module_10_res), .A2(
        n_majority7_module_91__or_module_11_res), .ZN(
        n_majority7_module_91_res) );
  DFF_X1 u_reg_module_92__cini_mul_v000_reg ( .D(n_majority7_module_91_res), 
        .CK(clock_5), .Q(n_reg_module_92_res), .QN() );
  BUF_X1 u_majority7_module_92_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_92_n7) );
  BUF_X1 u_majority7_module_92_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_92_n6) );
  BUF_X1 u_majority7_module_92_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_92_n5) );
  BUF_X1 u_majority7_module_92_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_92_n4) );
  BUF_X1 u_majority7_module_92_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_92_n3) );
  BUF_X1 u_majority7_module_92_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_92_n2) );
  BUF_X1 u_majority7_module_92_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_92_n1) );
  AND2_X1 u_majority7_module_92__and_module_1_U1 ( .A1(
        n_majority7_module_92_n7), .A2(n_majority7_module_92_n1), .ZN(
        n_majority7_module_92__and_module_1_res) );
  OR2_X1 u_majority7_module_92__or_module_1_U1 ( .A1(n_majority7_module_92_n1), 
        .A2(n_majority7_module_92_n7), .ZN(
        n_majority7_module_92__or_module_1_res) );
  AND2_X1 u_majority7_module_92__and_module_2_U1 ( .A1(
        n_majority7_module_92_n5), .A2(n_majority7_module_92_n3), .ZN(
        n_majority7_module_92__and_module_2_res) );
  OR2_X1 u_majority7_module_92__or_module_2_U1 ( .A1(n_majority7_module_92_n3), 
        .A2(n_majority7_module_92_n5), .ZN(
        n_majority7_module_92__or_module_2_res) );
  AND2_X1 u_majority7_module_92__and_module_3_U1 ( .A1(
        n_majority7_module_92_n6), .A2(n_majority7_module_92_n4), .ZN(
        n_majority7_module_92__and_module_3_res) );
  OR2_X1 u_majority7_module_92__or_module_3_U1 ( .A1(n_majority7_module_92_n4), 
        .A2(n_majority7_module_92_n6), .ZN(
        n_majority7_module_92__or_module_3_res) );
  AND2_X1 u_majority7_module_92__and_module_4_U1 ( .A1(
        n_majority7_module_92__and_module_2_res), .A2(
        n_majority7_module_92__and_module_1_res), .ZN(
        n_majority7_module_92__and_module_4_res) );
  OR2_X1 u_majority7_module_92__or_module_4_U1 ( .A1(
        n_majority7_module_92__and_module_1_res), .A2(
        n_majority7_module_92__and_module_2_res), .ZN(
        n_majority7_module_92__or_module_4_res) );
  AND2_X1 u_majority7_module_92__and_module_5_U1 ( .A1(
        n_majority7_module_92__and_module_3_res), .A2(n_majority7_module_92_n2), .ZN(n_majority7_module_92__and_module_5_res) );
  OR2_X1 u_majority7_module_92__or_module_5_U1 ( .A1(n_majority7_module_92_n2), 
        .A2(n_majority7_module_92__and_module_3_res), .ZN(
        n_majority7_module_92__or_module_5_res) );
  AND2_X1 u_majority7_module_92__and_module_6_U1 ( .A1(
        n_majority7_module_92__or_module_1_res), .A2(
        n_majority7_module_92__or_module_2_res), .ZN(
        n_majority7_module_92__and_module_6_res) );
  OR2_X1 u_majority7_module_92__or_module_6_U1 ( .A1(
        n_majority7_module_92__or_module_2_res), .A2(
        n_majority7_module_92__or_module_1_res), .ZN(
        n_majority7_module_92__or_module_6_res) );
  OR2_X1 u_majority7_module_92__or_module_7_U1 ( .A1(
        n_majority7_module_92__and_module_4_res), .A2(
        n_majority7_module_92__and_module_5_res), .ZN(
        n_majority7_module_92__or_module_7_res) );
  AND2_X1 u_majority7_module_92__and_module_7_U1 ( .A1(
        n_majority7_module_92__or_module_3_res), .A2(
        n_majority7_module_92__or_module_4_res), .ZN(
        n_majority7_module_92__and_module_7_res) );
  OR2_X1 u_majority7_module_92__or_module_8_U1 ( .A1(
        n_majority7_module_92__or_module_4_res), .A2(
        n_majority7_module_92__or_module_3_res), .ZN(
        n_majority7_module_92__or_module_8_res) );
  AND2_X1 u_majority7_module_92__and_module_8_U1 ( .A1(
        n_majority7_module_92__or_module_5_res), .A2(
        n_majority7_module_92__and_module_6_res), .ZN(
        n_majority7_module_92__and_module_8_res) );
  OR2_X1 u_majority7_module_92__or_module_9_U1 ( .A1(
        n_majority7_module_92__and_module_6_res), .A2(
        n_majority7_module_92__or_module_5_res), .ZN(
        n_majority7_module_92__or_module_9_res) );
  OR2_X1 u_majority7_module_92__or_module_10_U1 ( .A1(
        n_majority7_module_92__or_module_7_res), .A2(
        n_majority7_module_92__and_module_7_res), .ZN(
        n_majority7_module_92__or_module_10_res) );
  AND2_X1 u_majority7_module_92__and_module_9_U1 ( .A1(
        n_majority7_module_92__or_module_6_res), .A2(
        n_majority7_module_92__or_module_9_res), .ZN(
        n_majority7_module_92__and_module_9_res) );
  OR2_X1 u_majority7_module_92__or_module_11_U1 ( .A1(
        n_majority7_module_92__or_module_10_res), .A2(
        n_majority7_module_92__and_module_8_res), .ZN(
        n_majority7_module_92__or_module_11_res) );
  AND2_X1 u_majority7_module_92__and_module_10_U1 ( .A1(
        n_majority7_module_92__or_module_8_res), .A2(
        n_majority7_module_92__and_module_9_res), .ZN(
        n_majority7_module_92__and_module_10_res) );
  AND2_X1 u_majority7_module_92__and_module_11_U1 ( .A1(
        n_majority7_module_92__and_module_10_res), .A2(
        n_majority7_module_92__or_module_11_res), .ZN(
        n_majority7_module_92_res) );
  DFF_X1 u_reg_module_93__cini_mul_v000_reg ( .D(n_majority7_module_92_res), 
        .CK(clock_5), .Q(n_reg_module_93_res), .QN() );
  BUF_X1 u_majority7_module_93_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_93_n7) );
  BUF_X1 u_majority7_module_93_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_93_n6) );
  BUF_X1 u_majority7_module_93_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_93_n5) );
  BUF_X1 u_majority7_module_93_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_93_n4) );
  BUF_X1 u_majority7_module_93_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_93_n3) );
  BUF_X1 u_majority7_module_93_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_93_n2) );
  BUF_X1 u_majority7_module_93_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_93_n1) );
  AND2_X1 u_majority7_module_93__and_module_1_U1 ( .A1(
        n_majority7_module_93_n7), .A2(n_majority7_module_93_n1), .ZN(
        n_majority7_module_93__and_module_1_res) );
  OR2_X1 u_majority7_module_93__or_module_1_U1 ( .A1(n_majority7_module_93_n1), 
        .A2(n_majority7_module_93_n7), .ZN(
        n_majority7_module_93__or_module_1_res) );
  AND2_X1 u_majority7_module_93__and_module_2_U1 ( .A1(
        n_majority7_module_93_n5), .A2(n_majority7_module_93_n3), .ZN(
        n_majority7_module_93__and_module_2_res) );
  OR2_X1 u_majority7_module_93__or_module_2_U1 ( .A1(n_majority7_module_93_n3), 
        .A2(n_majority7_module_93_n5), .ZN(
        n_majority7_module_93__or_module_2_res) );
  AND2_X1 u_majority7_module_93__and_module_3_U1 ( .A1(
        n_majority7_module_93_n6), .A2(n_majority7_module_93_n4), .ZN(
        n_majority7_module_93__and_module_3_res) );
  OR2_X1 u_majority7_module_93__or_module_3_U1 ( .A1(n_majority7_module_93_n4), 
        .A2(n_majority7_module_93_n6), .ZN(
        n_majority7_module_93__or_module_3_res) );
  AND2_X1 u_majority7_module_93__and_module_4_U1 ( .A1(
        n_majority7_module_93__and_module_2_res), .A2(
        n_majority7_module_93__and_module_1_res), .ZN(
        n_majority7_module_93__and_module_4_res) );
  OR2_X1 u_majority7_module_93__or_module_4_U1 ( .A1(
        n_majority7_module_93__and_module_1_res), .A2(
        n_majority7_module_93__and_module_2_res), .ZN(
        n_majority7_module_93__or_module_4_res) );
  AND2_X1 u_majority7_module_93__and_module_5_U1 ( .A1(
        n_majority7_module_93__and_module_3_res), .A2(n_majority7_module_93_n2), .ZN(n_majority7_module_93__and_module_5_res) );
  OR2_X1 u_majority7_module_93__or_module_5_U1 ( .A1(n_majority7_module_93_n2), 
        .A2(n_majority7_module_93__and_module_3_res), .ZN(
        n_majority7_module_93__or_module_5_res) );
  AND2_X1 u_majority7_module_93__and_module_6_U1 ( .A1(
        n_majority7_module_93__or_module_1_res), .A2(
        n_majority7_module_93__or_module_2_res), .ZN(
        n_majority7_module_93__and_module_6_res) );
  OR2_X1 u_majority7_module_93__or_module_6_U1 ( .A1(
        n_majority7_module_93__or_module_2_res), .A2(
        n_majority7_module_93__or_module_1_res), .ZN(
        n_majority7_module_93__or_module_6_res) );
  OR2_X1 u_majority7_module_93__or_module_7_U1 ( .A1(
        n_majority7_module_93__and_module_4_res), .A2(
        n_majority7_module_93__and_module_5_res), .ZN(
        n_majority7_module_93__or_module_7_res) );
  AND2_X1 u_majority7_module_93__and_module_7_U1 ( .A1(
        n_majority7_module_93__or_module_3_res), .A2(
        n_majority7_module_93__or_module_4_res), .ZN(
        n_majority7_module_93__and_module_7_res) );
  OR2_X1 u_majority7_module_93__or_module_8_U1 ( .A1(
        n_majority7_module_93__or_module_4_res), .A2(
        n_majority7_module_93__or_module_3_res), .ZN(
        n_majority7_module_93__or_module_8_res) );
  AND2_X1 u_majority7_module_93__and_module_8_U1 ( .A1(
        n_majority7_module_93__or_module_5_res), .A2(
        n_majority7_module_93__and_module_6_res), .ZN(
        n_majority7_module_93__and_module_8_res) );
  OR2_X1 u_majority7_module_93__or_module_9_U1 ( .A1(
        n_majority7_module_93__and_module_6_res), .A2(
        n_majority7_module_93__or_module_5_res), .ZN(
        n_majority7_module_93__or_module_9_res) );
  OR2_X1 u_majority7_module_93__or_module_10_U1 ( .A1(
        n_majority7_module_93__or_module_7_res), .A2(
        n_majority7_module_93__and_module_7_res), .ZN(
        n_majority7_module_93__or_module_10_res) );
  AND2_X1 u_majority7_module_93__and_module_9_U1 ( .A1(
        n_majority7_module_93__or_module_6_res), .A2(
        n_majority7_module_93__or_module_9_res), .ZN(
        n_majority7_module_93__and_module_9_res) );
  OR2_X1 u_majority7_module_93__or_module_11_U1 ( .A1(
        n_majority7_module_93__or_module_10_res), .A2(
        n_majority7_module_93__and_module_8_res), .ZN(
        n_majority7_module_93__or_module_11_res) );
  AND2_X1 u_majority7_module_93__and_module_10_U1 ( .A1(
        n_majority7_module_93__or_module_8_res), .A2(
        n_majority7_module_93__and_module_9_res), .ZN(
        n_majority7_module_93__and_module_10_res) );
  AND2_X1 u_majority7_module_93__and_module_11_U1 ( .A1(
        n_majority7_module_93__and_module_10_res), .A2(
        n_majority7_module_93__or_module_11_res), .ZN(
        n_majority7_module_93_res) );
  DFF_X1 u_reg_module_94__cini_mul_v000_reg ( .D(n_majority7_module_93_res), 
        .CK(clock_5), .Q(n_reg_module_94_res), .QN() );
  BUF_X1 u_majority7_module_94_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_94_n7) );
  BUF_X1 u_majority7_module_94_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_94_n6) );
  BUF_X1 u_majority7_module_94_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_94_n5) );
  BUF_X1 u_majority7_module_94_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_94_n4) );
  BUF_X1 u_majority7_module_94_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_94_n3) );
  BUF_X1 u_majority7_module_94_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_94_n2) );
  BUF_X1 u_majority7_module_94_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_94_n1) );
  AND2_X1 u_majority7_module_94__and_module_1_U1 ( .A1(
        n_majority7_module_94_n7), .A2(n_majority7_module_94_n1), .ZN(
        n_majority7_module_94__and_module_1_res) );
  OR2_X1 u_majority7_module_94__or_module_1_U1 ( .A1(n_majority7_module_94_n1), 
        .A2(n_majority7_module_94_n7), .ZN(
        n_majority7_module_94__or_module_1_res) );
  AND2_X1 u_majority7_module_94__and_module_2_U1 ( .A1(
        n_majority7_module_94_n5), .A2(n_majority7_module_94_n3), .ZN(
        n_majority7_module_94__and_module_2_res) );
  OR2_X1 u_majority7_module_94__or_module_2_U1 ( .A1(n_majority7_module_94_n3), 
        .A2(n_majority7_module_94_n5), .ZN(
        n_majority7_module_94__or_module_2_res) );
  AND2_X1 u_majority7_module_94__and_module_3_U1 ( .A1(
        n_majority7_module_94_n6), .A2(n_majority7_module_94_n4), .ZN(
        n_majority7_module_94__and_module_3_res) );
  OR2_X1 u_majority7_module_94__or_module_3_U1 ( .A1(n_majority7_module_94_n4), 
        .A2(n_majority7_module_94_n6), .ZN(
        n_majority7_module_94__or_module_3_res) );
  AND2_X1 u_majority7_module_94__and_module_4_U1 ( .A1(
        n_majority7_module_94__and_module_2_res), .A2(
        n_majority7_module_94__and_module_1_res), .ZN(
        n_majority7_module_94__and_module_4_res) );
  OR2_X1 u_majority7_module_94__or_module_4_U1 ( .A1(
        n_majority7_module_94__and_module_1_res), .A2(
        n_majority7_module_94__and_module_2_res), .ZN(
        n_majority7_module_94__or_module_4_res) );
  AND2_X1 u_majority7_module_94__and_module_5_U1 ( .A1(
        n_majority7_module_94__and_module_3_res), .A2(n_majority7_module_94_n2), .ZN(n_majority7_module_94__and_module_5_res) );
  OR2_X1 u_majority7_module_94__or_module_5_U1 ( .A1(n_majority7_module_94_n2), 
        .A2(n_majority7_module_94__and_module_3_res), .ZN(
        n_majority7_module_94__or_module_5_res) );
  AND2_X1 u_majority7_module_94__and_module_6_U1 ( .A1(
        n_majority7_module_94__or_module_1_res), .A2(
        n_majority7_module_94__or_module_2_res), .ZN(
        n_majority7_module_94__and_module_6_res) );
  OR2_X1 u_majority7_module_94__or_module_6_U1 ( .A1(
        n_majority7_module_94__or_module_2_res), .A2(
        n_majority7_module_94__or_module_1_res), .ZN(
        n_majority7_module_94__or_module_6_res) );
  OR2_X1 u_majority7_module_94__or_module_7_U1 ( .A1(
        n_majority7_module_94__and_module_4_res), .A2(
        n_majority7_module_94__and_module_5_res), .ZN(
        n_majority7_module_94__or_module_7_res) );
  AND2_X1 u_majority7_module_94__and_module_7_U1 ( .A1(
        n_majority7_module_94__or_module_3_res), .A2(
        n_majority7_module_94__or_module_4_res), .ZN(
        n_majority7_module_94__and_module_7_res) );
  OR2_X1 u_majority7_module_94__or_module_8_U1 ( .A1(
        n_majority7_module_94__or_module_4_res), .A2(
        n_majority7_module_94__or_module_3_res), .ZN(
        n_majority7_module_94__or_module_8_res) );
  AND2_X1 u_majority7_module_94__and_module_8_U1 ( .A1(
        n_majority7_module_94__or_module_5_res), .A2(
        n_majority7_module_94__and_module_6_res), .ZN(
        n_majority7_module_94__and_module_8_res) );
  OR2_X1 u_majority7_module_94__or_module_9_U1 ( .A1(
        n_majority7_module_94__and_module_6_res), .A2(
        n_majority7_module_94__or_module_5_res), .ZN(
        n_majority7_module_94__or_module_9_res) );
  OR2_X1 u_majority7_module_94__or_module_10_U1 ( .A1(
        n_majority7_module_94__or_module_7_res), .A2(
        n_majority7_module_94__and_module_7_res), .ZN(
        n_majority7_module_94__or_module_10_res) );
  AND2_X1 u_majority7_module_94__and_module_9_U1 ( .A1(
        n_majority7_module_94__or_module_6_res), .A2(
        n_majority7_module_94__or_module_9_res), .ZN(
        n_majority7_module_94__and_module_9_res) );
  OR2_X1 u_majority7_module_94__or_module_11_U1 ( .A1(
        n_majority7_module_94__or_module_10_res), .A2(
        n_majority7_module_94__and_module_8_res), .ZN(
        n_majority7_module_94__or_module_11_res) );
  AND2_X1 u_majority7_module_94__and_module_10_U1 ( .A1(
        n_majority7_module_94__or_module_8_res), .A2(
        n_majority7_module_94__and_module_9_res), .ZN(
        n_majority7_module_94__and_module_10_res) );
  AND2_X1 u_majority7_module_94__and_module_11_U1 ( .A1(
        n_majority7_module_94__and_module_10_res), .A2(
        n_majority7_module_94__or_module_11_res), .ZN(
        n_majority7_module_94_res) );
  DFF_X1 u_reg_module_95__cini_mul_v000_reg ( .D(n_majority7_module_94_res), 
        .CK(clock_5), .Q(n_reg_module_95_res), .QN() );
  BUF_X1 u_majority7_module_95_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_95_n7) );
  BUF_X1 u_majority7_module_95_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_95_n6) );
  BUF_X1 u_majority7_module_95_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_95_n5) );
  BUF_X1 u_majority7_module_95_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_95_n4) );
  BUF_X1 u_majority7_module_95_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_95_n3) );
  BUF_X1 u_majority7_module_95_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_95_n2) );
  BUF_X1 u_majority7_module_95_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_95_n1) );
  AND2_X1 u_majority7_module_95__and_module_1_U1 ( .A1(
        n_majority7_module_95_n7), .A2(n_majority7_module_95_n1), .ZN(
        n_majority7_module_95__and_module_1_res) );
  OR2_X1 u_majority7_module_95__or_module_1_U1 ( .A1(n_majority7_module_95_n1), 
        .A2(n_majority7_module_95_n7), .ZN(
        n_majority7_module_95__or_module_1_res) );
  AND2_X1 u_majority7_module_95__and_module_2_U1 ( .A1(
        n_majority7_module_95_n5), .A2(n_majority7_module_95_n3), .ZN(
        n_majority7_module_95__and_module_2_res) );
  OR2_X1 u_majority7_module_95__or_module_2_U1 ( .A1(n_majority7_module_95_n3), 
        .A2(n_majority7_module_95_n5), .ZN(
        n_majority7_module_95__or_module_2_res) );
  AND2_X1 u_majority7_module_95__and_module_3_U1 ( .A1(
        n_majority7_module_95_n6), .A2(n_majority7_module_95_n4), .ZN(
        n_majority7_module_95__and_module_3_res) );
  OR2_X1 u_majority7_module_95__or_module_3_U1 ( .A1(n_majority7_module_95_n4), 
        .A2(n_majority7_module_95_n6), .ZN(
        n_majority7_module_95__or_module_3_res) );
  AND2_X1 u_majority7_module_95__and_module_4_U1 ( .A1(
        n_majority7_module_95__and_module_2_res), .A2(
        n_majority7_module_95__and_module_1_res), .ZN(
        n_majority7_module_95__and_module_4_res) );
  OR2_X1 u_majority7_module_95__or_module_4_U1 ( .A1(
        n_majority7_module_95__and_module_1_res), .A2(
        n_majority7_module_95__and_module_2_res), .ZN(
        n_majority7_module_95__or_module_4_res) );
  AND2_X1 u_majority7_module_95__and_module_5_U1 ( .A1(
        n_majority7_module_95__and_module_3_res), .A2(n_majority7_module_95_n2), .ZN(n_majority7_module_95__and_module_5_res) );
  OR2_X1 u_majority7_module_95__or_module_5_U1 ( .A1(n_majority7_module_95_n2), 
        .A2(n_majority7_module_95__and_module_3_res), .ZN(
        n_majority7_module_95__or_module_5_res) );
  AND2_X1 u_majority7_module_95__and_module_6_U1 ( .A1(
        n_majority7_module_95__or_module_1_res), .A2(
        n_majority7_module_95__or_module_2_res), .ZN(
        n_majority7_module_95__and_module_6_res) );
  OR2_X1 u_majority7_module_95__or_module_6_U1 ( .A1(
        n_majority7_module_95__or_module_2_res), .A2(
        n_majority7_module_95__or_module_1_res), .ZN(
        n_majority7_module_95__or_module_6_res) );
  OR2_X1 u_majority7_module_95__or_module_7_U1 ( .A1(
        n_majority7_module_95__and_module_4_res), .A2(
        n_majority7_module_95__and_module_5_res), .ZN(
        n_majority7_module_95__or_module_7_res) );
  AND2_X1 u_majority7_module_95__and_module_7_U1 ( .A1(
        n_majority7_module_95__or_module_3_res), .A2(
        n_majority7_module_95__or_module_4_res), .ZN(
        n_majority7_module_95__and_module_7_res) );
  OR2_X1 u_majority7_module_95__or_module_8_U1 ( .A1(
        n_majority7_module_95__or_module_4_res), .A2(
        n_majority7_module_95__or_module_3_res), .ZN(
        n_majority7_module_95__or_module_8_res) );
  AND2_X1 u_majority7_module_95__and_module_8_U1 ( .A1(
        n_majority7_module_95__or_module_5_res), .A2(
        n_majority7_module_95__and_module_6_res), .ZN(
        n_majority7_module_95__and_module_8_res) );
  OR2_X1 u_majority7_module_95__or_module_9_U1 ( .A1(
        n_majority7_module_95__and_module_6_res), .A2(
        n_majority7_module_95__or_module_5_res), .ZN(
        n_majority7_module_95__or_module_9_res) );
  OR2_X1 u_majority7_module_95__or_module_10_U1 ( .A1(
        n_majority7_module_95__or_module_7_res), .A2(
        n_majority7_module_95__and_module_7_res), .ZN(
        n_majority7_module_95__or_module_10_res) );
  AND2_X1 u_majority7_module_95__and_module_9_U1 ( .A1(
        n_majority7_module_95__or_module_6_res), .A2(
        n_majority7_module_95__or_module_9_res), .ZN(
        n_majority7_module_95__and_module_9_res) );
  OR2_X1 u_majority7_module_95__or_module_11_U1 ( .A1(
        n_majority7_module_95__or_module_10_res), .A2(
        n_majority7_module_95__and_module_8_res), .ZN(
        n_majority7_module_95__or_module_11_res) );
  AND2_X1 u_majority7_module_95__and_module_10_U1 ( .A1(
        n_majority7_module_95__or_module_8_res), .A2(
        n_majority7_module_95__and_module_9_res), .ZN(
        n_majority7_module_95__and_module_10_res) );
  AND2_X1 u_majority7_module_95__and_module_11_U1 ( .A1(
        n_majority7_module_95__and_module_10_res), .A2(
        n_majority7_module_95__or_module_11_res), .ZN(
        n_majority7_module_95_res) );
  DFF_X1 u_reg_module_96__cini_mul_v000_reg ( .D(n_majority7_module_95_res), 
        .CK(clock_5), .Q(n_reg_module_96_res), .QN() );
  BUF_X1 u_majority7_module_96_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_96_n7) );
  BUF_X1 u_majority7_module_96_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_96_n6) );
  BUF_X1 u_majority7_module_96_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_96_n5) );
  BUF_X1 u_majority7_module_96_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_96_n4) );
  BUF_X1 u_majority7_module_96_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_96_n3) );
  BUF_X1 u_majority7_module_96_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_96_n2) );
  BUF_X1 u_majority7_module_96_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_96_n1) );
  AND2_X1 u_majority7_module_96__and_module_1_U1 ( .A1(
        n_majority7_module_96_n7), .A2(n_majority7_module_96_n1), .ZN(
        n_majority7_module_96__and_module_1_res) );
  OR2_X1 u_majority7_module_96__or_module_1_U1 ( .A1(n_majority7_module_96_n1), 
        .A2(n_majority7_module_96_n7), .ZN(
        n_majority7_module_96__or_module_1_res) );
  AND2_X1 u_majority7_module_96__and_module_2_U1 ( .A1(
        n_majority7_module_96_n5), .A2(n_majority7_module_96_n3), .ZN(
        n_majority7_module_96__and_module_2_res) );
  OR2_X1 u_majority7_module_96__or_module_2_U1 ( .A1(n_majority7_module_96_n3), 
        .A2(n_majority7_module_96_n5), .ZN(
        n_majority7_module_96__or_module_2_res) );
  AND2_X1 u_majority7_module_96__and_module_3_U1 ( .A1(
        n_majority7_module_96_n6), .A2(n_majority7_module_96_n4), .ZN(
        n_majority7_module_96__and_module_3_res) );
  OR2_X1 u_majority7_module_96__or_module_3_U1 ( .A1(n_majority7_module_96_n4), 
        .A2(n_majority7_module_96_n6), .ZN(
        n_majority7_module_96__or_module_3_res) );
  AND2_X1 u_majority7_module_96__and_module_4_U1 ( .A1(
        n_majority7_module_96__and_module_2_res), .A2(
        n_majority7_module_96__and_module_1_res), .ZN(
        n_majority7_module_96__and_module_4_res) );
  OR2_X1 u_majority7_module_96__or_module_4_U1 ( .A1(
        n_majority7_module_96__and_module_1_res), .A2(
        n_majority7_module_96__and_module_2_res), .ZN(
        n_majority7_module_96__or_module_4_res) );
  AND2_X1 u_majority7_module_96__and_module_5_U1 ( .A1(
        n_majority7_module_96__and_module_3_res), .A2(n_majority7_module_96_n2), .ZN(n_majority7_module_96__and_module_5_res) );
  OR2_X1 u_majority7_module_96__or_module_5_U1 ( .A1(n_majority7_module_96_n2), 
        .A2(n_majority7_module_96__and_module_3_res), .ZN(
        n_majority7_module_96__or_module_5_res) );
  AND2_X1 u_majority7_module_96__and_module_6_U1 ( .A1(
        n_majority7_module_96__or_module_1_res), .A2(
        n_majority7_module_96__or_module_2_res), .ZN(
        n_majority7_module_96__and_module_6_res) );
  OR2_X1 u_majority7_module_96__or_module_6_U1 ( .A1(
        n_majority7_module_96__or_module_2_res), .A2(
        n_majority7_module_96__or_module_1_res), .ZN(
        n_majority7_module_96__or_module_6_res) );
  OR2_X1 u_majority7_module_96__or_module_7_U1 ( .A1(
        n_majority7_module_96__and_module_4_res), .A2(
        n_majority7_module_96__and_module_5_res), .ZN(
        n_majority7_module_96__or_module_7_res) );
  AND2_X1 u_majority7_module_96__and_module_7_U1 ( .A1(
        n_majority7_module_96__or_module_3_res), .A2(
        n_majority7_module_96__or_module_4_res), .ZN(
        n_majority7_module_96__and_module_7_res) );
  OR2_X1 u_majority7_module_96__or_module_8_U1 ( .A1(
        n_majority7_module_96__or_module_4_res), .A2(
        n_majority7_module_96__or_module_3_res), .ZN(
        n_majority7_module_96__or_module_8_res) );
  AND2_X1 u_majority7_module_96__and_module_8_U1 ( .A1(
        n_majority7_module_96__or_module_5_res), .A2(
        n_majority7_module_96__and_module_6_res), .ZN(
        n_majority7_module_96__and_module_8_res) );
  OR2_X1 u_majority7_module_96__or_module_9_U1 ( .A1(
        n_majority7_module_96__and_module_6_res), .A2(
        n_majority7_module_96__or_module_5_res), .ZN(
        n_majority7_module_96__or_module_9_res) );
  OR2_X1 u_majority7_module_96__or_module_10_U1 ( .A1(
        n_majority7_module_96__or_module_7_res), .A2(
        n_majority7_module_96__and_module_7_res), .ZN(
        n_majority7_module_96__or_module_10_res) );
  AND2_X1 u_majority7_module_96__and_module_9_U1 ( .A1(
        n_majority7_module_96__or_module_6_res), .A2(
        n_majority7_module_96__or_module_9_res), .ZN(
        n_majority7_module_96__and_module_9_res) );
  OR2_X1 u_majority7_module_96__or_module_11_U1 ( .A1(
        n_majority7_module_96__or_module_10_res), .A2(
        n_majority7_module_96__and_module_8_res), .ZN(
        n_majority7_module_96__or_module_11_res) );
  AND2_X1 u_majority7_module_96__and_module_10_U1 ( .A1(
        n_majority7_module_96__or_module_8_res), .A2(
        n_majority7_module_96__and_module_9_res), .ZN(
        n_majority7_module_96__and_module_10_res) );
  AND2_X1 u_majority7_module_96__and_module_11_U1 ( .A1(
        n_majority7_module_96__and_module_10_res), .A2(
        n_majority7_module_96__or_module_11_res), .ZN(
        n_majority7_module_96_res) );
  DFF_X1 u_reg_module_97__cini_mul_v000_reg ( .D(n_majority7_module_96_res), 
        .CK(clock_6), .Q(n_reg_module_97_res), .QN() );
  BUF_X1 u_majority7_module_97_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_97_n7) );
  BUF_X1 u_majority7_module_97_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_97_n6) );
  BUF_X1 u_majority7_module_97_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_97_n5) );
  BUF_X1 u_majority7_module_97_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_97_n4) );
  BUF_X1 u_majority7_module_97_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_97_n3) );
  BUF_X1 u_majority7_module_97_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_97_n2) );
  BUF_X1 u_majority7_module_97_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_97_n1) );
  AND2_X1 u_majority7_module_97__and_module_1_U1 ( .A1(
        n_majority7_module_97_n7), .A2(n_majority7_module_97_n1), .ZN(
        n_majority7_module_97__and_module_1_res) );
  OR2_X1 u_majority7_module_97__or_module_1_U1 ( .A1(n_majority7_module_97_n1), 
        .A2(n_majority7_module_97_n7), .ZN(
        n_majority7_module_97__or_module_1_res) );
  AND2_X1 u_majority7_module_97__and_module_2_U1 ( .A1(
        n_majority7_module_97_n5), .A2(n_majority7_module_97_n3), .ZN(
        n_majority7_module_97__and_module_2_res) );
  OR2_X1 u_majority7_module_97__or_module_2_U1 ( .A1(n_majority7_module_97_n3), 
        .A2(n_majority7_module_97_n5), .ZN(
        n_majority7_module_97__or_module_2_res) );
  AND2_X1 u_majority7_module_97__and_module_3_U1 ( .A1(
        n_majority7_module_97_n6), .A2(n_majority7_module_97_n4), .ZN(
        n_majority7_module_97__and_module_3_res) );
  OR2_X1 u_majority7_module_97__or_module_3_U1 ( .A1(n_majority7_module_97_n4), 
        .A2(n_majority7_module_97_n6), .ZN(
        n_majority7_module_97__or_module_3_res) );
  AND2_X1 u_majority7_module_97__and_module_4_U1 ( .A1(
        n_majority7_module_97__and_module_2_res), .A2(
        n_majority7_module_97__and_module_1_res), .ZN(
        n_majority7_module_97__and_module_4_res) );
  OR2_X1 u_majority7_module_97__or_module_4_U1 ( .A1(
        n_majority7_module_97__and_module_1_res), .A2(
        n_majority7_module_97__and_module_2_res), .ZN(
        n_majority7_module_97__or_module_4_res) );
  AND2_X1 u_majority7_module_97__and_module_5_U1 ( .A1(
        n_majority7_module_97__and_module_3_res), .A2(n_majority7_module_97_n2), .ZN(n_majority7_module_97__and_module_5_res) );
  OR2_X1 u_majority7_module_97__or_module_5_U1 ( .A1(n_majority7_module_97_n2), 
        .A2(n_majority7_module_97__and_module_3_res), .ZN(
        n_majority7_module_97__or_module_5_res) );
  AND2_X1 u_majority7_module_97__and_module_6_U1 ( .A1(
        n_majority7_module_97__or_module_1_res), .A2(
        n_majority7_module_97__or_module_2_res), .ZN(
        n_majority7_module_97__and_module_6_res) );
  OR2_X1 u_majority7_module_97__or_module_6_U1 ( .A1(
        n_majority7_module_97__or_module_2_res), .A2(
        n_majority7_module_97__or_module_1_res), .ZN(
        n_majority7_module_97__or_module_6_res) );
  OR2_X1 u_majority7_module_97__or_module_7_U1 ( .A1(
        n_majority7_module_97__and_module_4_res), .A2(
        n_majority7_module_97__and_module_5_res), .ZN(
        n_majority7_module_97__or_module_7_res) );
  AND2_X1 u_majority7_module_97__and_module_7_U1 ( .A1(
        n_majority7_module_97__or_module_3_res), .A2(
        n_majority7_module_97__or_module_4_res), .ZN(
        n_majority7_module_97__and_module_7_res) );
  OR2_X1 u_majority7_module_97__or_module_8_U1 ( .A1(
        n_majority7_module_97__or_module_4_res), .A2(
        n_majority7_module_97__or_module_3_res), .ZN(
        n_majority7_module_97__or_module_8_res) );
  AND2_X1 u_majority7_module_97__and_module_8_U1 ( .A1(
        n_majority7_module_97__or_module_5_res), .A2(
        n_majority7_module_97__and_module_6_res), .ZN(
        n_majority7_module_97__and_module_8_res) );
  OR2_X1 u_majority7_module_97__or_module_9_U1 ( .A1(
        n_majority7_module_97__and_module_6_res), .A2(
        n_majority7_module_97__or_module_5_res), .ZN(
        n_majority7_module_97__or_module_9_res) );
  OR2_X1 u_majority7_module_97__or_module_10_U1 ( .A1(
        n_majority7_module_97__or_module_7_res), .A2(
        n_majority7_module_97__and_module_7_res), .ZN(
        n_majority7_module_97__or_module_10_res) );
  AND2_X1 u_majority7_module_97__and_module_9_U1 ( .A1(
        n_majority7_module_97__or_module_6_res), .A2(
        n_majority7_module_97__or_module_9_res), .ZN(
        n_majority7_module_97__and_module_9_res) );
  OR2_X1 u_majority7_module_97__or_module_11_U1 ( .A1(
        n_majority7_module_97__or_module_10_res), .A2(
        n_majority7_module_97__and_module_8_res), .ZN(
        n_majority7_module_97__or_module_11_res) );
  AND2_X1 u_majority7_module_97__and_module_10_U1 ( .A1(
        n_majority7_module_97__or_module_8_res), .A2(
        n_majority7_module_97__and_module_9_res), .ZN(
        n_majority7_module_97__and_module_10_res) );
  AND2_X1 u_majority7_module_97__and_module_11_U1 ( .A1(
        n_majority7_module_97__and_module_10_res), .A2(
        n_majority7_module_97__or_module_11_res), .ZN(
        n_majority7_module_97_res) );
  DFF_X1 u_reg_module_98__cini_mul_v000_reg ( .D(n_majority7_module_97_res), 
        .CK(clock_6), .Q(n_reg_module_98_res), .QN() );
  BUF_X1 u_majority7_module_98_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_98_n7) );
  BUF_X1 u_majority7_module_98_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_98_n6) );
  BUF_X1 u_majority7_module_98_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_98_n5) );
  BUF_X1 u_majority7_module_98_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_98_n4) );
  BUF_X1 u_majority7_module_98_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_98_n3) );
  BUF_X1 u_majority7_module_98_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_98_n2) );
  BUF_X1 u_majority7_module_98_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_98_n1) );
  AND2_X1 u_majority7_module_98__and_module_1_U1 ( .A1(
        n_majority7_module_98_n7), .A2(n_majority7_module_98_n1), .ZN(
        n_majority7_module_98__and_module_1_res) );
  OR2_X1 u_majority7_module_98__or_module_1_U1 ( .A1(n_majority7_module_98_n1), 
        .A2(n_majority7_module_98_n7), .ZN(
        n_majority7_module_98__or_module_1_res) );
  AND2_X1 u_majority7_module_98__and_module_2_U1 ( .A1(
        n_majority7_module_98_n5), .A2(n_majority7_module_98_n3), .ZN(
        n_majority7_module_98__and_module_2_res) );
  OR2_X1 u_majority7_module_98__or_module_2_U1 ( .A1(n_majority7_module_98_n3), 
        .A2(n_majority7_module_98_n5), .ZN(
        n_majority7_module_98__or_module_2_res) );
  AND2_X1 u_majority7_module_98__and_module_3_U1 ( .A1(
        n_majority7_module_98_n6), .A2(n_majority7_module_98_n4), .ZN(
        n_majority7_module_98__and_module_3_res) );
  OR2_X1 u_majority7_module_98__or_module_3_U1 ( .A1(n_majority7_module_98_n4), 
        .A2(n_majority7_module_98_n6), .ZN(
        n_majority7_module_98__or_module_3_res) );
  AND2_X1 u_majority7_module_98__and_module_4_U1 ( .A1(
        n_majority7_module_98__and_module_2_res), .A2(
        n_majority7_module_98__and_module_1_res), .ZN(
        n_majority7_module_98__and_module_4_res) );
  OR2_X1 u_majority7_module_98__or_module_4_U1 ( .A1(
        n_majority7_module_98__and_module_1_res), .A2(
        n_majority7_module_98__and_module_2_res), .ZN(
        n_majority7_module_98__or_module_4_res) );
  AND2_X1 u_majority7_module_98__and_module_5_U1 ( .A1(
        n_majority7_module_98__and_module_3_res), .A2(n_majority7_module_98_n2), .ZN(n_majority7_module_98__and_module_5_res) );
  OR2_X1 u_majority7_module_98__or_module_5_U1 ( .A1(n_majority7_module_98_n2), 
        .A2(n_majority7_module_98__and_module_3_res), .ZN(
        n_majority7_module_98__or_module_5_res) );
  AND2_X1 u_majority7_module_98__and_module_6_U1 ( .A1(
        n_majority7_module_98__or_module_1_res), .A2(
        n_majority7_module_98__or_module_2_res), .ZN(
        n_majority7_module_98__and_module_6_res) );
  OR2_X1 u_majority7_module_98__or_module_6_U1 ( .A1(
        n_majority7_module_98__or_module_2_res), .A2(
        n_majority7_module_98__or_module_1_res), .ZN(
        n_majority7_module_98__or_module_6_res) );
  OR2_X1 u_majority7_module_98__or_module_7_U1 ( .A1(
        n_majority7_module_98__and_module_4_res), .A2(
        n_majority7_module_98__and_module_5_res), .ZN(
        n_majority7_module_98__or_module_7_res) );
  AND2_X1 u_majority7_module_98__and_module_7_U1 ( .A1(
        n_majority7_module_98__or_module_3_res), .A2(
        n_majority7_module_98__or_module_4_res), .ZN(
        n_majority7_module_98__and_module_7_res) );
  OR2_X1 u_majority7_module_98__or_module_8_U1 ( .A1(
        n_majority7_module_98__or_module_4_res), .A2(
        n_majority7_module_98__or_module_3_res), .ZN(
        n_majority7_module_98__or_module_8_res) );
  AND2_X1 u_majority7_module_98__and_module_8_U1 ( .A1(
        n_majority7_module_98__or_module_5_res), .A2(
        n_majority7_module_98__and_module_6_res), .ZN(
        n_majority7_module_98__and_module_8_res) );
  OR2_X1 u_majority7_module_98__or_module_9_U1 ( .A1(
        n_majority7_module_98__and_module_6_res), .A2(
        n_majority7_module_98__or_module_5_res), .ZN(
        n_majority7_module_98__or_module_9_res) );
  OR2_X1 u_majority7_module_98__or_module_10_U1 ( .A1(
        n_majority7_module_98__or_module_7_res), .A2(
        n_majority7_module_98__and_module_7_res), .ZN(
        n_majority7_module_98__or_module_10_res) );
  AND2_X1 u_majority7_module_98__and_module_9_U1 ( .A1(
        n_majority7_module_98__or_module_6_res), .A2(
        n_majority7_module_98__or_module_9_res), .ZN(
        n_majority7_module_98__and_module_9_res) );
  OR2_X1 u_majority7_module_98__or_module_11_U1 ( .A1(
        n_majority7_module_98__or_module_10_res), .A2(
        n_majority7_module_98__and_module_8_res), .ZN(
        n_majority7_module_98__or_module_11_res) );
  AND2_X1 u_majority7_module_98__and_module_10_U1 ( .A1(
        n_majority7_module_98__or_module_8_res), .A2(
        n_majority7_module_98__and_module_9_res), .ZN(
        n_majority7_module_98__and_module_10_res) );
  AND2_X1 u_majority7_module_98__and_module_11_U1 ( .A1(
        n_majority7_module_98__and_module_10_res), .A2(
        n_majority7_module_98__or_module_11_res), .ZN(
        n_majority7_module_98_res) );
  DFF_X1 u_reg_module_99__cini_mul_v000_reg ( .D(n_majority7_module_98_res), 
        .CK(clock_6), .Q(n_reg_module_99_res), .QN() );
  BUF_X1 u_majority7_module_99_U7 ( .A(n_xor_module_75_res), .Z(
        n_majority7_module_99_n7) );
  BUF_X1 u_majority7_module_99_U6 ( .A(n_xor_module_63_res), .Z(
        n_majority7_module_99_n6) );
  BUF_X1 u_majority7_module_99_U5 ( .A(n_xor_module_39_res), .Z(
        n_majority7_module_99_n5) );
  BUF_X1 u_majority7_module_99_U4 ( .A(n_xor_module_51_res), .Z(
        n_majority7_module_99_n4) );
  BUF_X1 u_majority7_module_99_U3 ( .A(n_xor_module_27_res), .Z(
        n_majority7_module_99_n3) );
  BUF_X1 u_majority7_module_99_U2 ( .A(n_xor_module_15_res), .Z(
        n_majority7_module_99_n2) );
  BUF_X1 u_majority7_module_99_U1 ( .A(n_xor_module_3_res), .Z(
        n_majority7_module_99_n1) );
  AND2_X1 u_majority7_module_99__and_module_1_U1 ( .A1(
        n_majority7_module_99_n7), .A2(n_majority7_module_99_n1), .ZN(
        n_majority7_module_99__and_module_1_res) );
  OR2_X1 u_majority7_module_99__or_module_1_U1 ( .A1(n_majority7_module_99_n1), 
        .A2(n_majority7_module_99_n7), .ZN(
        n_majority7_module_99__or_module_1_res) );
  AND2_X1 u_majority7_module_99__and_module_2_U1 ( .A1(
        n_majority7_module_99_n5), .A2(n_majority7_module_99_n3), .ZN(
        n_majority7_module_99__and_module_2_res) );
  OR2_X1 u_majority7_module_99__or_module_2_U1 ( .A1(n_majority7_module_99_n3), 
        .A2(n_majority7_module_99_n5), .ZN(
        n_majority7_module_99__or_module_2_res) );
  AND2_X1 u_majority7_module_99__and_module_3_U1 ( .A1(
        n_majority7_module_99_n6), .A2(n_majority7_module_99_n4), .ZN(
        n_majority7_module_99__and_module_3_res) );
  OR2_X1 u_majority7_module_99__or_module_3_U1 ( .A1(n_majority7_module_99_n4), 
        .A2(n_majority7_module_99_n6), .ZN(
        n_majority7_module_99__or_module_3_res) );
  AND2_X1 u_majority7_module_99__and_module_4_U1 ( .A1(
        n_majority7_module_99__and_module_2_res), .A2(
        n_majority7_module_99__and_module_1_res), .ZN(
        n_majority7_module_99__and_module_4_res) );
  OR2_X1 u_majority7_module_99__or_module_4_U1 ( .A1(
        n_majority7_module_99__and_module_1_res), .A2(
        n_majority7_module_99__and_module_2_res), .ZN(
        n_majority7_module_99__or_module_4_res) );
  AND2_X1 u_majority7_module_99__and_module_5_U1 ( .A1(
        n_majority7_module_99__and_module_3_res), .A2(n_majority7_module_99_n2), .ZN(n_majority7_module_99__and_module_5_res) );
  OR2_X1 u_majority7_module_99__or_module_5_U1 ( .A1(n_majority7_module_99_n2), 
        .A2(n_majority7_module_99__and_module_3_res), .ZN(
        n_majority7_module_99__or_module_5_res) );
  AND2_X1 u_majority7_module_99__and_module_6_U1 ( .A1(
        n_majority7_module_99__or_module_1_res), .A2(
        n_majority7_module_99__or_module_2_res), .ZN(
        n_majority7_module_99__and_module_6_res) );
  OR2_X1 u_majority7_module_99__or_module_6_U1 ( .A1(
        n_majority7_module_99__or_module_2_res), .A2(
        n_majority7_module_99__or_module_1_res), .ZN(
        n_majority7_module_99__or_module_6_res) );
  OR2_X1 u_majority7_module_99__or_module_7_U1 ( .A1(
        n_majority7_module_99__and_module_4_res), .A2(
        n_majority7_module_99__and_module_5_res), .ZN(
        n_majority7_module_99__or_module_7_res) );
  AND2_X1 u_majority7_module_99__and_module_7_U1 ( .A1(
        n_majority7_module_99__or_module_3_res), .A2(
        n_majority7_module_99__or_module_4_res), .ZN(
        n_majority7_module_99__and_module_7_res) );
  OR2_X1 u_majority7_module_99__or_module_8_U1 ( .A1(
        n_majority7_module_99__or_module_4_res), .A2(
        n_majority7_module_99__or_module_3_res), .ZN(
        n_majority7_module_99__or_module_8_res) );
  AND2_X1 u_majority7_module_99__and_module_8_U1 ( .A1(
        n_majority7_module_99__or_module_5_res), .A2(
        n_majority7_module_99__and_module_6_res), .ZN(
        n_majority7_module_99__and_module_8_res) );
  OR2_X1 u_majority7_module_99__or_module_9_U1 ( .A1(
        n_majority7_module_99__and_module_6_res), .A2(
        n_majority7_module_99__or_module_5_res), .ZN(
        n_majority7_module_99__or_module_9_res) );
  OR2_X1 u_majority7_module_99__or_module_10_U1 ( .A1(
        n_majority7_module_99__or_module_7_res), .A2(
        n_majority7_module_99__and_module_7_res), .ZN(
        n_majority7_module_99__or_module_10_res) );
  AND2_X1 u_majority7_module_99__and_module_9_U1 ( .A1(
        n_majority7_module_99__or_module_6_res), .A2(
        n_majority7_module_99__or_module_9_res), .ZN(
        n_majority7_module_99__and_module_9_res) );
  OR2_X1 u_majority7_module_99__or_module_11_U1 ( .A1(
        n_majority7_module_99__or_module_10_res), .A2(
        n_majority7_module_99__and_module_8_res), .ZN(
        n_majority7_module_99__or_module_11_res) );
  AND2_X1 u_majority7_module_99__and_module_10_U1 ( .A1(
        n_majority7_module_99__or_module_8_res), .A2(
        n_majority7_module_99__and_module_9_res), .ZN(
        n_majority7_module_99__and_module_10_res) );
  AND2_X1 u_majority7_module_99__and_module_11_U1 ( .A1(
        n_majority7_module_99__and_module_10_res), .A2(
        n_majority7_module_99__or_module_11_res), .ZN(
        n_majority7_module_99_res) );
  DFF_X1 u_reg_module_100__cini_mul_v000_reg ( .D(n_majority7_module_99_res), 
        .CK(clock_6), .Q(n_reg_module_100_res), .QN() );
  BUF_X1 u_majority7_module_100_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_100_n7) );
  BUF_X1 u_majority7_module_100_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_100_n6) );
  BUF_X1 u_majority7_module_100_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_100_n5) );
  BUF_X1 u_majority7_module_100_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_100_n4) );
  BUF_X1 u_majority7_module_100_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_100_n3) );
  BUF_X1 u_majority7_module_100_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_100_n2) );
  BUF_X1 u_majority7_module_100_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_100_n1) );
  AND2_X1 u_majority7_module_100__and_module_1_U1 ( .A1(
        n_majority7_module_100_n7), .A2(n_majority7_module_100_n1), .ZN(
        n_majority7_module_100__and_module_1_res) );
  OR2_X1 u_majority7_module_100__or_module_1_U1 ( .A1(
        n_majority7_module_100_n1), .A2(n_majority7_module_100_n7), .ZN(
        n_majority7_module_100__or_module_1_res) );
  AND2_X1 u_majority7_module_100__and_module_2_U1 ( .A1(
        n_majority7_module_100_n5), .A2(n_majority7_module_100_n3), .ZN(
        n_majority7_module_100__and_module_2_res) );
  OR2_X1 u_majority7_module_100__or_module_2_U1 ( .A1(
        n_majority7_module_100_n3), .A2(n_majority7_module_100_n5), .ZN(
        n_majority7_module_100__or_module_2_res) );
  AND2_X1 u_majority7_module_100__and_module_3_U1 ( .A1(
        n_majority7_module_100_n6), .A2(n_majority7_module_100_n4), .ZN(
        n_majority7_module_100__and_module_3_res) );
  OR2_X1 u_majority7_module_100__or_module_3_U1 ( .A1(
        n_majority7_module_100_n4), .A2(n_majority7_module_100_n6), .ZN(
        n_majority7_module_100__or_module_3_res) );
  AND2_X1 u_majority7_module_100__and_module_4_U1 ( .A1(
        n_majority7_module_100__and_module_2_res), .A2(
        n_majority7_module_100__and_module_1_res), .ZN(
        n_majority7_module_100__and_module_4_res) );
  OR2_X1 u_majority7_module_100__or_module_4_U1 ( .A1(
        n_majority7_module_100__and_module_1_res), .A2(
        n_majority7_module_100__and_module_2_res), .ZN(
        n_majority7_module_100__or_module_4_res) );
  AND2_X1 u_majority7_module_100__and_module_5_U1 ( .A1(
        n_majority7_module_100__and_module_3_res), .A2(
        n_majority7_module_100_n2), .ZN(
        n_majority7_module_100__and_module_5_res) );
  OR2_X1 u_majority7_module_100__or_module_5_U1 ( .A1(
        n_majority7_module_100_n2), .A2(
        n_majority7_module_100__and_module_3_res), .ZN(
        n_majority7_module_100__or_module_5_res) );
  AND2_X1 u_majority7_module_100__and_module_6_U1 ( .A1(
        n_majority7_module_100__or_module_1_res), .A2(
        n_majority7_module_100__or_module_2_res), .ZN(
        n_majority7_module_100__and_module_6_res) );
  OR2_X1 u_majority7_module_100__or_module_6_U1 ( .A1(
        n_majority7_module_100__or_module_2_res), .A2(
        n_majority7_module_100__or_module_1_res), .ZN(
        n_majority7_module_100__or_module_6_res) );
  OR2_X1 u_majority7_module_100__or_module_7_U1 ( .A1(
        n_majority7_module_100__and_module_4_res), .A2(
        n_majority7_module_100__and_module_5_res), .ZN(
        n_majority7_module_100__or_module_7_res) );
  AND2_X1 u_majority7_module_100__and_module_7_U1 ( .A1(
        n_majority7_module_100__or_module_3_res), .A2(
        n_majority7_module_100__or_module_4_res), .ZN(
        n_majority7_module_100__and_module_7_res) );
  OR2_X1 u_majority7_module_100__or_module_8_U1 ( .A1(
        n_majority7_module_100__or_module_4_res), .A2(
        n_majority7_module_100__or_module_3_res), .ZN(
        n_majority7_module_100__or_module_8_res) );
  AND2_X1 u_majority7_module_100__and_module_8_U1 ( .A1(
        n_majority7_module_100__or_module_5_res), .A2(
        n_majority7_module_100__and_module_6_res), .ZN(
        n_majority7_module_100__and_module_8_res) );
  OR2_X1 u_majority7_module_100__or_module_9_U1 ( .A1(
        n_majority7_module_100__and_module_6_res), .A2(
        n_majority7_module_100__or_module_5_res), .ZN(
        n_majority7_module_100__or_module_9_res) );
  OR2_X1 u_majority7_module_100__or_module_10_U1 ( .A1(
        n_majority7_module_100__or_module_7_res), .A2(
        n_majority7_module_100__and_module_7_res), .ZN(
        n_majority7_module_100__or_module_10_res) );
  AND2_X1 u_majority7_module_100__and_module_9_U1 ( .A1(
        n_majority7_module_100__or_module_6_res), .A2(
        n_majority7_module_100__or_module_9_res), .ZN(
        n_majority7_module_100__and_module_9_res) );
  OR2_X1 u_majority7_module_100__or_module_11_U1 ( .A1(
        n_majority7_module_100__or_module_10_res), .A2(
        n_majority7_module_100__and_module_8_res), .ZN(
        n_majority7_module_100__or_module_11_res) );
  AND2_X1 u_majority7_module_100__and_module_10_U1 ( .A1(
        n_majority7_module_100__or_module_8_res), .A2(
        n_majority7_module_100__and_module_9_res), .ZN(
        n_majority7_module_100__and_module_10_res) );
  AND2_X1 u_majority7_module_100__and_module_11_U1 ( .A1(
        n_majority7_module_100__and_module_10_res), .A2(
        n_majority7_module_100__or_module_11_res), .ZN(
        n_majority7_module_100_res) );
  DFF_X1 u_reg_module_101__cini_mul_v000_reg ( .D(n_majority7_module_100_res), 
        .CK(clock_6), .Q(n_reg_module_101_res), .QN() );
  BUF_X1 u_majority7_module_101_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_101_n7) );
  BUF_X1 u_majority7_module_101_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_101_n6) );
  BUF_X1 u_majority7_module_101_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_101_n5) );
  BUF_X1 u_majority7_module_101_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_101_n4) );
  BUF_X1 u_majority7_module_101_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_101_n3) );
  BUF_X1 u_majority7_module_101_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_101_n2) );
  BUF_X1 u_majority7_module_101_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_101_n1) );
  AND2_X1 u_majority7_module_101__and_module_1_U1 ( .A1(
        n_majority7_module_101_n7), .A2(n_majority7_module_101_n1), .ZN(
        n_majority7_module_101__and_module_1_res) );
  OR2_X1 u_majority7_module_101__or_module_1_U1 ( .A1(
        n_majority7_module_101_n1), .A2(n_majority7_module_101_n7), .ZN(
        n_majority7_module_101__or_module_1_res) );
  AND2_X1 u_majority7_module_101__and_module_2_U1 ( .A1(
        n_majority7_module_101_n5), .A2(n_majority7_module_101_n3), .ZN(
        n_majority7_module_101__and_module_2_res) );
  OR2_X1 u_majority7_module_101__or_module_2_U1 ( .A1(
        n_majority7_module_101_n3), .A2(n_majority7_module_101_n5), .ZN(
        n_majority7_module_101__or_module_2_res) );
  AND2_X1 u_majority7_module_101__and_module_3_U1 ( .A1(
        n_majority7_module_101_n6), .A2(n_majority7_module_101_n4), .ZN(
        n_majority7_module_101__and_module_3_res) );
  OR2_X1 u_majority7_module_101__or_module_3_U1 ( .A1(
        n_majority7_module_101_n4), .A2(n_majority7_module_101_n6), .ZN(
        n_majority7_module_101__or_module_3_res) );
  AND2_X1 u_majority7_module_101__and_module_4_U1 ( .A1(
        n_majority7_module_101__and_module_2_res), .A2(
        n_majority7_module_101__and_module_1_res), .ZN(
        n_majority7_module_101__and_module_4_res) );
  OR2_X1 u_majority7_module_101__or_module_4_U1 ( .A1(
        n_majority7_module_101__and_module_1_res), .A2(
        n_majority7_module_101__and_module_2_res), .ZN(
        n_majority7_module_101__or_module_4_res) );
  AND2_X1 u_majority7_module_101__and_module_5_U1 ( .A1(
        n_majority7_module_101__and_module_3_res), .A2(
        n_majority7_module_101_n2), .ZN(
        n_majority7_module_101__and_module_5_res) );
  OR2_X1 u_majority7_module_101__or_module_5_U1 ( .A1(
        n_majority7_module_101_n2), .A2(
        n_majority7_module_101__and_module_3_res), .ZN(
        n_majority7_module_101__or_module_5_res) );
  AND2_X1 u_majority7_module_101__and_module_6_U1 ( .A1(
        n_majority7_module_101__or_module_1_res), .A2(
        n_majority7_module_101__or_module_2_res), .ZN(
        n_majority7_module_101__and_module_6_res) );
  OR2_X1 u_majority7_module_101__or_module_6_U1 ( .A1(
        n_majority7_module_101__or_module_2_res), .A2(
        n_majority7_module_101__or_module_1_res), .ZN(
        n_majority7_module_101__or_module_6_res) );
  OR2_X1 u_majority7_module_101__or_module_7_U1 ( .A1(
        n_majority7_module_101__and_module_4_res), .A2(
        n_majority7_module_101__and_module_5_res), .ZN(
        n_majority7_module_101__or_module_7_res) );
  AND2_X1 u_majority7_module_101__and_module_7_U1 ( .A1(
        n_majority7_module_101__or_module_3_res), .A2(
        n_majority7_module_101__or_module_4_res), .ZN(
        n_majority7_module_101__and_module_7_res) );
  OR2_X1 u_majority7_module_101__or_module_8_U1 ( .A1(
        n_majority7_module_101__or_module_4_res), .A2(
        n_majority7_module_101__or_module_3_res), .ZN(
        n_majority7_module_101__or_module_8_res) );
  AND2_X1 u_majority7_module_101__and_module_8_U1 ( .A1(
        n_majority7_module_101__or_module_5_res), .A2(
        n_majority7_module_101__and_module_6_res), .ZN(
        n_majority7_module_101__and_module_8_res) );
  OR2_X1 u_majority7_module_101__or_module_9_U1 ( .A1(
        n_majority7_module_101__and_module_6_res), .A2(
        n_majority7_module_101__or_module_5_res), .ZN(
        n_majority7_module_101__or_module_9_res) );
  OR2_X1 u_majority7_module_101__or_module_10_U1 ( .A1(
        n_majority7_module_101__or_module_7_res), .A2(
        n_majority7_module_101__and_module_7_res), .ZN(
        n_majority7_module_101__or_module_10_res) );
  AND2_X1 u_majority7_module_101__and_module_9_U1 ( .A1(
        n_majority7_module_101__or_module_6_res), .A2(
        n_majority7_module_101__or_module_9_res), .ZN(
        n_majority7_module_101__and_module_9_res) );
  OR2_X1 u_majority7_module_101__or_module_11_U1 ( .A1(
        n_majority7_module_101__or_module_10_res), .A2(
        n_majority7_module_101__and_module_8_res), .ZN(
        n_majority7_module_101__or_module_11_res) );
  AND2_X1 u_majority7_module_101__and_module_10_U1 ( .A1(
        n_majority7_module_101__or_module_8_res), .A2(
        n_majority7_module_101__and_module_9_res), .ZN(
        n_majority7_module_101__and_module_10_res) );
  AND2_X1 u_majority7_module_101__and_module_11_U1 ( .A1(
        n_majority7_module_101__and_module_10_res), .A2(
        n_majority7_module_101__or_module_11_res), .ZN(
        n_majority7_module_101_res) );
  DFF_X1 u_reg_module_102__cini_mul_v000_reg ( .D(n_majority7_module_101_res), 
        .CK(clock_6), .Q(n_reg_module_102_res), .QN() );
  BUF_X1 u_majority7_module_102_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_102_n7) );
  BUF_X1 u_majority7_module_102_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_102_n6) );
  BUF_X1 u_majority7_module_102_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_102_n5) );
  BUF_X1 u_majority7_module_102_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_102_n4) );
  BUF_X1 u_majority7_module_102_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_102_n3) );
  BUF_X1 u_majority7_module_102_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_102_n2) );
  BUF_X1 u_majority7_module_102_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_102_n1) );
  AND2_X1 u_majority7_module_102__and_module_1_U1 ( .A1(
        n_majority7_module_102_n7), .A2(n_majority7_module_102_n1), .ZN(
        n_majority7_module_102__and_module_1_res) );
  OR2_X1 u_majority7_module_102__or_module_1_U1 ( .A1(
        n_majority7_module_102_n1), .A2(n_majority7_module_102_n7), .ZN(
        n_majority7_module_102__or_module_1_res) );
  AND2_X1 u_majority7_module_102__and_module_2_U1 ( .A1(
        n_majority7_module_102_n5), .A2(n_majority7_module_102_n3), .ZN(
        n_majority7_module_102__and_module_2_res) );
  OR2_X1 u_majority7_module_102__or_module_2_U1 ( .A1(
        n_majority7_module_102_n3), .A2(n_majority7_module_102_n5), .ZN(
        n_majority7_module_102__or_module_2_res) );
  AND2_X1 u_majority7_module_102__and_module_3_U1 ( .A1(
        n_majority7_module_102_n6), .A2(n_majority7_module_102_n4), .ZN(
        n_majority7_module_102__and_module_3_res) );
  OR2_X1 u_majority7_module_102__or_module_3_U1 ( .A1(
        n_majority7_module_102_n4), .A2(n_majority7_module_102_n6), .ZN(
        n_majority7_module_102__or_module_3_res) );
  AND2_X1 u_majority7_module_102__and_module_4_U1 ( .A1(
        n_majority7_module_102__and_module_2_res), .A2(
        n_majority7_module_102__and_module_1_res), .ZN(
        n_majority7_module_102__and_module_4_res) );
  OR2_X1 u_majority7_module_102__or_module_4_U1 ( .A1(
        n_majority7_module_102__and_module_1_res), .A2(
        n_majority7_module_102__and_module_2_res), .ZN(
        n_majority7_module_102__or_module_4_res) );
  AND2_X1 u_majority7_module_102__and_module_5_U1 ( .A1(
        n_majority7_module_102__and_module_3_res), .A2(
        n_majority7_module_102_n2), .ZN(
        n_majority7_module_102__and_module_5_res) );
  OR2_X1 u_majority7_module_102__or_module_5_U1 ( .A1(
        n_majority7_module_102_n2), .A2(
        n_majority7_module_102__and_module_3_res), .ZN(
        n_majority7_module_102__or_module_5_res) );
  AND2_X1 u_majority7_module_102__and_module_6_U1 ( .A1(
        n_majority7_module_102__or_module_1_res), .A2(
        n_majority7_module_102__or_module_2_res), .ZN(
        n_majority7_module_102__and_module_6_res) );
  OR2_X1 u_majority7_module_102__or_module_6_U1 ( .A1(
        n_majority7_module_102__or_module_2_res), .A2(
        n_majority7_module_102__or_module_1_res), .ZN(
        n_majority7_module_102__or_module_6_res) );
  OR2_X1 u_majority7_module_102__or_module_7_U1 ( .A1(
        n_majority7_module_102__and_module_4_res), .A2(
        n_majority7_module_102__and_module_5_res), .ZN(
        n_majority7_module_102__or_module_7_res) );
  AND2_X1 u_majority7_module_102__and_module_7_U1 ( .A1(
        n_majority7_module_102__or_module_3_res), .A2(
        n_majority7_module_102__or_module_4_res), .ZN(
        n_majority7_module_102__and_module_7_res) );
  OR2_X1 u_majority7_module_102__or_module_8_U1 ( .A1(
        n_majority7_module_102__or_module_4_res), .A2(
        n_majority7_module_102__or_module_3_res), .ZN(
        n_majority7_module_102__or_module_8_res) );
  AND2_X1 u_majority7_module_102__and_module_8_U1 ( .A1(
        n_majority7_module_102__or_module_5_res), .A2(
        n_majority7_module_102__and_module_6_res), .ZN(
        n_majority7_module_102__and_module_8_res) );
  OR2_X1 u_majority7_module_102__or_module_9_U1 ( .A1(
        n_majority7_module_102__and_module_6_res), .A2(
        n_majority7_module_102__or_module_5_res), .ZN(
        n_majority7_module_102__or_module_9_res) );
  OR2_X1 u_majority7_module_102__or_module_10_U1 ( .A1(
        n_majority7_module_102__or_module_7_res), .A2(
        n_majority7_module_102__and_module_7_res), .ZN(
        n_majority7_module_102__or_module_10_res) );
  AND2_X1 u_majority7_module_102__and_module_9_U1 ( .A1(
        n_majority7_module_102__or_module_6_res), .A2(
        n_majority7_module_102__or_module_9_res), .ZN(
        n_majority7_module_102__and_module_9_res) );
  OR2_X1 u_majority7_module_102__or_module_11_U1 ( .A1(
        n_majority7_module_102__or_module_10_res), .A2(
        n_majority7_module_102__and_module_8_res), .ZN(
        n_majority7_module_102__or_module_11_res) );
  AND2_X1 u_majority7_module_102__and_module_10_U1 ( .A1(
        n_majority7_module_102__or_module_8_res), .A2(
        n_majority7_module_102__and_module_9_res), .ZN(
        n_majority7_module_102__and_module_10_res) );
  AND2_X1 u_majority7_module_102__and_module_11_U1 ( .A1(
        n_majority7_module_102__and_module_10_res), .A2(
        n_majority7_module_102__or_module_11_res), .ZN(
        n_majority7_module_102_res) );
  DFF_X1 u_reg_module_103__cini_mul_v000_reg ( .D(n_majority7_module_102_res), 
        .CK(clock_6), .Q(n_reg_module_103_res), .QN() );
  BUF_X1 u_majority7_module_103_U7 ( .A(n_xor_module_78_res), .Z(
        n_majority7_module_103_n7) );
  BUF_X1 u_majority7_module_103_U6 ( .A(n_xor_module_66_res), .Z(
        n_majority7_module_103_n6) );
  BUF_X1 u_majority7_module_103_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_103_n5) );
  BUF_X1 u_majority7_module_103_U4 ( .A(n_xor_module_54_res), .Z(
        n_majority7_module_103_n4) );
  BUF_X1 u_majority7_module_103_U3 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_103_n3) );
  BUF_X1 u_majority7_module_103_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_103_n2) );
  BUF_X1 u_majority7_module_103_U1 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_103_n1) );
  AND2_X1 u_majority7_module_103__and_module_1_U1 ( .A1(
        n_majority7_module_103_n7), .A2(n_majority7_module_103_n1), .ZN(
        n_majority7_module_103__and_module_1_res) );
  OR2_X1 u_majority7_module_103__or_module_1_U1 ( .A1(
        n_majority7_module_103_n1), .A2(n_majority7_module_103_n7), .ZN(
        n_majority7_module_103__or_module_1_res) );
  AND2_X1 u_majority7_module_103__and_module_2_U1 ( .A1(
        n_majority7_module_103_n5), .A2(n_majority7_module_103_n3), .ZN(
        n_majority7_module_103__and_module_2_res) );
  OR2_X1 u_majority7_module_103__or_module_2_U1 ( .A1(
        n_majority7_module_103_n3), .A2(n_majority7_module_103_n5), .ZN(
        n_majority7_module_103__or_module_2_res) );
  AND2_X1 u_majority7_module_103__and_module_3_U1 ( .A1(
        n_majority7_module_103_n6), .A2(n_majority7_module_103_n4), .ZN(
        n_majority7_module_103__and_module_3_res) );
  OR2_X1 u_majority7_module_103__or_module_3_U1 ( .A1(
        n_majority7_module_103_n4), .A2(n_majority7_module_103_n6), .ZN(
        n_majority7_module_103__or_module_3_res) );
  AND2_X1 u_majority7_module_103__and_module_4_U1 ( .A1(
        n_majority7_module_103__and_module_2_res), .A2(
        n_majority7_module_103__and_module_1_res), .ZN(
        n_majority7_module_103__and_module_4_res) );
  OR2_X1 u_majority7_module_103__or_module_4_U1 ( .A1(
        n_majority7_module_103__and_module_1_res), .A2(
        n_majority7_module_103__and_module_2_res), .ZN(
        n_majority7_module_103__or_module_4_res) );
  AND2_X1 u_majority7_module_103__and_module_5_U1 ( .A1(
        n_majority7_module_103__and_module_3_res), .A2(
        n_majority7_module_103_n2), .ZN(
        n_majority7_module_103__and_module_5_res) );
  OR2_X1 u_majority7_module_103__or_module_5_U1 ( .A1(
        n_majority7_module_103_n2), .A2(
        n_majority7_module_103__and_module_3_res), .ZN(
        n_majority7_module_103__or_module_5_res) );
  AND2_X1 u_majority7_module_103__and_module_6_U1 ( .A1(
        n_majority7_module_103__or_module_1_res), .A2(
        n_majority7_module_103__or_module_2_res), .ZN(
        n_majority7_module_103__and_module_6_res) );
  OR2_X1 u_majority7_module_103__or_module_6_U1 ( .A1(
        n_majority7_module_103__or_module_2_res), .A2(
        n_majority7_module_103__or_module_1_res), .ZN(
        n_majority7_module_103__or_module_6_res) );
  OR2_X1 u_majority7_module_103__or_module_7_U1 ( .A1(
        n_majority7_module_103__and_module_4_res), .A2(
        n_majority7_module_103__and_module_5_res), .ZN(
        n_majority7_module_103__or_module_7_res) );
  AND2_X1 u_majority7_module_103__and_module_7_U1 ( .A1(
        n_majority7_module_103__or_module_3_res), .A2(
        n_majority7_module_103__or_module_4_res), .ZN(
        n_majority7_module_103__and_module_7_res) );
  OR2_X1 u_majority7_module_103__or_module_8_U1 ( .A1(
        n_majority7_module_103__or_module_4_res), .A2(
        n_majority7_module_103__or_module_3_res), .ZN(
        n_majority7_module_103__or_module_8_res) );
  AND2_X1 u_majority7_module_103__and_module_8_U1 ( .A1(
        n_majority7_module_103__or_module_5_res), .A2(
        n_majority7_module_103__and_module_6_res), .ZN(
        n_majority7_module_103__and_module_8_res) );
  OR2_X1 u_majority7_module_103__or_module_9_U1 ( .A1(
        n_majority7_module_103__and_module_6_res), .A2(
        n_majority7_module_103__or_module_5_res), .ZN(
        n_majority7_module_103__or_module_9_res) );
  OR2_X1 u_majority7_module_103__or_module_10_U1 ( .A1(
        n_majority7_module_103__or_module_7_res), .A2(
        n_majority7_module_103__and_module_7_res), .ZN(
        n_majority7_module_103__or_module_10_res) );
  AND2_X1 u_majority7_module_103__and_module_9_U1 ( .A1(
        n_majority7_module_103__or_module_6_res), .A2(
        n_majority7_module_103__or_module_9_res), .ZN(
        n_majority7_module_103__and_module_9_res) );
  OR2_X1 u_majority7_module_103__or_module_11_U1 ( .A1(
        n_majority7_module_103__or_module_10_res), .A2(
        n_majority7_module_103__and_module_8_res), .ZN(
        n_majority7_module_103__or_module_11_res) );
  AND2_X1 u_majority7_module_103__and_module_10_U1 ( .A1(
        n_majority7_module_103__or_module_8_res), .A2(
        n_majority7_module_103__and_module_9_res), .ZN(
        n_majority7_module_103__and_module_10_res) );
  AND2_X1 u_majority7_module_103__and_module_11_U1 ( .A1(
        n_majority7_module_103__and_module_10_res), .A2(
        n_majority7_module_103__or_module_11_res), .ZN(
        n_majority7_module_103_res) );
  DFF_X1 u_reg_module_104__cini_mul_v000_reg ( .D(n_majority7_module_103_res), 
        .CK(clock_6), .Q(n_reg_module_104_res), .QN() );
  BUF_X1 u_majority7_module_104_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_104_n7) );
  BUF_X1 u_majority7_module_104_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_104_n6) );
  BUF_X1 u_majority7_module_104_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_104_n5) );
  BUF_X1 u_majority7_module_104_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_104_n4) );
  BUF_X1 u_majority7_module_104_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_104_n3) );
  BUF_X1 u_majority7_module_104_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_104_n2) );
  BUF_X1 u_majority7_module_104_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_104_n1) );
  AND2_X1 u_majority7_module_104__and_module_1_U1 ( .A1(
        n_majority7_module_104_n7), .A2(n_majority7_module_104_n1), .ZN(
        n_majority7_module_104__and_module_1_res) );
  OR2_X1 u_majority7_module_104__or_module_1_U1 ( .A1(
        n_majority7_module_104_n1), .A2(n_majority7_module_104_n7), .ZN(
        n_majority7_module_104__or_module_1_res) );
  AND2_X1 u_majority7_module_104__and_module_2_U1 ( .A1(
        n_majority7_module_104_n5), .A2(n_majority7_module_104_n3), .ZN(
        n_majority7_module_104__and_module_2_res) );
  OR2_X1 u_majority7_module_104__or_module_2_U1 ( .A1(
        n_majority7_module_104_n3), .A2(n_majority7_module_104_n5), .ZN(
        n_majority7_module_104__or_module_2_res) );
  AND2_X1 u_majority7_module_104__and_module_3_U1 ( .A1(
        n_majority7_module_104_n6), .A2(n_majority7_module_104_n4), .ZN(
        n_majority7_module_104__and_module_3_res) );
  OR2_X1 u_majority7_module_104__or_module_3_U1 ( .A1(
        n_majority7_module_104_n4), .A2(n_majority7_module_104_n6), .ZN(
        n_majority7_module_104__or_module_3_res) );
  AND2_X1 u_majority7_module_104__and_module_4_U1 ( .A1(
        n_majority7_module_104__and_module_2_res), .A2(
        n_majority7_module_104__and_module_1_res), .ZN(
        n_majority7_module_104__and_module_4_res) );
  OR2_X1 u_majority7_module_104__or_module_4_U1 ( .A1(
        n_majority7_module_104__and_module_1_res), .A2(
        n_majority7_module_104__and_module_2_res), .ZN(
        n_majority7_module_104__or_module_4_res) );
  AND2_X1 u_majority7_module_104__and_module_5_U1 ( .A1(
        n_majority7_module_104__and_module_3_res), .A2(
        n_majority7_module_104_n2), .ZN(
        n_majority7_module_104__and_module_5_res) );
  OR2_X1 u_majority7_module_104__or_module_5_U1 ( .A1(
        n_majority7_module_104_n2), .A2(
        n_majority7_module_104__and_module_3_res), .ZN(
        n_majority7_module_104__or_module_5_res) );
  AND2_X1 u_majority7_module_104__and_module_6_U1 ( .A1(
        n_majority7_module_104__or_module_1_res), .A2(
        n_majority7_module_104__or_module_2_res), .ZN(
        n_majority7_module_104__and_module_6_res) );
  OR2_X1 u_majority7_module_104__or_module_6_U1 ( .A1(
        n_majority7_module_104__or_module_2_res), .A2(
        n_majority7_module_104__or_module_1_res), .ZN(
        n_majority7_module_104__or_module_6_res) );
  OR2_X1 u_majority7_module_104__or_module_7_U1 ( .A1(
        n_majority7_module_104__and_module_4_res), .A2(
        n_majority7_module_104__and_module_5_res), .ZN(
        n_majority7_module_104__or_module_7_res) );
  AND2_X1 u_majority7_module_104__and_module_7_U1 ( .A1(
        n_majority7_module_104__or_module_3_res), .A2(
        n_majority7_module_104__or_module_4_res), .ZN(
        n_majority7_module_104__and_module_7_res) );
  OR2_X1 u_majority7_module_104__or_module_8_U1 ( .A1(
        n_majority7_module_104__or_module_4_res), .A2(
        n_majority7_module_104__or_module_3_res), .ZN(
        n_majority7_module_104__or_module_8_res) );
  AND2_X1 u_majority7_module_104__and_module_8_U1 ( .A1(
        n_majority7_module_104__or_module_5_res), .A2(
        n_majority7_module_104__and_module_6_res), .ZN(
        n_majority7_module_104__and_module_8_res) );
  OR2_X1 u_majority7_module_104__or_module_9_U1 ( .A1(
        n_majority7_module_104__and_module_6_res), .A2(
        n_majority7_module_104__or_module_5_res), .ZN(
        n_majority7_module_104__or_module_9_res) );
  OR2_X1 u_majority7_module_104__or_module_10_U1 ( .A1(
        n_majority7_module_104__or_module_7_res), .A2(
        n_majority7_module_104__and_module_7_res), .ZN(
        n_majority7_module_104__or_module_10_res) );
  AND2_X1 u_majority7_module_104__and_module_9_U1 ( .A1(
        n_majority7_module_104__or_module_6_res), .A2(
        n_majority7_module_104__or_module_9_res), .ZN(
        n_majority7_module_104__and_module_9_res) );
  OR2_X1 u_majority7_module_104__or_module_11_U1 ( .A1(
        n_majority7_module_104__or_module_10_res), .A2(
        n_majority7_module_104__and_module_8_res), .ZN(
        n_majority7_module_104__or_module_11_res) );
  AND2_X1 u_majority7_module_104__and_module_10_U1 ( .A1(
        n_majority7_module_104__or_module_8_res), .A2(
        n_majority7_module_104__and_module_9_res), .ZN(
        n_majority7_module_104__and_module_10_res) );
  AND2_X1 u_majority7_module_104__and_module_11_U1 ( .A1(
        n_majority7_module_104__and_module_10_res), .A2(
        n_majority7_module_104__or_module_11_res), .ZN(
        n_majority7_module_104_res) );
  DFF_X1 u_reg_module_105__cini_mul_v000_reg ( .D(n_majority7_module_104_res), 
        .CK(clock_6), .Q(n_reg_module_105_res), .QN() );
  BUF_X1 u_majority7_module_105_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_105_n7) );
  BUF_X1 u_majority7_module_105_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_105_n6) );
  BUF_X1 u_majority7_module_105_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_105_n5) );
  BUF_X1 u_majority7_module_105_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_105_n4) );
  BUF_X1 u_majority7_module_105_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_105_n3) );
  BUF_X1 u_majority7_module_105_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_105_n2) );
  BUF_X1 u_majority7_module_105_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_105_n1) );
  AND2_X1 u_majority7_module_105__and_module_1_U1 ( .A1(
        n_majority7_module_105_n7), .A2(n_majority7_module_105_n1), .ZN(
        n_majority7_module_105__and_module_1_res) );
  OR2_X1 u_majority7_module_105__or_module_1_U1 ( .A1(
        n_majority7_module_105_n1), .A2(n_majority7_module_105_n7), .ZN(
        n_majority7_module_105__or_module_1_res) );
  AND2_X1 u_majority7_module_105__and_module_2_U1 ( .A1(
        n_majority7_module_105_n5), .A2(n_majority7_module_105_n3), .ZN(
        n_majority7_module_105__and_module_2_res) );
  OR2_X1 u_majority7_module_105__or_module_2_U1 ( .A1(
        n_majority7_module_105_n3), .A2(n_majority7_module_105_n5), .ZN(
        n_majority7_module_105__or_module_2_res) );
  AND2_X1 u_majority7_module_105__and_module_3_U1 ( .A1(
        n_majority7_module_105_n6), .A2(n_majority7_module_105_n4), .ZN(
        n_majority7_module_105__and_module_3_res) );
  OR2_X1 u_majority7_module_105__or_module_3_U1 ( .A1(
        n_majority7_module_105_n4), .A2(n_majority7_module_105_n6), .ZN(
        n_majority7_module_105__or_module_3_res) );
  AND2_X1 u_majority7_module_105__and_module_4_U1 ( .A1(
        n_majority7_module_105__and_module_2_res), .A2(
        n_majority7_module_105__and_module_1_res), .ZN(
        n_majority7_module_105__and_module_4_res) );
  OR2_X1 u_majority7_module_105__or_module_4_U1 ( .A1(
        n_majority7_module_105__and_module_1_res), .A2(
        n_majority7_module_105__and_module_2_res), .ZN(
        n_majority7_module_105__or_module_4_res) );
  AND2_X1 u_majority7_module_105__and_module_5_U1 ( .A1(
        n_majority7_module_105__and_module_3_res), .A2(
        n_majority7_module_105_n2), .ZN(
        n_majority7_module_105__and_module_5_res) );
  OR2_X1 u_majority7_module_105__or_module_5_U1 ( .A1(
        n_majority7_module_105_n2), .A2(
        n_majority7_module_105__and_module_3_res), .ZN(
        n_majority7_module_105__or_module_5_res) );
  AND2_X1 u_majority7_module_105__and_module_6_U1 ( .A1(
        n_majority7_module_105__or_module_1_res), .A2(
        n_majority7_module_105__or_module_2_res), .ZN(
        n_majority7_module_105__and_module_6_res) );
  OR2_X1 u_majority7_module_105__or_module_6_U1 ( .A1(
        n_majority7_module_105__or_module_2_res), .A2(
        n_majority7_module_105__or_module_1_res), .ZN(
        n_majority7_module_105__or_module_6_res) );
  OR2_X1 u_majority7_module_105__or_module_7_U1 ( .A1(
        n_majority7_module_105__and_module_4_res), .A2(
        n_majority7_module_105__and_module_5_res), .ZN(
        n_majority7_module_105__or_module_7_res) );
  AND2_X1 u_majority7_module_105__and_module_7_U1 ( .A1(
        n_majority7_module_105__or_module_3_res), .A2(
        n_majority7_module_105__or_module_4_res), .ZN(
        n_majority7_module_105__and_module_7_res) );
  OR2_X1 u_majority7_module_105__or_module_8_U1 ( .A1(
        n_majority7_module_105__or_module_4_res), .A2(
        n_majority7_module_105__or_module_3_res), .ZN(
        n_majority7_module_105__or_module_8_res) );
  AND2_X1 u_majority7_module_105__and_module_8_U1 ( .A1(
        n_majority7_module_105__or_module_5_res), .A2(
        n_majority7_module_105__and_module_6_res), .ZN(
        n_majority7_module_105__and_module_8_res) );
  OR2_X1 u_majority7_module_105__or_module_9_U1 ( .A1(
        n_majority7_module_105__and_module_6_res), .A2(
        n_majority7_module_105__or_module_5_res), .ZN(
        n_majority7_module_105__or_module_9_res) );
  OR2_X1 u_majority7_module_105__or_module_10_U1 ( .A1(
        n_majority7_module_105__or_module_7_res), .A2(
        n_majority7_module_105__and_module_7_res), .ZN(
        n_majority7_module_105__or_module_10_res) );
  AND2_X1 u_majority7_module_105__and_module_9_U1 ( .A1(
        n_majority7_module_105__or_module_6_res), .A2(
        n_majority7_module_105__or_module_9_res), .ZN(
        n_majority7_module_105__and_module_9_res) );
  OR2_X1 u_majority7_module_105__or_module_11_U1 ( .A1(
        n_majority7_module_105__or_module_10_res), .A2(
        n_majority7_module_105__and_module_8_res), .ZN(
        n_majority7_module_105__or_module_11_res) );
  AND2_X1 u_majority7_module_105__and_module_10_U1 ( .A1(
        n_majority7_module_105__or_module_8_res), .A2(
        n_majority7_module_105__and_module_9_res), .ZN(
        n_majority7_module_105__and_module_10_res) );
  AND2_X1 u_majority7_module_105__and_module_11_U1 ( .A1(
        n_majority7_module_105__and_module_10_res), .A2(
        n_majority7_module_105__or_module_11_res), .ZN(
        n_majority7_module_105_res) );
  DFF_X1 u_reg_module_106__cini_mul_v000_reg ( .D(n_majority7_module_105_res), 
        .CK(clock_6), .Q(n_reg_module_106_res), .QN() );
  BUF_X1 u_majority7_module_106_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_106_n7) );
  BUF_X1 u_majority7_module_106_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_106_n6) );
  BUF_X1 u_majority7_module_106_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_106_n5) );
  BUF_X1 u_majority7_module_106_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_106_n4) );
  BUF_X1 u_majority7_module_106_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_106_n3) );
  BUF_X1 u_majority7_module_106_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_106_n2) );
  BUF_X1 u_majority7_module_106_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_106_n1) );
  AND2_X1 u_majority7_module_106__and_module_1_U1 ( .A1(
        n_majority7_module_106_n7), .A2(n_majority7_module_106_n1), .ZN(
        n_majority7_module_106__and_module_1_res) );
  OR2_X1 u_majority7_module_106__or_module_1_U1 ( .A1(
        n_majority7_module_106_n1), .A2(n_majority7_module_106_n7), .ZN(
        n_majority7_module_106__or_module_1_res) );
  AND2_X1 u_majority7_module_106__and_module_2_U1 ( .A1(
        n_majority7_module_106_n5), .A2(n_majority7_module_106_n3), .ZN(
        n_majority7_module_106__and_module_2_res) );
  OR2_X1 u_majority7_module_106__or_module_2_U1 ( .A1(
        n_majority7_module_106_n3), .A2(n_majority7_module_106_n5), .ZN(
        n_majority7_module_106__or_module_2_res) );
  AND2_X1 u_majority7_module_106__and_module_3_U1 ( .A1(
        n_majority7_module_106_n6), .A2(n_majority7_module_106_n4), .ZN(
        n_majority7_module_106__and_module_3_res) );
  OR2_X1 u_majority7_module_106__or_module_3_U1 ( .A1(
        n_majority7_module_106_n4), .A2(n_majority7_module_106_n6), .ZN(
        n_majority7_module_106__or_module_3_res) );
  AND2_X1 u_majority7_module_106__and_module_4_U1 ( .A1(
        n_majority7_module_106__and_module_2_res), .A2(
        n_majority7_module_106__and_module_1_res), .ZN(
        n_majority7_module_106__and_module_4_res) );
  OR2_X1 u_majority7_module_106__or_module_4_U1 ( .A1(
        n_majority7_module_106__and_module_1_res), .A2(
        n_majority7_module_106__and_module_2_res), .ZN(
        n_majority7_module_106__or_module_4_res) );
  AND2_X1 u_majority7_module_106__and_module_5_U1 ( .A1(
        n_majority7_module_106__and_module_3_res), .A2(
        n_majority7_module_106_n2), .ZN(
        n_majority7_module_106__and_module_5_res) );
  OR2_X1 u_majority7_module_106__or_module_5_U1 ( .A1(
        n_majority7_module_106_n2), .A2(
        n_majority7_module_106__and_module_3_res), .ZN(
        n_majority7_module_106__or_module_5_res) );
  AND2_X1 u_majority7_module_106__and_module_6_U1 ( .A1(
        n_majority7_module_106__or_module_1_res), .A2(
        n_majority7_module_106__or_module_2_res), .ZN(
        n_majority7_module_106__and_module_6_res) );
  OR2_X1 u_majority7_module_106__or_module_6_U1 ( .A1(
        n_majority7_module_106__or_module_2_res), .A2(
        n_majority7_module_106__or_module_1_res), .ZN(
        n_majority7_module_106__or_module_6_res) );
  OR2_X1 u_majority7_module_106__or_module_7_U1 ( .A1(
        n_majority7_module_106__and_module_4_res), .A2(
        n_majority7_module_106__and_module_5_res), .ZN(
        n_majority7_module_106__or_module_7_res) );
  AND2_X1 u_majority7_module_106__and_module_7_U1 ( .A1(
        n_majority7_module_106__or_module_3_res), .A2(
        n_majority7_module_106__or_module_4_res), .ZN(
        n_majority7_module_106__and_module_7_res) );
  OR2_X1 u_majority7_module_106__or_module_8_U1 ( .A1(
        n_majority7_module_106__or_module_4_res), .A2(
        n_majority7_module_106__or_module_3_res), .ZN(
        n_majority7_module_106__or_module_8_res) );
  AND2_X1 u_majority7_module_106__and_module_8_U1 ( .A1(
        n_majority7_module_106__or_module_5_res), .A2(
        n_majority7_module_106__and_module_6_res), .ZN(
        n_majority7_module_106__and_module_8_res) );
  OR2_X1 u_majority7_module_106__or_module_9_U1 ( .A1(
        n_majority7_module_106__and_module_6_res), .A2(
        n_majority7_module_106__or_module_5_res), .ZN(
        n_majority7_module_106__or_module_9_res) );
  OR2_X1 u_majority7_module_106__or_module_10_U1 ( .A1(
        n_majority7_module_106__or_module_7_res), .A2(
        n_majority7_module_106__and_module_7_res), .ZN(
        n_majority7_module_106__or_module_10_res) );
  AND2_X1 u_majority7_module_106__and_module_9_U1 ( .A1(
        n_majority7_module_106__or_module_6_res), .A2(
        n_majority7_module_106__or_module_9_res), .ZN(
        n_majority7_module_106__and_module_9_res) );
  OR2_X1 u_majority7_module_106__or_module_11_U1 ( .A1(
        n_majority7_module_106__or_module_10_res), .A2(
        n_majority7_module_106__and_module_8_res), .ZN(
        n_majority7_module_106__or_module_11_res) );
  AND2_X1 u_majority7_module_106__and_module_10_U1 ( .A1(
        n_majority7_module_106__or_module_8_res), .A2(
        n_majority7_module_106__and_module_9_res), .ZN(
        n_majority7_module_106__and_module_10_res) );
  AND2_X1 u_majority7_module_106__and_module_11_U1 ( .A1(
        n_majority7_module_106__and_module_10_res), .A2(
        n_majority7_module_106__or_module_11_res), .ZN(
        n_majority7_module_106_res) );
  DFF_X1 u_reg_module_107__cini_mul_v000_reg ( .D(n_majority7_module_106_res), 
        .CK(clock_6), .Q(n_reg_module_107_res), .QN() );
  BUF_X1 u_majority7_module_107_U7 ( .A(n_xor_module_81_res), .Z(
        n_majority7_module_107_n7) );
  BUF_X1 u_majority7_module_107_U6 ( .A(n_xor_module_69_res), .Z(
        n_majority7_module_107_n6) );
  BUF_X1 u_majority7_module_107_U5 ( .A(n_xor_module_45_res), .Z(
        n_majority7_module_107_n5) );
  BUF_X1 u_majority7_module_107_U4 ( .A(n_xor_module_57_res), .Z(
        n_majority7_module_107_n4) );
  BUF_X1 u_majority7_module_107_U3 ( .A(n_xor_module_33_res), .Z(
        n_majority7_module_107_n3) );
  BUF_X1 u_majority7_module_107_U2 ( .A(n_xor_module_21_res), .Z(
        n_majority7_module_107_n2) );
  BUF_X1 u_majority7_module_107_U1 ( .A(n_xor_module_9_res), .Z(
        n_majority7_module_107_n1) );
  AND2_X1 u_majority7_module_107__and_module_1_U1 ( .A1(
        n_majority7_module_107_n7), .A2(n_majority7_module_107_n1), .ZN(
        n_majority7_module_107__and_module_1_res) );
  OR2_X1 u_majority7_module_107__or_module_1_U1 ( .A1(
        n_majority7_module_107_n1), .A2(n_majority7_module_107_n7), .ZN(
        n_majority7_module_107__or_module_1_res) );
  AND2_X1 u_majority7_module_107__and_module_2_U1 ( .A1(
        n_majority7_module_107_n5), .A2(n_majority7_module_107_n3), .ZN(
        n_majority7_module_107__and_module_2_res) );
  OR2_X1 u_majority7_module_107__or_module_2_U1 ( .A1(
        n_majority7_module_107_n3), .A2(n_majority7_module_107_n5), .ZN(
        n_majority7_module_107__or_module_2_res) );
  AND2_X1 u_majority7_module_107__and_module_3_U1 ( .A1(
        n_majority7_module_107_n6), .A2(n_majority7_module_107_n4), .ZN(
        n_majority7_module_107__and_module_3_res) );
  OR2_X1 u_majority7_module_107__or_module_3_U1 ( .A1(
        n_majority7_module_107_n4), .A2(n_majority7_module_107_n6), .ZN(
        n_majority7_module_107__or_module_3_res) );
  AND2_X1 u_majority7_module_107__and_module_4_U1 ( .A1(
        n_majority7_module_107__and_module_2_res), .A2(
        n_majority7_module_107__and_module_1_res), .ZN(
        n_majority7_module_107__and_module_4_res) );
  OR2_X1 u_majority7_module_107__or_module_4_U1 ( .A1(
        n_majority7_module_107__and_module_1_res), .A2(
        n_majority7_module_107__and_module_2_res), .ZN(
        n_majority7_module_107__or_module_4_res) );
  AND2_X1 u_majority7_module_107__and_module_5_U1 ( .A1(
        n_majority7_module_107__and_module_3_res), .A2(
        n_majority7_module_107_n2), .ZN(
        n_majority7_module_107__and_module_5_res) );
  OR2_X1 u_majority7_module_107__or_module_5_U1 ( .A1(
        n_majority7_module_107_n2), .A2(
        n_majority7_module_107__and_module_3_res), .ZN(
        n_majority7_module_107__or_module_5_res) );
  AND2_X1 u_majority7_module_107__and_module_6_U1 ( .A1(
        n_majority7_module_107__or_module_1_res), .A2(
        n_majority7_module_107__or_module_2_res), .ZN(
        n_majority7_module_107__and_module_6_res) );
  OR2_X1 u_majority7_module_107__or_module_6_U1 ( .A1(
        n_majority7_module_107__or_module_2_res), .A2(
        n_majority7_module_107__or_module_1_res), .ZN(
        n_majority7_module_107__or_module_6_res) );
  OR2_X1 u_majority7_module_107__or_module_7_U1 ( .A1(
        n_majority7_module_107__and_module_4_res), .A2(
        n_majority7_module_107__and_module_5_res), .ZN(
        n_majority7_module_107__or_module_7_res) );
  AND2_X1 u_majority7_module_107__and_module_7_U1 ( .A1(
        n_majority7_module_107__or_module_3_res), .A2(
        n_majority7_module_107__or_module_4_res), .ZN(
        n_majority7_module_107__and_module_7_res) );
  OR2_X1 u_majority7_module_107__or_module_8_U1 ( .A1(
        n_majority7_module_107__or_module_4_res), .A2(
        n_majority7_module_107__or_module_3_res), .ZN(
        n_majority7_module_107__or_module_8_res) );
  AND2_X1 u_majority7_module_107__and_module_8_U1 ( .A1(
        n_majority7_module_107__or_module_5_res), .A2(
        n_majority7_module_107__and_module_6_res), .ZN(
        n_majority7_module_107__and_module_8_res) );
  OR2_X1 u_majority7_module_107__or_module_9_U1 ( .A1(
        n_majority7_module_107__and_module_6_res), .A2(
        n_majority7_module_107__or_module_5_res), .ZN(
        n_majority7_module_107__or_module_9_res) );
  OR2_X1 u_majority7_module_107__or_module_10_U1 ( .A1(
        n_majority7_module_107__or_module_7_res), .A2(
        n_majority7_module_107__and_module_7_res), .ZN(
        n_majority7_module_107__or_module_10_res) );
  AND2_X1 u_majority7_module_107__and_module_9_U1 ( .A1(
        n_majority7_module_107__or_module_6_res), .A2(
        n_majority7_module_107__or_module_9_res), .ZN(
        n_majority7_module_107__and_module_9_res) );
  OR2_X1 u_majority7_module_107__or_module_11_U1 ( .A1(
        n_majority7_module_107__or_module_10_res), .A2(
        n_majority7_module_107__and_module_8_res), .ZN(
        n_majority7_module_107__or_module_11_res) );
  AND2_X1 u_majority7_module_107__and_module_10_U1 ( .A1(
        n_majority7_module_107__or_module_8_res), .A2(
        n_majority7_module_107__and_module_9_res), .ZN(
        n_majority7_module_107__and_module_10_res) );
  AND2_X1 u_majority7_module_107__and_module_11_U1 ( .A1(
        n_majority7_module_107__and_module_10_res), .A2(
        n_majority7_module_107__or_module_11_res), .ZN(
        n_majority7_module_107_res) );
  DFF_X1 u_reg_module_108__cini_mul_v000_reg ( .D(n_majority7_module_107_res), 
        .CK(clock_6), .Q(n_reg_module_108_res), .QN() );
  BUF_X1 u_majority7_module_108_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_108_n7) );
  BUF_X1 u_majority7_module_108_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_108_n6) );
  BUF_X1 u_majority7_module_108_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_108_n5) );
  BUF_X1 u_majority7_module_108_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_108_n4) );
  BUF_X1 u_majority7_module_108_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_108_n3) );
  BUF_X1 u_majority7_module_108_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_108_n2) );
  BUF_X1 u_majority7_module_108_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_108_n1) );
  AND2_X1 u_majority7_module_108__and_module_1_U1 ( .A1(
        n_majority7_module_108_n7), .A2(n_majority7_module_108_n1), .ZN(
        n_majority7_module_108__and_module_1_res) );
  OR2_X1 u_majority7_module_108__or_module_1_U1 ( .A1(
        n_majority7_module_108_n1), .A2(n_majority7_module_108_n7), .ZN(
        n_majority7_module_108__or_module_1_res) );
  AND2_X1 u_majority7_module_108__and_module_2_U1 ( .A1(
        n_majority7_module_108_n5), .A2(n_majority7_module_108_n3), .ZN(
        n_majority7_module_108__and_module_2_res) );
  OR2_X1 u_majority7_module_108__or_module_2_U1 ( .A1(
        n_majority7_module_108_n3), .A2(n_majority7_module_108_n5), .ZN(
        n_majority7_module_108__or_module_2_res) );
  AND2_X1 u_majority7_module_108__and_module_3_U1 ( .A1(
        n_majority7_module_108_n6), .A2(n_majority7_module_108_n4), .ZN(
        n_majority7_module_108__and_module_3_res) );
  OR2_X1 u_majority7_module_108__or_module_3_U1 ( .A1(
        n_majority7_module_108_n4), .A2(n_majority7_module_108_n6), .ZN(
        n_majority7_module_108__or_module_3_res) );
  AND2_X1 u_majority7_module_108__and_module_4_U1 ( .A1(
        n_majority7_module_108__and_module_2_res), .A2(
        n_majority7_module_108__and_module_1_res), .ZN(
        n_majority7_module_108__and_module_4_res) );
  OR2_X1 u_majority7_module_108__or_module_4_U1 ( .A1(
        n_majority7_module_108__and_module_1_res), .A2(
        n_majority7_module_108__and_module_2_res), .ZN(
        n_majority7_module_108__or_module_4_res) );
  AND2_X1 u_majority7_module_108__and_module_5_U1 ( .A1(
        n_majority7_module_108__and_module_3_res), .A2(
        n_majority7_module_108_n2), .ZN(
        n_majority7_module_108__and_module_5_res) );
  OR2_X1 u_majority7_module_108__or_module_5_U1 ( .A1(
        n_majority7_module_108_n2), .A2(
        n_majority7_module_108__and_module_3_res), .ZN(
        n_majority7_module_108__or_module_5_res) );
  AND2_X1 u_majority7_module_108__and_module_6_U1 ( .A1(
        n_majority7_module_108__or_module_1_res), .A2(
        n_majority7_module_108__or_module_2_res), .ZN(
        n_majority7_module_108__and_module_6_res) );
  OR2_X1 u_majority7_module_108__or_module_6_U1 ( .A1(
        n_majority7_module_108__or_module_2_res), .A2(
        n_majority7_module_108__or_module_1_res), .ZN(
        n_majority7_module_108__or_module_6_res) );
  OR2_X1 u_majority7_module_108__or_module_7_U1 ( .A1(
        n_majority7_module_108__and_module_4_res), .A2(
        n_majority7_module_108__and_module_5_res), .ZN(
        n_majority7_module_108__or_module_7_res) );
  AND2_X1 u_majority7_module_108__and_module_7_U1 ( .A1(
        n_majority7_module_108__or_module_3_res), .A2(
        n_majority7_module_108__or_module_4_res), .ZN(
        n_majority7_module_108__and_module_7_res) );
  OR2_X1 u_majority7_module_108__or_module_8_U1 ( .A1(
        n_majority7_module_108__or_module_4_res), .A2(
        n_majority7_module_108__or_module_3_res), .ZN(
        n_majority7_module_108__or_module_8_res) );
  AND2_X1 u_majority7_module_108__and_module_8_U1 ( .A1(
        n_majority7_module_108__or_module_5_res), .A2(
        n_majority7_module_108__and_module_6_res), .ZN(
        n_majority7_module_108__and_module_8_res) );
  OR2_X1 u_majority7_module_108__or_module_9_U1 ( .A1(
        n_majority7_module_108__and_module_6_res), .A2(
        n_majority7_module_108__or_module_5_res), .ZN(
        n_majority7_module_108__or_module_9_res) );
  OR2_X1 u_majority7_module_108__or_module_10_U1 ( .A1(
        n_majority7_module_108__or_module_7_res), .A2(
        n_majority7_module_108__and_module_7_res), .ZN(
        n_majority7_module_108__or_module_10_res) );
  AND2_X1 u_majority7_module_108__and_module_9_U1 ( .A1(
        n_majority7_module_108__or_module_6_res), .A2(
        n_majority7_module_108__or_module_9_res), .ZN(
        n_majority7_module_108__and_module_9_res) );
  OR2_X1 u_majority7_module_108__or_module_11_U1 ( .A1(
        n_majority7_module_108__or_module_10_res), .A2(
        n_majority7_module_108__and_module_8_res), .ZN(
        n_majority7_module_108__or_module_11_res) );
  AND2_X1 u_majority7_module_108__and_module_10_U1 ( .A1(
        n_majority7_module_108__or_module_8_res), .A2(
        n_majority7_module_108__and_module_9_res), .ZN(
        n_majority7_module_108__and_module_10_res) );
  AND2_X1 u_majority7_module_108__and_module_11_U1 ( .A1(
        n_majority7_module_108__and_module_10_res), .A2(
        n_majority7_module_108__or_module_11_res), .ZN(
        n_majority7_module_108_res) );
  DFF_X1 u_reg_module_109__cini_mul_v000_reg ( .D(n_majority7_module_108_res), 
        .CK(clock_6), .Q(n_reg_module_109_res), .QN() );
  BUF_X1 u_majority7_module_109_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_109_n7) );
  BUF_X1 u_majority7_module_109_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_109_n6) );
  BUF_X1 u_majority7_module_109_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_109_n5) );
  BUF_X1 u_majority7_module_109_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_109_n4) );
  BUF_X1 u_majority7_module_109_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_109_n3) );
  BUF_X1 u_majority7_module_109_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_109_n2) );
  BUF_X1 u_majority7_module_109_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_109_n1) );
  AND2_X1 u_majority7_module_109__and_module_1_U1 ( .A1(
        n_majority7_module_109_n7), .A2(n_majority7_module_109_n1), .ZN(
        n_majority7_module_109__and_module_1_res) );
  OR2_X1 u_majority7_module_109__or_module_1_U1 ( .A1(
        n_majority7_module_109_n1), .A2(n_majority7_module_109_n7), .ZN(
        n_majority7_module_109__or_module_1_res) );
  AND2_X1 u_majority7_module_109__and_module_2_U1 ( .A1(
        n_majority7_module_109_n5), .A2(n_majority7_module_109_n3), .ZN(
        n_majority7_module_109__and_module_2_res) );
  OR2_X1 u_majority7_module_109__or_module_2_U1 ( .A1(
        n_majority7_module_109_n3), .A2(n_majority7_module_109_n5), .ZN(
        n_majority7_module_109__or_module_2_res) );
  AND2_X1 u_majority7_module_109__and_module_3_U1 ( .A1(
        n_majority7_module_109_n6), .A2(n_majority7_module_109_n4), .ZN(
        n_majority7_module_109__and_module_3_res) );
  OR2_X1 u_majority7_module_109__or_module_3_U1 ( .A1(
        n_majority7_module_109_n4), .A2(n_majority7_module_109_n6), .ZN(
        n_majority7_module_109__or_module_3_res) );
  AND2_X1 u_majority7_module_109__and_module_4_U1 ( .A1(
        n_majority7_module_109__and_module_2_res), .A2(
        n_majority7_module_109__and_module_1_res), .ZN(
        n_majority7_module_109__and_module_4_res) );
  OR2_X1 u_majority7_module_109__or_module_4_U1 ( .A1(
        n_majority7_module_109__and_module_1_res), .A2(
        n_majority7_module_109__and_module_2_res), .ZN(
        n_majority7_module_109__or_module_4_res) );
  AND2_X1 u_majority7_module_109__and_module_5_U1 ( .A1(
        n_majority7_module_109__and_module_3_res), .A2(
        n_majority7_module_109_n2), .ZN(
        n_majority7_module_109__and_module_5_res) );
  OR2_X1 u_majority7_module_109__or_module_5_U1 ( .A1(
        n_majority7_module_109_n2), .A2(
        n_majority7_module_109__and_module_3_res), .ZN(
        n_majority7_module_109__or_module_5_res) );
  AND2_X1 u_majority7_module_109__and_module_6_U1 ( .A1(
        n_majority7_module_109__or_module_1_res), .A2(
        n_majority7_module_109__or_module_2_res), .ZN(
        n_majority7_module_109__and_module_6_res) );
  OR2_X1 u_majority7_module_109__or_module_6_U1 ( .A1(
        n_majority7_module_109__or_module_2_res), .A2(
        n_majority7_module_109__or_module_1_res), .ZN(
        n_majority7_module_109__or_module_6_res) );
  OR2_X1 u_majority7_module_109__or_module_7_U1 ( .A1(
        n_majority7_module_109__and_module_4_res), .A2(
        n_majority7_module_109__and_module_5_res), .ZN(
        n_majority7_module_109__or_module_7_res) );
  AND2_X1 u_majority7_module_109__and_module_7_U1 ( .A1(
        n_majority7_module_109__or_module_3_res), .A2(
        n_majority7_module_109__or_module_4_res), .ZN(
        n_majority7_module_109__and_module_7_res) );
  OR2_X1 u_majority7_module_109__or_module_8_U1 ( .A1(
        n_majority7_module_109__or_module_4_res), .A2(
        n_majority7_module_109__or_module_3_res), .ZN(
        n_majority7_module_109__or_module_8_res) );
  AND2_X1 u_majority7_module_109__and_module_8_U1 ( .A1(
        n_majority7_module_109__or_module_5_res), .A2(
        n_majority7_module_109__and_module_6_res), .ZN(
        n_majority7_module_109__and_module_8_res) );
  OR2_X1 u_majority7_module_109__or_module_9_U1 ( .A1(
        n_majority7_module_109__and_module_6_res), .A2(
        n_majority7_module_109__or_module_5_res), .ZN(
        n_majority7_module_109__or_module_9_res) );
  OR2_X1 u_majority7_module_109__or_module_10_U1 ( .A1(
        n_majority7_module_109__or_module_7_res), .A2(
        n_majority7_module_109__and_module_7_res), .ZN(
        n_majority7_module_109__or_module_10_res) );
  AND2_X1 u_majority7_module_109__and_module_9_U1 ( .A1(
        n_majority7_module_109__or_module_6_res), .A2(
        n_majority7_module_109__or_module_9_res), .ZN(
        n_majority7_module_109__and_module_9_res) );
  OR2_X1 u_majority7_module_109__or_module_11_U1 ( .A1(
        n_majority7_module_109__or_module_10_res), .A2(
        n_majority7_module_109__and_module_8_res), .ZN(
        n_majority7_module_109__or_module_11_res) );
  AND2_X1 u_majority7_module_109__and_module_10_U1 ( .A1(
        n_majority7_module_109__or_module_8_res), .A2(
        n_majority7_module_109__and_module_9_res), .ZN(
        n_majority7_module_109__and_module_10_res) );
  AND2_X1 u_majority7_module_109__and_module_11_U1 ( .A1(
        n_majority7_module_109__and_module_10_res), .A2(
        n_majority7_module_109__or_module_11_res), .ZN(
        n_majority7_module_109_res) );
  DFF_X1 u_reg_module_110__cini_mul_v000_reg ( .D(n_majority7_module_109_res), 
        .CK(clock_6), .Q(n_reg_module_110_res), .QN() );
  BUF_X1 u_majority7_module_110_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_110_n7) );
  BUF_X1 u_majority7_module_110_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_110_n6) );
  BUF_X1 u_majority7_module_110_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_110_n5) );
  BUF_X1 u_majority7_module_110_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_110_n4) );
  BUF_X1 u_majority7_module_110_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_110_n3) );
  BUF_X1 u_majority7_module_110_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_110_n2) );
  BUF_X1 u_majority7_module_110_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_110_n1) );
  AND2_X1 u_majority7_module_110__and_module_1_U1 ( .A1(
        n_majority7_module_110_n7), .A2(n_majority7_module_110_n1), .ZN(
        n_majority7_module_110__and_module_1_res) );
  OR2_X1 u_majority7_module_110__or_module_1_U1 ( .A1(
        n_majority7_module_110_n1), .A2(n_majority7_module_110_n7), .ZN(
        n_majority7_module_110__or_module_1_res) );
  AND2_X1 u_majority7_module_110__and_module_2_U1 ( .A1(
        n_majority7_module_110_n5), .A2(n_majority7_module_110_n3), .ZN(
        n_majority7_module_110__and_module_2_res) );
  OR2_X1 u_majority7_module_110__or_module_2_U1 ( .A1(
        n_majority7_module_110_n3), .A2(n_majority7_module_110_n5), .ZN(
        n_majority7_module_110__or_module_2_res) );
  AND2_X1 u_majority7_module_110__and_module_3_U1 ( .A1(
        n_majority7_module_110_n6), .A2(n_majority7_module_110_n4), .ZN(
        n_majority7_module_110__and_module_3_res) );
  OR2_X1 u_majority7_module_110__or_module_3_U1 ( .A1(
        n_majority7_module_110_n4), .A2(n_majority7_module_110_n6), .ZN(
        n_majority7_module_110__or_module_3_res) );
  AND2_X1 u_majority7_module_110__and_module_4_U1 ( .A1(
        n_majority7_module_110__and_module_2_res), .A2(
        n_majority7_module_110__and_module_1_res), .ZN(
        n_majority7_module_110__and_module_4_res) );
  OR2_X1 u_majority7_module_110__or_module_4_U1 ( .A1(
        n_majority7_module_110__and_module_1_res), .A2(
        n_majority7_module_110__and_module_2_res), .ZN(
        n_majority7_module_110__or_module_4_res) );
  AND2_X1 u_majority7_module_110__and_module_5_U1 ( .A1(
        n_majority7_module_110__and_module_3_res), .A2(
        n_majority7_module_110_n2), .ZN(
        n_majority7_module_110__and_module_5_res) );
  OR2_X1 u_majority7_module_110__or_module_5_U1 ( .A1(
        n_majority7_module_110_n2), .A2(
        n_majority7_module_110__and_module_3_res), .ZN(
        n_majority7_module_110__or_module_5_res) );
  AND2_X1 u_majority7_module_110__and_module_6_U1 ( .A1(
        n_majority7_module_110__or_module_1_res), .A2(
        n_majority7_module_110__or_module_2_res), .ZN(
        n_majority7_module_110__and_module_6_res) );
  OR2_X1 u_majority7_module_110__or_module_6_U1 ( .A1(
        n_majority7_module_110__or_module_2_res), .A2(
        n_majority7_module_110__or_module_1_res), .ZN(
        n_majority7_module_110__or_module_6_res) );
  OR2_X1 u_majority7_module_110__or_module_7_U1 ( .A1(
        n_majority7_module_110__and_module_4_res), .A2(
        n_majority7_module_110__and_module_5_res), .ZN(
        n_majority7_module_110__or_module_7_res) );
  AND2_X1 u_majority7_module_110__and_module_7_U1 ( .A1(
        n_majority7_module_110__or_module_3_res), .A2(
        n_majority7_module_110__or_module_4_res), .ZN(
        n_majority7_module_110__and_module_7_res) );
  OR2_X1 u_majority7_module_110__or_module_8_U1 ( .A1(
        n_majority7_module_110__or_module_4_res), .A2(
        n_majority7_module_110__or_module_3_res), .ZN(
        n_majority7_module_110__or_module_8_res) );
  AND2_X1 u_majority7_module_110__and_module_8_U1 ( .A1(
        n_majority7_module_110__or_module_5_res), .A2(
        n_majority7_module_110__and_module_6_res), .ZN(
        n_majority7_module_110__and_module_8_res) );
  OR2_X1 u_majority7_module_110__or_module_9_U1 ( .A1(
        n_majority7_module_110__and_module_6_res), .A2(
        n_majority7_module_110__or_module_5_res), .ZN(
        n_majority7_module_110__or_module_9_res) );
  OR2_X1 u_majority7_module_110__or_module_10_U1 ( .A1(
        n_majority7_module_110__or_module_7_res), .A2(
        n_majority7_module_110__and_module_7_res), .ZN(
        n_majority7_module_110__or_module_10_res) );
  AND2_X1 u_majority7_module_110__and_module_9_U1 ( .A1(
        n_majority7_module_110__or_module_6_res), .A2(
        n_majority7_module_110__or_module_9_res), .ZN(
        n_majority7_module_110__and_module_9_res) );
  OR2_X1 u_majority7_module_110__or_module_11_U1 ( .A1(
        n_majority7_module_110__or_module_10_res), .A2(
        n_majority7_module_110__and_module_8_res), .ZN(
        n_majority7_module_110__or_module_11_res) );
  AND2_X1 u_majority7_module_110__and_module_10_U1 ( .A1(
        n_majority7_module_110__or_module_8_res), .A2(
        n_majority7_module_110__and_module_9_res), .ZN(
        n_majority7_module_110__and_module_10_res) );
  AND2_X1 u_majority7_module_110__and_module_11_U1 ( .A1(
        n_majority7_module_110__and_module_10_res), .A2(
        n_majority7_module_110__or_module_11_res), .ZN(
        n_majority7_module_110_res) );
  DFF_X1 u_reg_module_111__cini_mul_v000_reg ( .D(n_majority7_module_110_res), 
        .CK(clock_6), .Q(n_reg_module_111_res), .QN() );
  BUF_X1 u_majority7_module_111_U7 ( .A(n_xor_module_84_res), .Z(
        n_majority7_module_111_n7) );
  BUF_X1 u_majority7_module_111_U6 ( .A(n_xor_module_72_res), .Z(
        n_majority7_module_111_n6) );
  BUF_X1 u_majority7_module_111_U5 ( .A(n_xor_module_48_res), .Z(
        n_majority7_module_111_n5) );
  BUF_X1 u_majority7_module_111_U4 ( .A(n_xor_module_60_res), .Z(
        n_majority7_module_111_n4) );
  BUF_X1 u_majority7_module_111_U3 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_111_n3) );
  BUF_X1 u_majority7_module_111_U2 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_111_n2) );
  BUF_X1 u_majority7_module_111_U1 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_111_n1) );
  AND2_X1 u_majority7_module_111__and_module_1_U1 ( .A1(
        n_majority7_module_111_n7), .A2(n_majority7_module_111_n1), .ZN(
        n_majority7_module_111__and_module_1_res) );
  OR2_X1 u_majority7_module_111__or_module_1_U1 ( .A1(
        n_majority7_module_111_n1), .A2(n_majority7_module_111_n7), .ZN(
        n_majority7_module_111__or_module_1_res) );
  AND2_X1 u_majority7_module_111__and_module_2_U1 ( .A1(
        n_majority7_module_111_n5), .A2(n_majority7_module_111_n3), .ZN(
        n_majority7_module_111__and_module_2_res) );
  OR2_X1 u_majority7_module_111__or_module_2_U1 ( .A1(
        n_majority7_module_111_n3), .A2(n_majority7_module_111_n5), .ZN(
        n_majority7_module_111__or_module_2_res) );
  AND2_X1 u_majority7_module_111__and_module_3_U1 ( .A1(
        n_majority7_module_111_n6), .A2(n_majority7_module_111_n4), .ZN(
        n_majority7_module_111__and_module_3_res) );
  OR2_X1 u_majority7_module_111__or_module_3_U1 ( .A1(
        n_majority7_module_111_n4), .A2(n_majority7_module_111_n6), .ZN(
        n_majority7_module_111__or_module_3_res) );
  AND2_X1 u_majority7_module_111__and_module_4_U1 ( .A1(
        n_majority7_module_111__and_module_2_res), .A2(
        n_majority7_module_111__and_module_1_res), .ZN(
        n_majority7_module_111__and_module_4_res) );
  OR2_X1 u_majority7_module_111__or_module_4_U1 ( .A1(
        n_majority7_module_111__and_module_1_res), .A2(
        n_majority7_module_111__and_module_2_res), .ZN(
        n_majority7_module_111__or_module_4_res) );
  AND2_X1 u_majority7_module_111__and_module_5_U1 ( .A1(
        n_majority7_module_111__and_module_3_res), .A2(
        n_majority7_module_111_n2), .ZN(
        n_majority7_module_111__and_module_5_res) );
  OR2_X1 u_majority7_module_111__or_module_5_U1 ( .A1(
        n_majority7_module_111_n2), .A2(
        n_majority7_module_111__and_module_3_res), .ZN(
        n_majority7_module_111__or_module_5_res) );
  AND2_X1 u_majority7_module_111__and_module_6_U1 ( .A1(
        n_majority7_module_111__or_module_1_res), .A2(
        n_majority7_module_111__or_module_2_res), .ZN(
        n_majority7_module_111__and_module_6_res) );
  OR2_X1 u_majority7_module_111__or_module_6_U1 ( .A1(
        n_majority7_module_111__or_module_2_res), .A2(
        n_majority7_module_111__or_module_1_res), .ZN(
        n_majority7_module_111__or_module_6_res) );
  OR2_X1 u_majority7_module_111__or_module_7_U1 ( .A1(
        n_majority7_module_111__and_module_4_res), .A2(
        n_majority7_module_111__and_module_5_res), .ZN(
        n_majority7_module_111__or_module_7_res) );
  AND2_X1 u_majority7_module_111__and_module_7_U1 ( .A1(
        n_majority7_module_111__or_module_3_res), .A2(
        n_majority7_module_111__or_module_4_res), .ZN(
        n_majority7_module_111__and_module_7_res) );
  OR2_X1 u_majority7_module_111__or_module_8_U1 ( .A1(
        n_majority7_module_111__or_module_4_res), .A2(
        n_majority7_module_111__or_module_3_res), .ZN(
        n_majority7_module_111__or_module_8_res) );
  AND2_X1 u_majority7_module_111__and_module_8_U1 ( .A1(
        n_majority7_module_111__or_module_5_res), .A2(
        n_majority7_module_111__and_module_6_res), .ZN(
        n_majority7_module_111__and_module_8_res) );
  OR2_X1 u_majority7_module_111__or_module_9_U1 ( .A1(
        n_majority7_module_111__and_module_6_res), .A2(
        n_majority7_module_111__or_module_5_res), .ZN(
        n_majority7_module_111__or_module_9_res) );
  OR2_X1 u_majority7_module_111__or_module_10_U1 ( .A1(
        n_majority7_module_111__or_module_7_res), .A2(
        n_majority7_module_111__and_module_7_res), .ZN(
        n_majority7_module_111__or_module_10_res) );
  AND2_X1 u_majority7_module_111__and_module_9_U1 ( .A1(
        n_majority7_module_111__or_module_6_res), .A2(
        n_majority7_module_111__or_module_9_res), .ZN(
        n_majority7_module_111__and_module_9_res) );
  OR2_X1 u_majority7_module_111__or_module_11_U1 ( .A1(
        n_majority7_module_111__or_module_10_res), .A2(
        n_majority7_module_111__and_module_8_res), .ZN(
        n_majority7_module_111__or_module_11_res) );
  AND2_X1 u_majority7_module_111__and_module_10_U1 ( .A1(
        n_majority7_module_111__or_module_8_res), .A2(
        n_majority7_module_111__and_module_9_res), .ZN(
        n_majority7_module_111__and_module_10_res) );
  AND2_X1 u_majority7_module_111__and_module_11_U1 ( .A1(
        n_majority7_module_111__and_module_10_res), .A2(
        n_majority7_module_111__or_module_11_res), .ZN(
        n_majority7_module_111_res) );
  DFF_X1 u_reg_module_112__cini_mul_v000_reg ( .D(n_majority7_module_111_res), 
        .CK(clock_6), .Q(n_reg_module_112_res), .QN() );
  AND2_X1 u_and_module_1_U1 ( .A1(n_reg_module_1_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_1_res) );
  DFF_X1 u_reg_module_113__cini_mul_v000_reg ( .D(n_and_module_1_res), .CK(
        clock_0), .Q(n_reg_module_113_res), .QN() );
  AND2_X1 u_and_module_2_U1 ( .A1(n_reg_module_5_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_2_res) );
  XOR2_X1 u_xor_module_85_U1 ( .A(p_rand_6), .B(n_and_module_2_res), .Z(
        n_xor_module_85_res) );
  DFF_X1 u_reg_module_114__cini_mul_v000_reg ( .D(n_xor_module_85_res), .CK(
        clock_0), .Q(n_reg_module_114_res), .QN() );
  AND2_X1 u_and_module_3_U1 ( .A1(n_reg_module_9_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_3_res) );
  XOR2_X1 u_xor_module_86_U1 ( .A(p_rand_7), .B(n_and_module_3_res), .Z(
        n_xor_module_86_res) );
  DFF_X1 u_reg_module_115__cini_mul_v000_reg ( .D(n_xor_module_86_res), .CK(
        clock_0), .Q(n_reg_module_115_res), .QN() );
  AND2_X1 u_and_module_4_U1 ( .A1(n_reg_module_13_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_4_res) );
  XOR2_X1 u_xor_module_87_U1 ( .A(p_rand_8), .B(n_and_module_4_res), .Z(
        n_xor_module_87_res) );
  DFF_X1 u_reg_module_116__cini_mul_v000_reg ( .D(n_xor_module_87_res), .CK(
        clock_0), .Q(n_reg_module_116_res), .QN() );
  AND2_X1 u_and_module_5_U1 ( .A1(n_reg_module_2_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_5_res) );
  XOR2_X1 u_xor_module_88_U1 ( .A(p_rand_6), .B(n_and_module_5_res), .Z(
        n_xor_module_88_res) );
  DFF_X1 u_reg_module_117__cini_mul_v000_reg ( .D(n_xor_module_88_res), .CK(
        clock_0), .Q(n_reg_module_117_res), .QN() );
  AND2_X1 u_and_module_6_U1 ( .A1(n_reg_module_6_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_6_res) );
  DFF_X1 u_reg_module_118__cini_mul_v000_reg ( .D(n_and_module_6_res), .CK(
        clock_0), .Q(n_reg_module_118_res), .QN() );
  AND2_X1 u_and_module_7_U1 ( .A1(n_reg_module_10_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_7_res) );
  XOR2_X1 u_xor_module_89_U1 ( .A(p_rand_9), .B(n_and_module_7_res), .Z(
        n_xor_module_89_res) );
  DFF_X1 u_reg_module_119__cini_mul_v000_reg ( .D(n_xor_module_89_res), .CK(
        clock_0), .Q(n_reg_module_119_res), .QN() );
  AND2_X1 u_and_module_8_U1 ( .A1(n_reg_module_14_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_8_res) );
  XOR2_X1 u_xor_module_90_U1 ( .A(p_rand_10), .B(n_and_module_8_res), .Z(
        n_xor_module_90_res) );
  DFF_X1 u_reg_module_120__cini_mul_v000_reg ( .D(n_xor_module_90_res), .CK(
        clock_0), .Q(n_reg_module_120_res), .QN() );
  AND2_X1 u_and_module_9_U1 ( .A1(n_reg_module_3_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_9_res) );
  XOR2_X1 u_xor_module_91_U1 ( .A(p_rand_7), .B(n_and_module_9_res), .Z(
        n_xor_module_91_res) );
  DFF_X1 u_reg_module_121__cini_mul_v000_reg ( .D(n_xor_module_91_res), .CK(
        clock_0), .Q(n_reg_module_121_res), .QN() );
  AND2_X1 u_and_module_10_U1 ( .A1(n_reg_module_7_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_10_res) );
  XOR2_X1 u_xor_module_92_U1 ( .A(p_rand_9), .B(n_and_module_10_res), .Z(
        n_xor_module_92_res) );
  DFF_X1 u_reg_module_122__cini_mul_v000_reg ( .D(n_xor_module_92_res), .CK(
        clock_0), .Q(n_reg_module_122_res), .QN() );
  AND2_X1 u_and_module_11_U1 ( .A1(n_reg_module_11_res), .A2(io_i0_s2_d0), 
        .ZN(n_and_module_11_res) );
  DFF_X1 u_reg_module_123__cini_mul_v000_reg ( .D(n_and_module_11_res), .CK(
        clock_0), .Q(n_reg_module_123_res), .QN() );
  AND2_X1 u_and_module_12_U1 ( .A1(n_reg_module_15_res), .A2(io_i0_s2_d0), 
        .ZN(n_and_module_12_res) );
  XOR2_X1 u_xor_module_93_U1 ( .A(p_rand_11), .B(n_and_module_12_res), .Z(
        n_xor_module_93_res) );
  DFF_X1 u_reg_module_124__cini_mul_v000_reg ( .D(n_xor_module_93_res), .CK(
        clock_0), .Q(n_reg_module_124_res), .QN() );
  AND2_X1 u_and_module_13_U1 ( .A1(n_reg_module_4_res), .A2(io_i0_s3_d0), .ZN(
        n_and_module_13_res) );
  XOR2_X1 u_xor_module_94_U1 ( .A(p_rand_8), .B(n_and_module_13_res), .Z(
        n_xor_module_94_res) );
  DFF_X1 u_reg_module_125__cini_mul_v000_reg ( .D(n_xor_module_94_res), .CK(
        clock_0), .Q(n_reg_module_125_res), .QN() );
  AND2_X1 u_and_module_14_U1 ( .A1(n_reg_module_8_res), .A2(io_i0_s3_d0), .ZN(
        n_and_module_14_res) );
  XOR2_X1 u_xor_module_95_U1 ( .A(p_rand_10), .B(n_and_module_14_res), .Z(
        n_xor_module_95_res) );
  DFF_X1 u_reg_module_126__cini_mul_v000_reg ( .D(n_xor_module_95_res), .CK(
        clock_0), .Q(n_reg_module_126_res), .QN() );
  AND2_X1 u_and_module_15_U1 ( .A1(n_reg_module_12_res), .A2(io_i0_s3_d0), 
        .ZN(n_and_module_15_res) );
  XOR2_X1 u_xor_module_96_U1 ( .A(p_rand_11), .B(n_and_module_15_res), .Z(
        n_xor_module_96_res) );
  DFF_X1 u_reg_module_127__cini_mul_v000_reg ( .D(n_xor_module_96_res), .CK(
        clock_0), .Q(n_reg_module_127_res), .QN() );
  AND2_X1 u_and_module_16_U1 ( .A1(n_reg_module_16_res), .A2(io_i0_s3_d0), 
        .ZN(n_and_module_16_res) );
  DFF_X1 u_reg_module_128__cini_mul_v000_reg ( .D(n_and_module_16_res), .CK(
        clock_0), .Q(n_reg_module_128_res), .QN() );
  AND2_X1 u_and_module_17_U1 ( .A1(n_reg_module_17_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_17_res) );
  DFF_X1 u_reg_module_129__cini_mul_v000_reg ( .D(n_and_module_17_res), .CK(
        clock_1), .Q(n_reg_module_129_res), .QN() );
  AND2_X1 u_and_module_18_U1 ( .A1(n_reg_module_21_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_18_res) );
  XOR2_X1 u_xor_module_97_U1 ( .A(p_rand_6), .B(n_and_module_18_res), .Z(
        n_xor_module_97_res) );
  DFF_X1 u_reg_module_130__cini_mul_v000_reg ( .D(n_xor_module_97_res), .CK(
        clock_1), .Q(n_reg_module_130_res), .QN() );
  AND2_X1 u_and_module_19_U1 ( .A1(n_reg_module_25_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_19_res) );
  XOR2_X1 u_xor_module_98_U1 ( .A(p_rand_7), .B(n_and_module_19_res), .Z(
        n_xor_module_98_res) );
  DFF_X1 u_reg_module_131__cini_mul_v000_reg ( .D(n_xor_module_98_res), .CK(
        clock_1), .Q(n_reg_module_131_res), .QN() );
  AND2_X1 u_and_module_20_U1 ( .A1(n_reg_module_29_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_20_res) );
  XOR2_X1 u_xor_module_99_U1 ( .A(p_rand_8), .B(n_and_module_20_res), .Z(
        n_xor_module_99_res) );
  DFF_X1 u_reg_module_132__cini_mul_v000_reg ( .D(n_xor_module_99_res), .CK(
        clock_1), .Q(n_reg_module_132_res), .QN() );
  AND2_X1 u_and_module_21_U1 ( .A1(n_reg_module_18_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_21_res) );
  XOR2_X1 u_xor_module_100_U1 ( .A(p_rand_6), .B(n_and_module_21_res), .Z(
        n_xor_module_100_res) );
  DFF_X1 u_reg_module_133__cini_mul_v000_reg ( .D(n_xor_module_100_res), .CK(
        clock_1), .Q(n_reg_module_133_res), .QN() );
  AND2_X1 u_and_module_22_U1 ( .A1(n_reg_module_22_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_22_res) );
  DFF_X1 u_reg_module_134__cini_mul_v000_reg ( .D(n_and_module_22_res), .CK(
        clock_1), .Q(n_reg_module_134_res), .QN() );
  AND2_X1 u_and_module_23_U1 ( .A1(n_reg_module_26_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_23_res) );
  XOR2_X1 u_xor_module_101_U1 ( .A(p_rand_9), .B(n_and_module_23_res), .Z(
        n_xor_module_101_res) );
  DFF_X1 u_reg_module_135__cini_mul_v000_reg ( .D(n_xor_module_101_res), .CK(
        clock_1), .Q(n_reg_module_135_res), .QN() );
  AND2_X1 u_and_module_24_U1 ( .A1(n_reg_module_30_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_24_res) );
  XOR2_X1 u_xor_module_102_U1 ( .A(p_rand_10), .B(n_and_module_24_res), .Z(
        n_xor_module_102_res) );
  DFF_X1 u_reg_module_136__cini_mul_v000_reg ( .D(n_xor_module_102_res), .CK(
        clock_1), .Q(n_reg_module_136_res), .QN() );
  AND2_X1 u_and_module_25_U1 ( .A1(n_reg_module_19_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_25_res) );
  XOR2_X1 u_xor_module_103_U1 ( .A(p_rand_7), .B(n_and_module_25_res), .Z(
        n_xor_module_103_res) );
  DFF_X1 u_reg_module_137__cini_mul_v000_reg ( .D(n_xor_module_103_res), .CK(
        clock_1), .Q(n_reg_module_137_res), .QN() );
  AND2_X1 u_and_module_26_U1 ( .A1(n_reg_module_23_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_26_res) );
  XOR2_X1 u_xor_module_104_U1 ( .A(p_rand_9), .B(n_and_module_26_res), .Z(
        n_xor_module_104_res) );
  DFF_X1 u_reg_module_138__cini_mul_v000_reg ( .D(n_xor_module_104_res), .CK(
        clock_1), .Q(n_reg_module_138_res), .QN() );
  AND2_X1 u_and_module_27_U1 ( .A1(n_reg_module_27_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_27_res) );
  DFF_X1 u_reg_module_139__cini_mul_v000_reg ( .D(n_and_module_27_res), .CK(
        clock_1), .Q(n_reg_module_139_res), .QN() );
  AND2_X1 u_and_module_28_U1 ( .A1(n_reg_module_31_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_28_res) );
  XOR2_X1 u_xor_module_105_U1 ( .A(p_rand_11), .B(n_and_module_28_res), .Z(
        n_xor_module_105_res) );
  DFF_X1 u_reg_module_140__cini_mul_v000_reg ( .D(n_xor_module_105_res), .CK(
        clock_1), .Q(n_reg_module_140_res), .QN() );
  AND2_X1 u_and_module_29_U1 ( .A1(n_reg_module_20_res), .A2(io_i0_s3_d1), 
        .ZN(n_and_module_29_res) );
  XOR2_X1 u_xor_module_106_U1 ( .A(p_rand_8), .B(n_and_module_29_res), .Z(
        n_xor_module_106_res) );
  DFF_X1 u_reg_module_141__cini_mul_v000_reg ( .D(n_xor_module_106_res), .CK(
        clock_1), .Q(n_reg_module_141_res), .QN() );
  AND2_X1 u_and_module_30_U1 ( .A1(n_reg_module_24_res), .A2(io_i0_s3_d1), 
        .ZN(n_and_module_30_res) );
  XOR2_X1 u_xor_module_107_U1 ( .A(p_rand_10), .B(n_and_module_30_res), .Z(
        n_xor_module_107_res) );
  DFF_X1 u_reg_module_142__cini_mul_v000_reg ( .D(n_xor_module_107_res), .CK(
        clock_1), .Q(n_reg_module_142_res), .QN() );
  AND2_X1 u_and_module_31_U1 ( .A1(n_reg_module_28_res), .A2(io_i0_s3_d1), 
        .ZN(n_and_module_31_res) );
  XOR2_X1 u_xor_module_108_U1 ( .A(p_rand_11), .B(n_and_module_31_res), .Z(
        n_xor_module_108_res) );
  DFF_X1 u_reg_module_143__cini_mul_v000_reg ( .D(n_xor_module_108_res), .CK(
        clock_1), .Q(n_reg_module_143_res), .QN() );
  AND2_X1 u_and_module_32_U1 ( .A1(n_reg_module_32_res), .A2(io_i0_s3_d1), 
        .ZN(n_and_module_32_res) );
  DFF_X1 u_reg_module_144__cini_mul_v000_reg ( .D(n_and_module_32_res), .CK(
        clock_1), .Q(n_reg_module_144_res), .QN() );
  AND2_X1 u_and_module_33_U1 ( .A1(n_reg_module_33_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_33_res) );
  DFF_X1 u_reg_module_145__cini_mul_v000_reg ( .D(n_and_module_33_res), .CK(
        clock_2), .Q(n_reg_module_145_res), .QN() );
  AND2_X1 u_and_module_34_U1 ( .A1(n_reg_module_37_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_34_res) );
  XOR2_X1 u_xor_module_109_U1 ( .A(p_rand_6), .B(n_and_module_34_res), .Z(
        n_xor_module_109_res) );
  DFF_X1 u_reg_module_146__cini_mul_v000_reg ( .D(n_xor_module_109_res), .CK(
        clock_2), .Q(n_reg_module_146_res), .QN() );
  AND2_X1 u_and_module_35_U1 ( .A1(n_reg_module_41_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_35_res) );
  XOR2_X1 u_xor_module_110_U1 ( .A(p_rand_7), .B(n_and_module_35_res), .Z(
        n_xor_module_110_res) );
  DFF_X1 u_reg_module_147__cini_mul_v000_reg ( .D(n_xor_module_110_res), .CK(
        clock_2), .Q(n_reg_module_147_res), .QN() );
  AND2_X1 u_and_module_36_U1 ( .A1(n_reg_module_45_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_36_res) );
  XOR2_X1 u_xor_module_111_U1 ( .A(p_rand_8), .B(n_and_module_36_res), .Z(
        n_xor_module_111_res) );
  DFF_X1 u_reg_module_148__cini_mul_v000_reg ( .D(n_xor_module_111_res), .CK(
        clock_2), .Q(n_reg_module_148_res), .QN() );
  AND2_X1 u_and_module_37_U1 ( .A1(n_reg_module_34_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_37_res) );
  XOR2_X1 u_xor_module_112_U1 ( .A(p_rand_6), .B(n_and_module_37_res), .Z(
        n_xor_module_112_res) );
  DFF_X1 u_reg_module_149__cini_mul_v000_reg ( .D(n_xor_module_112_res), .CK(
        clock_2), .Q(n_reg_module_149_res), .QN() );
  AND2_X1 u_and_module_38_U1 ( .A1(n_reg_module_38_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_38_res) );
  DFF_X1 u_reg_module_150__cini_mul_v000_reg ( .D(n_and_module_38_res), .CK(
        clock_2), .Q(n_reg_module_150_res), .QN() );
  AND2_X1 u_and_module_39_U1 ( .A1(n_reg_module_42_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_39_res) );
  XOR2_X1 u_xor_module_113_U1 ( .A(p_rand_9), .B(n_and_module_39_res), .Z(
        n_xor_module_113_res) );
  DFF_X1 u_reg_module_151__cini_mul_v000_reg ( .D(n_xor_module_113_res), .CK(
        clock_2), .Q(n_reg_module_151_res), .QN() );
  AND2_X1 u_and_module_40_U1 ( .A1(n_reg_module_46_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_40_res) );
  XOR2_X1 u_xor_module_114_U1 ( .A(p_rand_10), .B(n_and_module_40_res), .Z(
        n_xor_module_114_res) );
  DFF_X1 u_reg_module_152__cini_mul_v000_reg ( .D(n_xor_module_114_res), .CK(
        clock_2), .Q(n_reg_module_152_res), .QN() );
  AND2_X1 u_and_module_41_U1 ( .A1(n_reg_module_35_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_41_res) );
  XOR2_X1 u_xor_module_115_U1 ( .A(p_rand_7), .B(n_and_module_41_res), .Z(
        n_xor_module_115_res) );
  DFF_X1 u_reg_module_153__cini_mul_v000_reg ( .D(n_xor_module_115_res), .CK(
        clock_2), .Q(n_reg_module_153_res), .QN() );
  AND2_X1 u_and_module_42_U1 ( .A1(n_reg_module_39_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_42_res) );
  XOR2_X1 u_xor_module_116_U1 ( .A(p_rand_9), .B(n_and_module_42_res), .Z(
        n_xor_module_116_res) );
  DFF_X1 u_reg_module_154__cini_mul_v000_reg ( .D(n_xor_module_116_res), .CK(
        clock_2), .Q(n_reg_module_154_res), .QN() );
  AND2_X1 u_and_module_43_U1 ( .A1(n_reg_module_43_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_43_res) );
  DFF_X1 u_reg_module_155__cini_mul_v000_reg ( .D(n_and_module_43_res), .CK(
        clock_2), .Q(n_reg_module_155_res), .QN() );
  AND2_X1 u_and_module_44_U1 ( .A1(n_reg_module_47_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_44_res) );
  XOR2_X1 u_xor_module_117_U1 ( .A(p_rand_11), .B(n_and_module_44_res), .Z(
        n_xor_module_117_res) );
  DFF_X1 u_reg_module_156__cini_mul_v000_reg ( .D(n_xor_module_117_res), .CK(
        clock_2), .Q(n_reg_module_156_res), .QN() );
  AND2_X1 u_and_module_45_U1 ( .A1(n_reg_module_36_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_45_res) );
  XOR2_X1 u_xor_module_118_U1 ( .A(p_rand_8), .B(n_and_module_45_res), .Z(
        n_xor_module_118_res) );
  DFF_X1 u_reg_module_157__cini_mul_v000_reg ( .D(n_xor_module_118_res), .CK(
        clock_2), .Q(n_reg_module_157_res), .QN() );
  AND2_X1 u_and_module_46_U1 ( .A1(n_reg_module_40_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_46_res) );
  XOR2_X1 u_xor_module_119_U1 ( .A(p_rand_10), .B(n_and_module_46_res), .Z(
        n_xor_module_119_res) );
  DFF_X1 u_reg_module_158__cini_mul_v000_reg ( .D(n_xor_module_119_res), .CK(
        clock_2), .Q(n_reg_module_158_res), .QN() );
  AND2_X1 u_and_module_47_U1 ( .A1(n_reg_module_44_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_47_res) );
  XOR2_X1 u_xor_module_120_U1 ( .A(p_rand_11), .B(n_and_module_47_res), .Z(
        n_xor_module_120_res) );
  DFF_X1 u_reg_module_159__cini_mul_v000_reg ( .D(n_xor_module_120_res), .CK(
        clock_2), .Q(n_reg_module_159_res), .QN() );
  AND2_X1 u_and_module_48_U1 ( .A1(n_reg_module_48_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_48_res) );
  DFF_X1 u_reg_module_160__cini_mul_v000_reg ( .D(n_and_module_48_res), .CK(
        clock_2), .Q(n_reg_module_160_res), .QN() );
  AND2_X1 u_and_module_49_U1 ( .A1(n_reg_module_49_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_49_res) );
  DFF_X1 u_reg_module_161__cini_mul_v000_reg ( .D(n_and_module_49_res), .CK(
        clock_3), .Q(n_reg_module_161_res), .QN() );
  AND2_X1 u_and_module_50_U1 ( .A1(n_reg_module_53_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_50_res) );
  XOR2_X1 u_xor_module_121_U1 ( .A(p_rand_6), .B(n_and_module_50_res), .Z(
        n_xor_module_121_res) );
  DFF_X1 u_reg_module_162__cini_mul_v000_reg ( .D(n_xor_module_121_res), .CK(
        clock_3), .Q(n_reg_module_162_res), .QN() );
  AND2_X1 u_and_module_51_U1 ( .A1(n_reg_module_57_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_51_res) );
  XOR2_X1 u_xor_module_122_U1 ( .A(p_rand_7), .B(n_and_module_51_res), .Z(
        n_xor_module_122_res) );
  DFF_X1 u_reg_module_163__cini_mul_v000_reg ( .D(n_xor_module_122_res), .CK(
        clock_3), .Q(n_reg_module_163_res), .QN() );
  AND2_X1 u_and_module_52_U1 ( .A1(n_reg_module_61_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_52_res) );
  XOR2_X1 u_xor_module_123_U1 ( .A(p_rand_8), .B(n_and_module_52_res), .Z(
        n_xor_module_123_res) );
  DFF_X1 u_reg_module_164__cini_mul_v000_reg ( .D(n_xor_module_123_res), .CK(
        clock_3), .Q(n_reg_module_164_res), .QN() );
  AND2_X1 u_and_module_53_U1 ( .A1(n_reg_module_50_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_53_res) );
  XOR2_X1 u_xor_module_124_U1 ( .A(p_rand_6), .B(n_and_module_53_res), .Z(
        n_xor_module_124_res) );
  DFF_X1 u_reg_module_165__cini_mul_v000_reg ( .D(n_xor_module_124_res), .CK(
        clock_3), .Q(n_reg_module_165_res), .QN() );
  AND2_X1 u_and_module_54_U1 ( .A1(n_reg_module_54_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_54_res) );
  DFF_X1 u_reg_module_166__cini_mul_v000_reg ( .D(n_and_module_54_res), .CK(
        clock_3), .Q(n_reg_module_166_res), .QN() );
  AND2_X1 u_and_module_55_U1 ( .A1(n_reg_module_58_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_55_res) );
  XOR2_X1 u_xor_module_125_U1 ( .A(p_rand_9), .B(n_and_module_55_res), .Z(
        n_xor_module_125_res) );
  DFF_X1 u_reg_module_167__cini_mul_v000_reg ( .D(n_xor_module_125_res), .CK(
        clock_3), .Q(n_reg_module_167_res), .QN() );
  AND2_X1 u_and_module_56_U1 ( .A1(n_reg_module_62_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_56_res) );
  XOR2_X1 u_xor_module_126_U1 ( .A(p_rand_10), .B(n_and_module_56_res), .Z(
        n_xor_module_126_res) );
  DFF_X1 u_reg_module_168__cini_mul_v000_reg ( .D(n_xor_module_126_res), .CK(
        clock_3), .Q(n_reg_module_168_res), .QN() );
  AND2_X1 u_and_module_57_U1 ( .A1(n_reg_module_51_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_57_res) );
  XOR2_X1 u_xor_module_127_U1 ( .A(p_rand_7), .B(n_and_module_57_res), .Z(
        n_xor_module_127_res) );
  DFF_X1 u_reg_module_169__cini_mul_v000_reg ( .D(n_xor_module_127_res), .CK(
        clock_3), .Q(n_reg_module_169_res), .QN() );
  AND2_X1 u_and_module_58_U1 ( .A1(n_reg_module_55_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_58_res) );
  XOR2_X1 u_xor_module_128_U1 ( .A(p_rand_9), .B(n_and_module_58_res), .Z(
        n_xor_module_128_res) );
  DFF_X1 u_reg_module_170__cini_mul_v000_reg ( .D(n_xor_module_128_res), .CK(
        clock_3), .Q(n_reg_module_170_res), .QN() );
  AND2_X1 u_and_module_59_U1 ( .A1(n_reg_module_59_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_59_res) );
  DFF_X1 u_reg_module_171__cini_mul_v000_reg ( .D(n_and_module_59_res), .CK(
        clock_3), .Q(n_reg_module_171_res), .QN() );
  AND2_X1 u_and_module_60_U1 ( .A1(n_reg_module_63_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_60_res) );
  XOR2_X1 u_xor_module_129_U1 ( .A(p_rand_11), .B(n_and_module_60_res), .Z(
        n_xor_module_129_res) );
  DFF_X1 u_reg_module_172__cini_mul_v000_reg ( .D(n_xor_module_129_res), .CK(
        clock_3), .Q(n_reg_module_172_res), .QN() );
  AND2_X1 u_and_module_61_U1 ( .A1(n_reg_module_52_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_61_res) );
  XOR2_X1 u_xor_module_130_U1 ( .A(p_rand_8), .B(n_and_module_61_res), .Z(
        n_xor_module_130_res) );
  DFF_X1 u_reg_module_173__cini_mul_v000_reg ( .D(n_xor_module_130_res), .CK(
        clock_3), .Q(n_reg_module_173_res), .QN() );
  AND2_X1 u_and_module_62_U1 ( .A1(n_reg_module_56_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_62_res) );
  XOR2_X1 u_xor_module_131_U1 ( .A(p_rand_10), .B(n_and_module_62_res), .Z(
        n_xor_module_131_res) );
  DFF_X1 u_reg_module_174__cini_mul_v000_reg ( .D(n_xor_module_131_res), .CK(
        clock_3), .Q(n_reg_module_174_res), .QN() );
  AND2_X1 u_and_module_63_U1 ( .A1(n_reg_module_60_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_63_res) );
  XOR2_X1 u_xor_module_132_U1 ( .A(p_rand_11), .B(n_and_module_63_res), .Z(
        n_xor_module_132_res) );
  DFF_X1 u_reg_module_175__cini_mul_v000_reg ( .D(n_xor_module_132_res), .CK(
        clock_3), .Q(n_reg_module_175_res), .QN() );
  AND2_X1 u_and_module_64_U1 ( .A1(n_reg_module_64_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_64_res) );
  DFF_X1 u_reg_module_176__cini_mul_v000_reg ( .D(n_and_module_64_res), .CK(
        clock_3), .Q(n_reg_module_176_res), .QN() );
  AND2_X1 u_and_module_65_U1 ( .A1(n_reg_module_65_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_65_res) );
  DFF_X1 u_reg_module_177__cini_mul_v000_reg ( .D(n_and_module_65_res), .CK(
        clock_4), .Q(n_reg_module_177_res), .QN() );
  AND2_X1 u_and_module_66_U1 ( .A1(n_reg_module_69_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_66_res) );
  XOR2_X1 u_xor_module_133_U1 ( .A(p_rand_6), .B(n_and_module_66_res), .Z(
        n_xor_module_133_res) );
  DFF_X1 u_reg_module_178__cini_mul_v000_reg ( .D(n_xor_module_133_res), .CK(
        clock_4), .Q(n_reg_module_178_res), .QN() );
  AND2_X1 u_and_module_67_U1 ( .A1(n_reg_module_73_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_67_res) );
  XOR2_X1 u_xor_module_134_U1 ( .A(p_rand_7), .B(n_and_module_67_res), .Z(
        n_xor_module_134_res) );
  DFF_X1 u_reg_module_179__cini_mul_v000_reg ( .D(n_xor_module_134_res), .CK(
        clock_4), .Q(n_reg_module_179_res), .QN() );
  AND2_X1 u_and_module_68_U1 ( .A1(n_reg_module_77_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_68_res) );
  XOR2_X1 u_xor_module_135_U1 ( .A(p_rand_8), .B(n_and_module_68_res), .Z(
        n_xor_module_135_res) );
  DFF_X1 u_reg_module_180__cini_mul_v000_reg ( .D(n_xor_module_135_res), .CK(
        clock_4), .Q(n_reg_module_180_res), .QN() );
  AND2_X1 u_and_module_69_U1 ( .A1(n_reg_module_66_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_69_res) );
  XOR2_X1 u_xor_module_136_U1 ( .A(p_rand_6), .B(n_and_module_69_res), .Z(
        n_xor_module_136_res) );
  DFF_X1 u_reg_module_181__cini_mul_v000_reg ( .D(n_xor_module_136_res), .CK(
        clock_4), .Q(n_reg_module_181_res), .QN() );
  AND2_X1 u_and_module_70_U1 ( .A1(n_reg_module_70_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_70_res) );
  DFF_X1 u_reg_module_182__cini_mul_v000_reg ( .D(n_and_module_70_res), .CK(
        clock_4), .Q(n_reg_module_182_res), .QN() );
  AND2_X1 u_and_module_71_U1 ( .A1(n_reg_module_74_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_71_res) );
  XOR2_X1 u_xor_module_137_U1 ( .A(p_rand_9), .B(n_and_module_71_res), .Z(
        n_xor_module_137_res) );
  DFF_X1 u_reg_module_183__cini_mul_v000_reg ( .D(n_xor_module_137_res), .CK(
        clock_4), .Q(n_reg_module_183_res), .QN() );
  AND2_X1 u_and_module_72_U1 ( .A1(n_reg_module_78_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_72_res) );
  XOR2_X1 u_xor_module_138_U1 ( .A(p_rand_10), .B(n_and_module_72_res), .Z(
        n_xor_module_138_res) );
  DFF_X1 u_reg_module_184__cini_mul_v000_reg ( .D(n_xor_module_138_res), .CK(
        clock_4), .Q(n_reg_module_184_res), .QN() );
  AND2_X1 u_and_module_73_U1 ( .A1(n_reg_module_67_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_73_res) );
  XOR2_X1 u_xor_module_139_U1 ( .A(p_rand_7), .B(n_and_module_73_res), .Z(
        n_xor_module_139_res) );
  DFF_X1 u_reg_module_185__cini_mul_v000_reg ( .D(n_xor_module_139_res), .CK(
        clock_4), .Q(n_reg_module_185_res), .QN() );
  AND2_X1 u_and_module_74_U1 ( .A1(n_reg_module_71_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_74_res) );
  XOR2_X1 u_xor_module_140_U1 ( .A(p_rand_9), .B(n_and_module_74_res), .Z(
        n_xor_module_140_res) );
  DFF_X1 u_reg_module_186__cini_mul_v000_reg ( .D(n_xor_module_140_res), .CK(
        clock_4), .Q(n_reg_module_186_res), .QN() );
  AND2_X1 u_and_module_75_U1 ( .A1(n_reg_module_75_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_75_res) );
  DFF_X1 u_reg_module_187__cini_mul_v000_reg ( .D(n_and_module_75_res), .CK(
        clock_4), .Q(n_reg_module_187_res), .QN() );
  AND2_X1 u_and_module_76_U1 ( .A1(n_reg_module_79_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_76_res) );
  XOR2_X1 u_xor_module_141_U1 ( .A(p_rand_11), .B(n_and_module_76_res), .Z(
        n_xor_module_141_res) );
  DFF_X1 u_reg_module_188__cini_mul_v000_reg ( .D(n_xor_module_141_res), .CK(
        clock_4), .Q(n_reg_module_188_res), .QN() );
  AND2_X1 u_and_module_77_U1 ( .A1(n_reg_module_68_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_77_res) );
  XOR2_X1 u_xor_module_142_U1 ( .A(p_rand_8), .B(n_and_module_77_res), .Z(
        n_xor_module_142_res) );
  DFF_X1 u_reg_module_189__cini_mul_v000_reg ( .D(n_xor_module_142_res), .CK(
        clock_4), .Q(n_reg_module_189_res), .QN() );
  AND2_X1 u_and_module_78_U1 ( .A1(n_reg_module_72_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_78_res) );
  XOR2_X1 u_xor_module_143_U1 ( .A(p_rand_10), .B(n_and_module_78_res), .Z(
        n_xor_module_143_res) );
  DFF_X1 u_reg_module_190__cini_mul_v000_reg ( .D(n_xor_module_143_res), .CK(
        clock_4), .Q(n_reg_module_190_res), .QN() );
  AND2_X1 u_and_module_79_U1 ( .A1(n_reg_module_76_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_79_res) );
  XOR2_X1 u_xor_module_144_U1 ( .A(p_rand_11), .B(n_and_module_79_res), .Z(
        n_xor_module_144_res) );
  DFF_X1 u_reg_module_191__cini_mul_v000_reg ( .D(n_xor_module_144_res), .CK(
        clock_4), .Q(n_reg_module_191_res), .QN() );
  AND2_X1 u_and_module_80_U1 ( .A1(n_reg_module_80_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_80_res) );
  DFF_X1 u_reg_module_192__cini_mul_v000_reg ( .D(n_and_module_80_res), .CK(
        clock_4), .Q(n_reg_module_192_res), .QN() );
  AND2_X1 u_and_module_81_U1 ( .A1(n_reg_module_81_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_81_res) );
  DFF_X1 u_reg_module_193__cini_mul_v000_reg ( .D(n_and_module_81_res), .CK(
        clock_5), .Q(n_reg_module_193_res), .QN() );
  AND2_X1 u_and_module_82_U1 ( .A1(n_reg_module_85_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_82_res) );
  XOR2_X1 u_xor_module_145_U1 ( .A(p_rand_6), .B(n_and_module_82_res), .Z(
        n_xor_module_145_res) );
  DFF_X1 u_reg_module_194__cini_mul_v000_reg ( .D(n_xor_module_145_res), .CK(
        clock_5), .Q(n_reg_module_194_res), .QN() );
  AND2_X1 u_and_module_83_U1 ( .A1(n_reg_module_89_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_83_res) );
  XOR2_X1 u_xor_module_146_U1 ( .A(p_rand_7), .B(n_and_module_83_res), .Z(
        n_xor_module_146_res) );
  DFF_X1 u_reg_module_195__cini_mul_v000_reg ( .D(n_xor_module_146_res), .CK(
        clock_5), .Q(n_reg_module_195_res), .QN() );
  AND2_X1 u_and_module_84_U1 ( .A1(n_reg_module_93_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_84_res) );
  XOR2_X1 u_xor_module_147_U1 ( .A(p_rand_8), .B(n_and_module_84_res), .Z(
        n_xor_module_147_res) );
  DFF_X1 u_reg_module_196__cini_mul_v000_reg ( .D(n_xor_module_147_res), .CK(
        clock_5), .Q(n_reg_module_196_res), .QN() );
  AND2_X1 u_and_module_85_U1 ( .A1(n_reg_module_82_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_85_res) );
  XOR2_X1 u_xor_module_148_U1 ( .A(p_rand_6), .B(n_and_module_85_res), .Z(
        n_xor_module_148_res) );
  DFF_X1 u_reg_module_197__cini_mul_v000_reg ( .D(n_xor_module_148_res), .CK(
        clock_5), .Q(n_reg_module_197_res), .QN() );
  AND2_X1 u_and_module_86_U1 ( .A1(n_reg_module_86_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_86_res) );
  DFF_X1 u_reg_module_198__cini_mul_v000_reg ( .D(n_and_module_86_res), .CK(
        clock_5), .Q(n_reg_module_198_res), .QN() );
  AND2_X1 u_and_module_87_U1 ( .A1(n_reg_module_90_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_87_res) );
  XOR2_X1 u_xor_module_149_U1 ( .A(p_rand_9), .B(n_and_module_87_res), .Z(
        n_xor_module_149_res) );
  DFF_X1 u_reg_module_199__cini_mul_v000_reg ( .D(n_xor_module_149_res), .CK(
        clock_5), .Q(n_reg_module_199_res), .QN() );
  AND2_X1 u_and_module_88_U1 ( .A1(n_reg_module_94_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_88_res) );
  XOR2_X1 u_xor_module_150_U1 ( .A(p_rand_10), .B(n_and_module_88_res), .Z(
        n_xor_module_150_res) );
  DFF_X1 u_reg_module_200__cini_mul_v000_reg ( .D(n_xor_module_150_res), .CK(
        clock_5), .Q(n_reg_module_200_res), .QN() );
  AND2_X1 u_and_module_89_U1 ( .A1(n_reg_module_83_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_89_res) );
  XOR2_X1 u_xor_module_151_U1 ( .A(p_rand_7), .B(n_and_module_89_res), .Z(
        n_xor_module_151_res) );
  DFF_X1 u_reg_module_201__cini_mul_v000_reg ( .D(n_xor_module_151_res), .CK(
        clock_5), .Q(n_reg_module_201_res), .QN() );
  AND2_X1 u_and_module_90_U1 ( .A1(n_reg_module_87_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_90_res) );
  XOR2_X1 u_xor_module_152_U1 ( .A(p_rand_9), .B(n_and_module_90_res), .Z(
        n_xor_module_152_res) );
  DFF_X1 u_reg_module_202__cini_mul_v000_reg ( .D(n_xor_module_152_res), .CK(
        clock_5), .Q(n_reg_module_202_res), .QN() );
  AND2_X1 u_and_module_91_U1 ( .A1(n_reg_module_91_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_91_res) );
  DFF_X1 u_reg_module_203__cini_mul_v000_reg ( .D(n_and_module_91_res), .CK(
        clock_5), .Q(n_reg_module_203_res), .QN() );
  AND2_X1 u_and_module_92_U1 ( .A1(n_reg_module_95_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_92_res) );
  XOR2_X1 u_xor_module_153_U1 ( .A(p_rand_11), .B(n_and_module_92_res), .Z(
        n_xor_module_153_res) );
  DFF_X1 u_reg_module_204__cini_mul_v000_reg ( .D(n_xor_module_153_res), .CK(
        clock_5), .Q(n_reg_module_204_res), .QN() );
  AND2_X1 u_and_module_93_U1 ( .A1(n_reg_module_84_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_93_res) );
  XOR2_X1 u_xor_module_154_U1 ( .A(p_rand_8), .B(n_and_module_93_res), .Z(
        n_xor_module_154_res) );
  DFF_X1 u_reg_module_205__cini_mul_v000_reg ( .D(n_xor_module_154_res), .CK(
        clock_5), .Q(n_reg_module_205_res), .QN() );
  AND2_X1 u_and_module_94_U1 ( .A1(n_reg_module_88_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_94_res) );
  XOR2_X1 u_xor_module_155_U1 ( .A(p_rand_10), .B(n_and_module_94_res), .Z(
        n_xor_module_155_res) );
  DFF_X1 u_reg_module_206__cini_mul_v000_reg ( .D(n_xor_module_155_res), .CK(
        clock_5), .Q(n_reg_module_206_res), .QN() );
  AND2_X1 u_and_module_95_U1 ( .A1(n_reg_module_92_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_95_res) );
  XOR2_X1 u_xor_module_156_U1 ( .A(p_rand_11), .B(n_and_module_95_res), .Z(
        n_xor_module_156_res) );
  DFF_X1 u_reg_module_207__cini_mul_v000_reg ( .D(n_xor_module_156_res), .CK(
        clock_5), .Q(n_reg_module_207_res), .QN() );
  AND2_X1 u_and_module_96_U1 ( .A1(n_reg_module_96_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_96_res) );
  DFF_X1 u_reg_module_208__cini_mul_v000_reg ( .D(n_and_module_96_res), .CK(
        clock_5), .Q(n_reg_module_208_res), .QN() );
  AND2_X1 u_and_module_97_U1 ( .A1(n_reg_module_97_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_97_res) );
  DFF_X1 u_reg_module_209__cini_mul_v000_reg ( .D(n_and_module_97_res), .CK(
        clock_6), .Q(n_reg_module_209_res), .QN() );
  AND2_X1 u_and_module_98_U1 ( .A1(n_reg_module_101_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_98_res) );
  XOR2_X1 u_xor_module_157_U1 ( .A(p_rand_6), .B(n_and_module_98_res), .Z(
        n_xor_module_157_res) );
  DFF_X1 u_reg_module_210__cini_mul_v000_reg ( .D(n_xor_module_157_res), .CK(
        clock_6), .Q(n_reg_module_210_res), .QN() );
  AND2_X1 u_and_module_99_U1 ( .A1(n_reg_module_105_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_99_res) );
  XOR2_X1 u_xor_module_158_U1 ( .A(p_rand_7), .B(n_and_module_99_res), .Z(
        n_xor_module_158_res) );
  DFF_X1 u_reg_module_211__cini_mul_v000_reg ( .D(n_xor_module_158_res), .CK(
        clock_6), .Q(n_reg_module_211_res), .QN() );
  AND2_X1 u_and_module_100_U1 ( .A1(n_reg_module_109_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_100_res) );
  XOR2_X1 u_xor_module_159_U1 ( .A(p_rand_8), .B(n_and_module_100_res), .Z(
        n_xor_module_159_res) );
  DFF_X1 u_reg_module_212__cini_mul_v000_reg ( .D(n_xor_module_159_res), .CK(
        clock_6), .Q(n_reg_module_212_res), .QN() );
  AND2_X1 u_and_module_101_U1 ( .A1(n_reg_module_98_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_101_res) );
  XOR2_X1 u_xor_module_160_U1 ( .A(p_rand_6), .B(n_and_module_101_res), .Z(
        n_xor_module_160_res) );
  DFF_X1 u_reg_module_213__cini_mul_v000_reg ( .D(n_xor_module_160_res), .CK(
        clock_6), .Q(n_reg_module_213_res), .QN() );
  AND2_X1 u_and_module_102_U1 ( .A1(n_reg_module_102_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_102_res) );
  DFF_X1 u_reg_module_214__cini_mul_v000_reg ( .D(n_and_module_102_res), .CK(
        clock_6), .Q(n_reg_module_214_res), .QN() );
  AND2_X1 u_and_module_103_U1 ( .A1(n_reg_module_106_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_103_res) );
  XOR2_X1 u_xor_module_161_U1 ( .A(p_rand_9), .B(n_and_module_103_res), .Z(
        n_xor_module_161_res) );
  DFF_X1 u_reg_module_215__cini_mul_v000_reg ( .D(n_xor_module_161_res), .CK(
        clock_6), .Q(n_reg_module_215_res), .QN() );
  AND2_X1 u_and_module_104_U1 ( .A1(n_reg_module_110_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_104_res) );
  XOR2_X1 u_xor_module_162_U1 ( .A(p_rand_10), .B(n_and_module_104_res), .Z(
        n_xor_module_162_res) );
  DFF_X1 u_reg_module_216__cini_mul_v000_reg ( .D(n_xor_module_162_res), .CK(
        clock_6), .Q(n_reg_module_216_res), .QN() );
  AND2_X1 u_and_module_105_U1 ( .A1(n_reg_module_99_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_105_res) );
  XOR2_X1 u_xor_module_163_U1 ( .A(p_rand_7), .B(n_and_module_105_res), .Z(
        n_xor_module_163_res) );
  DFF_X1 u_reg_module_217__cini_mul_v000_reg ( .D(n_xor_module_163_res), .CK(
        clock_6), .Q(n_reg_module_217_res), .QN() );
  AND2_X1 u_and_module_106_U1 ( .A1(n_reg_module_103_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_106_res) );
  XOR2_X1 u_xor_module_164_U1 ( .A(p_rand_9), .B(n_and_module_106_res), .Z(
        n_xor_module_164_res) );
  DFF_X1 u_reg_module_218__cini_mul_v000_reg ( .D(n_xor_module_164_res), .CK(
        clock_6), .Q(n_reg_module_218_res), .QN() );
  AND2_X1 u_and_module_107_U1 ( .A1(n_reg_module_107_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_107_res) );
  DFF_X1 u_reg_module_219__cini_mul_v000_reg ( .D(n_and_module_107_res), .CK(
        clock_6), .Q(n_reg_module_219_res), .QN() );
  AND2_X1 u_and_module_108_U1 ( .A1(n_reg_module_111_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_108_res) );
  XOR2_X1 u_xor_module_165_U1 ( .A(p_rand_11), .B(n_and_module_108_res), .Z(
        n_xor_module_165_res) );
  DFF_X1 u_reg_module_220__cini_mul_v000_reg ( .D(n_xor_module_165_res), .CK(
        clock_6), .Q(n_reg_module_220_res), .QN() );
  AND2_X1 u_and_module_109_U1 ( .A1(n_reg_module_100_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_109_res) );
  XOR2_X1 u_xor_module_166_U1 ( .A(p_rand_8), .B(n_and_module_109_res), .Z(
        n_xor_module_166_res) );
  DFF_X1 u_reg_module_221__cini_mul_v000_reg ( .D(n_xor_module_166_res), .CK(
        clock_6), .Q(n_reg_module_221_res), .QN() );
  AND2_X1 u_and_module_110_U1 ( .A1(n_reg_module_104_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_110_res) );
  XOR2_X1 u_xor_module_167_U1 ( .A(p_rand_10), .B(n_and_module_110_res), .Z(
        n_xor_module_167_res) );
  DFF_X1 u_reg_module_222__cini_mul_v000_reg ( .D(n_xor_module_167_res), .CK(
        clock_6), .Q(n_reg_module_222_res), .QN() );
  AND2_X1 u_and_module_111_U1 ( .A1(n_reg_module_108_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_111_res) );
  XOR2_X1 u_xor_module_168_U1 ( .A(p_rand_11), .B(n_and_module_111_res), .Z(
        n_xor_module_168_res) );
  DFF_X1 u_reg_module_223__cini_mul_v000_reg ( .D(n_xor_module_168_res), .CK(
        clock_6), .Q(n_reg_module_223_res), .QN() );
  AND2_X1 u_and_module_112_U1 ( .A1(n_reg_module_112_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_112_res) );
  DFF_X1 u_reg_module_224__cini_mul_v000_reg ( .D(n_and_module_112_res), .CK(
        clock_6), .Q(n_reg_module_224_res), .QN() );
  XOR2_X1 u_xor_module_169_U1 ( .A(n_reg_module_114_res), .B(
        n_reg_module_113_res), .Z(n_xor_module_169_res) );
  XOR2_X1 u_xor_module_170_U1 ( .A(n_reg_module_115_res), .B(
        n_xor_module_169_res), .Z(n_xor_module_170_res) );
  XOR2_X1 u_xor_module_171_U1 ( .A(n_reg_module_116_res), .B(
        n_xor_module_170_res), .Z(io_o0_s0_d0) );
  XOR2_X1 u_xor_module_172_U1 ( .A(n_reg_module_117_res), .B(
        n_reg_module_118_res), .Z(n_xor_module_172_res) );
  XOR2_X1 u_xor_module_173_U1 ( .A(n_reg_module_119_res), .B(
        n_xor_module_172_res), .Z(n_xor_module_173_res) );
  XOR2_X1 u_xor_module_174_U1 ( .A(n_reg_module_120_res), .B(
        n_xor_module_173_res), .Z(io_o0_s1_d0) );
  XOR2_X1 u_xor_module_175_U1 ( .A(n_reg_module_121_res), .B(
        n_reg_module_123_res), .Z(n_xor_module_175_res) );
  XOR2_X1 u_xor_module_176_U1 ( .A(n_reg_module_122_res), .B(
        n_xor_module_175_res), .Z(n_xor_module_176_res) );
  XOR2_X1 u_xor_module_177_U1 ( .A(n_reg_module_124_res), .B(
        n_xor_module_176_res), .Z(io_o0_s2_d0) );
  XOR2_X1 u_xor_module_178_U1 ( .A(n_reg_module_125_res), .B(
        n_reg_module_128_res), .Z(n_xor_module_178_res) );
  XOR2_X1 u_xor_module_179_U1 ( .A(n_reg_module_126_res), .B(
        n_xor_module_178_res), .Z(n_xor_module_179_res) );
  XOR2_X1 u_xor_module_180_U1 ( .A(n_reg_module_127_res), .B(
        n_xor_module_179_res), .Z(io_o0_s3_d0) );
  XOR2_X1 u_xor_module_181_U1 ( .A(n_reg_module_130_res), .B(
        n_reg_module_129_res), .Z(n_xor_module_181_res) );
  XOR2_X1 u_xor_module_182_U1 ( .A(n_reg_module_131_res), .B(
        n_xor_module_181_res), .Z(n_xor_module_182_res) );
  XOR2_X1 u_xor_module_183_U1 ( .A(n_reg_module_132_res), .B(
        n_xor_module_182_res), .Z(io_o0_s0_d1) );
  XOR2_X1 u_xor_module_184_U1 ( .A(n_reg_module_133_res), .B(
        n_reg_module_134_res), .Z(n_xor_module_184_res) );
  XOR2_X1 u_xor_module_185_U1 ( .A(n_reg_module_135_res), .B(
        n_xor_module_184_res), .Z(n_xor_module_185_res) );
  XOR2_X1 u_xor_module_186_U1 ( .A(n_reg_module_136_res), .B(
        n_xor_module_185_res), .Z(io_o0_s1_d1) );
  XOR2_X1 u_xor_module_187_U1 ( .A(n_reg_module_137_res), .B(
        n_reg_module_139_res), .Z(n_xor_module_187_res) );
  XOR2_X1 u_xor_module_188_U1 ( .A(n_reg_module_138_res), .B(
        n_xor_module_187_res), .Z(n_xor_module_188_res) );
  XOR2_X1 u_xor_module_189_U1 ( .A(n_reg_module_140_res), .B(
        n_xor_module_188_res), .Z(io_o0_s2_d1) );
  XOR2_X1 u_xor_module_190_U1 ( .A(n_reg_module_141_res), .B(
        n_reg_module_144_res), .Z(n_xor_module_190_res) );
  XOR2_X1 u_xor_module_191_U1 ( .A(n_reg_module_142_res), .B(
        n_xor_module_190_res), .Z(n_xor_module_191_res) );
  XOR2_X1 u_xor_module_192_U1 ( .A(n_reg_module_143_res), .B(
        n_xor_module_191_res), .Z(io_o0_s3_d1) );
  XOR2_X1 u_xor_module_193_U1 ( .A(n_reg_module_146_res), .B(
        n_reg_module_145_res), .Z(n_xor_module_193_res) );
  XOR2_X1 u_xor_module_194_U1 ( .A(n_reg_module_147_res), .B(
        n_xor_module_193_res), .Z(n_xor_module_194_res) );
  XOR2_X1 u_xor_module_195_U1 ( .A(n_reg_module_148_res), .B(
        n_xor_module_194_res), .Z(io_o0_s0_d2) );
  XOR2_X1 u_xor_module_196_U1 ( .A(n_reg_module_149_res), .B(
        n_reg_module_150_res), .Z(n_xor_module_196_res) );
  XOR2_X1 u_xor_module_197_U1 ( .A(n_reg_module_151_res), .B(
        n_xor_module_196_res), .Z(n_xor_module_197_res) );
  XOR2_X1 u_xor_module_198_U1 ( .A(n_reg_module_152_res), .B(
        n_xor_module_197_res), .Z(io_o0_s1_d2) );
  XOR2_X1 u_xor_module_199_U1 ( .A(n_reg_module_153_res), .B(
        n_reg_module_155_res), .Z(n_xor_module_199_res) );
  XOR2_X1 u_xor_module_200_U1 ( .A(n_reg_module_154_res), .B(
        n_xor_module_199_res), .Z(n_xor_module_200_res) );
  XOR2_X1 u_xor_module_201_U1 ( .A(n_reg_module_156_res), .B(
        n_xor_module_200_res), .Z(io_o0_s2_d2) );
  XOR2_X1 u_xor_module_202_U1 ( .A(n_reg_module_157_res), .B(
        n_reg_module_160_res), .Z(n_xor_module_202_res) );
  XOR2_X1 u_xor_module_203_U1 ( .A(n_reg_module_158_res), .B(
        n_xor_module_202_res), .Z(n_xor_module_203_res) );
  XOR2_X1 u_xor_module_204_U1 ( .A(n_reg_module_159_res), .B(
        n_xor_module_203_res), .Z(io_o0_s3_d2) );
  XOR2_X1 u_xor_module_205_U1 ( .A(n_reg_module_162_res), .B(
        n_reg_module_161_res), .Z(n_xor_module_205_res) );
  XOR2_X1 u_xor_module_206_U1 ( .A(n_reg_module_163_res), .B(
        n_xor_module_205_res), .Z(n_xor_module_206_res) );
  XOR2_X1 u_xor_module_207_U1 ( .A(n_reg_module_164_res), .B(
        n_xor_module_206_res), .Z(io_o0_s0_d3) );
  XOR2_X1 u_xor_module_208_U1 ( .A(n_reg_module_165_res), .B(
        n_reg_module_166_res), .Z(n_xor_module_208_res) );
  XOR2_X1 u_xor_module_209_U1 ( .A(n_reg_module_167_res), .B(
        n_xor_module_208_res), .Z(n_xor_module_209_res) );
  XOR2_X1 u_xor_module_210_U1 ( .A(n_reg_module_168_res), .B(
        n_xor_module_209_res), .Z(io_o0_s1_d3) );
  XOR2_X1 u_xor_module_211_U1 ( .A(n_reg_module_169_res), .B(
        n_reg_module_171_res), .Z(n_xor_module_211_res) );
  XOR2_X1 u_xor_module_212_U1 ( .A(n_reg_module_170_res), .B(
        n_xor_module_211_res), .Z(n_xor_module_212_res) );
  XOR2_X1 u_xor_module_213_U1 ( .A(n_reg_module_172_res), .B(
        n_xor_module_212_res), .Z(io_o0_s2_d3) );
  XOR2_X1 u_xor_module_214_U1 ( .A(n_reg_module_173_res), .B(
        n_reg_module_176_res), .Z(n_xor_module_214_res) );
  XOR2_X1 u_xor_module_215_U1 ( .A(n_reg_module_174_res), .B(
        n_xor_module_214_res), .Z(n_xor_module_215_res) );
  XOR2_X1 u_xor_module_216_U1 ( .A(n_reg_module_175_res), .B(
        n_xor_module_215_res), .Z(io_o0_s3_d3) );
  XOR2_X1 u_xor_module_217_U1 ( .A(n_reg_module_178_res), .B(
        n_reg_module_177_res), .Z(n_xor_module_217_res) );
  XOR2_X1 u_xor_module_218_U1 ( .A(n_reg_module_179_res), .B(
        n_xor_module_217_res), .Z(n_xor_module_218_res) );
  XOR2_X1 u_xor_module_219_U1 ( .A(n_reg_module_180_res), .B(
        n_xor_module_218_res), .Z(io_o0_s0_d4) );
  XOR2_X1 u_xor_module_220_U1 ( .A(n_reg_module_181_res), .B(
        n_reg_module_182_res), .Z(n_xor_module_220_res) );
  XOR2_X1 u_xor_module_221_U1 ( .A(n_reg_module_183_res), .B(
        n_xor_module_220_res), .Z(n_xor_module_221_res) );
  XOR2_X1 u_xor_module_222_U1 ( .A(n_reg_module_184_res), .B(
        n_xor_module_221_res), .Z(io_o0_s1_d4) );
  XOR2_X1 u_xor_module_223_U1 ( .A(n_reg_module_185_res), .B(
        n_reg_module_187_res), .Z(n_xor_module_223_res) );
  XOR2_X1 u_xor_module_224_U1 ( .A(n_reg_module_186_res), .B(
        n_xor_module_223_res), .Z(n_xor_module_224_res) );
  XOR2_X1 u_xor_module_225_U1 ( .A(n_reg_module_188_res), .B(
        n_xor_module_224_res), .Z(io_o0_s2_d4) );
  XOR2_X1 u_xor_module_226_U1 ( .A(n_reg_module_189_res), .B(
        n_reg_module_192_res), .Z(n_xor_module_226_res) );
  XOR2_X1 u_xor_module_227_U1 ( .A(n_reg_module_190_res), .B(
        n_xor_module_226_res), .Z(n_xor_module_227_res) );
  XOR2_X1 u_xor_module_228_U1 ( .A(n_reg_module_191_res), .B(
        n_xor_module_227_res), .Z(io_o0_s3_d4) );
  XOR2_X1 u_xor_module_229_U1 ( .A(n_reg_module_194_res), .B(
        n_reg_module_193_res), .Z(n_xor_module_229_res) );
  XOR2_X1 u_xor_module_230_U1 ( .A(n_reg_module_195_res), .B(
        n_xor_module_229_res), .Z(n_xor_module_230_res) );
  XOR2_X1 u_xor_module_231_U1 ( .A(n_reg_module_196_res), .B(
        n_xor_module_230_res), .Z(io_o0_s0_d5) );
  XOR2_X1 u_xor_module_232_U1 ( .A(n_reg_module_197_res), .B(
        n_reg_module_198_res), .Z(n_xor_module_232_res) );
  XOR2_X1 u_xor_module_233_U1 ( .A(n_reg_module_199_res), .B(
        n_xor_module_232_res), .Z(n_xor_module_233_res) );
  XOR2_X1 u_xor_module_234_U1 ( .A(n_reg_module_200_res), .B(
        n_xor_module_233_res), .Z(io_o0_s1_d5) );
  XOR2_X1 u_xor_module_235_U1 ( .A(n_reg_module_201_res), .B(
        n_reg_module_203_res), .Z(n_xor_module_235_res) );
  XOR2_X1 u_xor_module_236_U1 ( .A(n_reg_module_202_res), .B(
        n_xor_module_235_res), .Z(n_xor_module_236_res) );
  XOR2_X1 u_xor_module_237_U1 ( .A(n_reg_module_204_res), .B(
        n_xor_module_236_res), .Z(io_o0_s2_d5) );
  XOR2_X1 u_xor_module_238_U1 ( .A(n_reg_module_205_res), .B(
        n_reg_module_208_res), .Z(n_xor_module_238_res) );
  XOR2_X1 u_xor_module_239_U1 ( .A(n_reg_module_206_res), .B(
        n_xor_module_238_res), .Z(n_xor_module_239_res) );
  XOR2_X1 u_xor_module_240_U1 ( .A(n_reg_module_207_res), .B(
        n_xor_module_239_res), .Z(io_o0_s3_d5) );
  XOR2_X1 u_xor_module_241_U1 ( .A(n_reg_module_210_res), .B(
        n_reg_module_209_res), .Z(n_xor_module_241_res) );
  XOR2_X1 u_xor_module_242_U1 ( .A(n_reg_module_211_res), .B(
        n_xor_module_241_res), .Z(n_xor_module_242_res) );
  XOR2_X1 u_xor_module_243_U1 ( .A(n_reg_module_212_res), .B(
        n_xor_module_242_res), .Z(io_o0_s0_d6) );
  XOR2_X1 u_xor_module_244_U1 ( .A(n_reg_module_213_res), .B(
        n_reg_module_214_res), .Z(n_xor_module_244_res) );
  XOR2_X1 u_xor_module_245_U1 ( .A(n_reg_module_215_res), .B(
        n_xor_module_244_res), .Z(n_xor_module_245_res) );
  XOR2_X1 u_xor_module_246_U1 ( .A(n_reg_module_216_res), .B(
        n_xor_module_245_res), .Z(io_o0_s1_d6) );
  XOR2_X1 u_xor_module_247_U1 ( .A(n_reg_module_217_res), .B(
        n_reg_module_219_res), .Z(n_xor_module_247_res) );
  XOR2_X1 u_xor_module_248_U1 ( .A(n_reg_module_218_res), .B(
        n_xor_module_247_res), .Z(n_xor_module_248_res) );
  XOR2_X1 u_xor_module_249_U1 ( .A(n_reg_module_220_res), .B(
        n_xor_module_248_res), .Z(io_o0_s2_d6) );
  XOR2_X1 u_xor_module_250_U1 ( .A(n_reg_module_221_res), .B(
        n_reg_module_224_res), .Z(n_xor_module_250_res) );
  XOR2_X1 u_xor_module_251_U1 ( .A(n_reg_module_222_res), .B(
        n_xor_module_250_res), .Z(n_xor_module_251_res) );
  XOR2_X1 u_xor_module_252_U1 ( .A(n_reg_module_223_res), .B(
        n_xor_module_251_res), .Z(io_o0_s3_d6) );
endmodule

