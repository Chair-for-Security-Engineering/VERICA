
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i0_s5, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, 
        io_i1_s5, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, 
        p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, 
        p_rand_12, p_rand_13, p_rand_14, io_o0_s0, io_o0_s1, io_o0_s2, 
        io_o0_s3, io_o0_s4, io_o0_s5 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i0_s5, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, io_i1_s5,
         p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6,
         p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12,
         p_rand_13, p_rand_14;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5;
  wire   n_hpc2_0_n207, n_hpc2_0_n206, n_hpc2_0_n205, n_hpc2_0_n204,
         n_hpc2_0_n203, n_hpc2_0_n202, n_hpc2_0_n201, n_hpc2_0_n200,
         n_hpc2_0_n199, n_hpc2_0_n198, n_hpc2_0_n197, n_hpc2_0_n196,
         n_hpc2_0_n195, n_hpc2_0_n194, n_hpc2_0_n193, n_hpc2_0_n192,
         n_hpc2_0_n191, n_hpc2_0_n190, n_hpc2_0_n189, n_hpc2_0_n188,
         n_hpc2_0_n187, n_hpc2_0_n186, n_hpc2_0_n185, n_hpc2_0_n184,
         n_hpc2_0_n183, n_hpc2_0_n182, n_hpc2_0_n181, n_hpc2_0_n180,
         n_hpc2_0_n179, n_hpc2_0_n178, n_hpc2_0_n177, n_hpc2_0_n176,
         n_hpc2_0_n175, n_hpc2_0_n174, n_hpc2_0_n173, n_hpc2_0_n172,
         n_hpc2_0_n171, n_hpc2_0_n170, n_hpc2_0_n169, n_hpc2_0_n168,
         n_hpc2_0_n167, n_hpc2_0_n166, n_hpc2_0_n165, n_hpc2_0_n164,
         n_hpc2_0_n163, n_hpc2_0_n162, n_hpc2_0_n161, n_hpc2_0_n160,
         n_hpc2_0_n159, n_hpc2_0_n158, n_hpc2_0_n157, n_hpc2_0_n156,
         n_hpc2_0_n155, n_hpc2_0_n154, n_hpc2_0_n153, n_hpc2_0_n152,
         n_hpc2_0_n151, n_hpc2_0_n150, n_hpc2_0_n149, n_hpc2_0_n148,
         n_hpc2_0_n147, n_hpc2_0_n146, n_hpc2_0_n145, n_hpc2_0_n144,
         n_hpc2_0_n143, n_hpc2_0_n142, n_hpc2_0_n141, n_hpc2_0_n140,
         n_hpc2_0_n139, n_hpc2_0_n138, n_hpc2_0_n137, n_hpc2_0_n136,
         n_hpc2_0_n135, n_hpc2_0_n134, n_hpc2_0_n133, n_hpc2_0_n132,
         n_hpc2_0_n131, n_hpc2_0_n130, n_hpc2_0_n129, n_hpc2_0_n128,
         n_hpc2_0_n127, n_hpc2_0_n126, n_hpc2_0_n125, n_hpc2_0_n124,
         n_hpc2_0_n123, n_hpc2_0_n122, n_hpc2_0_n121, n_hpc2_0_n120,
         n_hpc2_0_n119, n_hpc2_0_n118, n_hpc2_0_n117, n_hpc2_0_n116,
         n_hpc2_0_n115, n_hpc2_0_n114, n_hpc2_0_n113, n_hpc2_0_n112,
         n_hpc2_0_n111, n_hpc2_0_n110, n_hpc2_0_n109, n_hpc2_0_n108,
         n_hpc2_0_n107, n_hpc2_0_n106, n_hpc2_0_n105, n_hpc2_0_n104,
         n_hpc2_0_n103, n_hpc2_0_n102, n_hpc2_0_n101, n_hpc2_0_n100,
         n_hpc2_0_n99, n_hpc2_0_n98, n_hpc2_0_n97, n_hpc2_0_n96, n_hpc2_0_n95,
         n_hpc2_0_n94, n_hpc2_0_n93, n_hpc2_0_n92, n_hpc2_0_n91, n_hpc2_0_n90,
         n_hpc2_0_n89, n_hpc2_0_n88, n_hpc2_0_n87, n_hpc2_0_n86, n_hpc2_0_n85,
         n_hpc2_0_n84, n_hpc2_0_n83, n_hpc2_0_n82, n_hpc2_0_n81, n_hpc2_0_n80,
         n_hpc2_0_n79, n_hpc2_0_n78, n_hpc2_0_n77, n_hpc2_0_n76, n_hpc2_0_n75,
         n_hpc2_0_n74, n_hpc2_0_n73, n_hpc2_0_n72, n_hpc2_0_n71, n_hpc2_0_n70,
         n_hpc2_0_n69, n_hpc2_0_n68, n_hpc2_0_n67, n_hpc2_0_n66, n_hpc2_0_n65,
         n_hpc2_0_n64, n_hpc2_0_n63, n_hpc2_0_n62, n_hpc2_0_n61, n_hpc2_0_n60,
         n_hpc2_0_n59, n_hpc2_0_n58, n_hpc2_0_n57, n_hpc2_0_n56, n_hpc2_0_n55,
         n_hpc2_0_n54, n_hpc2_0_n53, n_hpc2_0_n52, n_hpc2_0_n51, n_hpc2_0_n50,
         n_hpc2_0_n49, n_hpc2_0_n48, n_hpc2_0_n47, n_hpc2_0_n46, n_hpc2_0_n45,
         n_hpc2_0_n44, n_hpc2_0_n43, n_hpc2_0_n42, n_hpc2_0_n41, n_hpc2_0_n40,
         n_hpc2_0_n39, n_hpc2_0_n38, n_hpc2_0_n37, n_hpc2_0_n36, n_hpc2_0_n35,
         n_hpc2_0_n34, n_hpc2_0_n33, n_hpc2_0_n32, n_hpc2_0_n31, n_hpc2_0_n30,
         n_hpc2_0_n29, n_hpc2_0_n28, n_hpc2_0_n27, n_hpc2_0_n26, n_hpc2_0_n25,
         n_hpc2_0_n24, n_hpc2_0_n23, n_hpc2_0_n22, n_hpc2_0_n21, n_hpc2_0_n20,
         n_hpc2_0_n19, n_hpc2_0_n18, n_hpc2_0_n17, n_hpc2_0_n16, n_hpc2_0_n15,
         n_hpc2_0_n14, n_hpc2_0_n13, n_hpc2_0_n12, n_hpc2_0_n11, n_hpc2_0_n10,
         n_hpc2_0_n9, n_hpc2_0_n8, n_hpc2_0_n7, n_hpc2_0_n6, n_hpc2_0_n5,
         n_hpc2_0_n4, n_hpc2_0_n3, n_hpc2_0_n2, n_hpc2_0_n1, n_hpc2_0_N101,
         n_hpc2_0_N100, n_hpc2_0_N99, n_hpc2_0_N98, n_hpc2_0_N97, n_hpc2_0_N96,
         n_hpc2_0_N95, n_hpc2_0_N94, n_hpc2_0_N93, n_hpc2_0_N92, n_hpc2_0_N91,
         n_hpc2_0_N90, n_hpc2_0_N89, n_hpc2_0_N88, n_hpc2_0_N87, n_hpc2_0_N86,
         n_hpc2_0_N85, n_hpc2_0_N84, n_hpc2_0_N83, n_hpc2_0_N82, n_hpc2_0_N81,
         n_hpc2_0_N80, n_hpc2_0_N79, n_hpc2_0_N78, n_hpc2_0_N77, n_hpc2_0_N76,
         n_hpc2_0_N75, n_hpc2_0_N74, n_hpc2_0_N73, n_hpc2_0_N72, n_hpc2_0_N71,
         n_hpc2_0_N70, n_hpc2_0_N69, n_hpc2_0_N68, n_hpc2_0_N67, n_hpc2_0_N66,
         n_hpc2_0_N65, n_hpc2_0_N64, n_hpc2_0_N63, n_hpc2_0_N62, n_hpc2_0_N61,
         n_hpc2_0_N60, n_hpc2_0_N59, n_hpc2_0_N58, n_hpc2_0_N57, n_hpc2_0_N56,
         n_hpc2_0_N55, n_hpc2_0_N54, n_hpc2_0_N53, n_hpc2_0_N52, n_hpc2_0_N51,
         n_hpc2_0_N50, n_hpc2_0_N49, n_hpc2_0_N48, n_hpc2_0_N47, n_hpc2_0_N46,
         n_hpc2_0_N45, n_hpc2_0_N44, n_hpc2_0_N43, n_hpc2_0_N42, n_hpc2_0_N41,
         n_hpc2_0_N40, n_hpc2_0_N39, n_hpc2_0_N38, n_hpc2_0_N37, n_hpc2_0_N36,
         n_hpc2_0_N35, n_hpc2_0_N34, n_hpc2_0_N33, n_hpc2_0_N32, n_hpc2_0_N31,
         n_hpc2_0_N30, n_hpc2_0_N29, n_hpc2_0_N28, n_hpc2_0_N27, n_hpc2_0_N26,
         n_hpc2_0_N25, n_hpc2_0_N24, n_hpc2_0_N23, n_hpc2_0_N22, n_hpc2_0_N21,
         n_hpc2_0_N20, n_hpc2_0_N19, n_hpc2_0_N18, n_hpc2_0_N17, n_hpc2_0_N16,
         n_hpc2_0_N15, n_hpc2_0_N14, n_hpc2_0_N13, n_hpc2_0_N12, n_hpc2_0_N11,
         n_hpc2_0_N10, n_hpc2_0_N9, n_hpc2_0_N8, n_hpc2_0_N7, n_hpc2_0_N6,
         n_hpc2_0__hpc_u54, n_hpc2_0__hpc_u45, n_hpc2_0__hpc_u35,
         n_hpc2_0__hpc_u25, n_hpc2_0__hpc_u15, n_hpc2_0__hpc_u05;

  NOR2_X1 u_hpc2_0_U164 ( .A1(n_hpc2_0_n207), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N10) );
  XOR2_X1 u_hpc2_0_U163 ( .A(io_i1_s3), .B(p_rand_13), .Z(n_hpc2_0_N100) );
  XOR2_X1 u_hpc2_0_U162 ( .A(io_i1_s4), .B(p_rand_14), .Z(n_hpc2_0_N101) );
  NOR2_X1 u_hpc2_0_U161 ( .A1(n_hpc2_0_n206), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N11) );
  NOR2_X1 u_hpc2_0_U160 ( .A1(n_hpc2_0_n205), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N12) );
  NOR2_X1 u_hpc2_0_U159 ( .A1(n_hpc2_0_n204), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N13) );
  NOR2_X1 u_hpc2_0_U158 ( .A1(n_hpc2_0_n203), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N14) );
  NOR2_X1 u_hpc2_0_U157 ( .A1(n_hpc2_0_n202), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N15) );
  NOR2_X1 u_hpc2_0_U156 ( .A1(n_hpc2_0_n201), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N16) );
  NOR2_X1 u_hpc2_0_U155 ( .A1(n_hpc2_0_n200), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N17) );
  NOR2_X1 u_hpc2_0_U154 ( .A1(n_hpc2_0_n199), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N18) );
  NOR2_X1 u_hpc2_0_U153 ( .A1(n_hpc2_0_n198), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N19) );
  NOR2_X1 u_hpc2_0_U152 ( .A1(n_hpc2_0_n197), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N20) );
  NOR2_X1 u_hpc2_0_U151 ( .A1(n_hpc2_0_n196), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N21) );
  NOR2_X1 u_hpc2_0_U150 ( .A1(n_hpc2_0_n195), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N22) );
  NOR2_X1 u_hpc2_0_U149 ( .A1(n_hpc2_0_n194), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N23) );
  NOR2_X1 u_hpc2_0_U148 ( .A1(n_hpc2_0_n193), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N24) );
  NOR2_X1 u_hpc2_0_U147 ( .A1(n_hpc2_0_n192), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N25) );
  NOR2_X1 u_hpc2_0_U146 ( .A1(n_hpc2_0_n191), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N26) );
  NOR2_X1 u_hpc2_0_U145 ( .A1(n_hpc2_0_n190), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N27) );
  NOR2_X1 u_hpc2_0_U144 ( .A1(n_hpc2_0_n189), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N28) );
  NOR2_X1 u_hpc2_0_U143 ( .A1(n_hpc2_0_n188), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N29) );
  NOR2_X1 u_hpc2_0_U142 ( .A1(n_hpc2_0_n187), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N30) );
  NOR2_X1 u_hpc2_0_U141 ( .A1(n_hpc2_0_n186), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N31) );
  NOR2_X1 u_hpc2_0_U140 ( .A1(n_hpc2_0_n185), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N32) );
  NOR2_X1 u_hpc2_0_U139 ( .A1(n_hpc2_0_n184), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N33) );
  NOR2_X1 u_hpc2_0_U138 ( .A1(n_hpc2_0_n183), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N34) );
  NOR2_X1 u_hpc2_0_U137 ( .A1(n_hpc2_0_n182), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N35) );
  NOR2_X1 u_hpc2_0_U136 ( .A1(n_hpc2_0_n181), .A2(n_hpc2_0_n12), .ZN(
        n_hpc2_0_N36) );
  NOR2_X1 u_hpc2_0_U135 ( .A1(n_hpc2_0_n180), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N37) );
  NOR2_X1 u_hpc2_0_U134 ( .A1(n_hpc2_0_n179), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N38) );
  NOR2_X1 u_hpc2_0_U133 ( .A1(n_hpc2_0_n178), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N39) );
  NOR2_X1 u_hpc2_0_U132 ( .A1(n_hpc2_0_n177), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N40) );
  NOR2_X1 u_hpc2_0_U131 ( .A1(n_hpc2_0_n176), .A2(n_hpc2_0_n11), .ZN(
        n_hpc2_0_N41) );
  NOR2_X1 u_hpc2_0_U130 ( .A1(n_hpc2_0_n174), .A2(n_hpc2_0_n175), .ZN(
        n_hpc2_0_N42) );
  NOR2_X1 u_hpc2_0_U129 ( .A1(n_hpc2_0_n172), .A2(n_hpc2_0_n173), .ZN(
        n_hpc2_0_N43) );
  NOR2_X1 u_hpc2_0_U128 ( .A1(n_hpc2_0_n170), .A2(n_hpc2_0_n171), .ZN(
        n_hpc2_0_N44) );
  NOR2_X1 u_hpc2_0_U127 ( .A1(n_hpc2_0_n168), .A2(n_hpc2_0_n169), .ZN(
        n_hpc2_0_N45) );
  NOR2_X1 u_hpc2_0_U126 ( .A1(n_hpc2_0_n166), .A2(n_hpc2_0_n167), .ZN(
        n_hpc2_0_N46) );
  NOR2_X1 u_hpc2_0_U125 ( .A1(n_hpc2_0_n174), .A2(n_hpc2_0_n165), .ZN(
        n_hpc2_0_N47) );
  NOR2_X1 u_hpc2_0_U124 ( .A1(n_hpc2_0_n163), .A2(n_hpc2_0_n164), .ZN(
        n_hpc2_0_N48) );
  NOR2_X1 u_hpc2_0_U123 ( .A1(n_hpc2_0_n161), .A2(n_hpc2_0_n162), .ZN(
        n_hpc2_0_N49) );
  NOR2_X1 u_hpc2_0_U122 ( .A1(n_hpc2_0_n159), .A2(n_hpc2_0_n160), .ZN(
        n_hpc2_0_N50) );
  NOR2_X1 u_hpc2_0_U121 ( .A1(n_hpc2_0_n157), .A2(n_hpc2_0_n158), .ZN(
        n_hpc2_0_N51) );
  NOR2_X1 u_hpc2_0_U120 ( .A1(n_hpc2_0_n172), .A2(n_hpc2_0_n156), .ZN(
        n_hpc2_0_N52) );
  NOR2_X1 u_hpc2_0_U119 ( .A1(n_hpc2_0_n163), .A2(n_hpc2_0_n155), .ZN(
        n_hpc2_0_N53) );
  NOR2_X1 u_hpc2_0_U118 ( .A1(n_hpc2_0_n153), .A2(n_hpc2_0_n154), .ZN(
        n_hpc2_0_N54) );
  NOR2_X1 u_hpc2_0_U117 ( .A1(n_hpc2_0_n151), .A2(n_hpc2_0_n152), .ZN(
        n_hpc2_0_N55) );
  NOR2_X1 u_hpc2_0_U116 ( .A1(n_hpc2_0_n149), .A2(n_hpc2_0_n150), .ZN(
        n_hpc2_0_N56) );
  NOR2_X1 u_hpc2_0_U115 ( .A1(n_hpc2_0_n170), .A2(n_hpc2_0_n148), .ZN(
        n_hpc2_0_N57) );
  NOR2_X1 u_hpc2_0_U114 ( .A1(n_hpc2_0_n161), .A2(n_hpc2_0_n147), .ZN(
        n_hpc2_0_N58) );
  NOR2_X1 u_hpc2_0_U113 ( .A1(n_hpc2_0_n153), .A2(n_hpc2_0_n146), .ZN(
        n_hpc2_0_N59) );
  NOR2_X1 u_hpc2_0_U112 ( .A1(n_hpc2_0_n145), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N6) );
  NOR2_X1 u_hpc2_0_U111 ( .A1(n_hpc2_0_n143), .A2(n_hpc2_0_n144), .ZN(
        n_hpc2_0_N60) );
  NOR2_X1 u_hpc2_0_U110 ( .A1(n_hpc2_0_n141), .A2(n_hpc2_0_n142), .ZN(
        n_hpc2_0_N61) );
  NOR2_X1 u_hpc2_0_U109 ( .A1(n_hpc2_0_n168), .A2(n_hpc2_0_n140), .ZN(
        n_hpc2_0_N62) );
  NOR2_X1 u_hpc2_0_U108 ( .A1(n_hpc2_0_n159), .A2(n_hpc2_0_n139), .ZN(
        n_hpc2_0_N63) );
  NOR2_X1 u_hpc2_0_U107 ( .A1(n_hpc2_0_n151), .A2(n_hpc2_0_n138), .ZN(
        n_hpc2_0_N64) );
  NOR2_X1 u_hpc2_0_U106 ( .A1(n_hpc2_0_n143), .A2(n_hpc2_0_n137), .ZN(
        n_hpc2_0_N65) );
  NOR2_X1 u_hpc2_0_U105 ( .A1(n_hpc2_0_n135), .A2(n_hpc2_0_n136), .ZN(
        n_hpc2_0_N66) );
  NOR2_X1 u_hpc2_0_U104 ( .A1(n_hpc2_0_n166), .A2(n_hpc2_0_n134), .ZN(
        n_hpc2_0_N67) );
  NOR2_X1 u_hpc2_0_U103 ( .A1(n_hpc2_0_n157), .A2(n_hpc2_0_n133), .ZN(
        n_hpc2_0_N68) );
  NOR2_X1 u_hpc2_0_U102 ( .A1(n_hpc2_0_n149), .A2(n_hpc2_0_n132), .ZN(
        n_hpc2_0_N69) );
  NOR2_X1 u_hpc2_0_U101 ( .A1(n_hpc2_0_n131), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N7) );
  NOR2_X1 u_hpc2_0_U100 ( .A1(n_hpc2_0_n141), .A2(n_hpc2_0_n130), .ZN(
        n_hpc2_0_N70) );
  NOR2_X1 u_hpc2_0_U99 ( .A1(n_hpc2_0_n135), .A2(n_hpc2_0_n129), .ZN(
        n_hpc2_0_N71) );
  XOR2_X1 u_hpc2_0_U98 ( .A(io_i1_s1), .B(p_rand_0), .Z(n_hpc2_0_N72) );
  XOR2_X1 u_hpc2_0_U97 ( .A(io_i1_s2), .B(p_rand_1), .Z(n_hpc2_0_N73) );
  XOR2_X1 u_hpc2_0_U96 ( .A(io_i1_s3), .B(p_rand_2), .Z(n_hpc2_0_N74) );
  XOR2_X1 u_hpc2_0_U95 ( .A(io_i1_s4), .B(p_rand_3), .Z(n_hpc2_0_N75) );
  XOR2_X1 u_hpc2_0_U94 ( .A(io_i1_s5), .B(p_rand_4), .Z(n_hpc2_0_N76) );
  XOR2_X1 u_hpc2_0_U93 ( .A(io_i1_s0), .B(p_rand_0), .Z(n_hpc2_0_N77) );
  XOR2_X1 u_hpc2_0_U92 ( .A(io_i1_s2), .B(p_rand_5), .Z(n_hpc2_0_N78) );
  XOR2_X1 u_hpc2_0_U91 ( .A(io_i1_s3), .B(p_rand_6), .Z(n_hpc2_0_N79) );
  NOR2_X1 u_hpc2_0_U90 ( .A1(n_hpc2_0_n128), .A2(n_hpc2_0_n8), .ZN(n_hpc2_0_N8) );
  XOR2_X1 u_hpc2_0_U89 ( .A(io_i1_s4), .B(p_rand_7), .Z(n_hpc2_0_N80) );
  XOR2_X1 u_hpc2_0_U88 ( .A(io_i1_s5), .B(p_rand_8), .Z(n_hpc2_0_N81) );
  XOR2_X1 u_hpc2_0_U87 ( .A(io_i1_s0), .B(p_rand_1), .Z(n_hpc2_0_N82) );
  XOR2_X1 u_hpc2_0_U86 ( .A(io_i1_s1), .B(p_rand_5), .Z(n_hpc2_0_N83) );
  XOR2_X1 u_hpc2_0_U85 ( .A(io_i1_s3), .B(p_rand_9), .Z(n_hpc2_0_N84) );
  XOR2_X1 u_hpc2_0_U84 ( .A(io_i1_s4), .B(p_rand_10), .Z(n_hpc2_0_N85) );
  XOR2_X1 u_hpc2_0_U83 ( .A(io_i1_s5), .B(p_rand_11), .Z(n_hpc2_0_N86) );
  XOR2_X1 u_hpc2_0_U82 ( .A(io_i1_s0), .B(p_rand_2), .Z(n_hpc2_0_N87) );
  XOR2_X1 u_hpc2_0_U81 ( .A(io_i1_s1), .B(p_rand_6), .Z(n_hpc2_0_N88) );
  XOR2_X1 u_hpc2_0_U80 ( .A(io_i1_s2), .B(p_rand_9), .Z(n_hpc2_0_N89) );
  NOR2_X1 u_hpc2_0_U79 ( .A1(n_hpc2_0_n127), .A2(n_hpc2_0_n7), .ZN(n_hpc2_0_N9) );
  XOR2_X1 u_hpc2_0_U78 ( .A(io_i1_s4), .B(p_rand_12), .Z(n_hpc2_0_N90) );
  XOR2_X1 u_hpc2_0_U77 ( .A(io_i1_s5), .B(p_rand_13), .Z(n_hpc2_0_N91) );
  XOR2_X1 u_hpc2_0_U76 ( .A(io_i1_s0), .B(p_rand_3), .Z(n_hpc2_0_N92) );
  XOR2_X1 u_hpc2_0_U75 ( .A(io_i1_s1), .B(p_rand_7), .Z(n_hpc2_0_N93) );
  XOR2_X1 u_hpc2_0_U74 ( .A(io_i1_s2), .B(p_rand_10), .Z(n_hpc2_0_N94) );
  XOR2_X1 u_hpc2_0_U73 ( .A(io_i1_s3), .B(p_rand_12), .Z(n_hpc2_0_N95) );
  XOR2_X1 u_hpc2_0_U72 ( .A(io_i1_s5), .B(p_rand_14), .Z(n_hpc2_0_N96) );
  XOR2_X1 u_hpc2_0_U71 ( .A(io_i1_s0), .B(p_rand_4), .Z(n_hpc2_0_N97) );
  XOR2_X1 u_hpc2_0_U70 ( .A(io_i1_s1), .B(p_rand_8), .Z(n_hpc2_0_N98) );
  XOR2_X1 u_hpc2_0_U69 ( .A(io_i1_s2), .B(p_rand_11), .Z(n_hpc2_0_N99) );
  INV_X1 u_hpc2_0_U68 ( .A(io_i0_s0), .ZN(n_hpc2_0_n1) );
  INV_X1 u_hpc2_0_U67 ( .A(io_i0_s1), .ZN(n_hpc2_0_n2) );
  INV_X1 u_hpc2_0_U66 ( .A(io_i0_s2), .ZN(n_hpc2_0_n3) );
  INV_X1 u_hpc2_0_U65 ( .A(io_i0_s3), .ZN(n_hpc2_0_n4) );
  INV_X1 u_hpc2_0_U64 ( .A(io_i0_s4), .ZN(n_hpc2_0_n5) );
  INV_X1 u_hpc2_0_U63 ( .A(io_i0_s5), .ZN(n_hpc2_0_n6) );
  XOR2_X1 u_hpc2_0_U62 ( .A(n_hpc2_0__hpc_u05), .B(n_hpc2_0_n124), .Z(
        n_hpc2_0_n65) );
  XOR2_X1 u_hpc2_0_U61 ( .A(n_hpc2_0_n122), .B(n_hpc2_0_n123), .Z(n_hpc2_0_n66) );
  XOR2_X1 u_hpc2_0_U60 ( .A(n_hpc2_0_n65), .B(n_hpc2_0_n66), .Z(n_hpc2_0_n61)
         );
  XOR2_X1 u_hpc2_0_U59 ( .A(n_hpc2_0_n118), .B(n_hpc2_0_n119), .Z(n_hpc2_0_n63) );
  XOR2_X1 u_hpc2_0_U58 ( .A(n_hpc2_0_n120), .B(n_hpc2_0_n121), .Z(n_hpc2_0_n64) );
  XOR2_X1 u_hpc2_0_U57 ( .A(n_hpc2_0_n63), .B(n_hpc2_0_n64), .Z(n_hpc2_0_n62)
         );
  XOR2_X1 u_hpc2_0_U56 ( .A(n_hpc2_0_n61), .B(n_hpc2_0_n62), .Z(n_hpc2_0_n60)
         );
  XOR2_X1 u_hpc2_0_U55 ( .A(n_hpc2_0_n60), .B(n_hpc2_0_n126), .Z(n_hpc2_0_n58)
         );
  XOR2_X1 u_hpc2_0_U54 ( .A(n_hpc2_0_n117), .B(n_hpc2_0_n125), .Z(n_hpc2_0_n59) );
  XOR2_X1 u_hpc2_0_U53 ( .A(n_hpc2_0_n58), .B(n_hpc2_0_n59), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U52 ( .A(n_hpc2_0__hpc_u15), .B(n_hpc2_0_n114), .Z(
        n_hpc2_0_n56) );
  XOR2_X1 u_hpc2_0_U51 ( .A(n_hpc2_0_n112), .B(n_hpc2_0_n113), .Z(n_hpc2_0_n57) );
  XOR2_X1 u_hpc2_0_U50 ( .A(n_hpc2_0_n56), .B(n_hpc2_0_n57), .Z(n_hpc2_0_n52)
         );
  XOR2_X1 u_hpc2_0_U49 ( .A(n_hpc2_0_n108), .B(n_hpc2_0_n109), .Z(n_hpc2_0_n54) );
  XOR2_X1 u_hpc2_0_U48 ( .A(n_hpc2_0_n110), .B(n_hpc2_0_n111), .Z(n_hpc2_0_n55) );
  XOR2_X1 u_hpc2_0_U47 ( .A(n_hpc2_0_n54), .B(n_hpc2_0_n55), .Z(n_hpc2_0_n53)
         );
  XOR2_X1 u_hpc2_0_U46 ( .A(n_hpc2_0_n52), .B(n_hpc2_0_n53), .Z(n_hpc2_0_n51)
         );
  XOR2_X1 u_hpc2_0_U45 ( .A(n_hpc2_0_n51), .B(n_hpc2_0_n116), .Z(n_hpc2_0_n49)
         );
  XOR2_X1 u_hpc2_0_U44 ( .A(n_hpc2_0_n107), .B(n_hpc2_0_n115), .Z(n_hpc2_0_n50) );
  XOR2_X1 u_hpc2_0_U43 ( .A(n_hpc2_0_n49), .B(n_hpc2_0_n50), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U42 ( .A(n_hpc2_0__hpc_u25), .B(n_hpc2_0_n104), .Z(
        n_hpc2_0_n47) );
  XOR2_X1 u_hpc2_0_U41 ( .A(n_hpc2_0_n102), .B(n_hpc2_0_n103), .Z(n_hpc2_0_n48) );
  XOR2_X1 u_hpc2_0_U40 ( .A(n_hpc2_0_n47), .B(n_hpc2_0_n48), .Z(n_hpc2_0_n43)
         );
  XOR2_X1 u_hpc2_0_U39 ( .A(n_hpc2_0_n98), .B(n_hpc2_0_n99), .Z(n_hpc2_0_n45)
         );
  XOR2_X1 u_hpc2_0_U38 ( .A(n_hpc2_0_n100), .B(n_hpc2_0_n101), .Z(n_hpc2_0_n46) );
  XOR2_X1 u_hpc2_0_U37 ( .A(n_hpc2_0_n45), .B(n_hpc2_0_n46), .Z(n_hpc2_0_n44)
         );
  XOR2_X1 u_hpc2_0_U36 ( .A(n_hpc2_0_n43), .B(n_hpc2_0_n44), .Z(n_hpc2_0_n42)
         );
  XOR2_X1 u_hpc2_0_U35 ( .A(n_hpc2_0_n42), .B(n_hpc2_0_n106), .Z(n_hpc2_0_n40)
         );
  XOR2_X1 u_hpc2_0_U34 ( .A(n_hpc2_0_n97), .B(n_hpc2_0_n105), .Z(n_hpc2_0_n41)
         );
  XOR2_X1 u_hpc2_0_U33 ( .A(n_hpc2_0_n40), .B(n_hpc2_0_n41), .Z(io_o0_s2) );
  XOR2_X1 u_hpc2_0_U32 ( .A(n_hpc2_0__hpc_u35), .B(n_hpc2_0_n94), .Z(
        n_hpc2_0_n38) );
  XOR2_X1 u_hpc2_0_U31 ( .A(n_hpc2_0_n92), .B(n_hpc2_0_n93), .Z(n_hpc2_0_n39)
         );
  XOR2_X1 u_hpc2_0_U30 ( .A(n_hpc2_0_n38), .B(n_hpc2_0_n39), .Z(n_hpc2_0_n34)
         );
  XOR2_X1 u_hpc2_0_U29 ( .A(n_hpc2_0_n88), .B(n_hpc2_0_n89), .Z(n_hpc2_0_n36)
         );
  XOR2_X1 u_hpc2_0_U28 ( .A(n_hpc2_0_n90), .B(n_hpc2_0_n91), .Z(n_hpc2_0_n37)
         );
  XOR2_X1 u_hpc2_0_U27 ( .A(n_hpc2_0_n36), .B(n_hpc2_0_n37), .Z(n_hpc2_0_n35)
         );
  XOR2_X1 u_hpc2_0_U26 ( .A(n_hpc2_0_n34), .B(n_hpc2_0_n35), .Z(n_hpc2_0_n33)
         );
  XOR2_X1 u_hpc2_0_U25 ( .A(n_hpc2_0_n33), .B(n_hpc2_0_n96), .Z(n_hpc2_0_n31)
         );
  XOR2_X1 u_hpc2_0_U24 ( .A(n_hpc2_0_n87), .B(n_hpc2_0_n95), .Z(n_hpc2_0_n32)
         );
  XOR2_X1 u_hpc2_0_U23 ( .A(n_hpc2_0_n31), .B(n_hpc2_0_n32), .Z(io_o0_s3) );
  XOR2_X1 u_hpc2_0_U22 ( .A(n_hpc2_0__hpc_u45), .B(n_hpc2_0_n84), .Z(
        n_hpc2_0_n29) );
  XOR2_X1 u_hpc2_0_U21 ( .A(n_hpc2_0_n82), .B(n_hpc2_0_n83), .Z(n_hpc2_0_n30)
         );
  XOR2_X1 u_hpc2_0_U20 ( .A(n_hpc2_0_n29), .B(n_hpc2_0_n30), .Z(n_hpc2_0_n25)
         );
  XOR2_X1 u_hpc2_0_U19 ( .A(n_hpc2_0_n78), .B(n_hpc2_0_n79), .Z(n_hpc2_0_n27)
         );
  XOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0_n80), .B(n_hpc2_0_n81), .Z(n_hpc2_0_n28)
         );
  XOR2_X1 u_hpc2_0_U17 ( .A(n_hpc2_0_n27), .B(n_hpc2_0_n28), .Z(n_hpc2_0_n26)
         );
  XOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_n25), .B(n_hpc2_0_n26), .Z(n_hpc2_0_n24)
         );
  XOR2_X1 u_hpc2_0_U15 ( .A(n_hpc2_0_n24), .B(n_hpc2_0_n86), .Z(n_hpc2_0_n22)
         );
  XOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0_n77), .B(n_hpc2_0_n85), .Z(n_hpc2_0_n23)
         );
  XOR2_X1 u_hpc2_0_U13 ( .A(n_hpc2_0_n22), .B(n_hpc2_0_n23), .Z(io_o0_s4) );
  XOR2_X1 u_hpc2_0_U12 ( .A(n_hpc2_0__hpc_u54), .B(n_hpc2_0_n74), .Z(
        n_hpc2_0_n20) );
  XOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_n72), .B(n_hpc2_0_n73), .Z(n_hpc2_0_n21)
         );
  XOR2_X1 u_hpc2_0_U10 ( .A(n_hpc2_0_n20), .B(n_hpc2_0_n21), .Z(n_hpc2_0_n16)
         );
  XOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_n68), .B(n_hpc2_0_n69), .Z(n_hpc2_0_n18)
         );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0_n70), .B(n_hpc2_0_n71), .Z(n_hpc2_0_n19)
         );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0_n18), .B(n_hpc2_0_n19), .Z(n_hpc2_0_n17)
         );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0_n16), .B(n_hpc2_0_n17), .Z(n_hpc2_0_n15)
         );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0_n15), .B(n_hpc2_0_n76), .Z(n_hpc2_0_n13)
         );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0_n67), .B(n_hpc2_0_n75), .Z(n_hpc2_0_n14)
         );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n13), .B(n_hpc2_0_n14), .Z(io_o0_s5) );
  DFF_X1 u_hpc2_0__hpc_av51_reg ( .D(n_hpc2_0_N38), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n69) );
  DFF_X1 u_hpc2_0__hpc_v51_reg ( .D(n_hpc2_0_N98), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n179) );
  DFF_X1 u_hpc2_0__hpc_av50_reg ( .D(n_hpc2_0_N37), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n67) );
  DFF_X1 u_hpc2_0__hpc_v50_reg ( .D(n_hpc2_0_N97), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n180) );
  DFF_X1 u_hpc2_0__hpc_av45_reg ( .D(n_hpc2_0_N36), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n82) );
  DFF_X1 u_hpc2_0__hpc_v45_reg ( .D(n_hpc2_0_N96), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n181) );
  DFF_X1 u_hpc2_0__hpc_av43_reg ( .D(n_hpc2_0_N35), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n81) );
  DFF_X1 u_hpc2_0__hpc_v43_reg ( .D(n_hpc2_0_N95), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n182) );
  DFF_X1 u_hpc2_0__hpc_av42_reg ( .D(n_hpc2_0_N34), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n80) );
  DFF_X1 u_hpc2_0__hpc_v42_reg ( .D(n_hpc2_0_N94), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n183) );
  DFF_X1 u_hpc2_0__hpc_av41_reg ( .D(n_hpc2_0_N33), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n79) );
  DFF_X1 u_hpc2_0__hpc_v41_reg ( .D(n_hpc2_0_N93), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n184) );
  DFF_X1 u_hpc2_0__hpc_av40_reg ( .D(n_hpc2_0_N32), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n77) );
  DFF_X1 u_hpc2_0__hpc_v40_reg ( .D(n_hpc2_0_N92), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n185) );
  DFF_X1 u_hpc2_0__hpc_av35_reg ( .D(n_hpc2_0_N31), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n92) );
  DFF_X1 u_hpc2_0__hpc_v35_reg ( .D(n_hpc2_0_N91), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n186) );
  DFF_X1 u_hpc2_0__hpc_av34_reg ( .D(n_hpc2_0_N30), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n91) );
  DFF_X1 u_hpc2_0__hpc_v34_reg ( .D(n_hpc2_0_N90), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n187) );
  DFF_X1 u_hpc2_0__hpc_av32_reg ( .D(n_hpc2_0_N29), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n90) );
  DFF_X1 u_hpc2_0__hpc_v32_reg ( .D(n_hpc2_0_N89), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n188) );
  DFF_X1 u_hpc2_0__hpc_av31_reg ( .D(n_hpc2_0_N28), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n89) );
  DFF_X1 u_hpc2_0__hpc_v31_reg ( .D(n_hpc2_0_N88), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n189) );
  DFF_X1 u_hpc2_0__hpc_av30_reg ( .D(n_hpc2_0_N27), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n87) );
  DFF_X1 u_hpc2_0__hpc_v30_reg ( .D(n_hpc2_0_N87), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n190) );
  DFF_X1 u_hpc2_0__hpc_av25_reg ( .D(n_hpc2_0_N26), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n102) );
  DFF_X1 u_hpc2_0__hpc_v25_reg ( .D(n_hpc2_0_N86), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n191) );
  DFF_X1 u_hpc2_0__hpc_av24_reg ( .D(n_hpc2_0_N25), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n101) );
  DFF_X1 u_hpc2_0__hpc_v24_reg ( .D(n_hpc2_0_N85), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n192) );
  DFF_X1 u_hpc2_0__hpc_av23_reg ( .D(n_hpc2_0_N24), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n100) );
  DFF_X1 u_hpc2_0__hpc_v23_reg ( .D(n_hpc2_0_N84), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n193) );
  DFF_X1 u_hpc2_0__hpc_av21_reg ( .D(n_hpc2_0_N23), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n99) );
  DFF_X1 u_hpc2_0__hpc_v21_reg ( .D(n_hpc2_0_N83), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n194) );
  DFF_X1 u_hpc2_0__hpc_av20_reg ( .D(n_hpc2_0_N22), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n97) );
  DFF_X1 u_hpc2_0__hpc_v20_reg ( .D(n_hpc2_0_N82), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n195) );
  DFF_X1 u_hpc2_0__hpc_av15_reg ( .D(n_hpc2_0_N21), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n112) );
  DFF_X1 u_hpc2_0__hpc_v15_reg ( .D(n_hpc2_0_N81), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n196) );
  DFF_X1 u_hpc2_0__hpc_av14_reg ( .D(n_hpc2_0_N20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n111) );
  DFF_X1 u_hpc2_0__hpc_v14_reg ( .D(n_hpc2_0_N80), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n197) );
  DFF_X1 u_hpc2_0__hpc_av13_reg ( .D(n_hpc2_0_N19), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n110) );
  DFF_X1 u_hpc2_0__hpc_v13_reg ( .D(n_hpc2_0_N79), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n198) );
  DFF_X1 u_hpc2_0__hpc_av12_reg ( .D(n_hpc2_0_N18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n109) );
  DFF_X1 u_hpc2_0__hpc_v12_reg ( .D(n_hpc2_0_N78), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n199) );
  DFF_X1 u_hpc2_0__hpc_av10_reg ( .D(n_hpc2_0_N17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n107) );
  DFF_X1 u_hpc2_0__hpc_v10_reg ( .D(n_hpc2_0_N77), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n200) );
  DFF_X1 u_hpc2_0__hpc_av05_reg ( .D(n_hpc2_0_N16), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n122) );
  DFF_X1 u_hpc2_0__hpc_v05_reg ( .D(n_hpc2_0_N76), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n201) );
  DFF_X1 u_hpc2_0__hpc_av04_reg ( .D(n_hpc2_0_N15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n121) );
  DFF_X1 u_hpc2_0__hpc_v04_reg ( .D(n_hpc2_0_N75), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n202) );
  DFF_X1 u_hpc2_0__hpc_av03_reg ( .D(n_hpc2_0_N14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n120) );
  DFF_X1 u_hpc2_0__hpc_v03_reg ( .D(n_hpc2_0_N74), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n203) );
  DFF_X1 u_hpc2_0__hpc_av02_reg ( .D(n_hpc2_0_N13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n119) );
  DFF_X1 u_hpc2_0__hpc_v02_reg ( .D(n_hpc2_0_N73), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n204) );
  DFF_X1 u_hpc2_0__hpc_av01_reg ( .D(n_hpc2_0_N12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n117) );
  DFF_X1 u_hpc2_0__hpc_v01_reg ( .D(n_hpc2_0_N72), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n205) );
  DFF_X1 u_hpc2_0__hpc_u54_reg ( .D(n_hpc2_0_N71), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u54), .QN() );
  DFF_X1 u_hpc2_0__hpc_u53_reg ( .D(n_hpc2_0_N70), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n74) );
  DFF_X1 u_hpc2_0__hpc_u52_reg ( .D(n_hpc2_0_N69), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n73) );
  DFF_X1 u_hpc2_0__hpc_u51_reg ( .D(n_hpc2_0_N68), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n76) );
  DFF_X1 u_hpc2_0__hpc_u50_reg ( .D(n_hpc2_0_N67), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n75) );
  DFF_X1 u_hpc2_0__hpc_u45_reg ( .D(n_hpc2_0_N66), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u45), .QN() );
  DFF_X1 u_hpc2_0__hpc_u43_reg ( .D(n_hpc2_0_N65), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n84) );
  DFF_X1 u_hpc2_0__hpc_u42_reg ( .D(n_hpc2_0_N64), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n83) );
  DFF_X1 u_hpc2_0__hpc_u41_reg ( .D(n_hpc2_0_N63), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n86) );
  DFF_X1 u_hpc2_0__hpc_u40_reg ( .D(n_hpc2_0_N62), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n85) );
  DFF_X1 u_hpc2_0__hpc_u35_reg ( .D(n_hpc2_0_N61), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u35), .QN() );
  DFF_X1 u_hpc2_0__hpc_u34_reg ( .D(n_hpc2_0_N60), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n94) );
  DFF_X1 u_hpc2_0__hpc_u32_reg ( .D(n_hpc2_0_N59), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n93) );
  DFF_X1 u_hpc2_0__hpc_u31_reg ( .D(n_hpc2_0_N58), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n96) );
  DFF_X1 u_hpc2_0__hpc_u30_reg ( .D(n_hpc2_0_N57), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n95) );
  DFF_X1 u_hpc2_0__hpc_u25_reg ( .D(n_hpc2_0_N56), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u25), .QN() );
  DFF_X1 u_hpc2_0__hpc_u24_reg ( .D(n_hpc2_0_N55), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n104) );
  DFF_X1 u_hpc2_0__hpc_u23_reg ( .D(n_hpc2_0_N54), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n103) );
  DFF_X1 u_hpc2_0__hpc_u21_reg ( .D(n_hpc2_0_N53), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n106) );
  DFF_X1 u_hpc2_0__hpc_u20_reg ( .D(n_hpc2_0_N52), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n105) );
  DFF_X1 u_hpc2_0__hpc_u15_reg ( .D(n_hpc2_0_N51), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u15), .QN() );
  DFF_X1 u_hpc2_0__hpc_u14_reg ( .D(n_hpc2_0_N50), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n114) );
  DFF_X1 u_hpc2_0__hpc_u13_reg ( .D(n_hpc2_0_N49), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n113) );
  DFF_X1 u_hpc2_0__hpc_u12_reg ( .D(n_hpc2_0_N48), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n116) );
  DFF_X1 u_hpc2_0__hpc_u10_reg ( .D(n_hpc2_0_N47), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n115) );
  DFF_X1 u_hpc2_0__hpc_u05_reg ( .D(n_hpc2_0_N46), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u05), .QN() );
  DFF_X1 u_hpc2_0__hpc_u04_reg ( .D(n_hpc2_0_N45), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n124) );
  DFF_X1 u_hpc2_0__hpc_u03_reg ( .D(n_hpc2_0_N44), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n123) );
  DFF_X1 u_hpc2_0__hpc_u02_reg ( .D(n_hpc2_0_N43), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n126) );
  DFF_X1 u_hpc2_0__hpc_u01_reg ( .D(n_hpc2_0_N42), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n125) );
  DFF_X1 u_hpc2_0__hpc_ab5_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n68) );
  DFF_X1 u_hpc2_0__hpc_b5_reg ( .D(io_i1_s5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n206) );
  DFF_X1 u_hpc2_0__hpc_ab4_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n78) );
  DFF_X1 u_hpc2_0__hpc_b4_reg ( .D(io_i1_s4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n207) );
  DFF_X1 u_hpc2_0__hpc_ab3_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n88) );
  DFF_X1 u_hpc2_0__hpc_b3_reg ( .D(io_i1_s3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n127) );
  DFF_X1 u_hpc2_0__hpc_ab2_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n98) );
  DFF_X1 u_hpc2_0__hpc_b2_reg ( .D(io_i1_s2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n128) );
  DFF_X1 u_hpc2_0__hpc_ab1_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n108) );
  DFF_X1 u_hpc2_0__hpc_b1_reg ( .D(io_i1_s1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n131) );
  DFF_X1 u_hpc2_0__hpc_ab0_reg ( .D(n_hpc2_0_N6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n118) );
  DFF_X1 u_hpc2_0__hpc_b0_reg ( .D(io_i1_s0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n145) );
  DFF_X1 u_hpc2_0__hpc_av54_reg ( .D(n_hpc2_0_N41), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n72) );
  DFF_X1 u_hpc2_0__hpc_av53_reg ( .D(n_hpc2_0_N40), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n71) );
  DFF_X1 u_hpc2_0__hpc_av52_reg ( .D(n_hpc2_0_N39), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n70) );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n133) );
  DFF_X1 u_hpc2_0_reg_pipeline_21_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n162) );
  DFF_X1 u_hpc2_0_reg_pipeline_27_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n173) );
  DFF_X1 u_hpc2_0_reg_pipeline_26_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n171) );
  DFF_X1 u_hpc2_0_reg_pipeline_28_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n175) );
  DFF_X1 u_hpc2_0_reg_pipeline_24_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n167) );
  DFF_X1 u_hpc2_0_reg_pipeline_29_reg ( .D(io_i0_s0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n10) );
  DFF_X1 u_hpc2_0_reg_pipeline_23_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n165) );
  DFF_X1 u_hpc2_0_reg_pipeline_19_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n158) );
  DFF_X1 u_hpc2_0_reg_pipeline_22_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n164) );
  DFF_X1 u_hpc2_0_reg_pipeline_25_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n169) );
  DFF_X1 u_hpc2_0_reg_pipeline_20_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n160) );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n136) );
  DFF_X1 u_hpc2_0_reg_pipeline_5_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n137) );
  DFF_X1 u_hpc2_0_reg_pipeline_9_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n142) );
  DFF_X1 u_hpc2_0_reg_pipeline_6_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n138) );
  DFF_X1 u_hpc2_0__hpc_r9_reg ( .D(p_rand_9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n153) );
  DFF_X1 u_hpc2_0__hpc_r6_reg ( .D(p_rand_6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n161) );
  DFF_X1 u_hpc2_0_reg_pipeline_7_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n139) );
  DFF_X1 u_hpc2_0__hpc_r8_reg ( .D(p_rand_8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n157) );
  DFF_X1 u_hpc2_0__hpc_r5_reg ( .D(p_rand_5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n163) );
  DFF_X1 u_hpc2_0__hpc_r3_reg ( .D(p_rand_3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n168) );
  DFF_X1 u_hpc2_0_reg_pipeline_8_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n140) );
  DFF_X1 u_hpc2_0__hpc_r7_reg ( .D(p_rand_7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n159) );
  DFF_X1 u_hpc2_0__hpc_r4_reg ( .D(p_rand_4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n166) );
  DFF_X1 u_hpc2_0__hpc_r2_reg ( .D(p_rand_2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n170) );
  DFF_X1 u_hpc2_0__hpc_r14_reg ( .D(p_rand_14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n135) );
  DFF_X1 u_hpc2_0_reg_pipeline_18_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n156) );
  DFF_X1 u_hpc2_0_reg_pipeline_17_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n155) );
  DFF_X1 u_hpc2_0_reg_pipeline_16_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n154) );
  DFF_X1 u_hpc2_0_reg_pipeline_15_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n152) );
  DFF_X1 u_hpc2_0_reg_pipeline_14_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n150) );
  DFF_X1 u_hpc2_0_reg_pipeline_13_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n148) );
  DFF_X1 u_hpc2_0_reg_pipeline_12_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n147) );
  DFF_X1 u_hpc2_0_reg_pipeline_11_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n146) );
  DFF_X1 u_hpc2_0_reg_pipeline_10_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n144) );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n132) );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n130) );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n129) );
  DFF_X1 u_hpc2_0__hpc_v54_reg ( .D(n_hpc2_0_N101), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n176) );
  DFF_X1 u_hpc2_0__hpc_v53_reg ( .D(n_hpc2_0_N100), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n177) );
  DFF_X1 u_hpc2_0__hpc_v52_reg ( .D(n_hpc2_0_N99), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n178) );
  DFF_X1 u_hpc2_0_reg_pipeline_34_reg ( .D(io_i0_s5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n11) );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(n_hpc2_0_n6), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n134) );
  DFF_X1 u_hpc2_0_reg_pipeline_30_reg ( .D(io_i0_s1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n9) );
  DFF_X1 u_hpc2_0_reg_pipeline_31_reg ( .D(io_i0_s2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n8) );
  DFF_X1 u_hpc2_0_reg_pipeline_32_reg ( .D(io_i0_s3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n7) );
  DFF_X1 u_hpc2_0_reg_pipeline_33_reg ( .D(io_i0_s4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n12) );
  DFF_X1 u_hpc2_0__hpc_r13_reg ( .D(p_rand_13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n141) );
  DFF_X1 u_hpc2_0__hpc_r12_reg ( .D(p_rand_12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n143) );
  DFF_X1 u_hpc2_0__hpc_r11_reg ( .D(p_rand_11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n149) );
  DFF_X1 u_hpc2_0__hpc_r10_reg ( .D(p_rand_10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n151) );
  DFF_X1 u_hpc2_0__hpc_r1_reg ( .D(p_rand_1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n172) );
  DFF_X1 u_hpc2_0__hpc_r0_reg ( .D(p_rand_0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n174) );
endmodule

