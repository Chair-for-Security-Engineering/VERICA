
module CINI ( io_a_0, io_a_1, io_a_2, io_b_0, io_b_1, io_b_2, io_c_0, io_c_1, 
        io_c_2, io_rand, clk, reset );
  input [4:0] io_a_0;
  input [4:0] io_a_1;
  input [4:0] io_a_2;
  input [4:0] io_b_0;
  input [4:0] io_b_1;
  input [4:0] io_b_2;
  output [4:0] io_c_0;
  output [4:0] io_c_1;
  output [4:0] io_c_2;
  input [2:0] io_rand;
  input clk, reset;
  wire   simpleNot_30_port_z, simpleNot_31_port_z, simpleNot_32_port_z,
         simpleNot_33_port_z, simpleNot_34_port_z, simpleNot_35_port_z,
         simpleNot_36_port_z, simpleNot_37_port_z, simpleNot_38_port_z,
         simpleNot_39_port_z, simpleNot_40_port_z, simpleNot_41_port_z,
         simpleNot_42_port_z, simpleNot_43_port_z, simpleNot_44_port_z,
         simpleNot_45_port_z, simpleNot_46_port_z, simpleNot_47_port_z,
         simpleNot_48_port_z, simpleNot_49_port_z, simpleNot_50_port_z,
         simpleNot_51_port_z, simpleNot_52_port_z, simpleNot_53_port_z,
         simpleNot_54_port_z, simpleNot_55_port_z, simpleNot_56_port_z,
         simpleNot_57_port_z, simpleNot_58_port_z, simpleNot_59_port_z,
         simpleXor_30_port_z, simpleXor_31_port_z, simpleXor_32_port_z,
         simpleXor_33_port_z, simpleXor_34_port_z, simpleXor_35_port_z,
         simpleXor_36_port_z, simpleXor_37_port_z, simpleXor_38_port_z,
         simpleXor_39_port_z, simpleXor_40_port_z, simpleXor_41_port_z,
         simpleXor_42_port_z, simpleXor_43_port_z, simpleXor_44_port_z,
         simpleXor_45_port_z, simpleXor_46_port_z, simpleXor_47_port_z,
         simpleXor_48_port_z, simpleXor_49_port_z, simpleXor_50_port_z,
         simpleXor_51_port_z, simpleXor_52_port_z, simpleXor_53_port_z,
         simpleXor_54_port_z, simpleXor_55_port_z, simpleXor_56_port_z,
         simpleXor_57_port_z, simpleXor_58_port_z, simpleXor_59_port_z,
         n_zz_io_c_0_0_, n_zz_io_c_1_0_, n_zz_io_c_2_0_, n_zz_io_c_0_4_0_,
         n_zz_io_c_1_4_0_, n_zz_io_c_2_4_0_, n_zz_io_c_0_8_0_,
         n_zz_io_c_1_8_0_, n_zz_io_c_2_8_0_, n_zz_io_c_0_12_0_,
         n_zz_io_c_1_12_0_, n_zz_io_c_2_12_0_, n_zz_io_c_0_16_0_,
         n_zz_io_c_1_16_0_, n_zz_io_c_2_16_0_, N0, N1, N2, N3, N4, N5, N6, N7,
         N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, cor_maj_59_port_o,
         cor_maj_58_port_o, cor_maj_57_port_o, cor_maj_56_port_o,
         cor_maj_55_port_o, cor_maj_54_port_o, cor_maj_53_port_o,
         cor_maj_52_port_o, cor_maj_51_port_o, cor_maj_50_port_o,
         cor_maj_49_port_o, cor_maj_48_port_o, cor_maj_47_port_o,
         cor_maj_46_port_o, cor_maj_45_port_o, cor_maj_44_port_o,
         cor_maj_43_port_o, cor_maj_42_port_o, cor_maj_41_port_o,
         cor_maj_40_port_o, cor_maj_39_port_o, cor_maj_38_port_o,
         cor_maj_37_port_o, cor_maj_36_port_o, cor_maj_35_port_o,
         cor_maj_34_port_o, cor_maj_33_port_o, cor_maj_32_port_o,
         cor_maj_31_port_o, cor_maj_30_port_o, cor_maj_30_n13, cor_maj_30_n12,
         cor_maj_30_n11, cor_maj_30_n10, cor_maj_30_n9, cor_maj_30_n8,
         cor_maj_30_n7, cor_maj_30_n6, cor_maj_30_n5, cor_maj_30_n4,
         cor_maj_30_n3, cor_maj_30_n2, cor_maj_30_n1, cor_maj_31_n26,
         cor_maj_31_n25, cor_maj_31_n24, cor_maj_31_n23, cor_maj_31_n22,
         cor_maj_31_n21, cor_maj_31_n20, cor_maj_31_n19, cor_maj_31_n18,
         cor_maj_31_n17, cor_maj_31_n16, cor_maj_31_n15, cor_maj_31_n14,
         cor_maj_32_n26, cor_maj_32_n25, cor_maj_32_n24, cor_maj_32_n23,
         cor_maj_32_n22, cor_maj_32_n21, cor_maj_32_n20, cor_maj_32_n19,
         cor_maj_32_n18, cor_maj_32_n17, cor_maj_32_n16, cor_maj_32_n15,
         cor_maj_32_n14, cor_maj_33_n26, cor_maj_33_n25, cor_maj_33_n24,
         cor_maj_33_n23, cor_maj_33_n22, cor_maj_33_n21, cor_maj_33_n20,
         cor_maj_33_n19, cor_maj_33_n18, cor_maj_33_n17, cor_maj_33_n16,
         cor_maj_33_n15, cor_maj_33_n14, cor_maj_34_n26, cor_maj_34_n25,
         cor_maj_34_n24, cor_maj_34_n23, cor_maj_34_n22, cor_maj_34_n21,
         cor_maj_34_n20, cor_maj_34_n19, cor_maj_34_n18, cor_maj_34_n17,
         cor_maj_34_n16, cor_maj_34_n15, cor_maj_34_n14, cor_maj_35_n26,
         cor_maj_35_n25, cor_maj_35_n24, cor_maj_35_n23, cor_maj_35_n22,
         cor_maj_35_n21, cor_maj_35_n20, cor_maj_35_n19, cor_maj_35_n18,
         cor_maj_35_n17, cor_maj_35_n16, cor_maj_35_n15, cor_maj_35_n14,
         cor_maj_36_n26, cor_maj_36_n25, cor_maj_36_n24, cor_maj_36_n23,
         cor_maj_36_n22, cor_maj_36_n21, cor_maj_36_n20, cor_maj_36_n19,
         cor_maj_36_n18, cor_maj_36_n17, cor_maj_36_n16, cor_maj_36_n15,
         cor_maj_36_n14, cor_maj_37_n26, cor_maj_37_n25, cor_maj_37_n24,
         cor_maj_37_n23, cor_maj_37_n22, cor_maj_37_n21, cor_maj_37_n20,
         cor_maj_37_n19, cor_maj_37_n18, cor_maj_37_n17, cor_maj_37_n16,
         cor_maj_37_n15, cor_maj_37_n14, cor_maj_38_n26, cor_maj_38_n25,
         cor_maj_38_n24, cor_maj_38_n23, cor_maj_38_n22, cor_maj_38_n21,
         cor_maj_38_n20, cor_maj_38_n19, cor_maj_38_n18, cor_maj_38_n17,
         cor_maj_38_n16, cor_maj_38_n15, cor_maj_38_n14, cor_maj_39_n26,
         cor_maj_39_n25, cor_maj_39_n24, cor_maj_39_n23, cor_maj_39_n22,
         cor_maj_39_n21, cor_maj_39_n20, cor_maj_39_n19, cor_maj_39_n18,
         cor_maj_39_n17, cor_maj_39_n16, cor_maj_39_n15, cor_maj_39_n14,
         cor_maj_40_n26, cor_maj_40_n25, cor_maj_40_n24, cor_maj_40_n23,
         cor_maj_40_n22, cor_maj_40_n21, cor_maj_40_n20, cor_maj_40_n19,
         cor_maj_40_n18, cor_maj_40_n17, cor_maj_40_n16, cor_maj_40_n15,
         cor_maj_40_n14, cor_maj_41_n26, cor_maj_41_n25, cor_maj_41_n24,
         cor_maj_41_n23, cor_maj_41_n22, cor_maj_41_n21, cor_maj_41_n20,
         cor_maj_41_n19, cor_maj_41_n18, cor_maj_41_n17, cor_maj_41_n16,
         cor_maj_41_n15, cor_maj_41_n14, cor_maj_42_n26, cor_maj_42_n25,
         cor_maj_42_n24, cor_maj_42_n23, cor_maj_42_n22, cor_maj_42_n21,
         cor_maj_42_n20, cor_maj_42_n19, cor_maj_42_n18, cor_maj_42_n17,
         cor_maj_42_n16, cor_maj_42_n15, cor_maj_42_n14, cor_maj_43_n26,
         cor_maj_43_n25, cor_maj_43_n24, cor_maj_43_n23, cor_maj_43_n22,
         cor_maj_43_n21, cor_maj_43_n20, cor_maj_43_n19, cor_maj_43_n18,
         cor_maj_43_n17, cor_maj_43_n16, cor_maj_43_n15, cor_maj_43_n14,
         cor_maj_44_n26, cor_maj_44_n25, cor_maj_44_n24, cor_maj_44_n23,
         cor_maj_44_n22, cor_maj_44_n21, cor_maj_44_n20, cor_maj_44_n19,
         cor_maj_44_n18, cor_maj_44_n17, cor_maj_44_n16, cor_maj_44_n15,
         cor_maj_44_n14, cor_maj_45_n26, cor_maj_45_n25, cor_maj_45_n24,
         cor_maj_45_n23, cor_maj_45_n22, cor_maj_45_n21, cor_maj_45_n20,
         cor_maj_45_n19, cor_maj_45_n18, cor_maj_45_n17, cor_maj_45_n16,
         cor_maj_45_n15, cor_maj_45_n14, cor_maj_46_n26, cor_maj_46_n25,
         cor_maj_46_n24, cor_maj_46_n23, cor_maj_46_n22, cor_maj_46_n21,
         cor_maj_46_n20, cor_maj_46_n19, cor_maj_46_n18, cor_maj_46_n17,
         cor_maj_46_n16, cor_maj_46_n15, cor_maj_46_n14, cor_maj_47_n26,
         cor_maj_47_n25, cor_maj_47_n24, cor_maj_47_n23, cor_maj_47_n22,
         cor_maj_47_n21, cor_maj_47_n20, cor_maj_47_n19, cor_maj_47_n18,
         cor_maj_47_n17, cor_maj_47_n16, cor_maj_47_n15, cor_maj_47_n14,
         cor_maj_48_n26, cor_maj_48_n25, cor_maj_48_n24, cor_maj_48_n23,
         cor_maj_48_n22, cor_maj_48_n21, cor_maj_48_n20, cor_maj_48_n19,
         cor_maj_48_n18, cor_maj_48_n17, cor_maj_48_n16, cor_maj_48_n15,
         cor_maj_48_n14, cor_maj_49_n26, cor_maj_49_n25, cor_maj_49_n24,
         cor_maj_49_n23, cor_maj_49_n22, cor_maj_49_n21, cor_maj_49_n20,
         cor_maj_49_n19, cor_maj_49_n18, cor_maj_49_n17, cor_maj_49_n16,
         cor_maj_49_n15, cor_maj_49_n14, cor_maj_50_n26, cor_maj_50_n25,
         cor_maj_50_n24, cor_maj_50_n23, cor_maj_50_n22, cor_maj_50_n21,
         cor_maj_50_n20, cor_maj_50_n19, cor_maj_50_n18, cor_maj_50_n17,
         cor_maj_50_n16, cor_maj_50_n15, cor_maj_50_n14, cor_maj_51_n26,
         cor_maj_51_n25, cor_maj_51_n24, cor_maj_51_n23, cor_maj_51_n22,
         cor_maj_51_n21, cor_maj_51_n20, cor_maj_51_n19, cor_maj_51_n18,
         cor_maj_51_n17, cor_maj_51_n16, cor_maj_51_n15, cor_maj_51_n14,
         cor_maj_52_n26, cor_maj_52_n25, cor_maj_52_n24, cor_maj_52_n23,
         cor_maj_52_n22, cor_maj_52_n21, cor_maj_52_n20, cor_maj_52_n19,
         cor_maj_52_n18, cor_maj_52_n17, cor_maj_52_n16, cor_maj_52_n15,
         cor_maj_52_n14, cor_maj_53_n26, cor_maj_53_n25, cor_maj_53_n24,
         cor_maj_53_n23, cor_maj_53_n22, cor_maj_53_n21, cor_maj_53_n20,
         cor_maj_53_n19, cor_maj_53_n18, cor_maj_53_n17, cor_maj_53_n16,
         cor_maj_53_n15, cor_maj_53_n14, cor_maj_54_n26, cor_maj_54_n25,
         cor_maj_54_n24, cor_maj_54_n23, cor_maj_54_n22, cor_maj_54_n21,
         cor_maj_54_n20, cor_maj_54_n19, cor_maj_54_n18, cor_maj_54_n17,
         cor_maj_54_n16, cor_maj_54_n15, cor_maj_54_n14, cor_maj_55_n26,
         cor_maj_55_n25, cor_maj_55_n24, cor_maj_55_n23, cor_maj_55_n22,
         cor_maj_55_n21, cor_maj_55_n20, cor_maj_55_n19, cor_maj_55_n18,
         cor_maj_55_n17, cor_maj_55_n16, cor_maj_55_n15, cor_maj_55_n14,
         cor_maj_56_n26, cor_maj_56_n25, cor_maj_56_n24, cor_maj_56_n23,
         cor_maj_56_n22, cor_maj_56_n21, cor_maj_56_n20, cor_maj_56_n19,
         cor_maj_56_n18, cor_maj_56_n17, cor_maj_56_n16, cor_maj_56_n15,
         cor_maj_56_n14, cor_maj_57_n26, cor_maj_57_n25, cor_maj_57_n24,
         cor_maj_57_n23, cor_maj_57_n22, cor_maj_57_n21, cor_maj_57_n20,
         cor_maj_57_n19, cor_maj_57_n18, cor_maj_57_n17, cor_maj_57_n16,
         cor_maj_57_n15, cor_maj_57_n14, cor_maj_58_n26, cor_maj_58_n25,
         cor_maj_58_n24, cor_maj_58_n23, cor_maj_58_n22, cor_maj_58_n21,
         cor_maj_58_n20, cor_maj_58_n19, cor_maj_58_n18, cor_maj_58_n17,
         cor_maj_58_n16, cor_maj_58_n15, cor_maj_58_n14, cor_maj_59_n26,
         cor_maj_59_n25, cor_maj_59_n24, cor_maj_59_n23, cor_maj_59_n22,
         cor_maj_59_n21, cor_maj_59_n20, cor_maj_59_n19, cor_maj_59_n18,
         cor_maj_59_n17, cor_maj_59_n16, cor_maj_59_n15, cor_maj_59_n14;
  wire   [4:0] v_1_0_1;
  wire   [4:0] v_1_0_2;
  wire   [4:0] v_1_1_0;
  wire   [4:0] v_1_1_2;
  wire   [4:0] v_1_2_0;
  wire   [4:0] v_1_2_1;
  wire   [4:0] cor_port_v_0_1;
  wire   [4:0] cor_port_v_0_2;
  wire   [4:0] cor_port_v_1_0;
  wire   [4:0] cor_port_v_1_2;
  wire   [4:0] cor_port_v_2_0;
  wire   [4:0] cor_port_v_2_1;
  wire   [2:1] n_zz_io_c_0_3;
  wire   [4:0] u_0_1;
  wire   [4:0] u_0_2;
  wire   [2:1] n_zz_io_c_1_3;
  wire   [4:0] u_1_0;
  wire   [4:0] u_1_2;
  wire   [2:1] n_zz_io_c_2_3;
  wire   [4:0] u_2_0;
  wire   [4:0] u_2_1;
  wire   [2:1] n_zz_io_c_0_7;
  wire   [2:1] n_zz_io_c_1_7;
  wire   [2:1] n_zz_io_c_2_7;
  wire   [2:1] n_zz_io_c_0_11;
  wire   [2:1] n_zz_io_c_1_11;
  wire   [2:1] n_zz_io_c_2_11;
  wire   [2:1] n_zz_io_c_0_15;
  wire   [2:1] n_zz_io_c_1_15;
  wire   [2:1] n_zz_io_c_2_15;
  wire   [2:1] n_zz_io_c_0_19;
  wire   [2:1] n_zz_io_c_1_19;
  wire   [2:1] n_zz_io_c_2_19;
  wire   [4:0] rand_reg_0;
  wire   [4:0] rand_reg_1;
  wire   [4:0] rand_reg_3;
  wire   [4:0] rand_reg_2;
  wire   [4:0] rand_reg_4;
  wire   [4:0] rand_reg_5;
  wire   [4:0] b_reg_0;
  wire   [4:0] b_reg_1;
  wire   [4:0] b_reg_2;

  DFF_X1 rand_reg_2_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[4]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[3]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[2]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[1]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[0]), 
        .QN() );
  DFF_X1 b_reg_1_reg_4_ ( .D(io_b_1[4]), .CK(clk), .Q(b_reg_1[4]), .QN() );
  DFF_X1 b_reg_1_reg_3_ ( .D(io_b_1[3]), .CK(clk), .Q(b_reg_1[3]), .QN() );
  DFF_X1 b_reg_1_reg_2_ ( .D(io_b_1[2]), .CK(clk), .Q(b_reg_1[2]), .QN() );
  DFF_X1 b_reg_1_reg_1_ ( .D(io_b_1[1]), .CK(clk), .Q(b_reg_1[1]), .QN() );
  DFF_X1 b_reg_1_reg_0_ ( .D(io_b_1[0]), .CK(clk), .Q(b_reg_1[0]), .QN() );
  DFF_X1 b_reg_2_reg_4_ ( .D(io_b_2[4]), .CK(clk), .Q(b_reg_2[4]), .QN() );
  DFF_X1 b_reg_2_reg_3_ ( .D(io_b_2[3]), .CK(clk), .Q(b_reg_2[3]), .QN() );
  DFF_X1 b_reg_2_reg_2_ ( .D(io_b_2[2]), .CK(clk), .Q(b_reg_2[2]), .QN() );
  DFF_X1 b_reg_2_reg_1_ ( .D(io_b_2[1]), .CK(clk), .Q(b_reg_2[1]), .QN() );
  DFF_X1 b_reg_2_reg_0_ ( .D(io_b_2[0]), .CK(clk), .Q(b_reg_2[0]), .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_2_ ( .D(N74), .CK(clk), .Q(n_zz_io_c_2_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_1_ ( .D(N73), .CK(clk), .Q(n_zz_io_c_2_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_0_ ( .D(N72), .CK(clk), .Q(n_zz_io_c_2_16_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_2_ ( .D(N71), .CK(clk), .Q(n_zz_io_c_1_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_1_ ( .D(N70), .CK(clk), .Q(n_zz_io_c_1_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_0_ ( .D(N69), .CK(clk), .Q(n_zz_io_c_1_16_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_2_ ( .D(N68), .CK(clk), .Q(n_zz_io_c_0_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_1_ ( .D(N67), .CK(clk), .Q(n_zz_io_c_0_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_15_reg_2_ ( .D(N65), .CK(clk), .Q(n_zz_io_c_2_15[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_15_reg_1_ ( .D(N64), .CK(clk), .Q(n_zz_io_c_2_15[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_15_reg_0_ ( .D(N63), .CK(clk), .Q(n_zz_io_c_2_12_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_15_reg_2_ ( .D(N62), .CK(clk), .Q(n_zz_io_c_1_15[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_15_reg_1_ ( .D(N61), .CK(clk), .Q(n_zz_io_c_1_15[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_15_reg_0_ ( .D(N60), .CK(clk), .Q(n_zz_io_c_1_12_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_15_reg_2_ ( .D(N59), .CK(clk), .Q(n_zz_io_c_0_15[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_15_reg_1_ ( .D(N58), .CK(clk), .Q(n_zz_io_c_0_15[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_11_reg_2_ ( .D(N56), .CK(clk), .Q(n_zz_io_c_2_11[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_11_reg_1_ ( .D(N55), .CK(clk), .Q(n_zz_io_c_2_11[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_11_reg_0_ ( .D(N54), .CK(clk), .Q(n_zz_io_c_2_8_0_), 
        .QN() );
  DFF_X1 rand_reg_5_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[4]), 
        .QN() );
  DFF_X1 u_2_1_reg_4_ ( .D(N29), .CK(clk), .Q(u_2_1[4]), .QN() );
  DFF_X1 rand_reg_5_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[3]), 
        .QN() );
  DFF_X1 u_2_1_reg_3_ ( .D(N23), .CK(clk), .Q(u_2_1[3]), .QN() );
  DFF_X1 rand_reg_5_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[2]), 
        .QN() );
  DFF_X1 u_2_1_reg_2_ ( .D(N17), .CK(clk), .Q(u_2_1[2]), .QN() );
  DFF_X1 rand_reg_5_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[1]), 
        .QN() );
  DFF_X1 u_2_1_reg_1_ ( .D(N11), .CK(clk), .Q(u_2_1[1]), .QN() );
  DFF_X1 rand_reg_5_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[0]), 
        .QN() );
  DFF_X1 u_2_1_reg_0_ ( .D(N5), .CK(clk), .Q(u_2_1[0]), .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_2_ ( .D(N53), .CK(clk), .Q(n_zz_io_c_1_11[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_1_ ( .D(N52), .CK(clk), .Q(n_zz_io_c_1_11[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_0_ ( .D(N51), .CK(clk), .Q(n_zz_io_c_1_8_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_2_ ( .D(N50), .CK(clk), .Q(n_zz_io_c_0_11[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_1_ ( .D(N49), .CK(clk), .Q(n_zz_io_c_0_11[1]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[4]), 
        .QN() );
  DFF_X1 u_0_1_reg_4_ ( .D(N24), .CK(clk), .Q(u_0_1[4]), .QN() );
  DFF_X1 rand_reg_0_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[3]), 
        .QN() );
  DFF_X1 u_0_1_reg_3_ ( .D(N18), .CK(clk), .Q(u_0_1[3]), .QN() );
  DFF_X1 rand_reg_0_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[2]), 
        .QN() );
  DFF_X1 u_0_1_reg_2_ ( .D(N12), .CK(clk), .Q(u_0_1[2]), .QN() );
  DFF_X1 rand_reg_0_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[1]), 
        .QN() );
  DFF_X1 u_0_1_reg_1_ ( .D(N6), .CK(clk), .Q(u_0_1[1]), .QN() );
  DFF_X1 rand_reg_0_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[0]), 
        .QN() );
  DFF_X1 u_0_1_reg_0_ ( .D(N0), .CK(clk), .Q(u_0_1[0]), .QN() );
  DFF_X1 rand_reg_3_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[4]), 
        .QN() );
  DFF_X1 u_1_0_reg_4_ ( .D(N26), .CK(clk), .Q(u_1_0[4]), .QN() );
  DFF_X1 rand_reg_3_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[3]), 
        .QN() );
  DFF_X1 u_1_0_reg_3_ ( .D(N20), .CK(clk), .Q(u_1_0[3]), .QN() );
  DFF_X1 rand_reg_3_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[2]), 
        .QN() );
  DFF_X1 u_1_0_reg_2_ ( .D(N14), .CK(clk), .Q(u_1_0[2]), .QN() );
  DFF_X1 rand_reg_3_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[1]), 
        .QN() );
  DFF_X1 u_1_0_reg_1_ ( .D(N8), .CK(clk), .Q(u_1_0[1]), .QN() );
  DFF_X1 rand_reg_3_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[0]), 
        .QN() );
  DFF_X1 u_1_0_reg_0_ ( .D(N2), .CK(clk), .Q(u_1_0[0]), .QN() );
  DFF_X1 u_1_2_reg_4_ ( .D(N27), .CK(clk), .Q(u_1_2[4]), .QN() );
  DFF_X1 u_1_2_reg_3_ ( .D(N21), .CK(clk), .Q(u_1_2[3]), .QN() );
  DFF_X1 u_1_2_reg_2_ ( .D(N15), .CK(clk), .Q(u_1_2[2]), .QN() );
  DFF_X1 u_1_2_reg_1_ ( .D(N9), .CK(clk), .Q(u_1_2[1]), .QN() );
  DFF_X1 u_1_2_reg_0_ ( .D(N3), .CK(clk), .Q(u_1_2[0]), .QN() );
  DFF_X1 u_zz_io_c_2_7_reg_2_ ( .D(N47), .CK(clk), .Q(n_zz_io_c_2_7[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_7_reg_1_ ( .D(N46), .CK(clk), .Q(n_zz_io_c_2_7[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_7_reg_0_ ( .D(N45), .CK(clk), .Q(n_zz_io_c_2_4_0_), .QN()
         );
  DFF_X1 rand_reg_1_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[4]), 
        .QN() );
  DFF_X1 u_0_2_reg_4_ ( .D(N25), .CK(clk), .Q(u_0_2[4]), .QN() );
  DFF_X1 rand_reg_1_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[3]), 
        .QN() );
  DFF_X1 u_0_2_reg_3_ ( .D(N19), .CK(clk), .Q(u_0_2[3]), .QN() );
  DFF_X1 rand_reg_1_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[2]), 
        .QN() );
  DFF_X1 u_0_2_reg_2_ ( .D(N13), .CK(clk), .Q(u_0_2[2]), .QN() );
  DFF_X1 rand_reg_1_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[1]), 
        .QN() );
  DFF_X1 u_0_2_reg_1_ ( .D(N7), .CK(clk), .Q(u_0_2[1]), .QN() );
  DFF_X1 rand_reg_1_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[0]), 
        .QN() );
  DFF_X1 u_0_2_reg_0_ ( .D(N1), .CK(clk), .Q(u_0_2[0]), .QN() );
  DFF_X1 rand_reg_4_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[4]), 
        .QN() );
  DFF_X1 u_2_0_reg_4_ ( .D(N28), .CK(clk), .Q(u_2_0[4]), .QN() );
  DFF_X1 rand_reg_4_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[3]), 
        .QN() );
  DFF_X1 u_2_0_reg_3_ ( .D(N22), .CK(clk), .Q(u_2_0[3]), .QN() );
  DFF_X1 rand_reg_4_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[2]), 
        .QN() );
  DFF_X1 u_2_0_reg_2_ ( .D(N16), .CK(clk), .Q(u_2_0[2]), .QN() );
  DFF_X1 rand_reg_4_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[1]), 
        .QN() );
  DFF_X1 u_2_0_reg_1_ ( .D(N10), .CK(clk), .Q(u_2_0[1]), .QN() );
  DFF_X1 rand_reg_4_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[0]), 
        .QN() );
  DFF_X1 u_2_0_reg_0_ ( .D(N4), .CK(clk), .Q(u_2_0[0]), .QN() );
  DFF_X1 b_reg_0_reg_4_ ( .D(io_b_0[4]), .CK(clk), .Q(b_reg_0[4]), .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_0_ ( .D(N66), .CK(clk), .Q(n_zz_io_c_0_16_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_3_ ( .D(io_b_0[3]), .CK(clk), .Q(b_reg_0[3]), .QN() );
  DFF_X1 u_zz_io_c_0_15_reg_0_ ( .D(N57), .CK(clk), .Q(n_zz_io_c_0_12_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_2_ ( .D(io_b_0[2]), .CK(clk), .Q(b_reg_0[2]), .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_0_ ( .D(N48), .CK(clk), .Q(n_zz_io_c_0_8_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_1_ ( .D(io_b_0[1]), .CK(clk), .Q(b_reg_0[1]), .QN() );
  DFF_X1 b_reg_0_reg_0_ ( .D(io_b_0[0]), .CK(clk), .Q(b_reg_0[0]), .QN() );
  DFF_X1 u_zz_io_c_1_7_reg_2_ ( .D(N44), .CK(clk), .Q(n_zz_io_c_1_7[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_7_reg_1_ ( .D(N43), .CK(clk), .Q(n_zz_io_c_1_7[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_7_reg_0_ ( .D(N42), .CK(clk), .Q(n_zz_io_c_1_4_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_7_reg_2_ ( .D(N41), .CK(clk), .Q(n_zz_io_c_0_7[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_7_reg_1_ ( .D(N40), .CK(clk), .Q(n_zz_io_c_0_7[1]), .QN()
         );
  DFF_X1 u_zz_io_c_0_7_reg_0_ ( .D(N39), .CK(clk), .Q(n_zz_io_c_0_4_0_), .QN()
         );
  DFF_X1 u_zz_io_c_2_3_reg_2_ ( .D(N38), .CK(clk), .Q(n_zz_io_c_2_3[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_3_reg_1_ ( .D(N37), .CK(clk), .Q(n_zz_io_c_2_3[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_3_reg_0_ ( .D(N36), .CK(clk), .Q(n_zz_io_c_2_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_3_reg_2_ ( .D(N35), .CK(clk), .Q(n_zz_io_c_1_3[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_3_reg_1_ ( .D(N34), .CK(clk), .Q(n_zz_io_c_1_3[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_3_reg_0_ ( .D(N33), .CK(clk), .Q(n_zz_io_c_1_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_3_reg_2_ ( .D(N32), .CK(clk), .Q(n_zz_io_c_0_3[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_3_reg_1_ ( .D(N31), .CK(clk), .Q(n_zz_io_c_0_3[1]), .QN()
         );
  DFF_X1 u_zz_io_c_0_3_reg_0_ ( .D(N30), .CK(clk), .Q(n_zz_io_c_0_0_), .QN()
         );
  XOR2_X2 U3 ( .A(io_rand[2]), .B(io_b_1[4]), .Z(v_1_2_1[4]) );
  XOR2_X2 U4 ( .A(io_rand[2]), .B(io_b_1[3]), .Z(v_1_2_1[3]) );
  XOR2_X2 U5 ( .A(io_rand[2]), .B(io_b_1[2]), .Z(v_1_2_1[2]) );
  XOR2_X2 U6 ( .A(io_rand[2]), .B(io_b_1[1]), .Z(v_1_2_1[1]) );
  XOR2_X2 U7 ( .A(io_rand[2]), .B(io_b_1[0]), .Z(v_1_2_1[0]) );
  XOR2_X2 U8 ( .A(io_rand[1]), .B(io_b_0[4]), .Z(v_1_2_0[4]) );
  XOR2_X2 U9 ( .A(io_rand[1]), .B(io_b_0[3]), .Z(v_1_2_0[3]) );
  XOR2_X2 U10 ( .A(io_rand[1]), .B(io_b_0[2]), .Z(v_1_2_0[2]) );
  XOR2_X2 U11 ( .A(io_rand[1]), .B(io_b_0[1]), .Z(v_1_2_0[1]) );
  XOR2_X2 U12 ( .A(io_rand[1]), .B(io_b_0[0]), .Z(v_1_2_0[0]) );
  XOR2_X2 U13 ( .A(io_rand[2]), .B(io_b_2[4]), .Z(v_1_1_2[4]) );
  XOR2_X2 U14 ( .A(io_rand[2]), .B(io_b_2[3]), .Z(v_1_1_2[3]) );
  XOR2_X2 U15 ( .A(io_rand[2]), .B(io_b_2[2]), .Z(v_1_1_2[2]) );
  XOR2_X2 U16 ( .A(io_rand[2]), .B(io_b_2[1]), .Z(v_1_1_2[1]) );
  XOR2_X2 U17 ( .A(io_rand[2]), .B(io_b_2[0]), .Z(v_1_1_2[0]) );
  XOR2_X2 U18 ( .A(io_rand[0]), .B(io_b_0[4]), .Z(v_1_1_0[4]) );
  XOR2_X2 U19 ( .A(io_rand[0]), .B(io_b_0[3]), .Z(v_1_1_0[3]) );
  XOR2_X2 U20 ( .A(io_rand[0]), .B(io_b_0[2]), .Z(v_1_1_0[2]) );
  XOR2_X2 U21 ( .A(io_rand[0]), .B(io_b_0[1]), .Z(v_1_1_0[1]) );
  XOR2_X2 U22 ( .A(io_rand[0]), .B(io_b_0[0]), .Z(v_1_1_0[0]) );
  XOR2_X2 U23 ( .A(io_rand[1]), .B(io_b_2[4]), .Z(v_1_0_2[4]) );
  XOR2_X2 U24 ( .A(io_rand[1]), .B(io_b_2[3]), .Z(v_1_0_2[3]) );
  XOR2_X2 U25 ( .A(io_rand[1]), .B(io_b_2[2]), .Z(v_1_0_2[2]) );
  XOR2_X2 U26 ( .A(io_rand[1]), .B(io_b_2[1]), .Z(v_1_0_2[1]) );
  XOR2_X2 U27 ( .A(io_rand[1]), .B(io_b_2[0]), .Z(v_1_0_2[0]) );
  XOR2_X2 U28 ( .A(io_rand[0]), .B(io_b_1[4]), .Z(v_1_0_1[4]) );
  XOR2_X2 U29 ( .A(io_rand[0]), .B(io_b_1[3]), .Z(v_1_0_1[3]) );
  XOR2_X2 U30 ( .A(io_rand[0]), .B(io_b_1[2]), .Z(v_1_0_1[2]) );
  XOR2_X2 U31 ( .A(io_rand[0]), .B(io_b_1[1]), .Z(v_1_0_1[1]) );
  XOR2_X2 U32 ( .A(io_rand[0]), .B(io_b_1[0]), .Z(v_1_0_1[0]) );
  AND2_X1 U138 ( .A1(b_reg_0[0]), .A2(io_a_0[0]), .ZN(N30) );
  AND2_X1 U139 ( .A1(cor_port_v_0_1[0]), .A2(io_a_0[0]), .ZN(N31) );
  AND2_X1 U140 ( .A1(b_reg_1[0]), .A2(io_a_1[0]), .ZN(N33) );
  AND2_X1 U141 ( .A1(cor_port_v_1_0[0]), .A2(io_a_1[0]), .ZN(N34) );
  AND2_X1 U142 ( .A1(b_reg_2[0]), .A2(io_a_2[0]), .ZN(N36) );
  AND2_X1 U143 ( .A1(cor_port_v_2_0[0]), .A2(io_a_2[0]), .ZN(N37) );
  AND2_X1 U144 ( .A1(b_reg_0[1]), .A2(io_a_0[1]), .ZN(N39) );
  AND2_X1 U145 ( .A1(cor_port_v_0_1[1]), .A2(io_a_0[1]), .ZN(N40) );
  AND2_X1 U146 ( .A1(b_reg_1[1]), .A2(io_a_1[1]), .ZN(N42) );
  AND2_X1 U147 ( .A1(cor_port_v_1_0[1]), .A2(io_a_1[1]), .ZN(N43) );
  AND2_X1 U148 ( .A1(b_reg_0[2]), .A2(io_a_0[2]), .ZN(N48) );
  AND2_X1 U149 ( .A1(b_reg_0[3]), .A2(io_a_0[3]), .ZN(N57) );
  AND2_X1 U150 ( .A1(b_reg_0[4]), .A2(io_a_0[4]), .ZN(N66) );
  AND2_X1 U151 ( .A1(b_reg_2[1]), .A2(io_a_2[1]), .ZN(N45) );
  AND2_X1 U152 ( .A1(cor_port_v_2_0[1]), .A2(io_a_2[1]), .ZN(N46) );
  AND2_X1 U153 ( .A1(cor_port_v_0_1[2]), .A2(io_a_0[2]), .ZN(N49) );
  AND2_X1 U154 ( .A1(b_reg_1[2]), .A2(io_a_1[2]), .ZN(N51) );
  AND2_X1 U155 ( .A1(cor_port_v_1_0[2]), .A2(io_a_1[2]), .ZN(N52) );
  AND2_X1 U156 ( .A1(b_reg_2[2]), .A2(io_a_2[2]), .ZN(N54) );
  AND2_X1 U157 ( .A1(cor_port_v_2_0[2]), .A2(io_a_2[2]), .ZN(N55) );
  AND2_X1 U158 ( .A1(cor_port_v_0_1[3]), .A2(io_a_0[3]), .ZN(N58) );
  AND2_X1 U159 ( .A1(b_reg_1[3]), .A2(io_a_1[3]), .ZN(N60) );
  AND2_X1 U160 ( .A1(cor_port_v_1_0[3]), .A2(io_a_1[3]), .ZN(N61) );
  AND2_X1 U161 ( .A1(b_reg_2[3]), .A2(io_a_2[3]), .ZN(N63) );
  AND2_X1 U162 ( .A1(cor_port_v_2_0[3]), .A2(io_a_2[3]), .ZN(N64) );
  AND2_X1 U163 ( .A1(cor_port_v_0_1[4]), .A2(io_a_0[4]), .ZN(N67) );
  AND2_X1 U164 ( .A1(b_reg_1[4]), .A2(io_a_1[4]), .ZN(N69) );
  AND2_X1 U165 ( .A1(cor_port_v_1_0[4]), .A2(io_a_1[4]), .ZN(N70) );
  AND2_X1 U166 ( .A1(b_reg_2[4]), .A2(io_a_2[4]), .ZN(N72) );
  AND2_X1 U167 ( .A1(cor_port_v_2_0[4]), .A2(io_a_2[4]), .ZN(N73) );
  AND2_X1 U168 ( .A1(io_a_0[0]), .A2(cor_port_v_0_2[0]), .ZN(N32) );
  AND2_X1 U169 ( .A1(io_a_1[0]), .A2(cor_port_v_1_2[0]), .ZN(N35) );
  AND2_X1 U170 ( .A1(io_a_2[0]), .A2(cor_port_v_2_1[0]), .ZN(N38) );
  AND2_X1 U171 ( .A1(io_a_0[1]), .A2(cor_port_v_0_2[1]), .ZN(N41) );
  AND2_X1 U172 ( .A1(io_a_1[1]), .A2(cor_port_v_1_2[1]), .ZN(N44) );
  AND2_X1 U173 ( .A1(simpleNot_34_port_z), .A2(rand_reg_4[0]), .ZN(N4) );
  AND2_X1 U174 ( .A1(simpleNot_40_port_z), .A2(rand_reg_4[1]), .ZN(N10) );
  AND2_X1 U175 ( .A1(simpleNot_46_port_z), .A2(rand_reg_4[2]), .ZN(N16) );
  AND2_X1 U176 ( .A1(simpleNot_52_port_z), .A2(rand_reg_4[3]), .ZN(N22) );
  AND2_X1 U177 ( .A1(simpleNot_58_port_z), .A2(rand_reg_4[4]), .ZN(N28) );
  AND2_X1 U178 ( .A1(simpleNot_31_port_z), .A2(rand_reg_1[0]), .ZN(N1) );
  AND2_X1 U179 ( .A1(simpleNot_37_port_z), .A2(rand_reg_1[1]), .ZN(N7) );
  AND2_X1 U180 ( .A1(simpleNot_43_port_z), .A2(rand_reg_1[2]), .ZN(N13) );
  AND2_X1 U181 ( .A1(simpleNot_49_port_z), .A2(rand_reg_1[3]), .ZN(N19) );
  AND2_X1 U182 ( .A1(simpleNot_55_port_z), .A2(rand_reg_1[4]), .ZN(N25) );
  AND2_X1 U183 ( .A1(io_a_2[1]), .A2(cor_port_v_2_1[1]), .ZN(N47) );
  AND2_X1 U184 ( .A1(simpleNot_33_port_z), .A2(rand_reg_2[0]), .ZN(N3) );
  AND2_X1 U185 ( .A1(simpleNot_39_port_z), .A2(rand_reg_2[1]), .ZN(N9) );
  AND2_X1 U186 ( .A1(simpleNot_45_port_z), .A2(rand_reg_2[2]), .ZN(N15) );
  AND2_X1 U187 ( .A1(simpleNot_51_port_z), .A2(rand_reg_2[3]), .ZN(N21) );
  AND2_X1 U188 ( .A1(simpleNot_57_port_z), .A2(rand_reg_2[4]), .ZN(N27) );
  AND2_X1 U189 ( .A1(simpleNot_32_port_z), .A2(rand_reg_3[0]), .ZN(N2) );
  AND2_X1 U190 ( .A1(simpleNot_38_port_z), .A2(rand_reg_3[1]), .ZN(N8) );
  AND2_X1 U191 ( .A1(simpleNot_44_port_z), .A2(rand_reg_3[2]), .ZN(N14) );
  AND2_X1 U192 ( .A1(simpleNot_50_port_z), .A2(rand_reg_3[3]), .ZN(N20) );
  AND2_X1 U193 ( .A1(simpleNot_56_port_z), .A2(rand_reg_3[4]), .ZN(N26) );
  AND2_X1 U194 ( .A1(simpleNot_30_port_z), .A2(rand_reg_0[0]), .ZN(N0) );
  AND2_X1 U195 ( .A1(simpleNot_36_port_z), .A2(rand_reg_0[1]), .ZN(N6) );
  AND2_X1 U196 ( .A1(simpleNot_42_port_z), .A2(rand_reg_0[2]), .ZN(N12) );
  AND2_X1 U197 ( .A1(simpleNot_48_port_z), .A2(rand_reg_0[3]), .ZN(N18) );
  AND2_X1 U198 ( .A1(simpleNot_54_port_z), .A2(rand_reg_0[4]), .ZN(N24) );
  AND2_X1 U199 ( .A1(io_a_0[2]), .A2(cor_port_v_0_2[2]), .ZN(N50) );
  AND2_X1 U200 ( .A1(io_a_1[2]), .A2(cor_port_v_1_2[2]), .ZN(N53) );
  AND2_X1 U201 ( .A1(simpleNot_35_port_z), .A2(rand_reg_5[0]), .ZN(N5) );
  AND2_X1 U202 ( .A1(simpleNot_41_port_z), .A2(rand_reg_5[1]), .ZN(N11) );
  AND2_X1 U203 ( .A1(simpleNot_47_port_z), .A2(rand_reg_5[2]), .ZN(N17) );
  AND2_X1 U204 ( .A1(simpleNot_53_port_z), .A2(rand_reg_5[3]), .ZN(N23) );
  AND2_X1 U205 ( .A1(simpleNot_59_port_z), .A2(rand_reg_5[4]), .ZN(N29) );
  AND2_X1 U206 ( .A1(io_a_2[2]), .A2(cor_port_v_2_1[2]), .ZN(N56) );
  AND2_X1 U207 ( .A1(io_a_0[3]), .A2(cor_port_v_0_2[3]), .ZN(N59) );
  AND2_X1 U208 ( .A1(io_a_1[3]), .A2(cor_port_v_1_2[3]), .ZN(N62) );
  AND2_X1 U209 ( .A1(io_a_2[3]), .A2(cor_port_v_2_1[3]), .ZN(N65) );
  AND2_X1 U210 ( .A1(io_a_0[4]), .A2(cor_port_v_0_2[4]), .ZN(N68) );
  AND2_X1 U211 ( .A1(io_a_1[4]), .A2(cor_port_v_1_2[4]), .ZN(N71) );
  AND2_X1 U212 ( .A1(io_a_2[4]), .A2(cor_port_v_2_1[4]), .ZN(N74) );
  XOR2_X1 U213 ( .A(n_zz_io_c_2_0_), .B(n5), .Z(io_c_2[0]) );
  XOR2_X1 U214 ( .A(simpleXor_35_port_z), .B(simpleXor_34_port_z), .Z(n5) );
  XOR2_X1 U215 ( .A(n_zz_io_c_2_4_0_), .B(n4), .Z(io_c_2[1]) );
  XOR2_X1 U216 ( .A(simpleXor_41_port_z), .B(simpleXor_40_port_z), .Z(n4) );
  XOR2_X1 U217 ( .A(n_zz_io_c_2_8_0_), .B(n3), .Z(io_c_2[2]) );
  XOR2_X1 U218 ( .A(simpleXor_47_port_z), .B(simpleXor_46_port_z), .Z(n3) );
  XOR2_X1 U219 ( .A(n_zz_io_c_2_12_0_), .B(n2), .Z(io_c_2[3]) );
  XOR2_X1 U220 ( .A(simpleXor_53_port_z), .B(simpleXor_52_port_z), .Z(n2) );
  XOR2_X1 U221 ( .A(n_zz_io_c_2_16_0_), .B(n1), .Z(io_c_2[4]) );
  XOR2_X1 U222 ( .A(simpleXor_59_port_z), .B(simpleXor_58_port_z), .Z(n1) );
  XOR2_X1 U223 ( .A(n_zz_io_c_1_0_), .B(n10), .Z(io_c_1[0]) );
  XOR2_X1 U224 ( .A(simpleXor_33_port_z), .B(simpleXor_32_port_z), .Z(n10) );
  XOR2_X1 U225 ( .A(n_zz_io_c_1_4_0_), .B(n9), .Z(io_c_1[1]) );
  XOR2_X1 U226 ( .A(simpleXor_39_port_z), .B(simpleXor_38_port_z), .Z(n9) );
  XOR2_X1 U227 ( .A(n_zz_io_c_1_8_0_), .B(n8), .Z(io_c_1[2]) );
  XOR2_X1 U228 ( .A(simpleXor_45_port_z), .B(simpleXor_44_port_z), .Z(n8) );
  XOR2_X1 U229 ( .A(n_zz_io_c_1_12_0_), .B(n7), .Z(io_c_1[3]) );
  XOR2_X1 U230 ( .A(simpleXor_51_port_z), .B(simpleXor_50_port_z), .Z(n7) );
  XOR2_X1 U231 ( .A(n_zz_io_c_1_16_0_), .B(n6), .Z(io_c_1[4]) );
  XOR2_X1 U232 ( .A(simpleXor_57_port_z), .B(simpleXor_56_port_z), .Z(n6) );
  XOR2_X1 U233 ( .A(n_zz_io_c_0_0_), .B(n15), .Z(io_c_0[0]) );
  XOR2_X1 U234 ( .A(simpleXor_31_port_z), .B(simpleXor_30_port_z), .Z(n15) );
  XOR2_X1 U235 ( .A(n_zz_io_c_0_4_0_), .B(n14), .Z(io_c_0[1]) );
  XOR2_X1 U236 ( .A(simpleXor_37_port_z), .B(simpleXor_36_port_z), .Z(n14) );
  XOR2_X1 U237 ( .A(n_zz_io_c_0_8_0_), .B(n13), .Z(io_c_0[2]) );
  XOR2_X1 U238 ( .A(simpleXor_43_port_z), .B(simpleXor_42_port_z), .Z(n13) );
  XOR2_X1 U239 ( .A(n_zz_io_c_0_12_0_), .B(n12), .Z(io_c_0[3]) );
  XOR2_X1 U240 ( .A(simpleXor_49_port_z), .B(simpleXor_48_port_z), .Z(n12) );
  XOR2_X1 U241 ( .A(n_zz_io_c_0_16_0_), .B(n11), .Z(io_c_0[4]) );
  XOR2_X1 U242 ( .A(simpleXor_55_port_z), .B(simpleXor_54_port_z), .Z(n11) );
  INV_X1 simpleNot_30_U1 ( .A(io_a_0[0]), .ZN(simpleNot_30_port_z) );
  INV_X1 simpleNot_31_U1 ( .A(io_a_0[0]), .ZN(simpleNot_31_port_z) );
  INV_X1 simpleNot_32_U1 ( .A(io_a_1[0]), .ZN(simpleNot_32_port_z) );
  INV_X1 simpleNot_33_U1 ( .A(io_a_1[0]), .ZN(simpleNot_33_port_z) );
  INV_X1 simpleNot_34_U1 ( .A(io_a_2[0]), .ZN(simpleNot_34_port_z) );
  INV_X1 simpleNot_35_U1 ( .A(io_a_2[0]), .ZN(simpleNot_35_port_z) );
  INV_X1 simpleNot_36_U1 ( .A(io_a_0[1]), .ZN(simpleNot_36_port_z) );
  INV_X1 simpleNot_37_U1 ( .A(io_a_0[1]), .ZN(simpleNot_37_port_z) );
  INV_X1 simpleNot_38_U1 ( .A(io_a_1[1]), .ZN(simpleNot_38_port_z) );
  INV_X1 simpleNot_39_U1 ( .A(io_a_1[1]), .ZN(simpleNot_39_port_z) );
  INV_X1 simpleNot_40_U1 ( .A(io_a_2[1]), .ZN(simpleNot_40_port_z) );
  INV_X1 simpleNot_41_U1 ( .A(io_a_2[1]), .ZN(simpleNot_41_port_z) );
  INV_X1 simpleNot_42_U1 ( .A(io_a_0[2]), .ZN(simpleNot_42_port_z) );
  INV_X1 simpleNot_43_U1 ( .A(io_a_0[2]), .ZN(simpleNot_43_port_z) );
  INV_X1 simpleNot_44_U1 ( .A(io_a_1[2]), .ZN(simpleNot_44_port_z) );
  INV_X1 simpleNot_45_U1 ( .A(io_a_1[2]), .ZN(simpleNot_45_port_z) );
  INV_X1 simpleNot_46_U1 ( .A(io_a_2[2]), .ZN(simpleNot_46_port_z) );
  INV_X1 simpleNot_47_U1 ( .A(io_a_2[2]), .ZN(simpleNot_47_port_z) );
  INV_X1 simpleNot_48_U1 ( .A(io_a_0[3]), .ZN(simpleNot_48_port_z) );
  INV_X1 simpleNot_49_U1 ( .A(io_a_0[3]), .ZN(simpleNot_49_port_z) );
  INV_X1 simpleNot_50_U1 ( .A(io_a_1[3]), .ZN(simpleNot_50_port_z) );
  INV_X1 simpleNot_51_U1 ( .A(io_a_1[3]), .ZN(simpleNot_51_port_z) );
  INV_X1 simpleNot_52_U1 ( .A(io_a_2[3]), .ZN(simpleNot_52_port_z) );
  INV_X1 simpleNot_53_U1 ( .A(io_a_2[3]), .ZN(simpleNot_53_port_z) );
  INV_X1 simpleNot_54_U1 ( .A(io_a_0[4]), .ZN(simpleNot_54_port_z) );
  INV_X1 simpleNot_55_U1 ( .A(io_a_0[4]), .ZN(simpleNot_55_port_z) );
  INV_X1 simpleNot_56_U1 ( .A(io_a_1[4]), .ZN(simpleNot_56_port_z) );
  INV_X1 simpleNot_57_U1 ( .A(io_a_1[4]), .ZN(simpleNot_57_port_z) );
  INV_X1 simpleNot_58_U1 ( .A(io_a_2[4]), .ZN(simpleNot_58_port_z) );
  INV_X1 simpleNot_59_U1 ( .A(io_a_2[4]), .ZN(simpleNot_59_port_z) );
  DFF_X1 cor_m_2_1_reg_0_ ( .D(cor_maj_55_port_o), .CK(clk), .Q(
        cor_port_v_2_1[0]), .QN() );
  DFF_X1 cor_m_2_1_reg_1_ ( .D(cor_maj_56_port_o), .CK(clk), .Q(
        cor_port_v_2_1[1]), .QN() );
  DFF_X1 cor_m_2_1_reg_2_ ( .D(cor_maj_57_port_o), .CK(clk), .Q(
        cor_port_v_2_1[2]), .QN() );
  DFF_X1 cor_m_2_1_reg_3_ ( .D(cor_maj_58_port_o), .CK(clk), .Q(
        cor_port_v_2_1[3]), .QN() );
  DFF_X1 cor_m_2_1_reg_4_ ( .D(cor_maj_59_port_o), .CK(clk), .Q(
        cor_port_v_2_1[4]), .QN() );
  DFF_X1 cor_m_2_0_reg_0_ ( .D(cor_maj_50_port_o), .CK(clk), .Q(
        cor_port_v_2_0[0]), .QN() );
  DFF_X1 cor_m_2_0_reg_1_ ( .D(cor_maj_51_port_o), .CK(clk), .Q(
        cor_port_v_2_0[1]), .QN() );
  DFF_X1 cor_m_2_0_reg_2_ ( .D(cor_maj_52_port_o), .CK(clk), .Q(
        cor_port_v_2_0[2]), .QN() );
  DFF_X1 cor_m_2_0_reg_3_ ( .D(cor_maj_53_port_o), .CK(clk), .Q(
        cor_port_v_2_0[3]), .QN() );
  DFF_X1 cor_m_2_0_reg_4_ ( .D(cor_maj_54_port_o), .CK(clk), .Q(
        cor_port_v_2_0[4]), .QN() );
  DFF_X1 cor_m_1_2_reg_0_ ( .D(cor_maj_45_port_o), .CK(clk), .Q(
        cor_port_v_1_2[0]), .QN() );
  DFF_X1 cor_m_1_2_reg_1_ ( .D(cor_maj_46_port_o), .CK(clk), .Q(
        cor_port_v_1_2[1]), .QN() );
  DFF_X1 cor_m_1_2_reg_2_ ( .D(cor_maj_47_port_o), .CK(clk), .Q(
        cor_port_v_1_2[2]), .QN() );
  DFF_X1 cor_m_1_2_reg_3_ ( .D(cor_maj_48_port_o), .CK(clk), .Q(
        cor_port_v_1_2[3]), .QN() );
  DFF_X1 cor_m_1_2_reg_4_ ( .D(cor_maj_49_port_o), .CK(clk), .Q(
        cor_port_v_1_2[4]), .QN() );
  DFF_X1 cor_m_1_0_reg_0_ ( .D(cor_maj_40_port_o), .CK(clk), .Q(
        cor_port_v_1_0[0]), .QN() );
  DFF_X1 cor_m_1_0_reg_1_ ( .D(cor_maj_41_port_o), .CK(clk), .Q(
        cor_port_v_1_0[1]), .QN() );
  DFF_X1 cor_m_1_0_reg_2_ ( .D(cor_maj_42_port_o), .CK(clk), .Q(
        cor_port_v_1_0[2]), .QN() );
  DFF_X1 cor_m_1_0_reg_3_ ( .D(cor_maj_43_port_o), .CK(clk), .Q(
        cor_port_v_1_0[3]), .QN() );
  DFF_X1 cor_m_1_0_reg_4_ ( .D(cor_maj_44_port_o), .CK(clk), .Q(
        cor_port_v_1_0[4]), .QN() );
  DFF_X1 cor_m_0_2_reg_0_ ( .D(cor_maj_35_port_o), .CK(clk), .Q(
        cor_port_v_0_2[0]), .QN() );
  DFF_X1 cor_m_0_2_reg_1_ ( .D(cor_maj_36_port_o), .CK(clk), .Q(
        cor_port_v_0_2[1]), .QN() );
  DFF_X1 cor_m_0_2_reg_2_ ( .D(cor_maj_37_port_o), .CK(clk), .Q(
        cor_port_v_0_2[2]), .QN() );
  DFF_X1 cor_m_0_2_reg_3_ ( .D(cor_maj_38_port_o), .CK(clk), .Q(
        cor_port_v_0_2[3]), .QN() );
  DFF_X1 cor_m_0_2_reg_4_ ( .D(cor_maj_39_port_o), .CK(clk), .Q(
        cor_port_v_0_2[4]), .QN() );
  DFF_X1 cor_m_0_1_reg_0_ ( .D(cor_maj_30_port_o), .CK(clk), .Q(
        cor_port_v_0_1[0]), .QN() );
  DFF_X1 cor_m_0_1_reg_1_ ( .D(cor_maj_31_port_o), .CK(clk), .Q(
        cor_port_v_0_1[1]), .QN() );
  DFF_X1 cor_m_0_1_reg_2_ ( .D(cor_maj_32_port_o), .CK(clk), .Q(
        cor_port_v_0_1[2]), .QN() );
  DFF_X1 cor_m_0_1_reg_3_ ( .D(cor_maj_33_port_o), .CK(clk), .Q(
        cor_port_v_0_1[3]), .QN() );
  DFF_X1 cor_m_0_1_reg_4_ ( .D(cor_maj_34_port_o), .CK(clk), .Q(
        cor_port_v_0_1[4]), .QN() );
  NAND2_X1 cor_maj_30_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_30_n9) );
  NAND2_X1 cor_maj_30_U14 ( .A1(cor_maj_30_n6), .A2(cor_maj_30_n5), .ZN(
        cor_maj_30_n10) );
  NAND2_X1 cor_maj_30_U13 ( .A1(cor_maj_30_n9), .A2(cor_maj_30_n10), .ZN(
        cor_maj_30_n8) );
  NAND2_X1 cor_maj_30_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_30_n11), .ZN(
        cor_maj_30_n13) );
  NAND2_X1 cor_maj_30_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_30_n12) );
  NAND2_X1 cor_maj_30_U10 ( .A1(cor_maj_30_n12), .A2(cor_maj_30_n13), .ZN(
        cor_maj_30_n7) );
  XOR2_X1 cor_maj_30_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_30_n5) );
  XOR2_X1 cor_maj_30_U8 ( .A(v_1_0_1[2]), .B(cor_maj_30_n11), .Z(cor_maj_30_n6) );
  XOR2_X1 cor_maj_30_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_30_n11)
         );
  OR2_X1 cor_maj_30_U6 ( .A1(cor_maj_30_n7), .A2(cor_maj_30_n8), .ZN(
        cor_maj_30_n3) );
  NAND2_X1 cor_maj_30_U5 ( .A1(cor_maj_30_n3), .A2(cor_maj_30_n4), .ZN(
        cor_maj_30_n2) );
  NAND2_X1 cor_maj_30_U4 ( .A1(cor_maj_30_n7), .A2(cor_maj_30_n8), .ZN(
        cor_maj_30_n1) );
  NAND2_X1 cor_maj_30_U3 ( .A1(cor_maj_30_n1), .A2(cor_maj_30_n2), .ZN(
        cor_maj_30_port_o) );
  XOR2_X1 cor_maj_30_U2 ( .A(cor_maj_30_n5), .B(cor_maj_30_n6), .Z(
        cor_maj_30_n4) );
  NAND2_X1 cor_maj_31_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_31_n18) );
  NAND2_X1 cor_maj_31_U14 ( .A1(cor_maj_31_n21), .A2(cor_maj_31_n22), .ZN(
        cor_maj_31_n17) );
  NAND2_X1 cor_maj_31_U13 ( .A1(cor_maj_31_n18), .A2(cor_maj_31_n17), .ZN(
        cor_maj_31_n19) );
  NAND2_X1 cor_maj_31_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_31_n16), .ZN(
        cor_maj_31_n14) );
  NAND2_X1 cor_maj_31_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_31_n15) );
  NAND2_X1 cor_maj_31_U10 ( .A1(cor_maj_31_n15), .A2(cor_maj_31_n14), .ZN(
        cor_maj_31_n20) );
  XOR2_X1 cor_maj_31_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_31_n22)
         );
  XOR2_X1 cor_maj_31_U8 ( .A(v_1_0_1[2]), .B(cor_maj_31_n16), .Z(
        cor_maj_31_n21) );
  XOR2_X1 cor_maj_31_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_31_n16)
         );
  OR2_X1 cor_maj_31_U6 ( .A1(cor_maj_31_n20), .A2(cor_maj_31_n19), .ZN(
        cor_maj_31_n24) );
  NAND2_X1 cor_maj_31_U5 ( .A1(cor_maj_31_n24), .A2(cor_maj_31_n23), .ZN(
        cor_maj_31_n25) );
  NAND2_X1 cor_maj_31_U4 ( .A1(cor_maj_31_n20), .A2(cor_maj_31_n19), .ZN(
        cor_maj_31_n26) );
  NAND2_X1 cor_maj_31_U3 ( .A1(cor_maj_31_n26), .A2(cor_maj_31_n25), .ZN(
        cor_maj_31_port_o) );
  XOR2_X1 cor_maj_31_U2 ( .A(cor_maj_31_n22), .B(cor_maj_31_n21), .Z(
        cor_maj_31_n23) );
  NAND2_X1 cor_maj_32_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_32_n18) );
  NAND2_X1 cor_maj_32_U14 ( .A1(cor_maj_32_n21), .A2(cor_maj_32_n22), .ZN(
        cor_maj_32_n17) );
  NAND2_X1 cor_maj_32_U13 ( .A1(cor_maj_32_n18), .A2(cor_maj_32_n17), .ZN(
        cor_maj_32_n19) );
  NAND2_X1 cor_maj_32_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_32_n16), .ZN(
        cor_maj_32_n14) );
  NAND2_X1 cor_maj_32_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_32_n15) );
  NAND2_X1 cor_maj_32_U10 ( .A1(cor_maj_32_n15), .A2(cor_maj_32_n14), .ZN(
        cor_maj_32_n20) );
  XOR2_X1 cor_maj_32_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_32_n22)
         );
  XOR2_X1 cor_maj_32_U8 ( .A(v_1_0_1[2]), .B(cor_maj_32_n16), .Z(
        cor_maj_32_n21) );
  XOR2_X1 cor_maj_32_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_32_n16)
         );
  OR2_X1 cor_maj_32_U6 ( .A1(cor_maj_32_n20), .A2(cor_maj_32_n19), .ZN(
        cor_maj_32_n24) );
  NAND2_X1 cor_maj_32_U5 ( .A1(cor_maj_32_n24), .A2(cor_maj_32_n23), .ZN(
        cor_maj_32_n25) );
  NAND2_X1 cor_maj_32_U4 ( .A1(cor_maj_32_n20), .A2(cor_maj_32_n19), .ZN(
        cor_maj_32_n26) );
  NAND2_X1 cor_maj_32_U3 ( .A1(cor_maj_32_n26), .A2(cor_maj_32_n25), .ZN(
        cor_maj_32_port_o) );
  XOR2_X1 cor_maj_32_U2 ( .A(cor_maj_32_n22), .B(cor_maj_32_n21), .Z(
        cor_maj_32_n23) );
  NAND2_X1 cor_maj_33_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_33_n18) );
  NAND2_X1 cor_maj_33_U14 ( .A1(cor_maj_33_n21), .A2(cor_maj_33_n22), .ZN(
        cor_maj_33_n17) );
  NAND2_X1 cor_maj_33_U13 ( .A1(cor_maj_33_n18), .A2(cor_maj_33_n17), .ZN(
        cor_maj_33_n19) );
  NAND2_X1 cor_maj_33_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_33_n16), .ZN(
        cor_maj_33_n14) );
  NAND2_X1 cor_maj_33_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_33_n15) );
  NAND2_X1 cor_maj_33_U10 ( .A1(cor_maj_33_n15), .A2(cor_maj_33_n14), .ZN(
        cor_maj_33_n20) );
  XOR2_X1 cor_maj_33_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_33_n22)
         );
  XOR2_X1 cor_maj_33_U8 ( .A(v_1_0_1[2]), .B(cor_maj_33_n16), .Z(
        cor_maj_33_n21) );
  XOR2_X1 cor_maj_33_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_33_n16)
         );
  OR2_X1 cor_maj_33_U6 ( .A1(cor_maj_33_n20), .A2(cor_maj_33_n19), .ZN(
        cor_maj_33_n24) );
  NAND2_X1 cor_maj_33_U5 ( .A1(cor_maj_33_n24), .A2(cor_maj_33_n23), .ZN(
        cor_maj_33_n25) );
  NAND2_X1 cor_maj_33_U4 ( .A1(cor_maj_33_n20), .A2(cor_maj_33_n19), .ZN(
        cor_maj_33_n26) );
  NAND2_X1 cor_maj_33_U3 ( .A1(cor_maj_33_n26), .A2(cor_maj_33_n25), .ZN(
        cor_maj_33_port_o) );
  XOR2_X1 cor_maj_33_U2 ( .A(cor_maj_33_n22), .B(cor_maj_33_n21), .Z(
        cor_maj_33_n23) );
  NAND2_X1 cor_maj_34_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_34_n18) );
  NAND2_X1 cor_maj_34_U14 ( .A1(cor_maj_34_n21), .A2(cor_maj_34_n22), .ZN(
        cor_maj_34_n17) );
  NAND2_X1 cor_maj_34_U13 ( .A1(cor_maj_34_n18), .A2(cor_maj_34_n17), .ZN(
        cor_maj_34_n19) );
  NAND2_X1 cor_maj_34_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_34_n16), .ZN(
        cor_maj_34_n14) );
  NAND2_X1 cor_maj_34_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_34_n15) );
  NAND2_X1 cor_maj_34_U10 ( .A1(cor_maj_34_n15), .A2(cor_maj_34_n14), .ZN(
        cor_maj_34_n20) );
  XOR2_X1 cor_maj_34_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_34_n22)
         );
  XOR2_X1 cor_maj_34_U8 ( .A(v_1_0_1[2]), .B(cor_maj_34_n16), .Z(
        cor_maj_34_n21) );
  XOR2_X1 cor_maj_34_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_34_n16)
         );
  OR2_X1 cor_maj_34_U6 ( .A1(cor_maj_34_n20), .A2(cor_maj_34_n19), .ZN(
        cor_maj_34_n24) );
  NAND2_X1 cor_maj_34_U5 ( .A1(cor_maj_34_n24), .A2(cor_maj_34_n23), .ZN(
        cor_maj_34_n25) );
  NAND2_X1 cor_maj_34_U4 ( .A1(cor_maj_34_n20), .A2(cor_maj_34_n19), .ZN(
        cor_maj_34_n26) );
  NAND2_X1 cor_maj_34_U3 ( .A1(cor_maj_34_n26), .A2(cor_maj_34_n25), .ZN(
        cor_maj_34_port_o) );
  XOR2_X1 cor_maj_34_U2 ( .A(cor_maj_34_n22), .B(cor_maj_34_n21), .Z(
        cor_maj_34_n23) );
  NAND2_X1 cor_maj_35_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_35_n18) );
  NAND2_X1 cor_maj_35_U14 ( .A1(cor_maj_35_n21), .A2(cor_maj_35_n22), .ZN(
        cor_maj_35_n17) );
  NAND2_X1 cor_maj_35_U13 ( .A1(cor_maj_35_n18), .A2(cor_maj_35_n17), .ZN(
        cor_maj_35_n19) );
  NAND2_X1 cor_maj_35_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_35_n16), .ZN(
        cor_maj_35_n14) );
  NAND2_X1 cor_maj_35_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_35_n15) );
  NAND2_X1 cor_maj_35_U10 ( .A1(cor_maj_35_n15), .A2(cor_maj_35_n14), .ZN(
        cor_maj_35_n20) );
  XOR2_X1 cor_maj_35_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_35_n22)
         );
  XOR2_X1 cor_maj_35_U8 ( .A(v_1_0_2[2]), .B(cor_maj_35_n16), .Z(
        cor_maj_35_n21) );
  XOR2_X1 cor_maj_35_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_35_n16)
         );
  OR2_X1 cor_maj_35_U6 ( .A1(cor_maj_35_n20), .A2(cor_maj_35_n19), .ZN(
        cor_maj_35_n24) );
  NAND2_X1 cor_maj_35_U5 ( .A1(cor_maj_35_n24), .A2(cor_maj_35_n23), .ZN(
        cor_maj_35_n25) );
  NAND2_X1 cor_maj_35_U4 ( .A1(cor_maj_35_n20), .A2(cor_maj_35_n19), .ZN(
        cor_maj_35_n26) );
  NAND2_X1 cor_maj_35_U3 ( .A1(cor_maj_35_n26), .A2(cor_maj_35_n25), .ZN(
        cor_maj_35_port_o) );
  XOR2_X1 cor_maj_35_U2 ( .A(cor_maj_35_n22), .B(cor_maj_35_n21), .Z(
        cor_maj_35_n23) );
  NAND2_X1 cor_maj_36_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_36_n18) );
  NAND2_X1 cor_maj_36_U14 ( .A1(cor_maj_36_n21), .A2(cor_maj_36_n22), .ZN(
        cor_maj_36_n17) );
  NAND2_X1 cor_maj_36_U13 ( .A1(cor_maj_36_n18), .A2(cor_maj_36_n17), .ZN(
        cor_maj_36_n19) );
  NAND2_X1 cor_maj_36_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_36_n16), .ZN(
        cor_maj_36_n14) );
  NAND2_X1 cor_maj_36_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_36_n15) );
  NAND2_X1 cor_maj_36_U10 ( .A1(cor_maj_36_n15), .A2(cor_maj_36_n14), .ZN(
        cor_maj_36_n20) );
  XOR2_X1 cor_maj_36_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_36_n22)
         );
  XOR2_X1 cor_maj_36_U8 ( .A(v_1_0_2[2]), .B(cor_maj_36_n16), .Z(
        cor_maj_36_n21) );
  XOR2_X1 cor_maj_36_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_36_n16)
         );
  OR2_X1 cor_maj_36_U6 ( .A1(cor_maj_36_n20), .A2(cor_maj_36_n19), .ZN(
        cor_maj_36_n24) );
  NAND2_X1 cor_maj_36_U5 ( .A1(cor_maj_36_n24), .A2(cor_maj_36_n23), .ZN(
        cor_maj_36_n25) );
  NAND2_X1 cor_maj_36_U4 ( .A1(cor_maj_36_n20), .A2(cor_maj_36_n19), .ZN(
        cor_maj_36_n26) );
  NAND2_X1 cor_maj_36_U3 ( .A1(cor_maj_36_n26), .A2(cor_maj_36_n25), .ZN(
        cor_maj_36_port_o) );
  XOR2_X1 cor_maj_36_U2 ( .A(cor_maj_36_n22), .B(cor_maj_36_n21), .Z(
        cor_maj_36_n23) );
  NAND2_X1 cor_maj_37_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_37_n18) );
  NAND2_X1 cor_maj_37_U14 ( .A1(cor_maj_37_n21), .A2(cor_maj_37_n22), .ZN(
        cor_maj_37_n17) );
  NAND2_X1 cor_maj_37_U13 ( .A1(cor_maj_37_n18), .A2(cor_maj_37_n17), .ZN(
        cor_maj_37_n19) );
  NAND2_X1 cor_maj_37_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_37_n16), .ZN(
        cor_maj_37_n14) );
  NAND2_X1 cor_maj_37_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_37_n15) );
  NAND2_X1 cor_maj_37_U10 ( .A1(cor_maj_37_n15), .A2(cor_maj_37_n14), .ZN(
        cor_maj_37_n20) );
  XOR2_X1 cor_maj_37_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_37_n22)
         );
  XOR2_X1 cor_maj_37_U8 ( .A(v_1_0_2[2]), .B(cor_maj_37_n16), .Z(
        cor_maj_37_n21) );
  XOR2_X1 cor_maj_37_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_37_n16)
         );
  OR2_X1 cor_maj_37_U6 ( .A1(cor_maj_37_n20), .A2(cor_maj_37_n19), .ZN(
        cor_maj_37_n24) );
  NAND2_X1 cor_maj_37_U5 ( .A1(cor_maj_37_n24), .A2(cor_maj_37_n23), .ZN(
        cor_maj_37_n25) );
  NAND2_X1 cor_maj_37_U4 ( .A1(cor_maj_37_n20), .A2(cor_maj_37_n19), .ZN(
        cor_maj_37_n26) );
  NAND2_X1 cor_maj_37_U3 ( .A1(cor_maj_37_n26), .A2(cor_maj_37_n25), .ZN(
        cor_maj_37_port_o) );
  XOR2_X1 cor_maj_37_U2 ( .A(cor_maj_37_n22), .B(cor_maj_37_n21), .Z(
        cor_maj_37_n23) );
  NAND2_X1 cor_maj_38_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_38_n18) );
  NAND2_X1 cor_maj_38_U14 ( .A1(cor_maj_38_n21), .A2(cor_maj_38_n22), .ZN(
        cor_maj_38_n17) );
  NAND2_X1 cor_maj_38_U13 ( .A1(cor_maj_38_n18), .A2(cor_maj_38_n17), .ZN(
        cor_maj_38_n19) );
  NAND2_X1 cor_maj_38_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_38_n16), .ZN(
        cor_maj_38_n14) );
  NAND2_X1 cor_maj_38_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_38_n15) );
  NAND2_X1 cor_maj_38_U10 ( .A1(cor_maj_38_n15), .A2(cor_maj_38_n14), .ZN(
        cor_maj_38_n20) );
  XOR2_X1 cor_maj_38_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_38_n22)
         );
  XOR2_X1 cor_maj_38_U8 ( .A(v_1_0_2[2]), .B(cor_maj_38_n16), .Z(
        cor_maj_38_n21) );
  XOR2_X1 cor_maj_38_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_38_n16)
         );
  OR2_X1 cor_maj_38_U6 ( .A1(cor_maj_38_n20), .A2(cor_maj_38_n19), .ZN(
        cor_maj_38_n24) );
  NAND2_X1 cor_maj_38_U5 ( .A1(cor_maj_38_n24), .A2(cor_maj_38_n23), .ZN(
        cor_maj_38_n25) );
  NAND2_X1 cor_maj_38_U4 ( .A1(cor_maj_38_n20), .A2(cor_maj_38_n19), .ZN(
        cor_maj_38_n26) );
  NAND2_X1 cor_maj_38_U3 ( .A1(cor_maj_38_n26), .A2(cor_maj_38_n25), .ZN(
        cor_maj_38_port_o) );
  XOR2_X1 cor_maj_38_U2 ( .A(cor_maj_38_n22), .B(cor_maj_38_n21), .Z(
        cor_maj_38_n23) );
  NAND2_X1 cor_maj_39_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_39_n18) );
  NAND2_X1 cor_maj_39_U14 ( .A1(cor_maj_39_n21), .A2(cor_maj_39_n22), .ZN(
        cor_maj_39_n17) );
  NAND2_X1 cor_maj_39_U13 ( .A1(cor_maj_39_n18), .A2(cor_maj_39_n17), .ZN(
        cor_maj_39_n19) );
  NAND2_X1 cor_maj_39_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_39_n16), .ZN(
        cor_maj_39_n14) );
  NAND2_X1 cor_maj_39_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_39_n15) );
  NAND2_X1 cor_maj_39_U10 ( .A1(cor_maj_39_n15), .A2(cor_maj_39_n14), .ZN(
        cor_maj_39_n20) );
  XOR2_X1 cor_maj_39_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_39_n22)
         );
  XOR2_X1 cor_maj_39_U8 ( .A(v_1_0_2[2]), .B(cor_maj_39_n16), .Z(
        cor_maj_39_n21) );
  XOR2_X1 cor_maj_39_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_39_n16)
         );
  OR2_X1 cor_maj_39_U6 ( .A1(cor_maj_39_n20), .A2(cor_maj_39_n19), .ZN(
        cor_maj_39_n24) );
  NAND2_X1 cor_maj_39_U5 ( .A1(cor_maj_39_n24), .A2(cor_maj_39_n23), .ZN(
        cor_maj_39_n25) );
  NAND2_X1 cor_maj_39_U4 ( .A1(cor_maj_39_n20), .A2(cor_maj_39_n19), .ZN(
        cor_maj_39_n26) );
  NAND2_X1 cor_maj_39_U3 ( .A1(cor_maj_39_n26), .A2(cor_maj_39_n25), .ZN(
        cor_maj_39_port_o) );
  XOR2_X1 cor_maj_39_U2 ( .A(cor_maj_39_n22), .B(cor_maj_39_n21), .Z(
        cor_maj_39_n23) );
  NAND2_X1 cor_maj_40_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_40_n18) );
  NAND2_X1 cor_maj_40_U14 ( .A1(cor_maj_40_n21), .A2(cor_maj_40_n22), .ZN(
        cor_maj_40_n17) );
  NAND2_X1 cor_maj_40_U13 ( .A1(cor_maj_40_n18), .A2(cor_maj_40_n17), .ZN(
        cor_maj_40_n19) );
  NAND2_X1 cor_maj_40_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_40_n16), .ZN(
        cor_maj_40_n14) );
  NAND2_X1 cor_maj_40_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_40_n15) );
  NAND2_X1 cor_maj_40_U10 ( .A1(cor_maj_40_n15), .A2(cor_maj_40_n14), .ZN(
        cor_maj_40_n20) );
  XOR2_X1 cor_maj_40_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_40_n22)
         );
  XOR2_X1 cor_maj_40_U8 ( .A(v_1_1_0[2]), .B(cor_maj_40_n16), .Z(
        cor_maj_40_n21) );
  XOR2_X1 cor_maj_40_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_40_n16)
         );
  OR2_X1 cor_maj_40_U6 ( .A1(cor_maj_40_n20), .A2(cor_maj_40_n19), .ZN(
        cor_maj_40_n24) );
  NAND2_X1 cor_maj_40_U5 ( .A1(cor_maj_40_n24), .A2(cor_maj_40_n23), .ZN(
        cor_maj_40_n25) );
  NAND2_X1 cor_maj_40_U4 ( .A1(cor_maj_40_n20), .A2(cor_maj_40_n19), .ZN(
        cor_maj_40_n26) );
  NAND2_X1 cor_maj_40_U3 ( .A1(cor_maj_40_n26), .A2(cor_maj_40_n25), .ZN(
        cor_maj_40_port_o) );
  XOR2_X1 cor_maj_40_U2 ( .A(cor_maj_40_n22), .B(cor_maj_40_n21), .Z(
        cor_maj_40_n23) );
  NAND2_X1 cor_maj_41_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_41_n18) );
  NAND2_X1 cor_maj_41_U14 ( .A1(cor_maj_41_n21), .A2(cor_maj_41_n22), .ZN(
        cor_maj_41_n17) );
  NAND2_X1 cor_maj_41_U13 ( .A1(cor_maj_41_n18), .A2(cor_maj_41_n17), .ZN(
        cor_maj_41_n19) );
  NAND2_X1 cor_maj_41_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_41_n16), .ZN(
        cor_maj_41_n14) );
  NAND2_X1 cor_maj_41_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_41_n15) );
  NAND2_X1 cor_maj_41_U10 ( .A1(cor_maj_41_n15), .A2(cor_maj_41_n14), .ZN(
        cor_maj_41_n20) );
  XOR2_X1 cor_maj_41_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_41_n22)
         );
  XOR2_X1 cor_maj_41_U8 ( .A(v_1_1_0[2]), .B(cor_maj_41_n16), .Z(
        cor_maj_41_n21) );
  XOR2_X1 cor_maj_41_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_41_n16)
         );
  OR2_X1 cor_maj_41_U6 ( .A1(cor_maj_41_n20), .A2(cor_maj_41_n19), .ZN(
        cor_maj_41_n24) );
  NAND2_X1 cor_maj_41_U5 ( .A1(cor_maj_41_n24), .A2(cor_maj_41_n23), .ZN(
        cor_maj_41_n25) );
  NAND2_X1 cor_maj_41_U4 ( .A1(cor_maj_41_n20), .A2(cor_maj_41_n19), .ZN(
        cor_maj_41_n26) );
  NAND2_X1 cor_maj_41_U3 ( .A1(cor_maj_41_n26), .A2(cor_maj_41_n25), .ZN(
        cor_maj_41_port_o) );
  XOR2_X1 cor_maj_41_U2 ( .A(cor_maj_41_n22), .B(cor_maj_41_n21), .Z(
        cor_maj_41_n23) );
  NAND2_X1 cor_maj_42_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_42_n18) );
  NAND2_X1 cor_maj_42_U14 ( .A1(cor_maj_42_n21), .A2(cor_maj_42_n22), .ZN(
        cor_maj_42_n17) );
  NAND2_X1 cor_maj_42_U13 ( .A1(cor_maj_42_n18), .A2(cor_maj_42_n17), .ZN(
        cor_maj_42_n19) );
  NAND2_X1 cor_maj_42_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_42_n16), .ZN(
        cor_maj_42_n14) );
  NAND2_X1 cor_maj_42_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_42_n15) );
  NAND2_X1 cor_maj_42_U10 ( .A1(cor_maj_42_n15), .A2(cor_maj_42_n14), .ZN(
        cor_maj_42_n20) );
  XOR2_X1 cor_maj_42_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_42_n22)
         );
  XOR2_X1 cor_maj_42_U8 ( .A(v_1_1_0[2]), .B(cor_maj_42_n16), .Z(
        cor_maj_42_n21) );
  XOR2_X1 cor_maj_42_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_42_n16)
         );
  OR2_X1 cor_maj_42_U6 ( .A1(cor_maj_42_n20), .A2(cor_maj_42_n19), .ZN(
        cor_maj_42_n24) );
  NAND2_X1 cor_maj_42_U5 ( .A1(cor_maj_42_n24), .A2(cor_maj_42_n23), .ZN(
        cor_maj_42_n25) );
  NAND2_X1 cor_maj_42_U4 ( .A1(cor_maj_42_n20), .A2(cor_maj_42_n19), .ZN(
        cor_maj_42_n26) );
  NAND2_X1 cor_maj_42_U3 ( .A1(cor_maj_42_n26), .A2(cor_maj_42_n25), .ZN(
        cor_maj_42_port_o) );
  XOR2_X1 cor_maj_42_U2 ( .A(cor_maj_42_n22), .B(cor_maj_42_n21), .Z(
        cor_maj_42_n23) );
  NAND2_X1 cor_maj_43_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_43_n18) );
  NAND2_X1 cor_maj_43_U14 ( .A1(cor_maj_43_n21), .A2(cor_maj_43_n22), .ZN(
        cor_maj_43_n17) );
  NAND2_X1 cor_maj_43_U13 ( .A1(cor_maj_43_n18), .A2(cor_maj_43_n17), .ZN(
        cor_maj_43_n19) );
  NAND2_X1 cor_maj_43_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_43_n16), .ZN(
        cor_maj_43_n14) );
  NAND2_X1 cor_maj_43_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_43_n15) );
  NAND2_X1 cor_maj_43_U10 ( .A1(cor_maj_43_n15), .A2(cor_maj_43_n14), .ZN(
        cor_maj_43_n20) );
  XOR2_X1 cor_maj_43_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_43_n22)
         );
  XOR2_X1 cor_maj_43_U8 ( .A(v_1_1_0[2]), .B(cor_maj_43_n16), .Z(
        cor_maj_43_n21) );
  XOR2_X1 cor_maj_43_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_43_n16)
         );
  OR2_X1 cor_maj_43_U6 ( .A1(cor_maj_43_n20), .A2(cor_maj_43_n19), .ZN(
        cor_maj_43_n24) );
  NAND2_X1 cor_maj_43_U5 ( .A1(cor_maj_43_n24), .A2(cor_maj_43_n23), .ZN(
        cor_maj_43_n25) );
  NAND2_X1 cor_maj_43_U4 ( .A1(cor_maj_43_n20), .A2(cor_maj_43_n19), .ZN(
        cor_maj_43_n26) );
  NAND2_X1 cor_maj_43_U3 ( .A1(cor_maj_43_n26), .A2(cor_maj_43_n25), .ZN(
        cor_maj_43_port_o) );
  XOR2_X1 cor_maj_43_U2 ( .A(cor_maj_43_n22), .B(cor_maj_43_n21), .Z(
        cor_maj_43_n23) );
  NAND2_X1 cor_maj_44_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_44_n18) );
  NAND2_X1 cor_maj_44_U14 ( .A1(cor_maj_44_n21), .A2(cor_maj_44_n22), .ZN(
        cor_maj_44_n17) );
  NAND2_X1 cor_maj_44_U13 ( .A1(cor_maj_44_n18), .A2(cor_maj_44_n17), .ZN(
        cor_maj_44_n19) );
  NAND2_X1 cor_maj_44_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_44_n16), .ZN(
        cor_maj_44_n14) );
  NAND2_X1 cor_maj_44_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_44_n15) );
  NAND2_X1 cor_maj_44_U10 ( .A1(cor_maj_44_n15), .A2(cor_maj_44_n14), .ZN(
        cor_maj_44_n20) );
  XOR2_X1 cor_maj_44_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_44_n22)
         );
  XOR2_X1 cor_maj_44_U8 ( .A(v_1_1_0[2]), .B(cor_maj_44_n16), .Z(
        cor_maj_44_n21) );
  XOR2_X1 cor_maj_44_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_44_n16)
         );
  OR2_X1 cor_maj_44_U6 ( .A1(cor_maj_44_n20), .A2(cor_maj_44_n19), .ZN(
        cor_maj_44_n24) );
  NAND2_X1 cor_maj_44_U5 ( .A1(cor_maj_44_n24), .A2(cor_maj_44_n23), .ZN(
        cor_maj_44_n25) );
  NAND2_X1 cor_maj_44_U4 ( .A1(cor_maj_44_n20), .A2(cor_maj_44_n19), .ZN(
        cor_maj_44_n26) );
  NAND2_X1 cor_maj_44_U3 ( .A1(cor_maj_44_n26), .A2(cor_maj_44_n25), .ZN(
        cor_maj_44_port_o) );
  XOR2_X1 cor_maj_44_U2 ( .A(cor_maj_44_n22), .B(cor_maj_44_n21), .Z(
        cor_maj_44_n23) );
  NAND2_X1 cor_maj_45_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_45_n18) );
  NAND2_X1 cor_maj_45_U14 ( .A1(cor_maj_45_n21), .A2(cor_maj_45_n22), .ZN(
        cor_maj_45_n17) );
  NAND2_X1 cor_maj_45_U13 ( .A1(cor_maj_45_n18), .A2(cor_maj_45_n17), .ZN(
        cor_maj_45_n19) );
  NAND2_X1 cor_maj_45_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_45_n16), .ZN(
        cor_maj_45_n14) );
  NAND2_X1 cor_maj_45_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_45_n15) );
  NAND2_X1 cor_maj_45_U10 ( .A1(cor_maj_45_n15), .A2(cor_maj_45_n14), .ZN(
        cor_maj_45_n20) );
  XOR2_X1 cor_maj_45_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_45_n22)
         );
  XOR2_X1 cor_maj_45_U8 ( .A(v_1_1_2[2]), .B(cor_maj_45_n16), .Z(
        cor_maj_45_n21) );
  XOR2_X1 cor_maj_45_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_45_n16)
         );
  OR2_X1 cor_maj_45_U6 ( .A1(cor_maj_45_n20), .A2(cor_maj_45_n19), .ZN(
        cor_maj_45_n24) );
  NAND2_X1 cor_maj_45_U5 ( .A1(cor_maj_45_n24), .A2(cor_maj_45_n23), .ZN(
        cor_maj_45_n25) );
  NAND2_X1 cor_maj_45_U4 ( .A1(cor_maj_45_n20), .A2(cor_maj_45_n19), .ZN(
        cor_maj_45_n26) );
  NAND2_X1 cor_maj_45_U3 ( .A1(cor_maj_45_n26), .A2(cor_maj_45_n25), .ZN(
        cor_maj_45_port_o) );
  XOR2_X1 cor_maj_45_U2 ( .A(cor_maj_45_n22), .B(cor_maj_45_n21), .Z(
        cor_maj_45_n23) );
  NAND2_X1 cor_maj_46_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_46_n18) );
  NAND2_X1 cor_maj_46_U14 ( .A1(cor_maj_46_n21), .A2(cor_maj_46_n22), .ZN(
        cor_maj_46_n17) );
  NAND2_X1 cor_maj_46_U13 ( .A1(cor_maj_46_n18), .A2(cor_maj_46_n17), .ZN(
        cor_maj_46_n19) );
  NAND2_X1 cor_maj_46_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_46_n16), .ZN(
        cor_maj_46_n14) );
  NAND2_X1 cor_maj_46_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_46_n15) );
  NAND2_X1 cor_maj_46_U10 ( .A1(cor_maj_46_n15), .A2(cor_maj_46_n14), .ZN(
        cor_maj_46_n20) );
  XOR2_X1 cor_maj_46_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_46_n22)
         );
  XOR2_X1 cor_maj_46_U8 ( .A(v_1_1_2[2]), .B(cor_maj_46_n16), .Z(
        cor_maj_46_n21) );
  XOR2_X1 cor_maj_46_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_46_n16)
         );
  OR2_X1 cor_maj_46_U6 ( .A1(cor_maj_46_n20), .A2(cor_maj_46_n19), .ZN(
        cor_maj_46_n24) );
  NAND2_X1 cor_maj_46_U5 ( .A1(cor_maj_46_n24), .A2(cor_maj_46_n23), .ZN(
        cor_maj_46_n25) );
  NAND2_X1 cor_maj_46_U4 ( .A1(cor_maj_46_n20), .A2(cor_maj_46_n19), .ZN(
        cor_maj_46_n26) );
  NAND2_X1 cor_maj_46_U3 ( .A1(cor_maj_46_n26), .A2(cor_maj_46_n25), .ZN(
        cor_maj_46_port_o) );
  XOR2_X1 cor_maj_46_U2 ( .A(cor_maj_46_n22), .B(cor_maj_46_n21), .Z(
        cor_maj_46_n23) );
  NAND2_X1 cor_maj_47_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_47_n18) );
  NAND2_X1 cor_maj_47_U14 ( .A1(cor_maj_47_n21), .A2(cor_maj_47_n22), .ZN(
        cor_maj_47_n17) );
  NAND2_X1 cor_maj_47_U13 ( .A1(cor_maj_47_n18), .A2(cor_maj_47_n17), .ZN(
        cor_maj_47_n19) );
  NAND2_X1 cor_maj_47_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_47_n16), .ZN(
        cor_maj_47_n14) );
  NAND2_X1 cor_maj_47_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_47_n15) );
  NAND2_X1 cor_maj_47_U10 ( .A1(cor_maj_47_n15), .A2(cor_maj_47_n14), .ZN(
        cor_maj_47_n20) );
  XOR2_X1 cor_maj_47_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_47_n22)
         );
  XOR2_X1 cor_maj_47_U8 ( .A(v_1_1_2[2]), .B(cor_maj_47_n16), .Z(
        cor_maj_47_n21) );
  XOR2_X1 cor_maj_47_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_47_n16)
         );
  OR2_X1 cor_maj_47_U6 ( .A1(cor_maj_47_n20), .A2(cor_maj_47_n19), .ZN(
        cor_maj_47_n24) );
  NAND2_X1 cor_maj_47_U5 ( .A1(cor_maj_47_n24), .A2(cor_maj_47_n23), .ZN(
        cor_maj_47_n25) );
  NAND2_X1 cor_maj_47_U4 ( .A1(cor_maj_47_n20), .A2(cor_maj_47_n19), .ZN(
        cor_maj_47_n26) );
  NAND2_X1 cor_maj_47_U3 ( .A1(cor_maj_47_n26), .A2(cor_maj_47_n25), .ZN(
        cor_maj_47_port_o) );
  XOR2_X1 cor_maj_47_U2 ( .A(cor_maj_47_n22), .B(cor_maj_47_n21), .Z(
        cor_maj_47_n23) );
  NAND2_X1 cor_maj_48_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_48_n18) );
  NAND2_X1 cor_maj_48_U14 ( .A1(cor_maj_48_n21), .A2(cor_maj_48_n22), .ZN(
        cor_maj_48_n17) );
  NAND2_X1 cor_maj_48_U13 ( .A1(cor_maj_48_n18), .A2(cor_maj_48_n17), .ZN(
        cor_maj_48_n19) );
  NAND2_X1 cor_maj_48_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_48_n16), .ZN(
        cor_maj_48_n14) );
  NAND2_X1 cor_maj_48_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_48_n15) );
  NAND2_X1 cor_maj_48_U10 ( .A1(cor_maj_48_n15), .A2(cor_maj_48_n14), .ZN(
        cor_maj_48_n20) );
  XOR2_X1 cor_maj_48_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_48_n22)
         );
  XOR2_X1 cor_maj_48_U8 ( .A(v_1_1_2[2]), .B(cor_maj_48_n16), .Z(
        cor_maj_48_n21) );
  XOR2_X1 cor_maj_48_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_48_n16)
         );
  OR2_X1 cor_maj_48_U6 ( .A1(cor_maj_48_n20), .A2(cor_maj_48_n19), .ZN(
        cor_maj_48_n24) );
  NAND2_X1 cor_maj_48_U5 ( .A1(cor_maj_48_n24), .A2(cor_maj_48_n23), .ZN(
        cor_maj_48_n25) );
  NAND2_X1 cor_maj_48_U4 ( .A1(cor_maj_48_n20), .A2(cor_maj_48_n19), .ZN(
        cor_maj_48_n26) );
  NAND2_X1 cor_maj_48_U3 ( .A1(cor_maj_48_n26), .A2(cor_maj_48_n25), .ZN(
        cor_maj_48_port_o) );
  XOR2_X1 cor_maj_48_U2 ( .A(cor_maj_48_n22), .B(cor_maj_48_n21), .Z(
        cor_maj_48_n23) );
  NAND2_X1 cor_maj_49_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_49_n18) );
  NAND2_X1 cor_maj_49_U14 ( .A1(cor_maj_49_n21), .A2(cor_maj_49_n22), .ZN(
        cor_maj_49_n17) );
  NAND2_X1 cor_maj_49_U13 ( .A1(cor_maj_49_n18), .A2(cor_maj_49_n17), .ZN(
        cor_maj_49_n19) );
  NAND2_X1 cor_maj_49_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_49_n16), .ZN(
        cor_maj_49_n14) );
  NAND2_X1 cor_maj_49_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_49_n15) );
  NAND2_X1 cor_maj_49_U10 ( .A1(cor_maj_49_n15), .A2(cor_maj_49_n14), .ZN(
        cor_maj_49_n20) );
  XOR2_X1 cor_maj_49_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_49_n22)
         );
  XOR2_X1 cor_maj_49_U8 ( .A(v_1_1_2[2]), .B(cor_maj_49_n16), .Z(
        cor_maj_49_n21) );
  XOR2_X1 cor_maj_49_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_49_n16)
         );
  OR2_X1 cor_maj_49_U6 ( .A1(cor_maj_49_n20), .A2(cor_maj_49_n19), .ZN(
        cor_maj_49_n24) );
  NAND2_X1 cor_maj_49_U5 ( .A1(cor_maj_49_n24), .A2(cor_maj_49_n23), .ZN(
        cor_maj_49_n25) );
  NAND2_X1 cor_maj_49_U4 ( .A1(cor_maj_49_n20), .A2(cor_maj_49_n19), .ZN(
        cor_maj_49_n26) );
  NAND2_X1 cor_maj_49_U3 ( .A1(cor_maj_49_n26), .A2(cor_maj_49_n25), .ZN(
        cor_maj_49_port_o) );
  XOR2_X1 cor_maj_49_U2 ( .A(cor_maj_49_n22), .B(cor_maj_49_n21), .Z(
        cor_maj_49_n23) );
  NAND2_X1 cor_maj_50_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_50_n18) );
  NAND2_X1 cor_maj_50_U14 ( .A1(cor_maj_50_n21), .A2(cor_maj_50_n22), .ZN(
        cor_maj_50_n17) );
  NAND2_X1 cor_maj_50_U13 ( .A1(cor_maj_50_n18), .A2(cor_maj_50_n17), .ZN(
        cor_maj_50_n19) );
  NAND2_X1 cor_maj_50_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_50_n16), .ZN(
        cor_maj_50_n14) );
  NAND2_X1 cor_maj_50_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_50_n15) );
  NAND2_X1 cor_maj_50_U10 ( .A1(cor_maj_50_n15), .A2(cor_maj_50_n14), .ZN(
        cor_maj_50_n20) );
  XOR2_X1 cor_maj_50_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_50_n22)
         );
  XOR2_X1 cor_maj_50_U8 ( .A(v_1_2_0[2]), .B(cor_maj_50_n16), .Z(
        cor_maj_50_n21) );
  XOR2_X1 cor_maj_50_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_50_n16)
         );
  OR2_X1 cor_maj_50_U6 ( .A1(cor_maj_50_n20), .A2(cor_maj_50_n19), .ZN(
        cor_maj_50_n24) );
  NAND2_X1 cor_maj_50_U5 ( .A1(cor_maj_50_n24), .A2(cor_maj_50_n23), .ZN(
        cor_maj_50_n25) );
  NAND2_X1 cor_maj_50_U4 ( .A1(cor_maj_50_n20), .A2(cor_maj_50_n19), .ZN(
        cor_maj_50_n26) );
  NAND2_X1 cor_maj_50_U3 ( .A1(cor_maj_50_n26), .A2(cor_maj_50_n25), .ZN(
        cor_maj_50_port_o) );
  XOR2_X1 cor_maj_50_U2 ( .A(cor_maj_50_n22), .B(cor_maj_50_n21), .Z(
        cor_maj_50_n23) );
  NAND2_X1 cor_maj_51_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_51_n18) );
  NAND2_X1 cor_maj_51_U14 ( .A1(cor_maj_51_n21), .A2(cor_maj_51_n22), .ZN(
        cor_maj_51_n17) );
  NAND2_X1 cor_maj_51_U13 ( .A1(cor_maj_51_n18), .A2(cor_maj_51_n17), .ZN(
        cor_maj_51_n19) );
  NAND2_X1 cor_maj_51_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_51_n16), .ZN(
        cor_maj_51_n14) );
  NAND2_X1 cor_maj_51_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_51_n15) );
  NAND2_X1 cor_maj_51_U10 ( .A1(cor_maj_51_n15), .A2(cor_maj_51_n14), .ZN(
        cor_maj_51_n20) );
  XOR2_X1 cor_maj_51_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_51_n22)
         );
  XOR2_X1 cor_maj_51_U8 ( .A(v_1_2_0[2]), .B(cor_maj_51_n16), .Z(
        cor_maj_51_n21) );
  XOR2_X1 cor_maj_51_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_51_n16)
         );
  OR2_X1 cor_maj_51_U6 ( .A1(cor_maj_51_n20), .A2(cor_maj_51_n19), .ZN(
        cor_maj_51_n24) );
  NAND2_X1 cor_maj_51_U5 ( .A1(cor_maj_51_n24), .A2(cor_maj_51_n23), .ZN(
        cor_maj_51_n25) );
  NAND2_X1 cor_maj_51_U4 ( .A1(cor_maj_51_n20), .A2(cor_maj_51_n19), .ZN(
        cor_maj_51_n26) );
  NAND2_X1 cor_maj_51_U3 ( .A1(cor_maj_51_n26), .A2(cor_maj_51_n25), .ZN(
        cor_maj_51_port_o) );
  XOR2_X1 cor_maj_51_U2 ( .A(cor_maj_51_n22), .B(cor_maj_51_n21), .Z(
        cor_maj_51_n23) );
  NAND2_X1 cor_maj_52_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_52_n18) );
  NAND2_X1 cor_maj_52_U14 ( .A1(cor_maj_52_n21), .A2(cor_maj_52_n22), .ZN(
        cor_maj_52_n17) );
  NAND2_X1 cor_maj_52_U13 ( .A1(cor_maj_52_n18), .A2(cor_maj_52_n17), .ZN(
        cor_maj_52_n19) );
  NAND2_X1 cor_maj_52_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_52_n16), .ZN(
        cor_maj_52_n14) );
  NAND2_X1 cor_maj_52_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_52_n15) );
  NAND2_X1 cor_maj_52_U10 ( .A1(cor_maj_52_n15), .A2(cor_maj_52_n14), .ZN(
        cor_maj_52_n20) );
  XOR2_X1 cor_maj_52_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_52_n22)
         );
  XOR2_X1 cor_maj_52_U8 ( .A(v_1_2_0[2]), .B(cor_maj_52_n16), .Z(
        cor_maj_52_n21) );
  XOR2_X1 cor_maj_52_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_52_n16)
         );
  OR2_X1 cor_maj_52_U6 ( .A1(cor_maj_52_n20), .A2(cor_maj_52_n19), .ZN(
        cor_maj_52_n24) );
  NAND2_X1 cor_maj_52_U5 ( .A1(cor_maj_52_n24), .A2(cor_maj_52_n23), .ZN(
        cor_maj_52_n25) );
  NAND2_X1 cor_maj_52_U4 ( .A1(cor_maj_52_n20), .A2(cor_maj_52_n19), .ZN(
        cor_maj_52_n26) );
  NAND2_X1 cor_maj_52_U3 ( .A1(cor_maj_52_n26), .A2(cor_maj_52_n25), .ZN(
        cor_maj_52_port_o) );
  XOR2_X1 cor_maj_52_U2 ( .A(cor_maj_52_n22), .B(cor_maj_52_n21), .Z(
        cor_maj_52_n23) );
  NAND2_X1 cor_maj_53_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_53_n18) );
  NAND2_X1 cor_maj_53_U14 ( .A1(cor_maj_53_n21), .A2(cor_maj_53_n22), .ZN(
        cor_maj_53_n17) );
  NAND2_X1 cor_maj_53_U13 ( .A1(cor_maj_53_n18), .A2(cor_maj_53_n17), .ZN(
        cor_maj_53_n19) );
  NAND2_X1 cor_maj_53_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_53_n16), .ZN(
        cor_maj_53_n14) );
  NAND2_X1 cor_maj_53_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_53_n15) );
  NAND2_X1 cor_maj_53_U10 ( .A1(cor_maj_53_n15), .A2(cor_maj_53_n14), .ZN(
        cor_maj_53_n20) );
  XOR2_X1 cor_maj_53_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_53_n22)
         );
  XOR2_X1 cor_maj_53_U8 ( .A(v_1_2_0[2]), .B(cor_maj_53_n16), .Z(
        cor_maj_53_n21) );
  XOR2_X1 cor_maj_53_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_53_n16)
         );
  OR2_X1 cor_maj_53_U6 ( .A1(cor_maj_53_n20), .A2(cor_maj_53_n19), .ZN(
        cor_maj_53_n24) );
  NAND2_X1 cor_maj_53_U5 ( .A1(cor_maj_53_n24), .A2(cor_maj_53_n23), .ZN(
        cor_maj_53_n25) );
  NAND2_X1 cor_maj_53_U4 ( .A1(cor_maj_53_n20), .A2(cor_maj_53_n19), .ZN(
        cor_maj_53_n26) );
  NAND2_X1 cor_maj_53_U3 ( .A1(cor_maj_53_n26), .A2(cor_maj_53_n25), .ZN(
        cor_maj_53_port_o) );
  XOR2_X1 cor_maj_53_U2 ( .A(cor_maj_53_n22), .B(cor_maj_53_n21), .Z(
        cor_maj_53_n23) );
  NAND2_X1 cor_maj_54_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_54_n18) );
  NAND2_X1 cor_maj_54_U14 ( .A1(cor_maj_54_n21), .A2(cor_maj_54_n22), .ZN(
        cor_maj_54_n17) );
  NAND2_X1 cor_maj_54_U13 ( .A1(cor_maj_54_n18), .A2(cor_maj_54_n17), .ZN(
        cor_maj_54_n19) );
  NAND2_X1 cor_maj_54_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_54_n16), .ZN(
        cor_maj_54_n14) );
  NAND2_X1 cor_maj_54_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_54_n15) );
  NAND2_X1 cor_maj_54_U10 ( .A1(cor_maj_54_n15), .A2(cor_maj_54_n14), .ZN(
        cor_maj_54_n20) );
  XOR2_X1 cor_maj_54_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_54_n22)
         );
  XOR2_X1 cor_maj_54_U8 ( .A(v_1_2_0[2]), .B(cor_maj_54_n16), .Z(
        cor_maj_54_n21) );
  XOR2_X1 cor_maj_54_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_54_n16)
         );
  OR2_X1 cor_maj_54_U6 ( .A1(cor_maj_54_n20), .A2(cor_maj_54_n19), .ZN(
        cor_maj_54_n24) );
  NAND2_X1 cor_maj_54_U5 ( .A1(cor_maj_54_n24), .A2(cor_maj_54_n23), .ZN(
        cor_maj_54_n25) );
  NAND2_X1 cor_maj_54_U4 ( .A1(cor_maj_54_n20), .A2(cor_maj_54_n19), .ZN(
        cor_maj_54_n26) );
  NAND2_X1 cor_maj_54_U3 ( .A1(cor_maj_54_n26), .A2(cor_maj_54_n25), .ZN(
        cor_maj_54_port_o) );
  XOR2_X1 cor_maj_54_U2 ( .A(cor_maj_54_n22), .B(cor_maj_54_n21), .Z(
        cor_maj_54_n23) );
  NAND2_X1 cor_maj_55_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_55_n18) );
  NAND2_X1 cor_maj_55_U14 ( .A1(cor_maj_55_n21), .A2(cor_maj_55_n22), .ZN(
        cor_maj_55_n17) );
  NAND2_X1 cor_maj_55_U13 ( .A1(cor_maj_55_n18), .A2(cor_maj_55_n17), .ZN(
        cor_maj_55_n19) );
  NAND2_X1 cor_maj_55_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_55_n16), .ZN(
        cor_maj_55_n14) );
  NAND2_X1 cor_maj_55_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_55_n15) );
  NAND2_X1 cor_maj_55_U10 ( .A1(cor_maj_55_n15), .A2(cor_maj_55_n14), .ZN(
        cor_maj_55_n20) );
  XOR2_X1 cor_maj_55_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_55_n22)
         );
  XOR2_X1 cor_maj_55_U8 ( .A(v_1_2_1[2]), .B(cor_maj_55_n16), .Z(
        cor_maj_55_n21) );
  XOR2_X1 cor_maj_55_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_55_n16)
         );
  OR2_X1 cor_maj_55_U6 ( .A1(cor_maj_55_n20), .A2(cor_maj_55_n19), .ZN(
        cor_maj_55_n24) );
  NAND2_X1 cor_maj_55_U5 ( .A1(cor_maj_55_n24), .A2(cor_maj_55_n23), .ZN(
        cor_maj_55_n25) );
  NAND2_X1 cor_maj_55_U4 ( .A1(cor_maj_55_n20), .A2(cor_maj_55_n19), .ZN(
        cor_maj_55_n26) );
  NAND2_X1 cor_maj_55_U3 ( .A1(cor_maj_55_n26), .A2(cor_maj_55_n25), .ZN(
        cor_maj_55_port_o) );
  XOR2_X1 cor_maj_55_U2 ( .A(cor_maj_55_n22), .B(cor_maj_55_n21), .Z(
        cor_maj_55_n23) );
  NAND2_X1 cor_maj_56_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_56_n18) );
  NAND2_X1 cor_maj_56_U14 ( .A1(cor_maj_56_n21), .A2(cor_maj_56_n22), .ZN(
        cor_maj_56_n17) );
  NAND2_X1 cor_maj_56_U13 ( .A1(cor_maj_56_n18), .A2(cor_maj_56_n17), .ZN(
        cor_maj_56_n19) );
  NAND2_X1 cor_maj_56_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_56_n16), .ZN(
        cor_maj_56_n14) );
  NAND2_X1 cor_maj_56_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_56_n15) );
  NAND2_X1 cor_maj_56_U10 ( .A1(cor_maj_56_n15), .A2(cor_maj_56_n14), .ZN(
        cor_maj_56_n20) );
  XOR2_X1 cor_maj_56_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_56_n22)
         );
  XOR2_X1 cor_maj_56_U8 ( .A(v_1_2_1[2]), .B(cor_maj_56_n16), .Z(
        cor_maj_56_n21) );
  XOR2_X1 cor_maj_56_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_56_n16)
         );
  OR2_X1 cor_maj_56_U6 ( .A1(cor_maj_56_n20), .A2(cor_maj_56_n19), .ZN(
        cor_maj_56_n24) );
  NAND2_X1 cor_maj_56_U5 ( .A1(cor_maj_56_n24), .A2(cor_maj_56_n23), .ZN(
        cor_maj_56_n25) );
  NAND2_X1 cor_maj_56_U4 ( .A1(cor_maj_56_n20), .A2(cor_maj_56_n19), .ZN(
        cor_maj_56_n26) );
  NAND2_X1 cor_maj_56_U3 ( .A1(cor_maj_56_n26), .A2(cor_maj_56_n25), .ZN(
        cor_maj_56_port_o) );
  XOR2_X1 cor_maj_56_U2 ( .A(cor_maj_56_n22), .B(cor_maj_56_n21), .Z(
        cor_maj_56_n23) );
  NAND2_X1 cor_maj_57_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_57_n18) );
  NAND2_X1 cor_maj_57_U14 ( .A1(cor_maj_57_n21), .A2(cor_maj_57_n22), .ZN(
        cor_maj_57_n17) );
  NAND2_X1 cor_maj_57_U13 ( .A1(cor_maj_57_n18), .A2(cor_maj_57_n17), .ZN(
        cor_maj_57_n19) );
  NAND2_X1 cor_maj_57_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_57_n16), .ZN(
        cor_maj_57_n14) );
  NAND2_X1 cor_maj_57_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_57_n15) );
  NAND2_X1 cor_maj_57_U10 ( .A1(cor_maj_57_n15), .A2(cor_maj_57_n14), .ZN(
        cor_maj_57_n20) );
  XOR2_X1 cor_maj_57_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_57_n22)
         );
  XOR2_X1 cor_maj_57_U8 ( .A(v_1_2_1[2]), .B(cor_maj_57_n16), .Z(
        cor_maj_57_n21) );
  XOR2_X1 cor_maj_57_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_57_n16)
         );
  OR2_X1 cor_maj_57_U6 ( .A1(cor_maj_57_n20), .A2(cor_maj_57_n19), .ZN(
        cor_maj_57_n24) );
  NAND2_X1 cor_maj_57_U5 ( .A1(cor_maj_57_n24), .A2(cor_maj_57_n23), .ZN(
        cor_maj_57_n25) );
  NAND2_X1 cor_maj_57_U4 ( .A1(cor_maj_57_n20), .A2(cor_maj_57_n19), .ZN(
        cor_maj_57_n26) );
  NAND2_X1 cor_maj_57_U3 ( .A1(cor_maj_57_n26), .A2(cor_maj_57_n25), .ZN(
        cor_maj_57_port_o) );
  XOR2_X1 cor_maj_57_U2 ( .A(cor_maj_57_n22), .B(cor_maj_57_n21), .Z(
        cor_maj_57_n23) );
  NAND2_X1 cor_maj_58_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_58_n18) );
  NAND2_X1 cor_maj_58_U14 ( .A1(cor_maj_58_n21), .A2(cor_maj_58_n22), .ZN(
        cor_maj_58_n17) );
  NAND2_X1 cor_maj_58_U13 ( .A1(cor_maj_58_n18), .A2(cor_maj_58_n17), .ZN(
        cor_maj_58_n19) );
  NAND2_X1 cor_maj_58_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_58_n16), .ZN(
        cor_maj_58_n14) );
  NAND2_X1 cor_maj_58_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_58_n15) );
  NAND2_X1 cor_maj_58_U10 ( .A1(cor_maj_58_n15), .A2(cor_maj_58_n14), .ZN(
        cor_maj_58_n20) );
  XOR2_X1 cor_maj_58_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_58_n22)
         );
  XOR2_X1 cor_maj_58_U8 ( .A(v_1_2_1[2]), .B(cor_maj_58_n16), .Z(
        cor_maj_58_n21) );
  XOR2_X1 cor_maj_58_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_58_n16)
         );
  OR2_X1 cor_maj_58_U6 ( .A1(cor_maj_58_n20), .A2(cor_maj_58_n19), .ZN(
        cor_maj_58_n24) );
  NAND2_X1 cor_maj_58_U5 ( .A1(cor_maj_58_n24), .A2(cor_maj_58_n23), .ZN(
        cor_maj_58_n25) );
  NAND2_X1 cor_maj_58_U4 ( .A1(cor_maj_58_n20), .A2(cor_maj_58_n19), .ZN(
        cor_maj_58_n26) );
  NAND2_X1 cor_maj_58_U3 ( .A1(cor_maj_58_n26), .A2(cor_maj_58_n25), .ZN(
        cor_maj_58_port_o) );
  XOR2_X1 cor_maj_58_U2 ( .A(cor_maj_58_n22), .B(cor_maj_58_n21), .Z(
        cor_maj_58_n23) );
  NAND2_X1 cor_maj_59_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_59_n18) );
  NAND2_X1 cor_maj_59_U14 ( .A1(cor_maj_59_n21), .A2(cor_maj_59_n22), .ZN(
        cor_maj_59_n17) );
  NAND2_X1 cor_maj_59_U13 ( .A1(cor_maj_59_n18), .A2(cor_maj_59_n17), .ZN(
        cor_maj_59_n19) );
  NAND2_X1 cor_maj_59_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_59_n16), .ZN(
        cor_maj_59_n14) );
  NAND2_X1 cor_maj_59_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_59_n15) );
  NAND2_X1 cor_maj_59_U10 ( .A1(cor_maj_59_n15), .A2(cor_maj_59_n14), .ZN(
        cor_maj_59_n20) );
  XOR2_X1 cor_maj_59_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_59_n22)
         );
  XOR2_X1 cor_maj_59_U8 ( .A(v_1_2_1[2]), .B(cor_maj_59_n16), .Z(
        cor_maj_59_n21) );
  XOR2_X1 cor_maj_59_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_59_n16)
         );
  OR2_X1 cor_maj_59_U6 ( .A1(cor_maj_59_n20), .A2(cor_maj_59_n19), .ZN(
        cor_maj_59_n24) );
  NAND2_X1 cor_maj_59_U5 ( .A1(cor_maj_59_n24), .A2(cor_maj_59_n23), .ZN(
        cor_maj_59_n25) );
  NAND2_X1 cor_maj_59_U4 ( .A1(cor_maj_59_n20), .A2(cor_maj_59_n19), .ZN(
        cor_maj_59_n26) );
  NAND2_X1 cor_maj_59_U3 ( .A1(cor_maj_59_n26), .A2(cor_maj_59_n25), .ZN(
        cor_maj_59_port_o) );
  XOR2_X1 cor_maj_59_U2 ( .A(cor_maj_59_n22), .B(cor_maj_59_n21), .Z(
        cor_maj_59_n23) );
  XOR2_X1 simpleXor_30_U1 ( .A(n_zz_io_c_0_3[1]), .B(u_0_1[0]), .Z(
        simpleXor_30_port_z) );
  XOR2_X1 simpleXor_31_U1 ( .A(n_zz_io_c_0_3[2]), .B(u_0_2[0]), .Z(
        simpleXor_31_port_z) );
  XOR2_X1 simpleXor_32_U1 ( .A(n_zz_io_c_1_3[1]), .B(u_1_0[0]), .Z(
        simpleXor_32_port_z) );
  XOR2_X1 simpleXor_33_U1 ( .A(n_zz_io_c_1_3[2]), .B(u_1_2[0]), .Z(
        simpleXor_33_port_z) );
  XOR2_X1 simpleXor_34_U1 ( .A(n_zz_io_c_2_3[1]), .B(u_2_0[0]), .Z(
        simpleXor_34_port_z) );
  XOR2_X1 simpleXor_35_U1 ( .A(n_zz_io_c_2_3[2]), .B(u_2_1[0]), .Z(
        simpleXor_35_port_z) );
  XOR2_X1 simpleXor_36_U1 ( .A(n_zz_io_c_0_7[1]), .B(u_0_1[1]), .Z(
        simpleXor_36_port_z) );
  XOR2_X1 simpleXor_37_U1 ( .A(n_zz_io_c_0_7[2]), .B(u_0_2[1]), .Z(
        simpleXor_37_port_z) );
  XOR2_X1 simpleXor_38_U1 ( .A(n_zz_io_c_1_7[1]), .B(u_1_0[1]), .Z(
        simpleXor_38_port_z) );
  XOR2_X1 simpleXor_39_U1 ( .A(n_zz_io_c_1_7[2]), .B(u_1_2[1]), .Z(
        simpleXor_39_port_z) );
  XOR2_X1 simpleXor_40_U1 ( .A(n_zz_io_c_2_7[1]), .B(u_2_0[1]), .Z(
        simpleXor_40_port_z) );
  XOR2_X1 simpleXor_41_U1 ( .A(n_zz_io_c_2_7[2]), .B(u_2_1[1]), .Z(
        simpleXor_41_port_z) );
  XOR2_X1 simpleXor_42_U1 ( .A(n_zz_io_c_0_11[1]), .B(u_0_1[2]), .Z(
        simpleXor_42_port_z) );
  XOR2_X1 simpleXor_43_U1 ( .A(n_zz_io_c_0_11[2]), .B(u_0_2[2]), .Z(
        simpleXor_43_port_z) );
  XOR2_X1 simpleXor_44_U1 ( .A(n_zz_io_c_1_11[1]), .B(u_1_0[2]), .Z(
        simpleXor_44_port_z) );
  XOR2_X1 simpleXor_45_U1 ( .A(n_zz_io_c_1_11[2]), .B(u_1_2[2]), .Z(
        simpleXor_45_port_z) );
  XOR2_X1 simpleXor_46_U1 ( .A(n_zz_io_c_2_11[1]), .B(u_2_0[2]), .Z(
        simpleXor_46_port_z) );
  XOR2_X1 simpleXor_47_U1 ( .A(n_zz_io_c_2_11[2]), .B(u_2_1[2]), .Z(
        simpleXor_47_port_z) );
  XOR2_X1 simpleXor_48_U1 ( .A(n_zz_io_c_0_15[1]), .B(u_0_1[3]), .Z(
        simpleXor_48_port_z) );
  XOR2_X1 simpleXor_49_U1 ( .A(n_zz_io_c_0_15[2]), .B(u_0_2[3]), .Z(
        simpleXor_49_port_z) );
  XOR2_X1 simpleXor_50_U1 ( .A(n_zz_io_c_1_15[1]), .B(u_1_0[3]), .Z(
        simpleXor_50_port_z) );
  XOR2_X1 simpleXor_51_U1 ( .A(n_zz_io_c_1_15[2]), .B(u_1_2[3]), .Z(
        simpleXor_51_port_z) );
  XOR2_X1 simpleXor_52_U1 ( .A(n_zz_io_c_2_15[1]), .B(u_2_0[3]), .Z(
        simpleXor_52_port_z) );
  XOR2_X1 simpleXor_53_U1 ( .A(n_zz_io_c_2_15[2]), .B(u_2_1[3]), .Z(
        simpleXor_53_port_z) );
  XOR2_X1 simpleXor_54_U1 ( .A(n_zz_io_c_0_19[1]), .B(u_0_1[4]), .Z(
        simpleXor_54_port_z) );
  XOR2_X1 simpleXor_55_U1 ( .A(n_zz_io_c_0_19[2]), .B(u_0_2[4]), .Z(
        simpleXor_55_port_z) );
  XOR2_X1 simpleXor_56_U1 ( .A(n_zz_io_c_1_19[1]), .B(u_1_0[4]), .Z(
        simpleXor_56_port_z) );
  XOR2_X1 simpleXor_57_U1 ( .A(n_zz_io_c_1_19[2]), .B(u_1_2[4]), .Z(
        simpleXor_57_port_z) );
  XOR2_X1 simpleXor_58_U1 ( .A(n_zz_io_c_2_19[1]), .B(u_2_0[4]), .Z(
        simpleXor_58_port_z) );
  XOR2_X1 simpleXor_59_U1 ( .A(n_zz_io_c_2_19[2]), .B(u_2_1[4]), .Z(
        simpleXor_59_port_z) );
endmodule

