
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, p_rand_0, 
        p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7, 
        p_rand_8, p_rand_9, io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4
 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, p_rand_0, p_rand_1,
         p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7, p_rand_8,
         p_rand_9;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4;
  wire   n_dom_0_n45, n_dom_0_n44, n_dom_0_n43, n_dom_0_n42, n_dom_0_n41,
         n_dom_0_n40, n_dom_0_n39, n_dom_0_n38, n_dom_0_n37, n_dom_0_n36,
         n_dom_0_n35, n_dom_0_n34, n_dom_0_n33, n_dom_0_n32, n_dom_0_n31,
         n_dom_0_n30, n_dom_0_n29, n_dom_0_n28, n_dom_0_n27, n_dom_0_n26,
         n_dom_0_n25, n_dom_0_n24, n_dom_0_n23, n_dom_0_n22, n_dom_0_n21,
         n_dom_0_n20, n_dom_0_n19, n_dom_0_n18, n_dom_0_n17, n_dom_0_n16,
         n_dom_0_n15, n_dom_0_n14, n_dom_0_n13, n_dom_0_n12, n_dom_0_n11,
         n_dom_0_n10, n_dom_0_n9, n_dom_0_n8, n_dom_0_n7, n_dom_0_n6,
         n_dom_0_n5, n_dom_0_n4, n_dom_0_n3, n_dom_0_n2, n_dom_0_n1,
         n_dom_0_N29, n_dom_0_N28, n_dom_0_N27, n_dom_0_N26, n_dom_0_N25,
         n_dom_0_N24, n_dom_0__dom_inter4_2, n_dom_0__dom_inter4,
         n_dom_0_reg_pipeline, n_dom_0_N23, n_dom_0__dom_inter3_6,
         n_dom_0__dom_inter3, n_dom_0_reg_pipeline_3, n_dom_0_N22,
         n_dom_0__dom_inter2_9, n_dom_0__dom_inter2, n_dom_0_reg_pipeline_7,
         n_dom_0_N21, n_dom_0__dom_inter1_14, n_dom_0__dom_inter1,
         n_dom_0_reg_pipeline_11, n_dom_0_N20, n_dom_0__dom_inter0_18,
         n_dom_0__dom_inter0, n_dom_0_reg_pipeline_15, n_dom_0_N19,
         n_dom_0_N18, n_dom_0_N17, n_dom_0_N16, n_dom_0_N15, n_dom_0_N14,
         n_dom_0_N13, n_dom_0_N12, n_dom_0_N11, n_dom_0_N10, n_dom_0_N9,
         n_dom_0_N8, n_dom_0_N7, n_dom_0_N6, n_dom_0_N5, n_dom_0_N4,
         n_dom_0_N3, n_dom_0_N2, n_dom_0_N1, n_dom_0_N0;

  NAND2_X1 u_dom_0_U67 ( .A1(io_i0_s0), .A2(io_i1_s4), .ZN(n_dom_0_n35) );
  XNOR2_X1 u_dom_0_U66 ( .A(p_rand_3), .B(n_dom_0_n35), .ZN(n_dom_0_N0) );
  NAND2_X1 u_dom_0_U65 ( .A1(io_i0_s0), .A2(io_i1_s3), .ZN(n_dom_0_n34) );
  XNOR2_X1 u_dom_0_U64 ( .A(p_rand_2), .B(n_dom_0_n34), .ZN(n_dom_0_N1) );
  NAND2_X1 u_dom_0_U63 ( .A1(io_i1_s3), .A2(io_i0_s2), .ZN(n_dom_0_n33) );
  XNOR2_X1 u_dom_0_U62 ( .A(p_rand_7), .B(n_dom_0_n33), .ZN(n_dom_0_N10) );
  NAND2_X1 u_dom_0_U61 ( .A1(io_i1_s1), .A2(io_i0_s2), .ZN(n_dom_0_n32) );
  XNOR2_X1 u_dom_0_U60 ( .A(p_rand_4), .B(n_dom_0_n32), .ZN(n_dom_0_N11) );
  NAND2_X1 u_dom_0_U59 ( .A1(io_i0_s3), .A2(io_i1_s4), .ZN(n_dom_0_n31) );
  XNOR2_X1 u_dom_0_U58 ( .A(p_rand_9), .B(n_dom_0_n31), .ZN(n_dom_0_N12) );
  NAND2_X1 u_dom_0_U57 ( .A1(io_i0_s3), .A2(io_i1_s2), .ZN(n_dom_0_n30) );
  XNOR2_X1 u_dom_0_U56 ( .A(p_rand_7), .B(n_dom_0_n30), .ZN(n_dom_0_N13) );
  NAND2_X1 u_dom_0_U55 ( .A1(io_i0_s3), .A2(io_i1_s1), .ZN(n_dom_0_n29) );
  XNOR2_X1 u_dom_0_U54 ( .A(p_rand_5), .B(n_dom_0_n29), .ZN(n_dom_0_N14) );
  NAND2_X1 u_dom_0_U53 ( .A1(io_i0_s3), .A2(io_i1_s0), .ZN(n_dom_0_n28) );
  XNOR2_X1 u_dom_0_U52 ( .A(p_rand_2), .B(n_dom_0_n28), .ZN(n_dom_0_N15) );
  NAND2_X1 u_dom_0_U51 ( .A1(io_i0_s4), .A2(io_i1_s3), .ZN(n_dom_0_n27) );
  XNOR2_X1 u_dom_0_U50 ( .A(p_rand_9), .B(n_dom_0_n27), .ZN(n_dom_0_N16) );
  NAND2_X1 u_dom_0_U49 ( .A1(io_i0_s4), .A2(io_i1_s2), .ZN(n_dom_0_n26) );
  XNOR2_X1 u_dom_0_U48 ( .A(p_rand_8), .B(n_dom_0_n26), .ZN(n_dom_0_N17) );
  NAND2_X1 u_dom_0_U47 ( .A1(io_i0_s4), .A2(io_i1_s1), .ZN(n_dom_0_n25) );
  XNOR2_X1 u_dom_0_U46 ( .A(p_rand_6), .B(n_dom_0_n25), .ZN(n_dom_0_N18) );
  NAND2_X1 u_dom_0_U45 ( .A1(io_i0_s4), .A2(io_i1_s0), .ZN(n_dom_0_n24) );
  XNOR2_X1 u_dom_0_U44 ( .A(p_rand_3), .B(n_dom_0_n24), .ZN(n_dom_0_N19) );
  NAND2_X1 u_dom_0_U43 ( .A1(io_i0_s0), .A2(io_i1_s2), .ZN(n_dom_0_n23) );
  XNOR2_X1 u_dom_0_U42 ( .A(p_rand_1), .B(n_dom_0_n23), .ZN(n_dom_0_N2) );
  XOR2_X1 u_dom_0_U41 ( .A(n_dom_0__dom_inter0), .B(n_dom_0_reg_pipeline_15), 
        .Z(n_dom_0_n22) );
  XOR2_X1 u_dom_0_U40 ( .A(n_dom_0_n22), .B(n_dom_0_n44), .Z(n_dom_0_n20) );
  XOR2_X1 u_dom_0_U39 ( .A(n_dom_0__dom_inter0_18), .B(n_dom_0_n45), .Z(
        n_dom_0_n21) );
  XOR2_X1 u_dom_0_U38 ( .A(n_dom_0_n20), .B(n_dom_0_n21), .Z(n_dom_0_N20) );
  XOR2_X1 u_dom_0_U37 ( .A(n_dom_0__dom_inter1), .B(n_dom_0_reg_pipeline_11), 
        .Z(n_dom_0_n19) );
  XOR2_X1 u_dom_0_U36 ( .A(n_dom_0_n19), .B(n_dom_0_n42), .Z(n_dom_0_n17) );
  XOR2_X1 u_dom_0_U35 ( .A(n_dom_0__dom_inter1_14), .B(n_dom_0_n43), .Z(
        n_dom_0_n18) );
  XOR2_X1 u_dom_0_U34 ( .A(n_dom_0_n17), .B(n_dom_0_n18), .Z(n_dom_0_N21) );
  XOR2_X1 u_dom_0_U33 ( .A(n_dom_0__dom_inter2), .B(n_dom_0_reg_pipeline_7), 
        .Z(n_dom_0_n16) );
  XOR2_X1 u_dom_0_U32 ( .A(n_dom_0_n16), .B(n_dom_0_n40), .Z(n_dom_0_n14) );
  XOR2_X1 u_dom_0_U31 ( .A(n_dom_0__dom_inter2_9), .B(n_dom_0_n41), .Z(
        n_dom_0_n15) );
  XOR2_X1 u_dom_0_U30 ( .A(n_dom_0_n14), .B(n_dom_0_n15), .Z(n_dom_0_N22) );
  XOR2_X1 u_dom_0_U29 ( .A(n_dom_0__dom_inter3), .B(n_dom_0_reg_pipeline_3), 
        .Z(n_dom_0_n13) );
  XOR2_X1 u_dom_0_U28 ( .A(n_dom_0_n13), .B(n_dom_0_n38), .Z(n_dom_0_n11) );
  XOR2_X1 u_dom_0_U27 ( .A(n_dom_0__dom_inter3_6), .B(n_dom_0_n39), .Z(
        n_dom_0_n12) );
  XOR2_X1 u_dom_0_U26 ( .A(n_dom_0_n11), .B(n_dom_0_n12), .Z(n_dom_0_N23) );
  XOR2_X1 u_dom_0_U25 ( .A(n_dom_0__dom_inter4), .B(n_dom_0_reg_pipeline), .Z(
        n_dom_0_n10) );
  XOR2_X1 u_dom_0_U24 ( .A(n_dom_0_n10), .B(n_dom_0_n36), .Z(n_dom_0_n8) );
  XOR2_X1 u_dom_0_U23 ( .A(n_dom_0__dom_inter4_2), .B(n_dom_0_n37), .Z(
        n_dom_0_n9) );
  XOR2_X1 u_dom_0_U22 ( .A(n_dom_0_n8), .B(n_dom_0_n9), .Z(n_dom_0_N24) );
  AND2_X1 u_dom_0_U21 ( .A1(io_i1_s4), .A2(io_i0_s4), .ZN(n_dom_0_N25) );
  AND2_X1 u_dom_0_U20 ( .A1(io_i0_s1), .A2(io_i1_s1), .ZN(n_dom_0_N26) );
  AND2_X1 u_dom_0_U19 ( .A1(io_i1_s0), .A2(io_i0_s0), .ZN(n_dom_0_N27) );
  AND2_X1 u_dom_0_U18 ( .A1(io_i1_s3), .A2(io_i0_s3), .ZN(n_dom_0_N28) );
  AND2_X1 u_dom_0_U17 ( .A1(io_i0_s2), .A2(io_i1_s2), .ZN(n_dom_0_N29) );
  NAND2_X1 u_dom_0_U16 ( .A1(io_i1_s1), .A2(io_i0_s0), .ZN(n_dom_0_n7) );
  XNOR2_X1 u_dom_0_U15 ( .A(p_rand_0), .B(n_dom_0_n7), .ZN(n_dom_0_N3) );
  NAND2_X1 u_dom_0_U14 ( .A1(io_i0_s1), .A2(io_i1_s4), .ZN(n_dom_0_n6) );
  XNOR2_X1 u_dom_0_U13 ( .A(p_rand_6), .B(n_dom_0_n6), .ZN(n_dom_0_N4) );
  NAND2_X1 u_dom_0_U12 ( .A1(io_i1_s3), .A2(io_i0_s1), .ZN(n_dom_0_n5) );
  XNOR2_X1 u_dom_0_U11 ( .A(p_rand_5), .B(n_dom_0_n5), .ZN(n_dom_0_N5) );
  NAND2_X1 u_dom_0_U10 ( .A1(io_i1_s2), .A2(io_i0_s1), .ZN(n_dom_0_n4) );
  XNOR2_X1 u_dom_0_U9 ( .A(p_rand_4), .B(n_dom_0_n4), .ZN(n_dom_0_N6) );
  NAND2_X1 u_dom_0_U8 ( .A1(io_i0_s1), .A2(io_i1_s0), .ZN(n_dom_0_n3) );
  XNOR2_X1 u_dom_0_U7 ( .A(p_rand_0), .B(n_dom_0_n3), .ZN(n_dom_0_N7) );
  NAND2_X1 u_dom_0_U6 ( .A1(io_i1_s4), .A2(io_i0_s2), .ZN(n_dom_0_n2) );
  XNOR2_X1 u_dom_0_U5 ( .A(p_rand_8), .B(n_dom_0_n2), .ZN(n_dom_0_N8) );
  NAND2_X1 u_dom_0_U4 ( .A1(io_i1_s0), .A2(io_i0_s2), .ZN(n_dom_0_n1) );
  XNOR2_X1 u_dom_0_U3 ( .A(p_rand_1), .B(n_dom_0_n1), .ZN(n_dom_0_N9) );
  DFF_X1 u_dom_0_dom_out1_reg ( .D(n_dom_0_N21), .CK(clock_0), .Q(io_o0_s1), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter1_13_reg ( .D(n_dom_0_N6), .CK(clock_0), .Q(), .QN(
        n_dom_0_n43) );
  DFF_X1 u_dom_0_dom_out4_reg ( .D(n_dom_0_N24), .CK(clock_0), .Q(io_o0_s4), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter4_1_reg ( .D(n_dom_0_N18), .CK(clock_0), .Q(), .QN(
        n_dom_0_n37) );
  DFF_X1 u_dom_0__dom_inter4_2_reg ( .D(n_dom_0_N19), .CK(clock_0), .Q(
        n_dom_0__dom_inter4_2), .QN() );
  DFF_X1 u_dom_0_dom_out3_reg ( .D(n_dom_0_N23), .CK(clock_0), .Q(io_o0_s3), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter3_4_reg ( .D(n_dom_0_N13), .CK(clock_0), .Q(), .QN(
        n_dom_0_n38) );
  DFF_X1 u_dom_0_dom_out2_reg ( .D(n_dom_0_N22), .CK(clock_0), .Q(io_o0_s2), 
        .QN() );
  DFF_X1 u_dom_0_reg_pipeline_7_reg ( .D(n_dom_0_N29), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_7), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_3_reg ( .D(n_dom_0_N28), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_3), .QN() );
  DFF_X1 u_dom_0__dom_inter4_reg ( .D(n_dom_0_N16), .CK(clock_0), .Q(
        n_dom_0__dom_inter4), .QN() );
  DFF_X1 u_dom_0__dom_inter2_reg ( .D(n_dom_0_N8), .CK(clock_0), .Q(
        n_dom_0__dom_inter2), .QN() );
  DFF_X1 u_dom_0_dom_out0_reg ( .D(n_dom_0_N20), .CK(clock_0), .Q(io_o0_s0), 
        .QN() );
  DFF_X1 u_dom_0_reg_pipeline_15_reg ( .D(n_dom_0_N27), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_15), .QN() );
  DFF_X1 u_dom_0__dom_inter1_reg ( .D(n_dom_0_N4), .CK(clock_0), .Q(
        n_dom_0__dom_inter1), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_11_reg ( .D(n_dom_0_N26), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_11), .QN() );
  DFF_X1 u_dom_0__dom_inter3_reg ( .D(n_dom_0_N12), .CK(clock_0), .Q(
        n_dom_0__dom_inter3), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_reg ( .D(n_dom_0_N25), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline), .QN() );
  DFF_X1 u_dom_0__dom_inter0_reg ( .D(n_dom_0_N0), .CK(clock_0), .Q(
        n_dom_0__dom_inter0), .QN() );
  DFF_X1 u_dom_0__dom_inter4_0_reg ( .D(n_dom_0_N17), .CK(clock_0), .Q(), .QN(
        n_dom_0_n36) );
  DFF_X1 u_dom_0__dom_inter0_17_reg ( .D(n_dom_0_N2), .CK(clock_0), .Q(), .QN(
        n_dom_0_n45) );
  DFF_X1 u_dom_0__dom_inter2_8_reg ( .D(n_dom_0_N10), .CK(clock_0), .Q(), .QN(
        n_dom_0_n41) );
  DFF_X1 u_dom_0__dom_inter0_18_reg ( .D(n_dom_0_N3), .CK(clock_0), .Q(
        n_dom_0__dom_inter0_18), .QN() );
  DFF_X1 u_dom_0__dom_inter2_9_reg ( .D(n_dom_0_N11), .CK(clock_0), .Q(
        n_dom_0__dom_inter2_9), .QN() );
  DFF_X1 u_dom_0__dom_inter2_10_reg ( .D(n_dom_0_N9), .CK(clock_0), .Q(), .QN(
        n_dom_0_n40) );
  DFF_X1 u_dom_0__dom_inter3_5_reg ( .D(n_dom_0_N14), .CK(clock_0), .Q(), .QN(
        n_dom_0_n39) );
  DFF_X1 u_dom_0__dom_inter1_14_reg ( .D(n_dom_0_N7), .CK(clock_0), .Q(
        n_dom_0__dom_inter1_14), .QN() );
  DFF_X1 u_dom_0__dom_inter3_6_reg ( .D(n_dom_0_N15), .CK(clock_0), .Q(
        n_dom_0__dom_inter3_6), .QN() );
  DFF_X1 u_dom_0__dom_inter0_16_reg ( .D(n_dom_0_N1), .CK(clock_0), .Q(), .QN(
        n_dom_0_n44) );
  DFF_X1 u_dom_0__dom_inter1_12_reg ( .D(n_dom_0_N5), .CK(clock_0), .Q(), .QN(
        n_dom_0_n42) );
endmodule

