
module sharedSbox_PL ( clk, A, PRNGQ, Q );
  input [23:0] A;
  input [51:0] PRNGQ;
  output [23:0] Q;
  input clk;
  wire   Zl_f1_11_, Zl_f1_9_, Zl_f1_8_, Zl_f1_7_, Zl_f1_5_, Zl_f1_4_, Zl_f1_3_,
         Zl_f1_1_, Zl_f1_0_, Inst_f1_linearMapping_n32,
         Inst_f1_linearMapping_n31, Inst_f1_linearMapping_n30,
         Inst_f1_linearMapping_n29, Inst_f1_linearMapping_n28,
         Inst_f1_linearMapping_n27, Inst_f1_linearMapping_n26,
         Inst_f1_linearMapping_n25, Inst_f1_linearMapping_n24,
         Inst_f1_linearMapping_n23, Inst_f1_linearMapping_n22,
         Inst_f1_linearMapping_n21, Inst_f1_linearMapping_n20,
         Inst_f1_linearMapping_n19, Inst_f1_linearMapping_n18,
         Inst_f1_linearMapping_n17, Inst_f1_linearMapping_n16,
         Inst_f1_linearMapping_n15, Inst_f1_linearMapping_n14,
         Inst_f1_linearMapping_n13, Inst_f1_linearMapping_n12,
         Inst_f1_phpplmul_himul_n98, Inst_f1_phpplmul_himul_n97,
         Inst_f1_phpplmul_himul_n96, Inst_f1_phpplmul_himul_n95,
         Inst_f1_phpplmul_himul_n94, Inst_f1_phpplmul_himul_n93,
         Inst_f1_phpplmul_himul_n92, Inst_f1_phpplmul_himul_n91,
         Inst_f1_phpplmul_himul_n90, Inst_f1_phpplmul_himul_n89,
         Inst_f1_phpplmul_himul_n88, Inst_f1_phpplmul_himul_n87,
         Inst_f1_phpplmul_himul_n86, Inst_f1_phpplmul_himul_n85,
         Inst_f1_phpplmul_himul_n84, Inst_f1_phpplmul_himul_n83,
         Inst_f1_phpplmul_himul_n82, Inst_f1_phpplmul_himul_n81,
         Inst_f1_phpplmul_himul_n80, Inst_f1_phpplmul_himul_n79,
         Inst_f1_phpplmul_himul_n78, Inst_f1_phpplmul_himul_n77,
         Inst_f1_phpplmul_himul_n76, Inst_f1_phpplmul_himul_n75,
         Inst_f1_phpplmul_himul_n74, Inst_f1_phpplmul_himul_n73,
         Inst_f1_phpplmul_himul_n72, Inst_f1_phpplmul_himul_n71,
         Inst_f1_phpplmul_himul_n70, Inst_f1_phpplmul_himul_n69,
         Inst_f1_phpplmul_himul_n68, Inst_f1_phpplmul_himul_n67,
         Inst_f1_phpplmul_himul_n66, Inst_f1_phpplmul_himul_n65,
         Inst_f1_phpplmul_himul_n64, Inst_f1_phpplmul_himul_n63,
         Inst_f1_phpplmul_himul_n62, Inst_f1_phpplmul_himul_n61,
         Inst_f1_phpplmul_himul_n60, Inst_f1_phpplmul_himul_n59,
         Inst_f1_phpplmul_himul_n58, Inst_f1_phpplmul_himul_n57,
         Inst_f1_phpplmul_himul_n56, Inst_f1_phpplmul_himul_n55,
         Inst_f1_phpplmul_himul_n54, Inst_f1_phpplmul_himul_n53,
         Inst_f1_phpplmul_himul_n52, Inst_f1_phpplmul_himul_n51,
         Inst_f1_phpplmul_himul_n50, Inst_f1_phpplmul_himul_n49,
         Inst_f1_phpplmul_himul_n48, Inst_f1_phpplmul_himul_n47,
         Inst_f1_phpplmul_himul_n46, Inst_f1_phpplmul_himul_n45,
         Inst_f1_phpplmul_himul_n44, Inst_f1_phpplmul_himul_n43,
         Inst_f1_phpplmul_himul_n42, Inst_f1_phpplmul_himul_n41,
         Inst_f1_phpplmul_himul_n40, Inst_f1_phpplmul_himul_n39,
         Inst_f1_phpplmul_himul_n38, Inst_f1_phpplmul_himul_n37,
         Inst_f1_phpplmul_himul_n36, Inst_f1_phpplmul_himul_n35,
         Inst_f1_phpplmul_himul_n34, Inst_f1_phpplmul_himul_n33,
         Inst_f1_phpplmul_himul_n32, Inst_f1_phpplmul_himul_n31,
         Inst_f1_phpplmul_himul_n30, Inst_f1_phpplmul_himul_n29,
         Inst_f1_phpplmul_himul_n28, Inst_f1_phpplmul_himul_n27,
         Inst_f1_phpplmul_himul_n26, Inst_f1_phpplmul_himul_n25,
         Inst_f1_phpplmul_himul_n24, Inst_f1_phpplmul_himul_n23,
         Inst_f1_phpplmul_himul_n22, Inst_f1_phpplmul_himul_n21,
         Inst_f1_phpplmul_himul_n20, Inst_f1_phpplmul_himul_n19,
         Inst_f1_phpplmul_himul_n18, Inst_f1_phpplmul_himul_n17,
         Inst_f1_phpplmul_himul_n16, Inst_f1_phpplmul_himul_n15,
         Inst_f1_phpplmul_himul_n14, Inst_f1_phpplmul_himul_n13,
         Inst_f1_phpplmul_himul_n12, Inst_f1_phpplmul_himul_n11,
         Inst_f1_phpplmul_himul_n10, Inst_f1_phpplmul_himul_n9,
         Inst_f1_phpplmul_himul_n8, Inst_f1_phpplmul_himul_n7,
         Inst_f1_phpplmul_himul_n6, Inst_f1_phpplmul_himul_n5,
         Inst_f1_phpplmul_himul_n4, Inst_f1_phpplmul_himul_n3,
         Inst_f1_phpplmul_himul_n2, Inst_f1_phpplmul_himul_n1,
         Inst_f1_phpplmul_summul_n340, Inst_f1_phpplmul_summul_n339,
         Inst_f1_phpplmul_summul_n338, Inst_f1_phpplmul_summul_n337,
         Inst_f1_phpplmul_summul_n336, Inst_f1_phpplmul_summul_n335,
         Inst_f1_phpplmul_summul_n334, Inst_f1_phpplmul_summul_n333,
         Inst_f1_phpplmul_summul_n332, Inst_f1_phpplmul_summul_n331,
         Inst_f1_phpplmul_summul_n330, Inst_f1_phpplmul_summul_n329,
         Inst_f1_phpplmul_summul_n328, Inst_f1_phpplmul_summul_n327,
         Inst_f1_phpplmul_summul_n326, Inst_f1_phpplmul_summul_n325,
         Inst_f1_phpplmul_summul_n324, Inst_f1_phpplmul_summul_n323,
         Inst_f1_phpplmul_summul_n322, Inst_f1_phpplmul_summul_n321,
         Inst_f1_phpplmul_summul_n320, Inst_f1_phpplmul_summul_n319,
         Inst_f1_phpplmul_summul_n318, Inst_f1_phpplmul_summul_n317,
         Inst_f1_phpplmul_summul_n316, Inst_f1_phpplmul_summul_n315,
         Inst_f1_phpplmul_summul_n314, Inst_f1_phpplmul_summul_n313,
         Inst_f1_phpplmul_summul_n312, Inst_f1_phpplmul_summul_n311,
         Inst_f1_phpplmul_summul_n310, Inst_f1_phpplmul_summul_n309,
         Inst_f1_phpplmul_summul_n308, Inst_f1_phpplmul_summul_n307,
         Inst_f1_phpplmul_summul_n306, Inst_f1_phpplmul_summul_n305,
         Inst_f1_phpplmul_summul_n304, Inst_f1_phpplmul_summul_n303,
         Inst_f1_phpplmul_summul_n302, Inst_f1_phpplmul_summul_n301,
         Inst_f1_phpplmul_summul_n300, Inst_f1_phpplmul_summul_n299,
         Inst_f1_phpplmul_summul_n298, Inst_f1_phpplmul_summul_n297,
         Inst_f1_phpplmul_summul_n296, Inst_f1_phpplmul_summul_n295,
         Inst_f1_phpplmul_summul_n294, Inst_f1_phpplmul_summul_n293,
         Inst_f1_phpplmul_summul_n292, Inst_f1_phpplmul_summul_n291,
         Inst_f1_phpplmul_summul_n290, Inst_f1_phpplmul_summul_n289,
         Inst_f1_phpplmul_summul_n288, Inst_f1_phpplmul_summul_n287,
         Inst_f1_phpplmul_summul_n286, Inst_f1_phpplmul_summul_n285,
         Inst_f1_phpplmul_summul_n284, Inst_f1_phpplmul_summul_n283,
         Inst_f1_phpplmul_summul_n282, Inst_f1_phpplmul_summul_n281,
         Inst_f1_phpplmul_summul_n280, Inst_f1_phpplmul_summul_n279,
         Inst_f1_phpplmul_summul_n278, Inst_f1_phpplmul_summul_n277,
         Inst_f1_phpplmul_summul_n276, Inst_f1_phpplmul_summul_n275,
         Inst_f1_phpplmul_summul_n274, Inst_f1_phpplmul_summul_n273,
         Inst_f1_phpplmul_summul_n272, Inst_f1_phpplmul_summul_n271,
         Inst_f1_phpplmul_summul_n270, Inst_f1_phpplmul_summul_n269,
         Inst_f1_phpplmul_summul_n268, Inst_f1_phpplmul_summul_n267,
         Inst_f1_phpplmul_summul_n266, Inst_f1_phpplmul_summul_n265,
         Inst_f1_phpplmul_summul_n264, Inst_f1_phpplmul_summul_n263,
         Inst_f1_phpplmul_summul_n262, Inst_f1_phpplmul_summul_n261,
         Inst_f1_phpplmul_summul_n260, Inst_f1_phpplmul_summul_n259,
         Inst_f1_phpplmul_summul_n258, Inst_f1_phpplmul_summul_n257,
         Inst_f1_phpplmul_summul_n256, Inst_f1_phpplmul_summul_n255,
         Inst_f1_phpplmul_summul_n254, Inst_f1_phpplmul_summul_n253,
         Inst_f1_phpplmul_summul_n252, Inst_f1_phpplmul_summul_n251,
         Inst_f1_phpplmul_summul_n250, Inst_f1_phpplmul_summul_n249,
         Inst_f1_phpplmul_summul_n248, Inst_f1_phpplmul_summul_n247,
         Inst_f1_phpplmul_summul_n246, Inst_f1_phpplmul_summul_n245,
         Inst_f1_phpplmul_summul_n244, Inst_f1_phpplmul_summul_n243,
         Inst_f1_phpplmul_lowmul_n340, Inst_f1_phpplmul_lowmul_n339,
         Inst_f1_phpplmul_lowmul_n338, Inst_f1_phpplmul_lowmul_n337,
         Inst_f1_phpplmul_lowmul_n336, Inst_f1_phpplmul_lowmul_n335,
         Inst_f1_phpplmul_lowmul_n334, Inst_f1_phpplmul_lowmul_n333,
         Inst_f1_phpplmul_lowmul_n332, Inst_f1_phpplmul_lowmul_n331,
         Inst_f1_phpplmul_lowmul_n330, Inst_f1_phpplmul_lowmul_n329,
         Inst_f1_phpplmul_lowmul_n328, Inst_f1_phpplmul_lowmul_n327,
         Inst_f1_phpplmul_lowmul_n326, Inst_f1_phpplmul_lowmul_n325,
         Inst_f1_phpplmul_lowmul_n324, Inst_f1_phpplmul_lowmul_n323,
         Inst_f1_phpplmul_lowmul_n322, Inst_f1_phpplmul_lowmul_n321,
         Inst_f1_phpplmul_lowmul_n320, Inst_f1_phpplmul_lowmul_n319,
         Inst_f1_phpplmul_lowmul_n318, Inst_f1_phpplmul_lowmul_n317,
         Inst_f1_phpplmul_lowmul_n316, Inst_f1_phpplmul_lowmul_n315,
         Inst_f1_phpplmul_lowmul_n314, Inst_f1_phpplmul_lowmul_n313,
         Inst_f1_phpplmul_lowmul_n312, Inst_f1_phpplmul_lowmul_n311,
         Inst_f1_phpplmul_lowmul_n310, Inst_f1_phpplmul_lowmul_n309,
         Inst_f1_phpplmul_lowmul_n308, Inst_f1_phpplmul_lowmul_n307,
         Inst_f1_phpplmul_lowmul_n306, Inst_f1_phpplmul_lowmul_n305,
         Inst_f1_phpplmul_lowmul_n304, Inst_f1_phpplmul_lowmul_n303,
         Inst_f1_phpplmul_lowmul_n302, Inst_f1_phpplmul_lowmul_n301,
         Inst_f1_phpplmul_lowmul_n300, Inst_f1_phpplmul_lowmul_n299,
         Inst_f1_phpplmul_lowmul_n298, Inst_f1_phpplmul_lowmul_n297,
         Inst_f1_phpplmul_lowmul_n296, Inst_f1_phpplmul_lowmul_n295,
         Inst_f1_phpplmul_lowmul_n294, Inst_f1_phpplmul_lowmul_n293,
         Inst_f1_phpplmul_lowmul_n292, Inst_f1_phpplmul_lowmul_n291,
         Inst_f1_phpplmul_lowmul_n290, Inst_f1_phpplmul_lowmul_n289,
         Inst_f1_phpplmul_lowmul_n288, Inst_f1_phpplmul_lowmul_n287,
         Inst_f1_phpplmul_lowmul_n286, Inst_f1_phpplmul_lowmul_n285,
         Inst_f1_phpplmul_lowmul_n284, Inst_f1_phpplmul_lowmul_n283,
         Inst_f1_phpplmul_lowmul_n282, Inst_f1_phpplmul_lowmul_n281,
         Inst_f1_phpplmul_lowmul_n280, Inst_f1_phpplmul_lowmul_n279,
         Inst_f1_phpplmul_lowmul_n278, Inst_f1_phpplmul_lowmul_n277,
         Inst_f1_phpplmul_lowmul_n276, Inst_f1_phpplmul_lowmul_n275,
         Inst_f1_phpplmul_lowmul_n274, Inst_f1_phpplmul_lowmul_n273,
         Inst_f1_phpplmul_lowmul_n272, Inst_f1_phpplmul_lowmul_n271,
         Inst_f1_phpplmul_lowmul_n270, Inst_f1_phpplmul_lowmul_n269,
         Inst_f1_phpplmul_lowmul_n268, Inst_f1_phpplmul_lowmul_n267,
         Inst_f1_phpplmul_lowmul_n266, Inst_f1_phpplmul_lowmul_n265,
         Inst_f1_phpplmul_lowmul_n264, Inst_f1_phpplmul_lowmul_n263,
         Inst_f1_phpplmul_lowmul_n262, Inst_f1_phpplmul_lowmul_n261,
         Inst_f1_phpplmul_lowmul_n260, Inst_f1_phpplmul_lowmul_n259,
         Inst_f1_phpplmul_lowmul_n258, Inst_f1_phpplmul_lowmul_n257,
         Inst_f1_phpplmul_lowmul_n256, Inst_f1_phpplmul_lowmul_n255,
         Inst_f1_phpplmul_lowmul_n254, Inst_f1_phpplmul_lowmul_n253,
         Inst_f1_phpplmul_lowmul_n252, Inst_f1_phpplmul_lowmul_n251,
         Inst_f1_phpplmul_lowmul_n250, Inst_f1_phpplmul_lowmul_n249,
         Inst_f1_phpplmul_lowmul_n248, Inst_f1_phpplmul_lowmul_n247,
         Inst_f1_phpplmul_lowmul_n246, Inst_f1_phpplmul_lowmul_n245,
         Inst_f1_phpplmul_lowmul_n244, Inst_f1_phpplmul_lowmul_n243,
         Inst_f2_abmul_pw2_0_, Inst_f2_abmul_pw2_1_, Inst_f2_abmul_pw2_2_,
         Inst_f2_abmul_pw2_3_, Inst_f2_abmul_pw2_4_, Inst_f2_abmul_pw2_5_,
         Inst_f2_dinv_1_mul_n340, Inst_f2_dinv_1_mul_n339,
         Inst_f2_dinv_1_mul_n338, Inst_f2_dinv_1_mul_n337,
         Inst_f2_dinv_1_mul_n336, Inst_f2_dinv_1_mul_n335,
         Inst_f2_dinv_1_mul_n334, Inst_f2_dinv_1_mul_n333,
         Inst_f2_dinv_1_mul_n332, Inst_f2_dinv_1_mul_n331,
         Inst_f2_dinv_1_mul_n330, Inst_f2_dinv_1_mul_n329,
         Inst_f2_dinv_1_mul_n328, Inst_f2_dinv_1_mul_n327,
         Inst_f2_dinv_1_mul_n326, Inst_f2_dinv_1_mul_n325,
         Inst_f2_dinv_1_mul_n324, Inst_f2_dinv_1_mul_n323,
         Inst_f2_dinv_1_mul_n322, Inst_f2_dinv_1_mul_n321,
         Inst_f2_dinv_1_mul_n320, Inst_f2_dinv_1_mul_n319,
         Inst_f2_dinv_1_mul_n318, Inst_f2_dinv_1_mul_n317,
         Inst_f2_dinv_1_mul_n316, Inst_f2_dinv_1_mul_n315,
         Inst_f2_dinv_1_mul_n314, Inst_f2_dinv_1_mul_n313,
         Inst_f2_dinv_1_mul_n312, Inst_f2_dinv_1_mul_n311,
         Inst_f2_dinv_1_mul_n310, Inst_f2_dinv_1_mul_n309,
         Inst_f2_dinv_1_mul_n308, Inst_f2_dinv_1_mul_n307,
         Inst_f2_dinv_1_mul_n306, Inst_f2_dinv_1_mul_n305,
         Inst_f2_dinv_1_mul_n304, Inst_f2_dinv_1_mul_n303,
         Inst_f2_dinv_1_mul_n302, Inst_f2_dinv_1_mul_n301,
         Inst_f2_dinv_1_mul_n300, Inst_f2_dinv_1_mul_n299,
         Inst_f2_dinv_1_mul_n298, Inst_f2_dinv_1_mul_n297,
         Inst_f2_dinv_1_mul_n296, Inst_f2_dinv_1_mul_n295,
         Inst_f2_dinv_1_mul_n294, Inst_f2_dinv_1_mul_n293,
         Inst_f2_dinv_1_mul_n292, Inst_f2_dinv_1_mul_n291,
         Inst_f2_dinv_1_mul_n290, Inst_f2_dinv_1_mul_n289,
         Inst_f2_dinv_1_mul_n288, Inst_f2_dinv_1_mul_n287,
         Inst_f2_dinv_1_mul_n286, Inst_f2_dinv_1_mul_n285,
         Inst_f2_dinv_1_mul_n284, Inst_f2_dinv_1_mul_n283,
         Inst_f2_dinv_1_mul_n282, Inst_f2_dinv_1_mul_n281,
         Inst_f2_dinv_1_mul_n280, Inst_f2_dinv_1_mul_n279,
         Inst_f2_dinv_1_mul_n278, Inst_f2_dinv_1_mul_n277,
         Inst_f2_dinv_1_mul_n276, Inst_f2_dinv_1_mul_n275,
         Inst_f2_dinv_1_mul_n274, Inst_f2_dinv_1_mul_n273,
         Inst_f2_dinv_1_mul_n272, Inst_f2_dinv_1_mul_n271,
         Inst_f2_dinv_1_mul_n270, Inst_f2_dinv_1_mul_n269,
         Inst_f2_dinv_1_mul_n268, Inst_f2_dinv_1_mul_n267,
         Inst_f2_dinv_1_mul_n266, Inst_f2_dinv_1_mul_n265,
         Inst_f2_dinv_1_mul_n264, Inst_f2_dinv_1_mul_n263,
         Inst_f2_dinv_1_mul_n262, Inst_f2_dinv_1_mul_n261,
         Inst_f2_dinv_1_mul_n260, Inst_f2_dinv_1_mul_n259,
         Inst_f2_dinv_1_mul_n258, Inst_f2_dinv_1_mul_n257,
         Inst_f2_dinv_1_mul_n256, Inst_f2_dinv_1_mul_n255,
         Inst_f2_dinv_1_mul_n254, Inst_f2_dinv_1_mul_n253,
         Inst_f2_dinv_1_mul_n252, Inst_f2_dinv_1_mul_n251,
         Inst_f2_dinv_1_mul_n250, Inst_f2_dinv_1_mul_n249,
         Inst_f2_dinv_1_mul_n248, Inst_f2_dinv_1_mul_n247,
         Inst_f2_dinv_1_mul_n246, Inst_f2_dinv_1_mul_n245,
         Inst_f2_dinv_1_mul_n244, Inst_f2_dinv_1_mul_n243, Inst_f3_dinv_2_d_0_,
         Inst_f3_dinv_2_d_1_, Inst_f3_dinv_2_d_2_, Inst_f3_dinv_2_d_3_,
         Inst_f3_dinv_2_d_4_, Inst_f3_dinv_2_d_5_, Inst_f3_dinv_2_himul_n341,
         Inst_f3_dinv_2_himul_n340, Inst_f3_dinv_2_himul_n339,
         Inst_f3_dinv_2_himul_n338, Inst_f3_dinv_2_himul_n337,
         Inst_f3_dinv_2_himul_n336, Inst_f3_dinv_2_himul_n335,
         Inst_f3_dinv_2_himul_n334, Inst_f3_dinv_2_himul_n333,
         Inst_f3_dinv_2_himul_n332, Inst_f3_dinv_2_himul_n331,
         Inst_f3_dinv_2_himul_n330, Inst_f3_dinv_2_himul_n329,
         Inst_f3_dinv_2_himul_n328, Inst_f3_dinv_2_himul_n327,
         Inst_f3_dinv_2_himul_n326, Inst_f3_dinv_2_himul_n325,
         Inst_f3_dinv_2_himul_n324, Inst_f3_dinv_2_himul_n323,
         Inst_f3_dinv_2_himul_n322, Inst_f3_dinv_2_himul_n321,
         Inst_f3_dinv_2_himul_n320, Inst_f3_dinv_2_himul_n319,
         Inst_f3_dinv_2_himul_n318, Inst_f3_dinv_2_himul_n317,
         Inst_f3_dinv_2_himul_n316, Inst_f3_dinv_2_himul_n315,
         Inst_f3_dinv_2_himul_n314, Inst_f3_dinv_2_himul_n313,
         Inst_f3_dinv_2_himul_n312, Inst_f3_dinv_2_himul_n311,
         Inst_f3_dinv_2_himul_n310, Inst_f3_dinv_2_himul_n309,
         Inst_f3_dinv_2_himul_n308, Inst_f3_dinv_2_himul_n307,
         Inst_f3_dinv_2_himul_n306, Inst_f3_dinv_2_himul_n305,
         Inst_f3_dinv_2_himul_n304, Inst_f3_dinv_2_himul_n303,
         Inst_f3_dinv_2_himul_n302, Inst_f3_dinv_2_himul_n301,
         Inst_f3_dinv_2_himul_n300, Inst_f3_dinv_2_himul_n299,
         Inst_f3_dinv_2_himul_n298, Inst_f3_dinv_2_himul_n297,
         Inst_f3_dinv_2_himul_n296, Inst_f3_dinv_2_himul_n295,
         Inst_f3_dinv_2_himul_n294, Inst_f3_dinv_2_himul_n293,
         Inst_f3_dinv_2_himul_n292, Inst_f3_dinv_2_himul_n291,
         Inst_f3_dinv_2_himul_n290, Inst_f3_dinv_2_himul_n289,
         Inst_f3_dinv_2_himul_n288, Inst_f3_dinv_2_himul_n287,
         Inst_f3_dinv_2_himul_n286, Inst_f3_dinv_2_himul_n285,
         Inst_f3_dinv_2_himul_n284, Inst_f3_dinv_2_himul_n283,
         Inst_f3_dinv_2_himul_n282, Inst_f3_dinv_2_himul_n281,
         Inst_f3_dinv_2_himul_n280, Inst_f3_dinv_2_himul_n279,
         Inst_f3_dinv_2_himul_n278, Inst_f3_dinv_2_himul_n277,
         Inst_f3_dinv_2_himul_n276, Inst_f3_dinv_2_himul_n275,
         Inst_f3_dinv_2_himul_n274, Inst_f3_dinv_2_himul_n273,
         Inst_f3_dinv_2_himul_n272, Inst_f3_dinv_2_himul_n271,
         Inst_f3_dinv_2_himul_n270, Inst_f3_dinv_2_himul_n269,
         Inst_f3_dinv_2_himul_n268, Inst_f3_dinv_2_himul_n267,
         Inst_f3_dinv_2_himul_n266, Inst_f3_dinv_2_himul_n265,
         Inst_f3_dinv_2_himul_n264, Inst_f3_dinv_2_himul_n263,
         Inst_f3_dinv_2_himul_n262, Inst_f3_dinv_2_himul_n261,
         Inst_f3_dinv_2_himul_n260, Inst_f3_dinv_2_himul_n259,
         Inst_f3_dinv_2_himul_n258, Inst_f3_dinv_2_himul_n257,
         Inst_f3_dinv_2_himul_n256, Inst_f3_dinv_2_himul_n255,
         Inst_f3_dinv_2_himul_n254, Inst_f3_dinv_2_himul_n253,
         Inst_f3_dinv_2_himul_n252, Inst_f3_dinv_2_himul_n251,
         Inst_f3_dinv_2_himul_n250, Inst_f3_dinv_2_himul_n249,
         Inst_f3_dinv_2_himul_n248, Inst_f3_dinv_2_himul_n247,
         Inst_f3_dinv_2_himul_n246, Inst_f3_dinv_2_himul_n245,
         Inst_f3_dinv_2_himul_n244, Inst_f3_dinv_2_lowmul_n340,
         Inst_f3_dinv_2_lowmul_n339, Inst_f3_dinv_2_lowmul_n338,
         Inst_f3_dinv_2_lowmul_n337, Inst_f3_dinv_2_lowmul_n336,
         Inst_f3_dinv_2_lowmul_n335, Inst_f3_dinv_2_lowmul_n334,
         Inst_f3_dinv_2_lowmul_n333, Inst_f3_dinv_2_lowmul_n332,
         Inst_f3_dinv_2_lowmul_n331, Inst_f3_dinv_2_lowmul_n330,
         Inst_f3_dinv_2_lowmul_n329, Inst_f3_dinv_2_lowmul_n328,
         Inst_f3_dinv_2_lowmul_n327, Inst_f3_dinv_2_lowmul_n326,
         Inst_f3_dinv_2_lowmul_n325, Inst_f3_dinv_2_lowmul_n324,
         Inst_f3_dinv_2_lowmul_n323, Inst_f3_dinv_2_lowmul_n322,
         Inst_f3_dinv_2_lowmul_n321, Inst_f3_dinv_2_lowmul_n320,
         Inst_f3_dinv_2_lowmul_n319, Inst_f3_dinv_2_lowmul_n318,
         Inst_f3_dinv_2_lowmul_n317, Inst_f3_dinv_2_lowmul_n316,
         Inst_f3_dinv_2_lowmul_n315, Inst_f3_dinv_2_lowmul_n314,
         Inst_f3_dinv_2_lowmul_n313, Inst_f3_dinv_2_lowmul_n312,
         Inst_f3_dinv_2_lowmul_n311, Inst_f3_dinv_2_lowmul_n310,
         Inst_f3_dinv_2_lowmul_n309, Inst_f3_dinv_2_lowmul_n308,
         Inst_f3_dinv_2_lowmul_n307, Inst_f3_dinv_2_lowmul_n306,
         Inst_f3_dinv_2_lowmul_n305, Inst_f3_dinv_2_lowmul_n304,
         Inst_f3_dinv_2_lowmul_n303, Inst_f3_dinv_2_lowmul_n302,
         Inst_f3_dinv_2_lowmul_n301, Inst_f3_dinv_2_lowmul_n300,
         Inst_f3_dinv_2_lowmul_n299, Inst_f3_dinv_2_lowmul_n298,
         Inst_f3_dinv_2_lowmul_n297, Inst_f3_dinv_2_lowmul_n296,
         Inst_f3_dinv_2_lowmul_n295, Inst_f3_dinv_2_lowmul_n294,
         Inst_f3_dinv_2_lowmul_n293, Inst_f3_dinv_2_lowmul_n292,
         Inst_f3_dinv_2_lowmul_n291, Inst_f3_dinv_2_lowmul_n290,
         Inst_f3_dinv_2_lowmul_n289, Inst_f3_dinv_2_lowmul_n288,
         Inst_f3_dinv_2_lowmul_n287, Inst_f3_dinv_2_lowmul_n286,
         Inst_f3_dinv_2_lowmul_n285, Inst_f3_dinv_2_lowmul_n284,
         Inst_f3_dinv_2_lowmul_n283, Inst_f3_dinv_2_lowmul_n282,
         Inst_f3_dinv_2_lowmul_n281, Inst_f3_dinv_2_lowmul_n280,
         Inst_f3_dinv_2_lowmul_n279, Inst_f3_dinv_2_lowmul_n278,
         Inst_f3_dinv_2_lowmul_n277, Inst_f3_dinv_2_lowmul_n276,
         Inst_f3_dinv_2_lowmul_n275, Inst_f3_dinv_2_lowmul_n274,
         Inst_f3_dinv_2_lowmul_n273, Inst_f3_dinv_2_lowmul_n272,
         Inst_f3_dinv_2_lowmul_n271, Inst_f3_dinv_2_lowmul_n270,
         Inst_f3_dinv_2_lowmul_n269, Inst_f3_dinv_2_lowmul_n268,
         Inst_f3_dinv_2_lowmul_n267, Inst_f3_dinv_2_lowmul_n266,
         Inst_f3_dinv_2_lowmul_n265, Inst_f3_dinv_2_lowmul_n264,
         Inst_f3_dinv_2_lowmul_n263, Inst_f3_dinv_2_lowmul_n262,
         Inst_f3_dinv_2_lowmul_n261, Inst_f3_dinv_2_lowmul_n260,
         Inst_f3_dinv_2_lowmul_n259, Inst_f3_dinv_2_lowmul_n258,
         Inst_f3_dinv_2_lowmul_n257, Inst_f3_dinv_2_lowmul_n256,
         Inst_f3_dinv_2_lowmul_n255, Inst_f3_dinv_2_lowmul_n254,
         Inst_f3_dinv_2_lowmul_n253, Inst_f3_dinv_2_lowmul_n252,
         Inst_f3_dinv_2_lowmul_n251, Inst_f3_dinv_2_lowmul_n250,
         Inst_f3_dinv_2_lowmul_n249, Inst_f3_dinv_2_lowmul_n248,
         Inst_f3_dinv_2_lowmul_n247, Inst_f3_dinv_2_lowmul_n246,
         Inst_f3_dinv_2_lowmul_n245, Inst_f3_dinv_2_lowmul_n244,
         Inst_f3_dinv_2_lowmul_n243, Inst_f4_multd_L_himul_n340,
         Inst_f4_multd_L_himul_n339, Inst_f4_multd_L_himul_n338,
         Inst_f4_multd_L_himul_n337, Inst_f4_multd_L_himul_n336,
         Inst_f4_multd_L_himul_n335, Inst_f4_multd_L_himul_n334,
         Inst_f4_multd_L_himul_n333, Inst_f4_multd_L_himul_n332,
         Inst_f4_multd_L_himul_n331, Inst_f4_multd_L_himul_n330,
         Inst_f4_multd_L_himul_n329, Inst_f4_multd_L_himul_n328,
         Inst_f4_multd_L_himul_n327, Inst_f4_multd_L_himul_n326,
         Inst_f4_multd_L_himul_n325, Inst_f4_multd_L_himul_n324,
         Inst_f4_multd_L_himul_n323, Inst_f4_multd_L_himul_n322,
         Inst_f4_multd_L_himul_n321, Inst_f4_multd_L_himul_n320,
         Inst_f4_multd_L_himul_n319, Inst_f4_multd_L_himul_n318,
         Inst_f4_multd_L_himul_n317, Inst_f4_multd_L_himul_n316,
         Inst_f4_multd_L_himul_n315, Inst_f4_multd_L_himul_n314,
         Inst_f4_multd_L_himul_n313, Inst_f4_multd_L_himul_n312,
         Inst_f4_multd_L_himul_n311, Inst_f4_multd_L_himul_n310,
         Inst_f4_multd_L_himul_n309, Inst_f4_multd_L_himul_n308,
         Inst_f4_multd_L_himul_n307, Inst_f4_multd_L_himul_n306,
         Inst_f4_multd_L_himul_n305, Inst_f4_multd_L_himul_n304,
         Inst_f4_multd_L_himul_n303, Inst_f4_multd_L_himul_n302,
         Inst_f4_multd_L_himul_n301, Inst_f4_multd_L_himul_n300,
         Inst_f4_multd_L_himul_n299, Inst_f4_multd_L_himul_n298,
         Inst_f4_multd_L_himul_n297, Inst_f4_multd_L_himul_n296,
         Inst_f4_multd_L_himul_n295, Inst_f4_multd_L_himul_n294,
         Inst_f4_multd_L_himul_n293, Inst_f4_multd_L_himul_n292,
         Inst_f4_multd_L_himul_n291, Inst_f4_multd_L_himul_n290,
         Inst_f4_multd_L_himul_n289, Inst_f4_multd_L_himul_n288,
         Inst_f4_multd_L_himul_n287, Inst_f4_multd_L_himul_n286,
         Inst_f4_multd_L_himul_n285, Inst_f4_multd_L_himul_n284,
         Inst_f4_multd_L_himul_n283, Inst_f4_multd_L_himul_n282,
         Inst_f4_multd_L_himul_n281, Inst_f4_multd_L_himul_n280,
         Inst_f4_multd_L_himul_n279, Inst_f4_multd_L_himul_n278,
         Inst_f4_multd_L_himul_n277, Inst_f4_multd_L_himul_n276,
         Inst_f4_multd_L_himul_n275, Inst_f4_multd_L_himul_n274,
         Inst_f4_multd_L_himul_n273, Inst_f4_multd_L_himul_n272,
         Inst_f4_multd_L_himul_n271, Inst_f4_multd_L_himul_n270,
         Inst_f4_multd_L_himul_n269, Inst_f4_multd_L_himul_n268,
         Inst_f4_multd_L_himul_n267, Inst_f4_multd_L_himul_n266,
         Inst_f4_multd_L_himul_n265, Inst_f4_multd_L_himul_n264,
         Inst_f4_multd_L_himul_n263, Inst_f4_multd_L_himul_n262,
         Inst_f4_multd_L_himul_n261, Inst_f4_multd_L_himul_n260,
         Inst_f4_multd_L_himul_n259, Inst_f4_multd_L_himul_n258,
         Inst_f4_multd_L_himul_n257, Inst_f4_multd_L_himul_n256,
         Inst_f4_multd_L_himul_n255, Inst_f4_multd_L_himul_n254,
         Inst_f4_multd_L_himul_n253, Inst_f4_multd_L_himul_n252,
         Inst_f4_multd_L_himul_n251, Inst_f4_multd_L_himul_n250,
         Inst_f4_multd_L_himul_n249, Inst_f4_multd_L_himul_n248,
         Inst_f4_multd_L_himul_n247, Inst_f4_multd_L_himul_n246,
         Inst_f4_multd_L_himul_n245, Inst_f4_multd_L_himul_n244,
         Inst_f4_multd_L_himul_n243, Inst_f4_multd_L_summul_n340,
         Inst_f4_multd_L_summul_n339, Inst_f4_multd_L_summul_n338,
         Inst_f4_multd_L_summul_n337, Inst_f4_multd_L_summul_n336,
         Inst_f4_multd_L_summul_n335, Inst_f4_multd_L_summul_n334,
         Inst_f4_multd_L_summul_n333, Inst_f4_multd_L_summul_n332,
         Inst_f4_multd_L_summul_n331, Inst_f4_multd_L_summul_n330,
         Inst_f4_multd_L_summul_n329, Inst_f4_multd_L_summul_n328,
         Inst_f4_multd_L_summul_n327, Inst_f4_multd_L_summul_n326,
         Inst_f4_multd_L_summul_n325, Inst_f4_multd_L_summul_n324,
         Inst_f4_multd_L_summul_n323, Inst_f4_multd_L_summul_n322,
         Inst_f4_multd_L_summul_n321, Inst_f4_multd_L_summul_n320,
         Inst_f4_multd_L_summul_n319, Inst_f4_multd_L_summul_n318,
         Inst_f4_multd_L_summul_n317, Inst_f4_multd_L_summul_n316,
         Inst_f4_multd_L_summul_n315, Inst_f4_multd_L_summul_n314,
         Inst_f4_multd_L_summul_n313, Inst_f4_multd_L_summul_n312,
         Inst_f4_multd_L_summul_n311, Inst_f4_multd_L_summul_n310,
         Inst_f4_multd_L_summul_n309, Inst_f4_multd_L_summul_n308,
         Inst_f4_multd_L_summul_n307, Inst_f4_multd_L_summul_n306,
         Inst_f4_multd_L_summul_n305, Inst_f4_multd_L_summul_n304,
         Inst_f4_multd_L_summul_n303, Inst_f4_multd_L_summul_n302,
         Inst_f4_multd_L_summul_n301, Inst_f4_multd_L_summul_n300,
         Inst_f4_multd_L_summul_n299, Inst_f4_multd_L_summul_n298,
         Inst_f4_multd_L_summul_n297, Inst_f4_multd_L_summul_n296,
         Inst_f4_multd_L_summul_n295, Inst_f4_multd_L_summul_n294,
         Inst_f4_multd_L_summul_n293, Inst_f4_multd_L_summul_n292,
         Inst_f4_multd_L_summul_n291, Inst_f4_multd_L_summul_n290,
         Inst_f4_multd_L_summul_n289, Inst_f4_multd_L_summul_n288,
         Inst_f4_multd_L_summul_n287, Inst_f4_multd_L_summul_n286,
         Inst_f4_multd_L_summul_n285, Inst_f4_multd_L_summul_n284,
         Inst_f4_multd_L_summul_n283, Inst_f4_multd_L_summul_n282,
         Inst_f4_multd_L_summul_n281, Inst_f4_multd_L_summul_n280,
         Inst_f4_multd_L_summul_n279, Inst_f4_multd_L_summul_n278,
         Inst_f4_multd_L_summul_n277, Inst_f4_multd_L_summul_n276,
         Inst_f4_multd_L_summul_n275, Inst_f4_multd_L_summul_n274,
         Inst_f4_multd_L_summul_n273, Inst_f4_multd_L_summul_n272,
         Inst_f4_multd_L_summul_n271, Inst_f4_multd_L_summul_n270,
         Inst_f4_multd_L_summul_n269, Inst_f4_multd_L_summul_n268,
         Inst_f4_multd_L_summul_n267, Inst_f4_multd_L_summul_n266,
         Inst_f4_multd_L_summul_n265, Inst_f4_multd_L_summul_n264,
         Inst_f4_multd_L_summul_n263, Inst_f4_multd_L_summul_n262,
         Inst_f4_multd_L_summul_n261, Inst_f4_multd_L_summul_n260,
         Inst_f4_multd_L_summul_n259, Inst_f4_multd_L_summul_n258,
         Inst_f4_multd_L_summul_n257, Inst_f4_multd_L_summul_n256,
         Inst_f4_multd_L_summul_n255, Inst_f4_multd_L_summul_n254,
         Inst_f4_multd_L_summul_n253, Inst_f4_multd_L_summul_n252,
         Inst_f4_multd_L_summul_n251, Inst_f4_multd_L_summul_n250,
         Inst_f4_multd_L_summul_n249, Inst_f4_multd_L_summul_n248,
         Inst_f4_multd_L_summul_n247, Inst_f4_multd_L_summul_n246,
         Inst_f4_multd_L_summul_n245, Inst_f4_multd_L_summul_n244,
         Inst_f4_multd_L_summul_n243, Inst_f4_multd_L_lowmul_n340,
         Inst_f4_multd_L_lowmul_n339, Inst_f4_multd_L_lowmul_n338,
         Inst_f4_multd_L_lowmul_n337, Inst_f4_multd_L_lowmul_n336,
         Inst_f4_multd_L_lowmul_n335, Inst_f4_multd_L_lowmul_n334,
         Inst_f4_multd_L_lowmul_n333, Inst_f4_multd_L_lowmul_n332,
         Inst_f4_multd_L_lowmul_n331, Inst_f4_multd_L_lowmul_n330,
         Inst_f4_multd_L_lowmul_n329, Inst_f4_multd_L_lowmul_n328,
         Inst_f4_multd_L_lowmul_n327, Inst_f4_multd_L_lowmul_n326,
         Inst_f4_multd_L_lowmul_n325, Inst_f4_multd_L_lowmul_n324,
         Inst_f4_multd_L_lowmul_n323, Inst_f4_multd_L_lowmul_n322,
         Inst_f4_multd_L_lowmul_n321, Inst_f4_multd_L_lowmul_n320,
         Inst_f4_multd_L_lowmul_n319, Inst_f4_multd_L_lowmul_n318,
         Inst_f4_multd_L_lowmul_n317, Inst_f4_multd_L_lowmul_n316,
         Inst_f4_multd_L_lowmul_n315, Inst_f4_multd_L_lowmul_n314,
         Inst_f4_multd_L_lowmul_n313, Inst_f4_multd_L_lowmul_n312,
         Inst_f4_multd_L_lowmul_n311, Inst_f4_multd_L_lowmul_n310,
         Inst_f4_multd_L_lowmul_n309, Inst_f4_multd_L_lowmul_n308,
         Inst_f4_multd_L_lowmul_n307, Inst_f4_multd_L_lowmul_n306,
         Inst_f4_multd_L_lowmul_n305, Inst_f4_multd_L_lowmul_n304,
         Inst_f4_multd_L_lowmul_n303, Inst_f4_multd_L_lowmul_n302,
         Inst_f4_multd_L_lowmul_n301, Inst_f4_multd_L_lowmul_n300,
         Inst_f4_multd_L_lowmul_n299, Inst_f4_multd_L_lowmul_n298,
         Inst_f4_multd_L_lowmul_n297, Inst_f4_multd_L_lowmul_n296,
         Inst_f4_multd_L_lowmul_n295, Inst_f4_multd_L_lowmul_n294,
         Inst_f4_multd_L_lowmul_n293, Inst_f4_multd_L_lowmul_n292,
         Inst_f4_multd_L_lowmul_n291, Inst_f4_multd_L_lowmul_n290,
         Inst_f4_multd_L_lowmul_n289, Inst_f4_multd_L_lowmul_n288,
         Inst_f4_multd_L_lowmul_n287, Inst_f4_multd_L_lowmul_n286,
         Inst_f4_multd_L_lowmul_n285, Inst_f4_multd_L_lowmul_n284,
         Inst_f4_multd_L_lowmul_n283, Inst_f4_multd_L_lowmul_n282,
         Inst_f4_multd_L_lowmul_n281, Inst_f4_multd_L_lowmul_n280,
         Inst_f4_multd_L_lowmul_n279, Inst_f4_multd_L_lowmul_n278,
         Inst_f4_multd_L_lowmul_n277, Inst_f4_multd_L_lowmul_n276,
         Inst_f4_multd_L_lowmul_n275, Inst_f4_multd_L_lowmul_n274,
         Inst_f4_multd_L_lowmul_n273, Inst_f4_multd_L_lowmul_n272,
         Inst_f4_multd_L_lowmul_n271, Inst_f4_multd_L_lowmul_n270,
         Inst_f4_multd_L_lowmul_n269, Inst_f4_multd_L_lowmul_n268,
         Inst_f4_multd_L_lowmul_n267, Inst_f4_multd_L_lowmul_n266,
         Inst_f4_multd_L_lowmul_n265, Inst_f4_multd_L_lowmul_n264,
         Inst_f4_multd_L_lowmul_n263, Inst_f4_multd_L_lowmul_n262,
         Inst_f4_multd_L_lowmul_n261, Inst_f4_multd_L_lowmul_n260,
         Inst_f4_multd_L_lowmul_n259, Inst_f4_multd_L_lowmul_n258,
         Inst_f4_multd_L_lowmul_n257, Inst_f4_multd_L_lowmul_n256,
         Inst_f4_multd_L_lowmul_n255, Inst_f4_multd_L_lowmul_n254,
         Inst_f4_multd_L_lowmul_n253, Inst_f4_multd_L_lowmul_n252,
         Inst_f4_multd_L_lowmul_n251, Inst_f4_multd_L_lowmul_n250,
         Inst_f4_multd_L_lowmul_n249, Inst_f4_multd_L_lowmul_n248,
         Inst_f4_multd_L_lowmul_n247, Inst_f4_multd_L_lowmul_n246,
         Inst_f4_multd_L_lowmul_n245, Inst_f4_multd_L_lowmul_n244,
         Inst_f4_multd_L_lowmul_n243, Inst_f4_multd_H_himul_n340,
         Inst_f4_multd_H_himul_n339, Inst_f4_multd_H_himul_n338,
         Inst_f4_multd_H_himul_n337, Inst_f4_multd_H_himul_n336,
         Inst_f4_multd_H_himul_n335, Inst_f4_multd_H_himul_n334,
         Inst_f4_multd_H_himul_n333, Inst_f4_multd_H_himul_n332,
         Inst_f4_multd_H_himul_n331, Inst_f4_multd_H_himul_n330,
         Inst_f4_multd_H_himul_n329, Inst_f4_multd_H_himul_n328,
         Inst_f4_multd_H_himul_n327, Inst_f4_multd_H_himul_n326,
         Inst_f4_multd_H_himul_n325, Inst_f4_multd_H_himul_n324,
         Inst_f4_multd_H_himul_n323, Inst_f4_multd_H_himul_n322,
         Inst_f4_multd_H_himul_n321, Inst_f4_multd_H_himul_n320,
         Inst_f4_multd_H_himul_n319, Inst_f4_multd_H_himul_n318,
         Inst_f4_multd_H_himul_n317, Inst_f4_multd_H_himul_n316,
         Inst_f4_multd_H_himul_n315, Inst_f4_multd_H_himul_n314,
         Inst_f4_multd_H_himul_n313, Inst_f4_multd_H_himul_n312,
         Inst_f4_multd_H_himul_n311, Inst_f4_multd_H_himul_n310,
         Inst_f4_multd_H_himul_n309, Inst_f4_multd_H_himul_n308,
         Inst_f4_multd_H_himul_n307, Inst_f4_multd_H_himul_n306,
         Inst_f4_multd_H_himul_n305, Inst_f4_multd_H_himul_n304,
         Inst_f4_multd_H_himul_n303, Inst_f4_multd_H_himul_n302,
         Inst_f4_multd_H_himul_n301, Inst_f4_multd_H_himul_n300,
         Inst_f4_multd_H_himul_n299, Inst_f4_multd_H_himul_n298,
         Inst_f4_multd_H_himul_n297, Inst_f4_multd_H_himul_n296,
         Inst_f4_multd_H_himul_n295, Inst_f4_multd_H_himul_n294,
         Inst_f4_multd_H_himul_n293, Inst_f4_multd_H_himul_n292,
         Inst_f4_multd_H_himul_n291, Inst_f4_multd_H_himul_n290,
         Inst_f4_multd_H_himul_n289, Inst_f4_multd_H_himul_n288,
         Inst_f4_multd_H_himul_n287, Inst_f4_multd_H_himul_n286,
         Inst_f4_multd_H_himul_n285, Inst_f4_multd_H_himul_n284,
         Inst_f4_multd_H_himul_n283, Inst_f4_multd_H_himul_n282,
         Inst_f4_multd_H_himul_n281, Inst_f4_multd_H_himul_n280,
         Inst_f4_multd_H_himul_n279, Inst_f4_multd_H_himul_n278,
         Inst_f4_multd_H_himul_n277, Inst_f4_multd_H_himul_n276,
         Inst_f4_multd_H_himul_n275, Inst_f4_multd_H_himul_n274,
         Inst_f4_multd_H_himul_n273, Inst_f4_multd_H_himul_n272,
         Inst_f4_multd_H_himul_n271, Inst_f4_multd_H_himul_n270,
         Inst_f4_multd_H_himul_n269, Inst_f4_multd_H_himul_n268,
         Inst_f4_multd_H_himul_n267, Inst_f4_multd_H_himul_n266,
         Inst_f4_multd_H_himul_n265, Inst_f4_multd_H_himul_n264,
         Inst_f4_multd_H_himul_n263, Inst_f4_multd_H_himul_n262,
         Inst_f4_multd_H_himul_n261, Inst_f4_multd_H_himul_n260,
         Inst_f4_multd_H_himul_n259, Inst_f4_multd_H_himul_n258,
         Inst_f4_multd_H_himul_n257, Inst_f4_multd_H_himul_n256,
         Inst_f4_multd_H_himul_n255, Inst_f4_multd_H_himul_n254,
         Inst_f4_multd_H_himul_n253, Inst_f4_multd_H_himul_n252,
         Inst_f4_multd_H_himul_n251, Inst_f4_multd_H_himul_n250,
         Inst_f4_multd_H_himul_n249, Inst_f4_multd_H_himul_n248,
         Inst_f4_multd_H_himul_n247, Inst_f4_multd_H_himul_n246,
         Inst_f4_multd_H_himul_n245, Inst_f4_multd_H_himul_n244,
         Inst_f4_multd_H_himul_n243, Inst_f4_multd_H_summul_n340,
         Inst_f4_multd_H_summul_n339, Inst_f4_multd_H_summul_n338,
         Inst_f4_multd_H_summul_n337, Inst_f4_multd_H_summul_n336,
         Inst_f4_multd_H_summul_n335, Inst_f4_multd_H_summul_n334,
         Inst_f4_multd_H_summul_n333, Inst_f4_multd_H_summul_n332,
         Inst_f4_multd_H_summul_n331, Inst_f4_multd_H_summul_n330,
         Inst_f4_multd_H_summul_n329, Inst_f4_multd_H_summul_n328,
         Inst_f4_multd_H_summul_n327, Inst_f4_multd_H_summul_n326,
         Inst_f4_multd_H_summul_n325, Inst_f4_multd_H_summul_n324,
         Inst_f4_multd_H_summul_n323, Inst_f4_multd_H_summul_n322,
         Inst_f4_multd_H_summul_n321, Inst_f4_multd_H_summul_n320,
         Inst_f4_multd_H_summul_n319, Inst_f4_multd_H_summul_n318,
         Inst_f4_multd_H_summul_n317, Inst_f4_multd_H_summul_n316,
         Inst_f4_multd_H_summul_n315, Inst_f4_multd_H_summul_n314,
         Inst_f4_multd_H_summul_n313, Inst_f4_multd_H_summul_n312,
         Inst_f4_multd_H_summul_n311, Inst_f4_multd_H_summul_n310,
         Inst_f4_multd_H_summul_n309, Inst_f4_multd_H_summul_n308,
         Inst_f4_multd_H_summul_n307, Inst_f4_multd_H_summul_n306,
         Inst_f4_multd_H_summul_n305, Inst_f4_multd_H_summul_n304,
         Inst_f4_multd_H_summul_n303, Inst_f4_multd_H_summul_n302,
         Inst_f4_multd_H_summul_n301, Inst_f4_multd_H_summul_n300,
         Inst_f4_multd_H_summul_n299, Inst_f4_multd_H_summul_n298,
         Inst_f4_multd_H_summul_n297, Inst_f4_multd_H_summul_n296,
         Inst_f4_multd_H_summul_n295, Inst_f4_multd_H_summul_n294,
         Inst_f4_multd_H_summul_n293, Inst_f4_multd_H_summul_n292,
         Inst_f4_multd_H_summul_n291, Inst_f4_multd_H_summul_n290,
         Inst_f4_multd_H_summul_n289, Inst_f4_multd_H_summul_n288,
         Inst_f4_multd_H_summul_n287, Inst_f4_multd_H_summul_n286,
         Inst_f4_multd_H_summul_n285, Inst_f4_multd_H_summul_n284,
         Inst_f4_multd_H_summul_n283, Inst_f4_multd_H_summul_n282,
         Inst_f4_multd_H_summul_n281, Inst_f4_multd_H_summul_n280,
         Inst_f4_multd_H_summul_n279, Inst_f4_multd_H_summul_n278,
         Inst_f4_multd_H_summul_n277, Inst_f4_multd_H_summul_n276,
         Inst_f4_multd_H_summul_n275, Inst_f4_multd_H_summul_n274,
         Inst_f4_multd_H_summul_n273, Inst_f4_multd_H_summul_n272,
         Inst_f4_multd_H_summul_n271, Inst_f4_multd_H_summul_n270,
         Inst_f4_multd_H_summul_n269, Inst_f4_multd_H_summul_n268,
         Inst_f4_multd_H_summul_n267, Inst_f4_multd_H_summul_n266,
         Inst_f4_multd_H_summul_n265, Inst_f4_multd_H_summul_n264,
         Inst_f4_multd_H_summul_n263, Inst_f4_multd_H_summul_n262,
         Inst_f4_multd_H_summul_n261, Inst_f4_multd_H_summul_n260,
         Inst_f4_multd_H_summul_n259, Inst_f4_multd_H_summul_n258,
         Inst_f4_multd_H_summul_n257, Inst_f4_multd_H_summul_n256,
         Inst_f4_multd_H_summul_n255, Inst_f4_multd_H_summul_n254,
         Inst_f4_multd_H_summul_n253, Inst_f4_multd_H_summul_n252,
         Inst_f4_multd_H_summul_n251, Inst_f4_multd_H_summul_n250,
         Inst_f4_multd_H_summul_n249, Inst_f4_multd_H_summul_n248,
         Inst_f4_multd_H_summul_n247, Inst_f4_multd_H_summul_n246,
         Inst_f4_multd_H_summul_n245, Inst_f4_multd_H_summul_n244,
         Inst_f4_multd_H_summul_n243, Inst_f4_multd_H_lowmul_n340,
         Inst_f4_multd_H_lowmul_n339, Inst_f4_multd_H_lowmul_n338,
         Inst_f4_multd_H_lowmul_n337, Inst_f4_multd_H_lowmul_n336,
         Inst_f4_multd_H_lowmul_n335, Inst_f4_multd_H_lowmul_n334,
         Inst_f4_multd_H_lowmul_n333, Inst_f4_multd_H_lowmul_n332,
         Inst_f4_multd_H_lowmul_n331, Inst_f4_multd_H_lowmul_n330,
         Inst_f4_multd_H_lowmul_n329, Inst_f4_multd_H_lowmul_n328,
         Inst_f4_multd_H_lowmul_n327, Inst_f4_multd_H_lowmul_n326,
         Inst_f4_multd_H_lowmul_n325, Inst_f4_multd_H_lowmul_n324,
         Inst_f4_multd_H_lowmul_n323, Inst_f4_multd_H_lowmul_n322,
         Inst_f4_multd_H_lowmul_n321, Inst_f4_multd_H_lowmul_n320,
         Inst_f4_multd_H_lowmul_n319, Inst_f4_multd_H_lowmul_n318,
         Inst_f4_multd_H_lowmul_n317, Inst_f4_multd_H_lowmul_n316,
         Inst_f4_multd_H_lowmul_n315, Inst_f4_multd_H_lowmul_n314,
         Inst_f4_multd_H_lowmul_n313, Inst_f4_multd_H_lowmul_n312,
         Inst_f4_multd_H_lowmul_n311, Inst_f4_multd_H_lowmul_n310,
         Inst_f4_multd_H_lowmul_n309, Inst_f4_multd_H_lowmul_n308,
         Inst_f4_multd_H_lowmul_n307, Inst_f4_multd_H_lowmul_n306,
         Inst_f4_multd_H_lowmul_n305, Inst_f4_multd_H_lowmul_n304,
         Inst_f4_multd_H_lowmul_n303, Inst_f4_multd_H_lowmul_n302,
         Inst_f4_multd_H_lowmul_n301, Inst_f4_multd_H_lowmul_n300,
         Inst_f4_multd_H_lowmul_n299, Inst_f4_multd_H_lowmul_n298,
         Inst_f4_multd_H_lowmul_n297, Inst_f4_multd_H_lowmul_n296,
         Inst_f4_multd_H_lowmul_n295, Inst_f4_multd_H_lowmul_n294,
         Inst_f4_multd_H_lowmul_n293, Inst_f4_multd_H_lowmul_n292,
         Inst_f4_multd_H_lowmul_n291, Inst_f4_multd_H_lowmul_n290,
         Inst_f4_multd_H_lowmul_n289, Inst_f4_multd_H_lowmul_n288,
         Inst_f4_multd_H_lowmul_n287, Inst_f4_multd_H_lowmul_n286,
         Inst_f4_multd_H_lowmul_n285, Inst_f4_multd_H_lowmul_n284,
         Inst_f4_multd_H_lowmul_n283, Inst_f4_multd_H_lowmul_n282,
         Inst_f4_multd_H_lowmul_n281, Inst_f4_multd_H_lowmul_n280,
         Inst_f4_multd_H_lowmul_n279, Inst_f4_multd_H_lowmul_n278,
         Inst_f4_multd_H_lowmul_n277, Inst_f4_multd_H_lowmul_n276,
         Inst_f4_multd_H_lowmul_n275, Inst_f4_multd_H_lowmul_n274,
         Inst_f4_multd_H_lowmul_n273, Inst_f4_multd_H_lowmul_n272,
         Inst_f4_multd_H_lowmul_n271, Inst_f4_multd_H_lowmul_n270,
         Inst_f4_multd_H_lowmul_n269, Inst_f4_multd_H_lowmul_n268,
         Inst_f4_multd_H_lowmul_n267, Inst_f4_multd_H_lowmul_n266,
         Inst_f4_multd_H_lowmul_n265, Inst_f4_multd_H_lowmul_n264,
         Inst_f4_multd_H_lowmul_n263, Inst_f4_multd_H_lowmul_n262,
         Inst_f4_multd_H_lowmul_n261, Inst_f4_multd_H_lowmul_n260,
         Inst_f4_multd_H_lowmul_n259, Inst_f4_multd_H_lowmul_n258,
         Inst_f4_multd_H_lowmul_n257, Inst_f4_multd_H_lowmul_n256,
         Inst_f4_multd_H_lowmul_n255, Inst_f4_multd_H_lowmul_n254,
         Inst_f4_multd_H_lowmul_n253, Inst_f4_multd_H_lowmul_n252,
         Inst_f4_multd_H_lowmul_n251, Inst_f4_multd_H_lowmul_n250,
         Inst_f4_multd_H_lowmul_n249, Inst_f4_multd_H_lowmul_n248,
         Inst_f4_multd_H_lowmul_n247, Inst_f4_multd_H_lowmul_n246,
         Inst_f4_multd_H_lowmul_n245, Inst_f4_multd_H_lowmul_n244,
         Inst_f4_multd_H_lowmul_n243, Inst_f5_phwillwin_pw2_0_,
         Inst_f5_phwillwin_pw2_1_, Inst_f5_phwillwin_pw2_2_,
         Inst_f5_phwillwin_pw2_3_, Inst_f5_phwillwin_pw2_4_,
         Inst_f5_phwillwin_pw2_5_, Inst_f5_plwillwin_pw2_0_,
         Inst_f5_plwillwin_pw2_1_, Inst_f5_plwillwin_pw2_2_,
         Inst_f5_plwillwin_pw2_3_, Inst_f5_plwillwin_pw2_4_,
         Inst_f5_plwillwin_pw2_5_, Inst_f5_invlinearMapping_n9,
         Inst_f5_invlinearMapping_n8, Inst_f5_invlinearMapping_n7,
         Inst_f5_invlinearMapping_n6, Inst_f5_invlinearMapping_n5,
         Inst_f5_invlinearMapping_n4, Inst_f5_invlinearMapping_n3,
         Inst_f5_invlinearMapping_n2, Inst_f5_invlinearMapping_n1;
  wire   [11:0] Zh_f1;
  wire   [11:0] ab2;
  wire   [5:0] ph;
  wire   [5:0] p;
  wire   [5:0] pl;
  wire   [29:0] FF1_out;
  wire   [11:0] Zh_f2;
  wire   [11:0] Zl_f2;
  wire   [5:0] gamma1;
  wire   [5:0] sA2N;
  wire   [5:0] ab;
  wire   [5:0] gamma0;
  wire   [23:0] FF2_out;
  wire   [11:0] Zh_f3;
  wire   [11:0] Zl_f3;
  wire   [11:0] muld;
  wire   [35:0] FF3_out;
  wire   [5:0] ph_H;
  wire   [5:0] p_H;
  wire   [5:0] pl_H;
  wire   [5:0] ph_L;
  wire   [5:0] p_L;
  wire   [5:0] pl_L;
  wire   [35:0] FF4_out;
  wire   [11:1] Inst_f1_sZ;
  wire   [5:0] Inst_f1_phpplmul_Orig_pl;
  wire   [5:0] Inst_f1_phpplmul_Orig_p;
  wire   [5:0] Inst_f1_phpplmul_Orig_ph;
  wire   [5:0] Inst_f1_phpplmul_sB;
  wire   [5:0] Inst_f1_phpplmul_sA;
  wire   [1:0] Inst_f1_phpplmul_AddNewMaskph_MaskXOR;
  wire   [1:0] Inst_f1_phpplmul_AddNewMaskp_MaskXOR;
  wire   [1:0] Inst_f1_phpplmul_AddNewMaskpl_MaskXOR;
  wire   [11:0] Inst_f2_abin;
  wire   [5:0] Inst_f2_dinv_1_Orig_sA2N;
  wire   [5:1] Inst_f2_dinv_1_sA2;
  wire   [5:0] Inst_f2_dinv_1_Orig_ab;
  wire   [1:0] Inst_f2_dinv_1_AddNewMaskab_MaskXOR;
  wire   [1:0] Inst_f2_dinv_1_AddNewMasksA2N_MaskXOR;
  wire   [5:0] Inst_f3_dinv_2_ph;
  wire   [5:0] Inst_f3_dinv_2_pl;
  wire   [3:0] Inst_f3_dinv_2_AddNewMaskQ_MaskXOR;
  wire   [5:0] Inst_f4_multd_L_Orig_pl;
  wire   [5:0] Inst_f4_multd_L_Orig_p;
  wire   [5:0] Inst_f4_multd_L_Orig_ph;
  wire   [5:0] Inst_f4_multd_L_sB;
  wire   [5:0] Inst_f4_multd_L_sA;
  wire   [1:0] Inst_f4_multd_L_AddNewMaskph_MaskXOR;
  wire   [1:0] Inst_f4_multd_L_AddNewMaskp_MaskXOR;
  wire   [1:0] Inst_f4_multd_L_AddNewMaskpl_MaskXOR;
  wire   [5:0] Inst_f4_multd_H_Orig_pl;
  wire   [5:0] Inst_f4_multd_H_Orig_p;
  wire   [5:0] Inst_f4_multd_H_Orig_ph;
  wire   [5:0] Inst_f4_multd_H_sB;
  wire   [5:0] Inst_f4_multd_H_sA;
  wire   [1:0] Inst_f4_multd_H_AddNewMaskph_MaskXOR;
  wire   [1:0] Inst_f4_multd_H_AddNewMaskp_MaskXOR;
  wire   [1:0] Inst_f4_multd_H_AddNewMaskpl_MaskXOR;
  wire   [11:0] Inst_f5_pl;
  wire   [11:0] Inst_f5_ph;

  XOR2_X1 Inst_f1_U12 ( .A(Zh_f1[9]), .B(Zl_f1_9_), .Z(Inst_f1_sZ[9]) );
  XOR2_X1 Inst_f1_U11 ( .A(Zh_f1[8]), .B(Zl_f1_8_), .Z(ab2[8]) );
  XOR2_X1 Inst_f1_U10 ( .A(Zh_f1[7]), .B(Zl_f1_7_), .Z(Inst_f1_sZ[7]) );
  XOR2_X1 Inst_f1_U9 ( .A(Zh_f1[6]), .B(A[8]), .Z(Inst_f1_sZ[6]) );
  XOR2_X1 Inst_f1_U8 ( .A(Zh_f1[5]), .B(Zl_f1_5_), .Z(Inst_f1_sZ[5]) );
  XOR2_X1 Inst_f1_U7 ( .A(Zh_f1[4]), .B(Zl_f1_4_), .Z(ab2[4]) );
  XOR2_X1 Inst_f1_U6 ( .A(Zh_f1[3]), .B(Zl_f1_3_), .Z(Inst_f1_sZ[3]) );
  XOR2_X1 Inst_f1_U5 ( .A(Zh_f1[2]), .B(A[0]), .Z(Inst_f1_sZ[2]) );
  XOR2_X1 Inst_f1_U4 ( .A(Zh_f1[1]), .B(Zl_f1_1_), .Z(Inst_f1_sZ[1]) );
  XOR2_X1 Inst_f1_U3 ( .A(Zh_f1[11]), .B(Zl_f1_11_), .Z(Inst_f1_sZ[11]) );
  XOR2_X1 Inst_f1_U2 ( .A(Zh_f1[10]), .B(A[16]), .Z(Inst_f1_sZ[10]) );
  XOR2_X1 Inst_f1_U1 ( .A(Zh_f1[0]), .B(Zl_f1_0_), .Z(ab2[0]) );
  XNOR2_X1 Inst_f1_linearMapping_U42 ( .A(Inst_f1_linearMapping_n32), .B(
        Inst_f1_linearMapping_n31), .ZN(Zh_f1[11]) );
  XNOR2_X1 Inst_f1_linearMapping_U41 ( .A(Inst_f1_linearMapping_n30), .B(
        Inst_f1_linearMapping_n29), .ZN(Inst_f1_linearMapping_n31) );
  XNOR2_X1 Inst_f1_linearMapping_U40 ( .A(A[17]), .B(A[18]), .ZN(
        Inst_f1_linearMapping_n30) );
  XNOR2_X1 Inst_f1_linearMapping_U39 ( .A(Inst_f1_linearMapping_n28), .B(
        Inst_f1_linearMapping_n27), .ZN(Zh_f1[7]) );
  XNOR2_X1 Inst_f1_linearMapping_U38 ( .A(A[11]), .B(Inst_f1_linearMapping_n27), .ZN(Zl_f1_4_) );
  XNOR2_X1 Inst_f1_linearMapping_U37 ( .A(Inst_f1_linearMapping_n26), .B(
        Inst_f1_linearMapping_n25), .ZN(Inst_f1_linearMapping_n27) );
  XNOR2_X1 Inst_f1_linearMapping_U36 ( .A(A[9]), .B(A[10]), .ZN(
        Inst_f1_linearMapping_n26) );
  XNOR2_X1 Inst_f1_linearMapping_U35 ( .A(Inst_f1_linearMapping_n22), .B(
        Inst_f1_linearMapping_n21), .ZN(Inst_f1_linearMapping_n23) );
  XNOR2_X1 Inst_f1_linearMapping_U34 ( .A(A[1]), .B(A[2]), .ZN(
        Inst_f1_linearMapping_n22) );
  XOR2_X1 Inst_f1_linearMapping_U33 ( .A(A[1]), .B(Inst_f1_linearMapping_n20), 
        .Z(Zl_f1_3_) );
  XNOR2_X1 Inst_f1_linearMapping_U32 ( .A(Inst_f1_linearMapping_n19), .B(
        Inst_f1_linearMapping_n18), .ZN(Inst_f1_linearMapping_n20) );
  XNOR2_X1 Inst_f1_linearMapping_U31 ( .A(A[3]), .B(A[4]), .ZN(
        Inst_f1_linearMapping_n18) );
  XOR2_X1 Inst_f1_linearMapping_U30 ( .A(A[0]), .B(A[7]), .Z(
        Inst_f1_linearMapping_n19) );
  XNOR2_X1 Inst_f1_linearMapping_U29 ( .A(A[19]), .B(A[20]), .ZN(
        Inst_f1_linearMapping_n16) );
  XOR2_X1 Inst_f1_linearMapping_U28 ( .A(A[16]), .B(A[23]), .Z(
        Inst_f1_linearMapping_n17) );
  XOR2_X1 Inst_f1_linearMapping_U27 ( .A(A[9]), .B(Zl_f1_5_), .Z(Zh_f1[5]) );
  XOR2_X1 Inst_f1_linearMapping_U26 ( .A(A[9]), .B(Inst_f1_linearMapping_n15), 
        .Z(Zl_f1_7_) );
  XNOR2_X1 Inst_f1_linearMapping_U25 ( .A(Inst_f1_linearMapping_n14), .B(
        Inst_f1_linearMapping_n13), .ZN(Inst_f1_linearMapping_n15) );
  XNOR2_X1 Inst_f1_linearMapping_U24 ( .A(A[11]), .B(A[12]), .ZN(
        Inst_f1_linearMapping_n13) );
  XOR2_X1 Inst_f1_linearMapping_U23 ( .A(A[8]), .B(A[15]), .Z(
        Inst_f1_linearMapping_n14) );
  XOR2_X1 Inst_f1_linearMapping_U22 ( .A(A[15]), .B(A[13]), .Z(
        Inst_f1_linearMapping_n28) );
  XNOR2_X1 Inst_f1_linearMapping_U21 ( .A(A[8]), .B(A[14]), .ZN(
        Inst_f1_linearMapping_n25) );
  XOR2_X1 Inst_f1_linearMapping_U20 ( .A(A[23]), .B(A[21]), .Z(
        Inst_f1_linearMapping_n32) );
  XOR2_X1 Inst_f1_linearMapping_U19 ( .A(A[7]), .B(A[5]), .Z(
        Inst_f1_linearMapping_n24) );
  XNOR2_X1 Inst_f1_linearMapping_U18 ( .A(A[0]), .B(A[6]), .ZN(
        Inst_f1_linearMapping_n21) );
  XNOR2_X1 Inst_f1_linearMapping_U17 ( .A(A[16]), .B(A[22]), .ZN(
        Inst_f1_linearMapping_n29) );
  XNOR2_X2 Inst_f1_linearMapping_U16 ( .A(A[21]), .B(Inst_f1_linearMapping_n29), .ZN(Zl_f1_9_) );
  XOR2_X2 Inst_f1_linearMapping_U15 ( .A(A[17]), .B(Zl_f1_9_), .Z(Zh_f1[9]) );
  XOR2_X2 Inst_f1_linearMapping_U14 ( .A(A[20]), .B(Zl_f1_9_), .Z(Zh_f1[10])
         );
  XNOR2_X2 Inst_f1_linearMapping_U13 ( .A(A[5]), .B(Inst_f1_linearMapping_n21), 
        .ZN(Zl_f1_1_) );
  XOR2_X2 Inst_f1_linearMapping_U12 ( .A(A[1]), .B(Zl_f1_1_), .Z(Zh_f1[1]) );
  XOR2_X2 Inst_f1_linearMapping_U11 ( .A(A[4]), .B(Zl_f1_1_), .Z(Zh_f1[2]) );
  XNOR2_X2 Inst_f1_linearMapping_U10 ( .A(A[13]), .B(Inst_f1_linearMapping_n25), .ZN(Zl_f1_5_) );
  XOR2_X2 Inst_f1_linearMapping_U9 ( .A(A[12]), .B(Zl_f1_5_), .Z(Zh_f1[6]) );
  XNOR2_X2 Inst_f1_linearMapping_U8 ( .A(A[3]), .B(Inst_f1_linearMapping_n23), 
        .ZN(Zl_f1_0_) );
  XNOR2_X2 Inst_f1_linearMapping_U7 ( .A(Inst_f1_linearMapping_n32), .B(
        Inst_f1_linearMapping_n29), .ZN(Zh_f1[8]) );
  XNOR2_X2 Inst_f1_linearMapping_U6 ( .A(Inst_f1_linearMapping_n24), .B(
        Inst_f1_linearMapping_n21), .ZN(Zh_f1[0]) );
  XNOR2_X2 Inst_f1_linearMapping_U5 ( .A(Inst_f1_linearMapping_n28), .B(
        Inst_f1_linearMapping_n25), .ZN(Zh_f1[4]) );
  XNOR2_X2 Inst_f1_linearMapping_U4 ( .A(A[19]), .B(Inst_f1_linearMapping_n31), 
        .ZN(Zl_f1_8_) );
  XNOR2_X2 Inst_f1_linearMapping_U3 ( .A(Inst_f1_linearMapping_n24), .B(
        Inst_f1_linearMapping_n23), .ZN(Zh_f1[3]) );
  XOR2_X1 Inst_f1_linearMapping_U2 ( .A(Inst_f1_linearMapping_n17), .B(
        Inst_f1_linearMapping_n16), .Z(Inst_f1_linearMapping_n12) );
  XNOR2_X2 Inst_f1_linearMapping_U1 ( .A(A[17]), .B(Inst_f1_linearMapping_n12), 
        .ZN(Zl_f1_11_) );
  XOR2_X1 Inst_f1_abSQ_U6 ( .A(Inst_f1_sZ[11]), .B(Inst_f1_sZ[9]), .Z(ab2[10])
         );
  XOR2_X1 Inst_f1_abSQ_U5 ( .A(Inst_f1_sZ[10]), .B(ab2[8]), .Z(ab2[11]) );
  XOR2_X1 Inst_f1_abSQ_U4 ( .A(Inst_f1_sZ[5]), .B(Inst_f1_sZ[7]), .Z(ab2[6])
         );
  XOR2_X1 Inst_f1_abSQ_U3 ( .A(ab2[4]), .B(Inst_f1_sZ[6]), .Z(ab2[7]) );
  XOR2_X1 Inst_f1_abSQ_U2 ( .A(Inst_f1_sZ[1]), .B(Inst_f1_sZ[3]), .Z(ab2[2])
         );
  XOR2_X1 Inst_f1_abSQ_U1 ( .A(ab2[0]), .B(Inst_f1_sZ[2]), .Z(ab2[3]) );
  XOR2_X1 Inst_f1_abSQ_NxGamma_U3 ( .A(ab2[8]), .B(Inst_f1_sZ[9]), .Z(ab2[9])
         );
  XOR2_X1 Inst_f1_abSQ_NxGamma_U2 ( .A(ab2[4]), .B(Inst_f1_sZ[5]), .Z(ab2[5])
         );
  XOR2_X1 Inst_f1_abSQ_NxGamma_U1 ( .A(ab2[0]), .B(Inst_f1_sZ[1]), .Z(ab2[1])
         );
  XOR2_X1 Inst_f1_phpplmul_U12 ( .A(Zl_f1_11_), .B(Zl_f1_9_), .Z(
        Inst_f1_phpplmul_sB[5]) );
  XOR2_X1 Inst_f1_phpplmul_U11 ( .A(A[16]), .B(Zl_f1_8_), .Z(
        Inst_f1_phpplmul_sB[4]) );
  XOR2_X1 Inst_f1_phpplmul_U10 ( .A(Zl_f1_5_), .B(Zl_f1_7_), .Z(
        Inst_f1_phpplmul_sB[3]) );
  XOR2_X1 Inst_f1_phpplmul_U9 ( .A(Zl_f1_4_), .B(A[8]), .Z(
        Inst_f1_phpplmul_sB[2]) );
  XOR2_X1 Inst_f1_phpplmul_U8 ( .A(Zl_f1_1_), .B(Zl_f1_3_), .Z(
        Inst_f1_phpplmul_sB[1]) );
  XOR2_X1 Inst_f1_phpplmul_U7 ( .A(Zl_f1_0_), .B(A[0]), .Z(
        Inst_f1_phpplmul_sB[0]) );
  XOR2_X1 Inst_f1_phpplmul_U6 ( .A(Zh_f1[11]), .B(Zh_f1[9]), .Z(
        Inst_f1_phpplmul_sA[5]) );
  XOR2_X1 Inst_f1_phpplmul_U5 ( .A(Zh_f1[10]), .B(Zh_f1[8]), .Z(
        Inst_f1_phpplmul_sA[4]) );
  XOR2_X1 Inst_f1_phpplmul_U4 ( .A(Zh_f1[5]), .B(Zh_f1[7]), .Z(
        Inst_f1_phpplmul_sA[3]) );
  XOR2_X1 Inst_f1_phpplmul_U3 ( .A(Zh_f1[4]), .B(Zh_f1[6]), .Z(
        Inst_f1_phpplmul_sA[2]) );
  XOR2_X1 Inst_f1_phpplmul_U2 ( .A(Zh_f1[1]), .B(Zh_f1[3]), .Z(
        Inst_f1_phpplmul_sA[1]) );
  XOR2_X1 Inst_f1_phpplmul_U1 ( .A(Zh_f1[0]), .B(Zh_f1[2]), .Z(
        Inst_f1_phpplmul_sA[0]) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U104 ( .A(Inst_f1_phpplmul_himul_n94), .B(
        Inst_f1_phpplmul_himul_n93), .ZN(Inst_f1_phpplmul_Orig_ph[4]) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U103 ( .A(Inst_f1_phpplmul_himul_n92), .B(
        Inst_f1_phpplmul_himul_n91), .ZN(Inst_f1_phpplmul_himul_n93) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U102 ( .A(Inst_f1_phpplmul_himul_n90), .B(
        Inst_f1_phpplmul_himul_n89), .ZN(Inst_f1_phpplmul_himul_n91) );
  NAND2_X1 Inst_f1_phpplmul_himul_U101 ( .A1(Inst_f1_phpplmul_himul_n88), .A2(
        Zh_f1[6]), .ZN(Inst_f1_phpplmul_himul_n90) );
  NAND2_X1 Inst_f1_phpplmul_himul_U100 ( .A1(Inst_f1_phpplmul_himul_n87), .A2(
        Inst_f1_phpplmul_himul_n86), .ZN(Inst_f1_phpplmul_himul_n92) );
  NAND2_X1 Inst_f1_phpplmul_himul_U99 ( .A1(A[0]), .A2(
        Inst_f1_phpplmul_himul_n85), .ZN(Inst_f1_phpplmul_himul_n86) );
  OR2_X1 Inst_f1_phpplmul_himul_U98 ( .A1(Inst_f1_phpplmul_himul_n85), .A2(
        Inst_f1_phpplmul_himul_n95), .ZN(Inst_f1_phpplmul_himul_n87) );
  XOR2_X1 Inst_f1_phpplmul_himul_U97 ( .A(Zh_f1[3]), .B(
        Inst_f1_phpplmul_himul_n84), .Z(Inst_f1_phpplmul_himul_n85) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U96 ( .A(Inst_f1_phpplmul_himul_n83), .B(
        Inst_f1_phpplmul_himul_n97), .ZN(Inst_f1_phpplmul_himul_n94) );
  XOR2_X1 Inst_f1_phpplmul_himul_U95 ( .A(Inst_f1_phpplmul_himul_n82), .B(
        Inst_f1_phpplmul_himul_n81), .Z(Inst_f1_phpplmul_himul_n97) );
  NAND2_X1 Inst_f1_phpplmul_himul_U94 ( .A1(A[8]), .A2(Zh_f1[3]), .ZN(
        Inst_f1_phpplmul_himul_n81) );
  NOR2_X1 Inst_f1_phpplmul_himul_U93 ( .A1(Inst_f1_phpplmul_himul_n80), .A2(
        Inst_f1_phpplmul_himul_n95), .ZN(Inst_f1_phpplmul_himul_n82) );
  INV_X1 Inst_f1_phpplmul_himul_U92 ( .A(Zl_f1_3_), .ZN(
        Inst_f1_phpplmul_himul_n95) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U91 ( .A(Zh_f1[2]), .B(Zh_f1[6]), .ZN(
        Inst_f1_phpplmul_himul_n80) );
  NAND2_X1 Inst_f1_phpplmul_himul_U90 ( .A1(Inst_f1_phpplmul_himul_n79), .A2(
        Inst_f1_phpplmul_himul_n78), .ZN(Inst_f1_phpplmul_himul_n83) );
  NAND2_X1 Inst_f1_phpplmul_himul_U89 ( .A1(Zh_f1[3]), .A2(
        Inst_f1_phpplmul_himul_n77), .ZN(Inst_f1_phpplmul_himul_n78) );
  NAND2_X1 Inst_f1_phpplmul_himul_U88 ( .A1(Zh_f1[2]), .A2(Zl_f1_7_), .ZN(
        Inst_f1_phpplmul_himul_n79) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U87 ( .A(Inst_f1_phpplmul_himul_n76), .B(
        Inst_f1_phpplmul_himul_n75), .ZN(Inst_f1_phpplmul_Orig_ph[3]) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U86 ( .A(Inst_f1_phpplmul_himul_n74), .B(
        Inst_f1_phpplmul_himul_n73), .ZN(Inst_f1_phpplmul_himul_n75) );
  XOR2_X1 Inst_f1_phpplmul_himul_U85 ( .A(Inst_f1_phpplmul_himul_n72), .B(
        Inst_f1_phpplmul_himul_n71), .Z(Inst_f1_phpplmul_himul_n74) );
  NAND2_X1 Inst_f1_phpplmul_himul_U84 ( .A1(Zh_f1[10]), .A2(A[16]), .ZN(
        Inst_f1_phpplmul_himul_n71) );
  NAND2_X1 Inst_f1_phpplmul_himul_U83 ( .A1(Zh_f1[11]), .A2(Zl_f1_11_), .ZN(
        Inst_f1_phpplmul_himul_n72) );
  XOR2_X1 Inst_f1_phpplmul_himul_U82 ( .A(Inst_f1_phpplmul_himul_n70), .B(
        Inst_f1_phpplmul_himul_n69), .Z(Inst_f1_phpplmul_himul_n76) );
  XOR2_X1 Inst_f1_phpplmul_himul_U81 ( .A(Inst_f1_phpplmul_himul_n68), .B(
        Inst_f1_phpplmul_himul_n67), .Z(Inst_f1_phpplmul_himul_n69) );
  NAND2_X1 Inst_f1_phpplmul_himul_U80 ( .A1(Zh_f1[10]), .A2(
        Inst_f1_phpplmul_himul_n66), .ZN(Inst_f1_phpplmul_himul_n67) );
  NAND2_X1 Inst_f1_phpplmul_himul_U79 ( .A1(Zh_f1[2]), .A2(Zl_f1_11_), .ZN(
        Inst_f1_phpplmul_himul_n68) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U78 ( .A(Inst_f1_phpplmul_himul_n65), .B(
        Inst_f1_phpplmul_himul_n64), .ZN(Inst_f1_phpplmul_himul_n70) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U77 ( .A(Zh_f1[11]), .B(
        Inst_f1_phpplmul_himul_n63), .ZN(Inst_f1_phpplmul_himul_n64) );
  XOR2_X1 Inst_f1_phpplmul_himul_U76 ( .A(Inst_f1_phpplmul_himul_n62), .B(
        Inst_f1_phpplmul_himul_n61), .Z(Inst_f1_phpplmul_himul_n63) );
  NAND2_X1 Inst_f1_phpplmul_himul_U75 ( .A1(A[0]), .A2(Zh_f1[10]), .ZN(
        Inst_f1_phpplmul_himul_n61) );
  NOR2_X1 Inst_f1_phpplmul_himul_U74 ( .A1(Inst_f1_phpplmul_himul_n60), .A2(
        Zl_f1_3_), .ZN(Inst_f1_phpplmul_himul_n62) );
  NAND2_X1 Inst_f1_phpplmul_himul_U73 ( .A1(Inst_f1_phpplmul_himul_n59), .A2(
        A[16]), .ZN(Inst_f1_phpplmul_himul_n65) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U72 ( .A(Inst_f1_phpplmul_himul_n96), .B(
        Inst_f1_phpplmul_himul_n58), .ZN(Inst_f1_phpplmul_himul_n59) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U71 ( .A(Zh_f1[3]), .B(
        Inst_f1_phpplmul_himul_n57), .ZN(Inst_f1_phpplmul_himul_n58) );
  INV_X1 Inst_f1_phpplmul_himul_U70 ( .A(Zh_f1[2]), .ZN(
        Inst_f1_phpplmul_himul_n96) );
  XOR2_X1 Inst_f1_phpplmul_himul_U69 ( .A(Inst_f1_phpplmul_himul_n56), .B(
        Inst_f1_phpplmul_himul_n55), .Z(Inst_f1_phpplmul_Orig_ph[2]) );
  NAND2_X1 Inst_f1_phpplmul_himul_U68 ( .A1(Inst_f1_phpplmul_himul_n54), .A2(
        Inst_f1_phpplmul_himul_n53), .ZN(Inst_f1_phpplmul_himul_n55) );
  OR2_X1 Inst_f1_phpplmul_himul_U67 ( .A1(Zl_f1_11_), .A2(
        Inst_f1_phpplmul_himul_n60), .ZN(Inst_f1_phpplmul_himul_n53) );
  NAND2_X1 Inst_f1_phpplmul_himul_U66 ( .A1(Inst_f1_phpplmul_himul_n52), .A2(
        Zl_f1_11_), .ZN(Inst_f1_phpplmul_himul_n54) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U65 ( .A(Inst_f1_phpplmul_himul_n51), .B(
        Zh_f1[2]), .ZN(Inst_f1_phpplmul_himul_n52) );
  XOR2_X1 Inst_f1_phpplmul_himul_U64 ( .A(Inst_f1_phpplmul_himul_n50), .B(
        Inst_f1_phpplmul_himul_n49), .Z(Inst_f1_phpplmul_himul_n56) );
  NOR2_X1 Inst_f1_phpplmul_himul_U63 ( .A1(Inst_f1_phpplmul_himul_n57), .A2(
        Inst_f1_phpplmul_himul_n48), .ZN(Inst_f1_phpplmul_himul_n49) );
  XOR2_X1 Inst_f1_phpplmul_himul_U62 ( .A(Inst_f1_phpplmul_himul_n66), .B(
        Zl_f1_3_), .Z(Inst_f1_phpplmul_himul_n48) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U61 ( .A(Inst_f1_phpplmul_himul_n47), .B(
        Inst_f1_phpplmul_himul_n46), .ZN(Inst_f1_phpplmul_himul_n50) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U60 ( .A(A[0]), .B(
        Inst_f1_phpplmul_himul_n89), .ZN(Inst_f1_phpplmul_himul_n46) );
  XOR2_X1 Inst_f1_phpplmul_himul_U59 ( .A(Inst_f1_phpplmul_himul_n45), .B(
        Inst_f1_phpplmul_himul_n44), .Z(Inst_f1_phpplmul_himul_n89) );
  NAND2_X1 Inst_f1_phpplmul_himul_U58 ( .A1(Zh_f1[3]), .A2(A[0]), .ZN(
        Inst_f1_phpplmul_himul_n44) );
  NAND2_X1 Inst_f1_phpplmul_himul_U57 ( .A1(Zh_f1[2]), .A2(Zl_f1_3_), .ZN(
        Inst_f1_phpplmul_himul_n45) );
  XOR2_X1 Inst_f1_phpplmul_himul_U56 ( .A(Inst_f1_phpplmul_himul_n43), .B(
        Inst_f1_phpplmul_himul_n73), .Z(Inst_f1_phpplmul_himul_n47) );
  XOR2_X1 Inst_f1_phpplmul_himul_U55 ( .A(Inst_f1_phpplmul_himul_n42), .B(
        Inst_f1_phpplmul_himul_n41), .Z(Inst_f1_phpplmul_himul_n73) );
  NAND2_X1 Inst_f1_phpplmul_himul_U54 ( .A1(Zh_f1[10]), .A2(Zl_f1_3_), .ZN(
        Inst_f1_phpplmul_himul_n41) );
  NAND2_X1 Inst_f1_phpplmul_himul_U53 ( .A1(Zh_f1[11]), .A2(A[0]), .ZN(
        Inst_f1_phpplmul_himul_n42) );
  XOR2_X1 Inst_f1_phpplmul_himul_U52 ( .A(Inst_f1_phpplmul_himul_n40), .B(
        Inst_f1_phpplmul_himul_n39), .Z(Inst_f1_phpplmul_himul_n43) );
  NAND2_X1 Inst_f1_phpplmul_himul_U51 ( .A1(A[16]), .A2(
        Inst_f1_phpplmul_himul_n60), .ZN(Inst_f1_phpplmul_himul_n39) );
  INV_X1 Inst_f1_phpplmul_himul_U50 ( .A(Zh_f1[3]), .ZN(
        Inst_f1_phpplmul_himul_n60) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U49 ( .A(Inst_f1_phpplmul_himul_n38), .B(
        Inst_f1_phpplmul_himul_n37), .ZN(Inst_f1_phpplmul_Orig_ph[1]) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U48 ( .A(Inst_f1_phpplmul_himul_n36), .B(
        Inst_f1_phpplmul_himul_n35), .ZN(Inst_f1_phpplmul_himul_n38) );
  NAND2_X1 Inst_f1_phpplmul_himul_U47 ( .A1(Inst_f1_phpplmul_himul_n34), .A2(
        Zh_f1[6]), .ZN(Inst_f1_phpplmul_himul_n35) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U46 ( .A(A[8]), .B(
        Inst_f1_phpplmul_himul_n66), .ZN(Inst_f1_phpplmul_himul_n34) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U45 ( .A(Inst_f1_phpplmul_himul_n33), .B(
        Inst_f1_phpplmul_himul_n32), .ZN(Inst_f1_phpplmul_himul_n36) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U44 ( .A(Inst_f1_phpplmul_himul_n31), .B(
        Inst_f1_phpplmul_himul_n30), .ZN(Inst_f1_phpplmul_himul_n32) );
  NAND2_X1 Inst_f1_phpplmul_himul_U43 ( .A1(Inst_f1_phpplmul_himul_n29), .A2(
        Inst_f1_phpplmul_himul_n88), .ZN(Inst_f1_phpplmul_himul_n30) );
  XOR2_X1 Inst_f1_phpplmul_himul_U42 ( .A(A[8]), .B(Zl_f1_7_), .Z(
        Inst_f1_phpplmul_himul_n88) );
  XOR2_X1 Inst_f1_phpplmul_himul_U41 ( .A(Zh_f1[6]), .B(Zh_f1[10]), .Z(
        Inst_f1_phpplmul_himul_n29) );
  NAND2_X1 Inst_f1_phpplmul_himul_U40 ( .A1(Zh_f1[7]), .A2(A[16]), .ZN(
        Inst_f1_phpplmul_himul_n31) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U39 ( .A(Inst_f1_phpplmul_himul_n28), .B(
        Inst_f1_phpplmul_himul_n27), .ZN(Inst_f1_phpplmul_himul_n33) );
  XOR2_X1 Inst_f1_phpplmul_himul_U38 ( .A(Inst_f1_phpplmul_himul_n26), .B(
        Inst_f1_phpplmul_himul_n25), .Z(Inst_f1_phpplmul_himul_n28) );
  NOR2_X1 Inst_f1_phpplmul_himul_U37 ( .A1(Inst_f1_phpplmul_himul_n51), .A2(
        A[16]), .ZN(Inst_f1_phpplmul_himul_n25) );
  INV_X1 Inst_f1_phpplmul_himul_U36 ( .A(Zh_f1[10]), .ZN(
        Inst_f1_phpplmul_himul_n51) );
  NOR2_X1 Inst_f1_phpplmul_himul_U35 ( .A1(Inst_f1_phpplmul_himul_n57), .A2(
        Zl_f1_11_), .ZN(Inst_f1_phpplmul_himul_n26) );
  INV_X1 Inst_f1_phpplmul_himul_U34 ( .A(Zh_f1[11]), .ZN(
        Inst_f1_phpplmul_himul_n57) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U33 ( .A(Inst_f1_phpplmul_himul_n24), .B(
        Inst_f1_phpplmul_himul_n23), .ZN(Inst_f1_phpplmul_Orig_ph[0]) );
  NAND2_X1 Inst_f1_phpplmul_himul_U32 ( .A1(Zh_f1[6]), .A2(Zl_f1_11_), .ZN(
        Inst_f1_phpplmul_himul_n23) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U31 ( .A(Inst_f1_phpplmul_himul_n98), .B(
        Inst_f1_phpplmul_himul_n22), .ZN(Inst_f1_phpplmul_himul_n24) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U30 ( .A(Inst_f1_phpplmul_himul_n21), .B(
        Inst_f1_phpplmul_himul_n20), .ZN(Inst_f1_phpplmul_himul_n22) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U29 ( .A(Inst_f1_phpplmul_himul_n19), .B(
        Inst_f1_phpplmul_himul_n18), .ZN(Inst_f1_phpplmul_himul_n20) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U28 ( .A(Inst_f1_phpplmul_himul_n17), .B(
        Inst_f1_phpplmul_himul_n37), .ZN(Inst_f1_phpplmul_himul_n18) );
  NAND2_X1 Inst_f1_phpplmul_himul_U27 ( .A1(A[8]), .A2(
        Inst_f1_phpplmul_himul_n16), .ZN(Inst_f1_phpplmul_himul_n37) );
  XOR2_X1 Inst_f1_phpplmul_himul_U26 ( .A(Zh_f1[7]), .B(Zh_f1[11]), .Z(
        Inst_f1_phpplmul_himul_n16) );
  NOR2_X1 Inst_f1_phpplmul_himul_U25 ( .A1(Inst_f1_phpplmul_himul_n15), .A2(
        Inst_f1_phpplmul_himul_n77), .ZN(Inst_f1_phpplmul_himul_n17) );
  INV_X1 Inst_f1_phpplmul_himul_U24 ( .A(Zl_f1_7_), .ZN(
        Inst_f1_phpplmul_himul_n77) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U23 ( .A(Zh_f1[11]), .B(Zh_f1[10]), .ZN(
        Inst_f1_phpplmul_himul_n15) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U22 ( .A(Inst_f1_phpplmul_himul_n40), .B(
        A[16]), .ZN(Inst_f1_phpplmul_himul_n19) );
  NAND2_X1 Inst_f1_phpplmul_himul_U21 ( .A1(Zh_f1[10]), .A2(Zl_f1_11_), .ZN(
        Inst_f1_phpplmul_himul_n40) );
  NOR2_X1 Inst_f1_phpplmul_himul_U20 ( .A1(Inst_f1_phpplmul_himul_n84), .A2(
        Inst_f1_phpplmul_himul_n66), .ZN(Inst_f1_phpplmul_himul_n21) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U19 ( .A(A[16]), .B(Zl_f1_11_), .ZN(
        Inst_f1_phpplmul_himul_n66) );
  INV_X1 Inst_f1_phpplmul_himul_U18 ( .A(Zh_f1[7]), .ZN(
        Inst_f1_phpplmul_himul_n84) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U17 ( .A(Inst_f1_phpplmul_himul_n27), .B(
        Inst_f1_phpplmul_himul_n14), .ZN(Inst_f1_phpplmul_himul_n98) );
  NAND2_X1 Inst_f1_phpplmul_himul_U16 ( .A1(Zh_f1[6]), .A2(A[8]), .ZN(
        Inst_f1_phpplmul_himul_n14) );
  NAND2_X1 Inst_f1_phpplmul_himul_U15 ( .A1(Zl_f1_7_), .A2(Zh_f1[7]), .ZN(
        Inst_f1_phpplmul_himul_n27) );
  XOR2_X1 Inst_f1_phpplmul_himul_U14 ( .A(Inst_f1_phpplmul_himul_n98), .B(
        Inst_f1_phpplmul_himul_n13), .Z(Inst_f1_phpplmul_Orig_ph[5]) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U13 ( .A(Inst_f1_phpplmul_himul_n12), .B(
        Inst_f1_phpplmul_himul_n10), .ZN(Inst_f1_phpplmul_himul_n13) );
  NAND2_X1 Inst_f1_phpplmul_himul_U12 ( .A1(Inst_f1_phpplmul_himul_n11), .A2(
        Inst_f1_phpplmul_himul_n7), .ZN(Inst_f1_phpplmul_himul_n12) );
  NAND2_X1 Inst_f1_phpplmul_himul_U11 ( .A1(Inst_f1_phpplmul_himul_n1), .A2(
        Zl_f1_3_), .ZN(Inst_f1_phpplmul_himul_n11) );
  XOR2_X1 Inst_f1_phpplmul_himul_U10 ( .A(Inst_f1_phpplmul_himul_n97), .B(
        Inst_f1_phpplmul_himul_n9), .Z(Inst_f1_phpplmul_himul_n10) );
  NOR2_X1 Inst_f1_phpplmul_himul_U9 ( .A1(Inst_f1_phpplmul_himul_n96), .A2(
        Inst_f1_phpplmul_himul_n8), .ZN(Inst_f1_phpplmul_himul_n9) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U8 ( .A(A[8]), .B(Zl_f1_7_), .ZN(
        Inst_f1_phpplmul_himul_n8) );
  XOR2_X1 Inst_f1_phpplmul_himul_U7 ( .A(Inst_f1_phpplmul_himul_n4), .B(
        Inst_f1_phpplmul_himul_n6), .Z(Inst_f1_phpplmul_himul_n7) );
  NAND2_X1 Inst_f1_phpplmul_himul_U6 ( .A1(Inst_f1_phpplmul_himul_n5), .A2(
        Zh_f1[3]), .ZN(Inst_f1_phpplmul_himul_n6) );
  NAND2_X1 Inst_f1_phpplmul_himul_U5 ( .A1(A[0]), .A2(
        Inst_f1_phpplmul_himul_n95), .ZN(Inst_f1_phpplmul_himul_n5) );
  NAND2_X1 Inst_f1_phpplmul_himul_U4 ( .A1(A[0]), .A2(
        Inst_f1_phpplmul_himul_n3), .ZN(Inst_f1_phpplmul_himul_n4) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U3 ( .A(Inst_f1_phpplmul_himul_n2), .B(
        Zh_f1[7]), .ZN(Inst_f1_phpplmul_himul_n3) );
  XNOR2_X1 Inst_f1_phpplmul_himul_U2 ( .A(Zh_f1[2]), .B(Zh_f1[6]), .ZN(
        Inst_f1_phpplmul_himul_n2) );
  INV_X1 Inst_f1_phpplmul_himul_U1 ( .A(A[0]), .ZN(Inst_f1_phpplmul_himul_n1)
         );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_MaskXORInst_U2 ( .A(PRNGQ[0]), .B(
        PRNGQ[2]), .Z(Inst_f1_phpplmul_AddNewMaskph_MaskXOR[0]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_MaskXORInst_U1 ( .A(PRNGQ[1]), .B(
        PRNGQ[3]), .Z(Inst_f1_phpplmul_AddNewMaskph_MaskXOR[1]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_XORInst1_U2 ( .A(
        Inst_f1_phpplmul_Orig_ph[4]), .B(
        Inst_f1_phpplmul_AddNewMaskph_MaskXOR[0]), .Z(ph[4]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_XORInst1_U1 ( .A(
        Inst_f1_phpplmul_Orig_ph[5]), .B(
        Inst_f1_phpplmul_AddNewMaskph_MaskXOR[1]), .Z(ph[5]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_XORInst2_U4 ( .A(
        Inst_f1_phpplmul_Orig_ph[3]), .B(PRNGQ[3]), .Z(ph[3]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_XORInst2_U3 ( .A(
        Inst_f1_phpplmul_Orig_ph[2]), .B(PRNGQ[2]), .Z(ph[2]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_XORInst2_U2 ( .A(
        Inst_f1_phpplmul_Orig_ph[1]), .B(PRNGQ[1]), .Z(ph[1]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskph_XORInst2_U1 ( .A(
        Inst_f1_phpplmul_Orig_ph[0]), .B(PRNGQ[0]), .Z(ph[0]) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U104 ( .A(Inst_f1_phpplmul_summul_n336), 
        .B(Inst_f1_phpplmul_summul_n335), .ZN(Inst_f1_phpplmul_Orig_p[4]) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U103 ( .A(Inst_f1_phpplmul_summul_n334), 
        .B(Inst_f1_phpplmul_summul_n333), .ZN(Inst_f1_phpplmul_summul_n335) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U102 ( .A(Inst_f1_phpplmul_summul_n332), 
        .B(Inst_f1_phpplmul_summul_n331), .ZN(Inst_f1_phpplmul_summul_n333) );
  NAND2_X1 Inst_f1_phpplmul_summul_U101 ( .A1(Inst_f1_phpplmul_summul_n330), 
        .A2(Inst_f1_phpplmul_sA[2]), .ZN(Inst_f1_phpplmul_summul_n332) );
  NAND2_X1 Inst_f1_phpplmul_summul_U100 ( .A1(Inst_f1_phpplmul_summul_n329), 
        .A2(Inst_f1_phpplmul_summul_n328), .ZN(Inst_f1_phpplmul_summul_n334)
         );
  NAND2_X1 Inst_f1_phpplmul_summul_U99 ( .A1(Inst_f1_phpplmul_sB[0]), .A2(
        Inst_f1_phpplmul_summul_n327), .ZN(Inst_f1_phpplmul_summul_n328) );
  OR2_X1 Inst_f1_phpplmul_summul_U98 ( .A1(Inst_f1_phpplmul_summul_n327), .A2(
        Inst_f1_phpplmul_summul_n337), .ZN(Inst_f1_phpplmul_summul_n329) );
  XOR2_X1 Inst_f1_phpplmul_summul_U97 ( .A(Inst_f1_phpplmul_sA[1]), .B(
        Inst_f1_phpplmul_summul_n326), .Z(Inst_f1_phpplmul_summul_n327) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U96 ( .A(Inst_f1_phpplmul_summul_n325), .B(
        Inst_f1_phpplmul_summul_n339), .ZN(Inst_f1_phpplmul_summul_n336) );
  XOR2_X1 Inst_f1_phpplmul_summul_U95 ( .A(Inst_f1_phpplmul_summul_n324), .B(
        Inst_f1_phpplmul_summul_n323), .Z(Inst_f1_phpplmul_summul_n339) );
  NAND2_X1 Inst_f1_phpplmul_summul_U94 ( .A1(Inst_f1_phpplmul_sB[2]), .A2(
        Inst_f1_phpplmul_sA[1]), .ZN(Inst_f1_phpplmul_summul_n323) );
  NOR2_X1 Inst_f1_phpplmul_summul_U93 ( .A1(Inst_f1_phpplmul_summul_n322), 
        .A2(Inst_f1_phpplmul_summul_n337), .ZN(Inst_f1_phpplmul_summul_n324)
         );
  INV_X1 Inst_f1_phpplmul_summul_U92 ( .A(Inst_f1_phpplmul_sB[1]), .ZN(
        Inst_f1_phpplmul_summul_n337) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U91 ( .A(Inst_f1_phpplmul_sA[0]), .B(
        Inst_f1_phpplmul_sA[2]), .ZN(Inst_f1_phpplmul_summul_n322) );
  NAND2_X1 Inst_f1_phpplmul_summul_U90 ( .A1(Inst_f1_phpplmul_summul_n321), 
        .A2(Inst_f1_phpplmul_summul_n320), .ZN(Inst_f1_phpplmul_summul_n325)
         );
  NAND2_X1 Inst_f1_phpplmul_summul_U89 ( .A1(Inst_f1_phpplmul_sA[1]), .A2(
        Inst_f1_phpplmul_summul_n319), .ZN(Inst_f1_phpplmul_summul_n320) );
  NAND2_X1 Inst_f1_phpplmul_summul_U88 ( .A1(Inst_f1_phpplmul_sA[0]), .A2(
        Inst_f1_phpplmul_sB[3]), .ZN(Inst_f1_phpplmul_summul_n321) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U87 ( .A(Inst_f1_phpplmul_summul_n318), .B(
        Inst_f1_phpplmul_summul_n317), .ZN(Inst_f1_phpplmul_Orig_p[3]) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U86 ( .A(Inst_f1_phpplmul_summul_n316), .B(
        Inst_f1_phpplmul_summul_n315), .ZN(Inst_f1_phpplmul_summul_n317) );
  XOR2_X1 Inst_f1_phpplmul_summul_U85 ( .A(Inst_f1_phpplmul_summul_n314), .B(
        Inst_f1_phpplmul_summul_n313), .Z(Inst_f1_phpplmul_summul_n316) );
  NAND2_X1 Inst_f1_phpplmul_summul_U84 ( .A1(Inst_f1_phpplmul_sA[4]), .A2(
        Inst_f1_phpplmul_sB[4]), .ZN(Inst_f1_phpplmul_summul_n313) );
  NAND2_X1 Inst_f1_phpplmul_summul_U83 ( .A1(Inst_f1_phpplmul_sA[5]), .A2(
        Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n314) );
  XOR2_X1 Inst_f1_phpplmul_summul_U82 ( .A(Inst_f1_phpplmul_summul_n312), .B(
        Inst_f1_phpplmul_summul_n311), .Z(Inst_f1_phpplmul_summul_n318) );
  XOR2_X1 Inst_f1_phpplmul_summul_U81 ( .A(Inst_f1_phpplmul_summul_n310), .B(
        Inst_f1_phpplmul_summul_n309), .Z(Inst_f1_phpplmul_summul_n311) );
  NAND2_X1 Inst_f1_phpplmul_summul_U80 ( .A1(Inst_f1_phpplmul_sA[4]), .A2(
        Inst_f1_phpplmul_summul_n308), .ZN(Inst_f1_phpplmul_summul_n309) );
  NAND2_X1 Inst_f1_phpplmul_summul_U79 ( .A1(Inst_f1_phpplmul_sA[0]), .A2(
        Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n310) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U78 ( .A(Inst_f1_phpplmul_summul_n307), .B(
        Inst_f1_phpplmul_summul_n306), .ZN(Inst_f1_phpplmul_summul_n312) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U77 ( .A(Inst_f1_phpplmul_sA[5]), .B(
        Inst_f1_phpplmul_summul_n305), .ZN(Inst_f1_phpplmul_summul_n306) );
  XOR2_X1 Inst_f1_phpplmul_summul_U76 ( .A(Inst_f1_phpplmul_summul_n304), .B(
        Inst_f1_phpplmul_summul_n303), .Z(Inst_f1_phpplmul_summul_n305) );
  NAND2_X1 Inst_f1_phpplmul_summul_U75 ( .A1(Inst_f1_phpplmul_sB[0]), .A2(
        Inst_f1_phpplmul_sA[4]), .ZN(Inst_f1_phpplmul_summul_n303) );
  NOR2_X1 Inst_f1_phpplmul_summul_U74 ( .A1(Inst_f1_phpplmul_summul_n302), 
        .A2(Inst_f1_phpplmul_sB[1]), .ZN(Inst_f1_phpplmul_summul_n304) );
  NAND2_X1 Inst_f1_phpplmul_summul_U73 ( .A1(Inst_f1_phpplmul_summul_n301), 
        .A2(Inst_f1_phpplmul_sB[4]), .ZN(Inst_f1_phpplmul_summul_n307) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U72 ( .A(Inst_f1_phpplmul_summul_n338), .B(
        Inst_f1_phpplmul_summul_n300), .ZN(Inst_f1_phpplmul_summul_n301) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U71 ( .A(Inst_f1_phpplmul_sA[1]), .B(
        Inst_f1_phpplmul_summul_n299), .ZN(Inst_f1_phpplmul_summul_n300) );
  INV_X1 Inst_f1_phpplmul_summul_U70 ( .A(Inst_f1_phpplmul_sA[0]), .ZN(
        Inst_f1_phpplmul_summul_n338) );
  XOR2_X1 Inst_f1_phpplmul_summul_U69 ( .A(Inst_f1_phpplmul_summul_n298), .B(
        Inst_f1_phpplmul_summul_n297), .Z(Inst_f1_phpplmul_Orig_p[2]) );
  NAND2_X1 Inst_f1_phpplmul_summul_U68 ( .A1(Inst_f1_phpplmul_summul_n296), 
        .A2(Inst_f1_phpplmul_summul_n295), .ZN(Inst_f1_phpplmul_summul_n297)
         );
  OR2_X1 Inst_f1_phpplmul_summul_U67 ( .A1(Inst_f1_phpplmul_sB[5]), .A2(
        Inst_f1_phpplmul_summul_n302), .ZN(Inst_f1_phpplmul_summul_n295) );
  NAND2_X1 Inst_f1_phpplmul_summul_U66 ( .A1(Inst_f1_phpplmul_summul_n294), 
        .A2(Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n296) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U65 ( .A(Inst_f1_phpplmul_summul_n293), .B(
        Inst_f1_phpplmul_sA[0]), .ZN(Inst_f1_phpplmul_summul_n294) );
  XOR2_X1 Inst_f1_phpplmul_summul_U64 ( .A(Inst_f1_phpplmul_summul_n292), .B(
        Inst_f1_phpplmul_summul_n291), .Z(Inst_f1_phpplmul_summul_n298) );
  NOR2_X1 Inst_f1_phpplmul_summul_U63 ( .A1(Inst_f1_phpplmul_summul_n299), 
        .A2(Inst_f1_phpplmul_summul_n290), .ZN(Inst_f1_phpplmul_summul_n291)
         );
  XOR2_X1 Inst_f1_phpplmul_summul_U62 ( .A(Inst_f1_phpplmul_summul_n308), .B(
        Inst_f1_phpplmul_sB[1]), .Z(Inst_f1_phpplmul_summul_n290) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U61 ( .A(Inst_f1_phpplmul_summul_n289), .B(
        Inst_f1_phpplmul_summul_n288), .ZN(Inst_f1_phpplmul_summul_n292) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U60 ( .A(Inst_f1_phpplmul_sB[0]), .B(
        Inst_f1_phpplmul_summul_n331), .ZN(Inst_f1_phpplmul_summul_n288) );
  XOR2_X1 Inst_f1_phpplmul_summul_U59 ( .A(Inst_f1_phpplmul_summul_n287), .B(
        Inst_f1_phpplmul_summul_n286), .Z(Inst_f1_phpplmul_summul_n331) );
  NAND2_X1 Inst_f1_phpplmul_summul_U58 ( .A1(Inst_f1_phpplmul_sA[1]), .A2(
        Inst_f1_phpplmul_sB[0]), .ZN(Inst_f1_phpplmul_summul_n286) );
  NAND2_X1 Inst_f1_phpplmul_summul_U57 ( .A1(Inst_f1_phpplmul_sA[0]), .A2(
        Inst_f1_phpplmul_sB[1]), .ZN(Inst_f1_phpplmul_summul_n287) );
  XOR2_X1 Inst_f1_phpplmul_summul_U56 ( .A(Inst_f1_phpplmul_summul_n285), .B(
        Inst_f1_phpplmul_summul_n315), .Z(Inst_f1_phpplmul_summul_n289) );
  XOR2_X1 Inst_f1_phpplmul_summul_U55 ( .A(Inst_f1_phpplmul_summul_n284), .B(
        Inst_f1_phpplmul_summul_n283), .Z(Inst_f1_phpplmul_summul_n315) );
  NAND2_X1 Inst_f1_phpplmul_summul_U54 ( .A1(Inst_f1_phpplmul_sA[4]), .A2(
        Inst_f1_phpplmul_sB[1]), .ZN(Inst_f1_phpplmul_summul_n283) );
  NAND2_X1 Inst_f1_phpplmul_summul_U53 ( .A1(Inst_f1_phpplmul_sA[5]), .A2(
        Inst_f1_phpplmul_sB[0]), .ZN(Inst_f1_phpplmul_summul_n284) );
  XOR2_X1 Inst_f1_phpplmul_summul_U52 ( .A(Inst_f1_phpplmul_summul_n282), .B(
        Inst_f1_phpplmul_summul_n281), .Z(Inst_f1_phpplmul_summul_n285) );
  NAND2_X1 Inst_f1_phpplmul_summul_U51 ( .A1(Inst_f1_phpplmul_sB[4]), .A2(
        Inst_f1_phpplmul_summul_n302), .ZN(Inst_f1_phpplmul_summul_n281) );
  INV_X1 Inst_f1_phpplmul_summul_U50 ( .A(Inst_f1_phpplmul_sA[1]), .ZN(
        Inst_f1_phpplmul_summul_n302) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U49 ( .A(Inst_f1_phpplmul_summul_n280), .B(
        Inst_f1_phpplmul_summul_n279), .ZN(Inst_f1_phpplmul_Orig_p[1]) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U48 ( .A(Inst_f1_phpplmul_summul_n278), .B(
        Inst_f1_phpplmul_summul_n277), .ZN(Inst_f1_phpplmul_summul_n280) );
  NAND2_X1 Inst_f1_phpplmul_summul_U47 ( .A1(Inst_f1_phpplmul_summul_n276), 
        .A2(Inst_f1_phpplmul_sA[2]), .ZN(Inst_f1_phpplmul_summul_n277) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U46 ( .A(Inst_f1_phpplmul_sB[2]), .B(
        Inst_f1_phpplmul_summul_n308), .ZN(Inst_f1_phpplmul_summul_n276) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U45 ( .A(Inst_f1_phpplmul_summul_n275), .B(
        Inst_f1_phpplmul_summul_n274), .ZN(Inst_f1_phpplmul_summul_n278) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U44 ( .A(Inst_f1_phpplmul_summul_n273), .B(
        Inst_f1_phpplmul_summul_n272), .ZN(Inst_f1_phpplmul_summul_n274) );
  NAND2_X1 Inst_f1_phpplmul_summul_U43 ( .A1(Inst_f1_phpplmul_summul_n271), 
        .A2(Inst_f1_phpplmul_summul_n330), .ZN(Inst_f1_phpplmul_summul_n272)
         );
  XOR2_X1 Inst_f1_phpplmul_summul_U42 ( .A(Inst_f1_phpplmul_sB[2]), .B(
        Inst_f1_phpplmul_sB[3]), .Z(Inst_f1_phpplmul_summul_n330) );
  XOR2_X1 Inst_f1_phpplmul_summul_U41 ( .A(Inst_f1_phpplmul_sA[2]), .B(
        Inst_f1_phpplmul_sA[4]), .Z(Inst_f1_phpplmul_summul_n271) );
  NAND2_X1 Inst_f1_phpplmul_summul_U40 ( .A1(Inst_f1_phpplmul_sA[3]), .A2(
        Inst_f1_phpplmul_sB[4]), .ZN(Inst_f1_phpplmul_summul_n273) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U39 ( .A(Inst_f1_phpplmul_summul_n270), .B(
        Inst_f1_phpplmul_summul_n269), .ZN(Inst_f1_phpplmul_summul_n275) );
  XOR2_X1 Inst_f1_phpplmul_summul_U38 ( .A(Inst_f1_phpplmul_summul_n268), .B(
        Inst_f1_phpplmul_summul_n267), .Z(Inst_f1_phpplmul_summul_n270) );
  NOR2_X1 Inst_f1_phpplmul_summul_U37 ( .A1(Inst_f1_phpplmul_summul_n293), 
        .A2(Inst_f1_phpplmul_sB[4]), .ZN(Inst_f1_phpplmul_summul_n267) );
  INV_X1 Inst_f1_phpplmul_summul_U36 ( .A(Inst_f1_phpplmul_sA[4]), .ZN(
        Inst_f1_phpplmul_summul_n293) );
  NOR2_X1 Inst_f1_phpplmul_summul_U35 ( .A1(Inst_f1_phpplmul_summul_n299), 
        .A2(Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n268) );
  INV_X1 Inst_f1_phpplmul_summul_U34 ( .A(Inst_f1_phpplmul_sA[5]), .ZN(
        Inst_f1_phpplmul_summul_n299) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U33 ( .A(Inst_f1_phpplmul_summul_n266), .B(
        Inst_f1_phpplmul_summul_n265), .ZN(Inst_f1_phpplmul_Orig_p[0]) );
  NAND2_X1 Inst_f1_phpplmul_summul_U32 ( .A1(Inst_f1_phpplmul_sA[2]), .A2(
        Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n265) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U31 ( .A(Inst_f1_phpplmul_summul_n340), .B(
        Inst_f1_phpplmul_summul_n264), .ZN(Inst_f1_phpplmul_summul_n266) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U30 ( .A(Inst_f1_phpplmul_summul_n263), .B(
        Inst_f1_phpplmul_summul_n262), .ZN(Inst_f1_phpplmul_summul_n264) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U29 ( .A(Inst_f1_phpplmul_summul_n261), .B(
        Inst_f1_phpplmul_summul_n260), .ZN(Inst_f1_phpplmul_summul_n262) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U28 ( .A(Inst_f1_phpplmul_summul_n259), .B(
        Inst_f1_phpplmul_summul_n279), .ZN(Inst_f1_phpplmul_summul_n260) );
  NAND2_X1 Inst_f1_phpplmul_summul_U27 ( .A1(Inst_f1_phpplmul_sB[2]), .A2(
        Inst_f1_phpplmul_summul_n258), .ZN(Inst_f1_phpplmul_summul_n279) );
  XOR2_X1 Inst_f1_phpplmul_summul_U26 ( .A(Inst_f1_phpplmul_sA[3]), .B(
        Inst_f1_phpplmul_sA[5]), .Z(Inst_f1_phpplmul_summul_n258) );
  NOR2_X1 Inst_f1_phpplmul_summul_U25 ( .A1(Inst_f1_phpplmul_summul_n257), 
        .A2(Inst_f1_phpplmul_summul_n319), .ZN(Inst_f1_phpplmul_summul_n259)
         );
  INV_X1 Inst_f1_phpplmul_summul_U24 ( .A(Inst_f1_phpplmul_sB[3]), .ZN(
        Inst_f1_phpplmul_summul_n319) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U23 ( .A(Inst_f1_phpplmul_sA[5]), .B(
        Inst_f1_phpplmul_sA[4]), .ZN(Inst_f1_phpplmul_summul_n257) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U22 ( .A(Inst_f1_phpplmul_summul_n282), .B(
        Inst_f1_phpplmul_sB[4]), .ZN(Inst_f1_phpplmul_summul_n261) );
  NAND2_X1 Inst_f1_phpplmul_summul_U21 ( .A1(Inst_f1_phpplmul_sA[4]), .A2(
        Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n282) );
  NOR2_X1 Inst_f1_phpplmul_summul_U20 ( .A1(Inst_f1_phpplmul_summul_n326), 
        .A2(Inst_f1_phpplmul_summul_n308), .ZN(Inst_f1_phpplmul_summul_n263)
         );
  XNOR2_X1 Inst_f1_phpplmul_summul_U19 ( .A(Inst_f1_phpplmul_sB[4]), .B(
        Inst_f1_phpplmul_sB[5]), .ZN(Inst_f1_phpplmul_summul_n308) );
  INV_X1 Inst_f1_phpplmul_summul_U18 ( .A(Inst_f1_phpplmul_sA[3]), .ZN(
        Inst_f1_phpplmul_summul_n326) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U17 ( .A(Inst_f1_phpplmul_summul_n269), .B(
        Inst_f1_phpplmul_summul_n256), .ZN(Inst_f1_phpplmul_summul_n340) );
  NAND2_X1 Inst_f1_phpplmul_summul_U16 ( .A1(Inst_f1_phpplmul_sA[2]), .A2(
        Inst_f1_phpplmul_sB[2]), .ZN(Inst_f1_phpplmul_summul_n256) );
  NAND2_X1 Inst_f1_phpplmul_summul_U15 ( .A1(Inst_f1_phpplmul_sB[3]), .A2(
        Inst_f1_phpplmul_sA[3]), .ZN(Inst_f1_phpplmul_summul_n269) );
  XOR2_X1 Inst_f1_phpplmul_summul_U14 ( .A(Inst_f1_phpplmul_summul_n340), .B(
        Inst_f1_phpplmul_summul_n255), .Z(Inst_f1_phpplmul_Orig_p[5]) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U13 ( .A(Inst_f1_phpplmul_summul_n254), .B(
        Inst_f1_phpplmul_summul_n252), .ZN(Inst_f1_phpplmul_summul_n255) );
  NAND2_X1 Inst_f1_phpplmul_summul_U12 ( .A1(Inst_f1_phpplmul_summul_n253), 
        .A2(Inst_f1_phpplmul_summul_n249), .ZN(Inst_f1_phpplmul_summul_n254)
         );
  NAND2_X1 Inst_f1_phpplmul_summul_U11 ( .A1(Inst_f1_phpplmul_summul_n243), 
        .A2(Inst_f1_phpplmul_sB[1]), .ZN(Inst_f1_phpplmul_summul_n253) );
  XOR2_X1 Inst_f1_phpplmul_summul_U10 ( .A(Inst_f1_phpplmul_summul_n339), .B(
        Inst_f1_phpplmul_summul_n251), .Z(Inst_f1_phpplmul_summul_n252) );
  NOR2_X1 Inst_f1_phpplmul_summul_U9 ( .A1(Inst_f1_phpplmul_summul_n338), .A2(
        Inst_f1_phpplmul_summul_n250), .ZN(Inst_f1_phpplmul_summul_n251) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U8 ( .A(Inst_f1_phpplmul_sB[2]), .B(
        Inst_f1_phpplmul_sB[3]), .ZN(Inst_f1_phpplmul_summul_n250) );
  XOR2_X1 Inst_f1_phpplmul_summul_U7 ( .A(Inst_f1_phpplmul_summul_n246), .B(
        Inst_f1_phpplmul_summul_n248), .Z(Inst_f1_phpplmul_summul_n249) );
  NAND2_X1 Inst_f1_phpplmul_summul_U6 ( .A1(Inst_f1_phpplmul_summul_n247), 
        .A2(Inst_f1_phpplmul_sA[1]), .ZN(Inst_f1_phpplmul_summul_n248) );
  NAND2_X1 Inst_f1_phpplmul_summul_U5 ( .A1(Inst_f1_phpplmul_sB[0]), .A2(
        Inst_f1_phpplmul_summul_n337), .ZN(Inst_f1_phpplmul_summul_n247) );
  NAND2_X1 Inst_f1_phpplmul_summul_U4 ( .A1(Inst_f1_phpplmul_sB[0]), .A2(
        Inst_f1_phpplmul_summul_n245), .ZN(Inst_f1_phpplmul_summul_n246) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U3 ( .A(Inst_f1_phpplmul_summul_n244), .B(
        Inst_f1_phpplmul_sA[3]), .ZN(Inst_f1_phpplmul_summul_n245) );
  XNOR2_X1 Inst_f1_phpplmul_summul_U2 ( .A(Inst_f1_phpplmul_sA[0]), .B(
        Inst_f1_phpplmul_sA[2]), .ZN(Inst_f1_phpplmul_summul_n244) );
  INV_X1 Inst_f1_phpplmul_summul_U1 ( .A(Inst_f1_phpplmul_sB[0]), .ZN(
        Inst_f1_phpplmul_summul_n243) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_MaskXORInst_U2 ( .A(PRNGQ[4]), .B(
        PRNGQ[6]), .Z(Inst_f1_phpplmul_AddNewMaskp_MaskXOR[0]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_MaskXORInst_U1 ( .A(PRNGQ[5]), .B(
        PRNGQ[7]), .Z(Inst_f1_phpplmul_AddNewMaskp_MaskXOR[1]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_XORInst1_U2 ( .A(
        Inst_f1_phpplmul_Orig_p[4]), .B(
        Inst_f1_phpplmul_AddNewMaskp_MaskXOR[0]), .Z(p[4]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_XORInst1_U1 ( .A(
        Inst_f1_phpplmul_Orig_p[5]), .B(
        Inst_f1_phpplmul_AddNewMaskp_MaskXOR[1]), .Z(p[5]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_XORInst2_U4 ( .A(
        Inst_f1_phpplmul_Orig_p[3]), .B(PRNGQ[7]), .Z(p[3]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_XORInst2_U3 ( .A(
        Inst_f1_phpplmul_Orig_p[2]), .B(PRNGQ[6]), .Z(p[2]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_XORInst2_U2 ( .A(
        Inst_f1_phpplmul_Orig_p[1]), .B(PRNGQ[5]), .Z(p[1]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskp_XORInst2_U1 ( .A(
        Inst_f1_phpplmul_Orig_p[0]), .B(PRNGQ[4]), .Z(p[0]) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U104 ( .A(Inst_f1_phpplmul_lowmul_n336), 
        .B(Inst_f1_phpplmul_lowmul_n335), .ZN(Inst_f1_phpplmul_Orig_pl[4]) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U103 ( .A(Inst_f1_phpplmul_lowmul_n334), 
        .B(Inst_f1_phpplmul_lowmul_n333), .ZN(Inst_f1_phpplmul_lowmul_n335) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U102 ( .A(Inst_f1_phpplmul_lowmul_n332), 
        .B(Inst_f1_phpplmul_lowmul_n331), .ZN(Inst_f1_phpplmul_lowmul_n333) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U101 ( .A1(Inst_f1_phpplmul_lowmul_n330), 
        .A2(Zh_f1[4]), .ZN(Inst_f1_phpplmul_lowmul_n332) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U100 ( .A1(Inst_f1_phpplmul_lowmul_n329), 
        .A2(Inst_f1_phpplmul_lowmul_n328), .ZN(Inst_f1_phpplmul_lowmul_n334)
         );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U99 ( .A1(Zl_f1_0_), .A2(
        Inst_f1_phpplmul_lowmul_n327), .ZN(Inst_f1_phpplmul_lowmul_n328) );
  OR2_X1 Inst_f1_phpplmul_lowmul_U98 ( .A1(Inst_f1_phpplmul_lowmul_n327), .A2(
        Inst_f1_phpplmul_lowmul_n337), .ZN(Inst_f1_phpplmul_lowmul_n329) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U97 ( .A(Zh_f1[1]), .B(
        Inst_f1_phpplmul_lowmul_n326), .Z(Inst_f1_phpplmul_lowmul_n327) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U96 ( .A(Inst_f1_phpplmul_lowmul_n325), .B(
        Inst_f1_phpplmul_lowmul_n339), .ZN(Inst_f1_phpplmul_lowmul_n336) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U95 ( .A(Inst_f1_phpplmul_lowmul_n324), .B(
        Inst_f1_phpplmul_lowmul_n323), .Z(Inst_f1_phpplmul_lowmul_n339) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U94 ( .A1(Zl_f1_4_), .A2(Zh_f1[1]), .ZN(
        Inst_f1_phpplmul_lowmul_n323) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U93 ( .A1(Inst_f1_phpplmul_lowmul_n322), 
        .A2(Inst_f1_phpplmul_lowmul_n337), .ZN(Inst_f1_phpplmul_lowmul_n324)
         );
  INV_X1 Inst_f1_phpplmul_lowmul_U92 ( .A(Zl_f1_1_), .ZN(
        Inst_f1_phpplmul_lowmul_n337) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U91 ( .A(Zh_f1[0]), .B(Zh_f1[4]), .ZN(
        Inst_f1_phpplmul_lowmul_n322) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U90 ( .A1(Inst_f1_phpplmul_lowmul_n321), 
        .A2(Inst_f1_phpplmul_lowmul_n320), .ZN(Inst_f1_phpplmul_lowmul_n325)
         );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U89 ( .A1(Zh_f1[1]), .A2(
        Inst_f1_phpplmul_lowmul_n319), .ZN(Inst_f1_phpplmul_lowmul_n320) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U88 ( .A1(Zh_f1[0]), .A2(Zl_f1_5_), .ZN(
        Inst_f1_phpplmul_lowmul_n321) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U87 ( .A(Inst_f1_phpplmul_lowmul_n318), .B(
        Inst_f1_phpplmul_lowmul_n317), .ZN(Inst_f1_phpplmul_Orig_pl[3]) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U86 ( .A(Inst_f1_phpplmul_lowmul_n316), .B(
        Inst_f1_phpplmul_lowmul_n315), .ZN(Inst_f1_phpplmul_lowmul_n317) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U85 ( .A(Inst_f1_phpplmul_lowmul_n314), .B(
        Inst_f1_phpplmul_lowmul_n313), .Z(Inst_f1_phpplmul_lowmul_n316) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U84 ( .A1(Zh_f1[8]), .A2(Zl_f1_8_), .ZN(
        Inst_f1_phpplmul_lowmul_n313) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U83 ( .A1(Zh_f1[9]), .A2(Zl_f1_9_), .ZN(
        Inst_f1_phpplmul_lowmul_n314) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U82 ( .A(Inst_f1_phpplmul_lowmul_n312), .B(
        Inst_f1_phpplmul_lowmul_n311), .Z(Inst_f1_phpplmul_lowmul_n318) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U81 ( .A(Inst_f1_phpplmul_lowmul_n310), .B(
        Inst_f1_phpplmul_lowmul_n309), .Z(Inst_f1_phpplmul_lowmul_n311) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U80 ( .A1(Zh_f1[8]), .A2(
        Inst_f1_phpplmul_lowmul_n308), .ZN(Inst_f1_phpplmul_lowmul_n309) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U79 ( .A1(Zh_f1[0]), .A2(Zl_f1_9_), .ZN(
        Inst_f1_phpplmul_lowmul_n310) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U78 ( .A(Inst_f1_phpplmul_lowmul_n307), .B(
        Inst_f1_phpplmul_lowmul_n306), .ZN(Inst_f1_phpplmul_lowmul_n312) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U77 ( .A(Zh_f1[9]), .B(
        Inst_f1_phpplmul_lowmul_n305), .ZN(Inst_f1_phpplmul_lowmul_n306) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U76 ( .A(Inst_f1_phpplmul_lowmul_n304), .B(
        Inst_f1_phpplmul_lowmul_n303), .Z(Inst_f1_phpplmul_lowmul_n305) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U75 ( .A1(Zl_f1_0_), .A2(Zh_f1[8]), .ZN(
        Inst_f1_phpplmul_lowmul_n303) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U74 ( .A1(Inst_f1_phpplmul_lowmul_n302), 
        .A2(Zl_f1_1_), .ZN(Inst_f1_phpplmul_lowmul_n304) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U73 ( .A1(Inst_f1_phpplmul_lowmul_n301), 
        .A2(Zl_f1_8_), .ZN(Inst_f1_phpplmul_lowmul_n307) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U72 ( .A(Inst_f1_phpplmul_lowmul_n338), .B(
        Inst_f1_phpplmul_lowmul_n300), .ZN(Inst_f1_phpplmul_lowmul_n301) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U71 ( .A(Zh_f1[1]), .B(
        Inst_f1_phpplmul_lowmul_n299), .ZN(Inst_f1_phpplmul_lowmul_n300) );
  INV_X1 Inst_f1_phpplmul_lowmul_U70 ( .A(Zh_f1[0]), .ZN(
        Inst_f1_phpplmul_lowmul_n338) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U69 ( .A(Inst_f1_phpplmul_lowmul_n298), .B(
        Inst_f1_phpplmul_lowmul_n297), .Z(Inst_f1_phpplmul_Orig_pl[2]) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U68 ( .A1(Inst_f1_phpplmul_lowmul_n296), 
        .A2(Inst_f1_phpplmul_lowmul_n295), .ZN(Inst_f1_phpplmul_lowmul_n297)
         );
  OR2_X1 Inst_f1_phpplmul_lowmul_U67 ( .A1(Zl_f1_9_), .A2(
        Inst_f1_phpplmul_lowmul_n302), .ZN(Inst_f1_phpplmul_lowmul_n295) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U66 ( .A1(Inst_f1_phpplmul_lowmul_n294), 
        .A2(Zl_f1_9_), .ZN(Inst_f1_phpplmul_lowmul_n296) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U65 ( .A(Inst_f1_phpplmul_lowmul_n293), .B(
        Zh_f1[0]), .ZN(Inst_f1_phpplmul_lowmul_n294) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U64 ( .A(Inst_f1_phpplmul_lowmul_n292), .B(
        Inst_f1_phpplmul_lowmul_n291), .Z(Inst_f1_phpplmul_lowmul_n298) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U63 ( .A1(Inst_f1_phpplmul_lowmul_n299), 
        .A2(Inst_f1_phpplmul_lowmul_n290), .ZN(Inst_f1_phpplmul_lowmul_n291)
         );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U62 ( .A(Inst_f1_phpplmul_lowmul_n308), .B(
        Zl_f1_1_), .Z(Inst_f1_phpplmul_lowmul_n290) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U61 ( .A(Inst_f1_phpplmul_lowmul_n289), .B(
        Inst_f1_phpplmul_lowmul_n288), .ZN(Inst_f1_phpplmul_lowmul_n292) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U60 ( .A(Zl_f1_0_), .B(
        Inst_f1_phpplmul_lowmul_n331), .ZN(Inst_f1_phpplmul_lowmul_n288) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U59 ( .A(Inst_f1_phpplmul_lowmul_n287), .B(
        Inst_f1_phpplmul_lowmul_n286), .Z(Inst_f1_phpplmul_lowmul_n331) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U58 ( .A1(Zh_f1[1]), .A2(Zl_f1_0_), .ZN(
        Inst_f1_phpplmul_lowmul_n286) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U57 ( .A1(Zh_f1[0]), .A2(Zl_f1_1_), .ZN(
        Inst_f1_phpplmul_lowmul_n287) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U56 ( .A(Inst_f1_phpplmul_lowmul_n285), .B(
        Inst_f1_phpplmul_lowmul_n315), .Z(Inst_f1_phpplmul_lowmul_n289) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U55 ( .A(Inst_f1_phpplmul_lowmul_n284), .B(
        Inst_f1_phpplmul_lowmul_n283), .Z(Inst_f1_phpplmul_lowmul_n315) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U54 ( .A1(Zh_f1[8]), .A2(Zl_f1_1_), .ZN(
        Inst_f1_phpplmul_lowmul_n283) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U53 ( .A1(Zh_f1[9]), .A2(Zl_f1_0_), .ZN(
        Inst_f1_phpplmul_lowmul_n284) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U52 ( .A(Inst_f1_phpplmul_lowmul_n282), .B(
        Inst_f1_phpplmul_lowmul_n281), .Z(Inst_f1_phpplmul_lowmul_n285) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U51 ( .A1(Zl_f1_8_), .A2(
        Inst_f1_phpplmul_lowmul_n302), .ZN(Inst_f1_phpplmul_lowmul_n281) );
  INV_X1 Inst_f1_phpplmul_lowmul_U50 ( .A(Zh_f1[1]), .ZN(
        Inst_f1_phpplmul_lowmul_n302) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U49 ( .A(Inst_f1_phpplmul_lowmul_n280), .B(
        Inst_f1_phpplmul_lowmul_n279), .ZN(Inst_f1_phpplmul_Orig_pl[1]) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U48 ( .A(Inst_f1_phpplmul_lowmul_n278), .B(
        Inst_f1_phpplmul_lowmul_n277), .ZN(Inst_f1_phpplmul_lowmul_n280) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U47 ( .A1(Inst_f1_phpplmul_lowmul_n276), 
        .A2(Zh_f1[4]), .ZN(Inst_f1_phpplmul_lowmul_n277) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U46 ( .A(Zl_f1_4_), .B(
        Inst_f1_phpplmul_lowmul_n308), .ZN(Inst_f1_phpplmul_lowmul_n276) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U45 ( .A(Inst_f1_phpplmul_lowmul_n275), .B(
        Inst_f1_phpplmul_lowmul_n274), .ZN(Inst_f1_phpplmul_lowmul_n278) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U44 ( .A(Inst_f1_phpplmul_lowmul_n273), .B(
        Inst_f1_phpplmul_lowmul_n272), .ZN(Inst_f1_phpplmul_lowmul_n274) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U43 ( .A1(Inst_f1_phpplmul_lowmul_n271), 
        .A2(Inst_f1_phpplmul_lowmul_n330), .ZN(Inst_f1_phpplmul_lowmul_n272)
         );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U42 ( .A(Zl_f1_4_), .B(Zl_f1_5_), .Z(
        Inst_f1_phpplmul_lowmul_n330) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U41 ( .A(Zh_f1[4]), .B(Zh_f1[8]), .Z(
        Inst_f1_phpplmul_lowmul_n271) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U40 ( .A1(Zh_f1[5]), .A2(Zl_f1_8_), .ZN(
        Inst_f1_phpplmul_lowmul_n273) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U39 ( .A(Inst_f1_phpplmul_lowmul_n270), .B(
        Inst_f1_phpplmul_lowmul_n269), .ZN(Inst_f1_phpplmul_lowmul_n275) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U38 ( .A(Inst_f1_phpplmul_lowmul_n268), .B(
        Inst_f1_phpplmul_lowmul_n267), .Z(Inst_f1_phpplmul_lowmul_n270) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U37 ( .A1(Inst_f1_phpplmul_lowmul_n293), 
        .A2(Zl_f1_8_), .ZN(Inst_f1_phpplmul_lowmul_n267) );
  INV_X1 Inst_f1_phpplmul_lowmul_U36 ( .A(Zh_f1[8]), .ZN(
        Inst_f1_phpplmul_lowmul_n293) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U35 ( .A1(Inst_f1_phpplmul_lowmul_n299), 
        .A2(Zl_f1_9_), .ZN(Inst_f1_phpplmul_lowmul_n268) );
  INV_X1 Inst_f1_phpplmul_lowmul_U34 ( .A(Zh_f1[9]), .ZN(
        Inst_f1_phpplmul_lowmul_n299) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U33 ( .A(Inst_f1_phpplmul_lowmul_n266), .B(
        Inst_f1_phpplmul_lowmul_n265), .ZN(Inst_f1_phpplmul_Orig_pl[0]) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U32 ( .A1(Zh_f1[4]), .A2(Zl_f1_9_), .ZN(
        Inst_f1_phpplmul_lowmul_n265) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U31 ( .A(Inst_f1_phpplmul_lowmul_n340), .B(
        Inst_f1_phpplmul_lowmul_n264), .ZN(Inst_f1_phpplmul_lowmul_n266) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U30 ( .A(Inst_f1_phpplmul_lowmul_n263), .B(
        Inst_f1_phpplmul_lowmul_n262), .ZN(Inst_f1_phpplmul_lowmul_n264) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U29 ( .A(Inst_f1_phpplmul_lowmul_n261), .B(
        Inst_f1_phpplmul_lowmul_n260), .ZN(Inst_f1_phpplmul_lowmul_n262) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U28 ( .A(Inst_f1_phpplmul_lowmul_n259), .B(
        Inst_f1_phpplmul_lowmul_n279), .ZN(Inst_f1_phpplmul_lowmul_n260) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U27 ( .A1(Zl_f1_4_), .A2(
        Inst_f1_phpplmul_lowmul_n258), .ZN(Inst_f1_phpplmul_lowmul_n279) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U26 ( .A(Zh_f1[5]), .B(Zh_f1[9]), .Z(
        Inst_f1_phpplmul_lowmul_n258) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U25 ( .A1(Inst_f1_phpplmul_lowmul_n257), 
        .A2(Inst_f1_phpplmul_lowmul_n319), .ZN(Inst_f1_phpplmul_lowmul_n259)
         );
  INV_X1 Inst_f1_phpplmul_lowmul_U24 ( .A(Zl_f1_5_), .ZN(
        Inst_f1_phpplmul_lowmul_n319) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U23 ( .A(Zh_f1[9]), .B(Zh_f1[8]), .ZN(
        Inst_f1_phpplmul_lowmul_n257) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U22 ( .A(Inst_f1_phpplmul_lowmul_n282), .B(
        Zl_f1_8_), .ZN(Inst_f1_phpplmul_lowmul_n261) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U21 ( .A1(Zh_f1[8]), .A2(Zl_f1_9_), .ZN(
        Inst_f1_phpplmul_lowmul_n282) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U20 ( .A1(Inst_f1_phpplmul_lowmul_n326), 
        .A2(Inst_f1_phpplmul_lowmul_n308), .ZN(Inst_f1_phpplmul_lowmul_n263)
         );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U19 ( .A(Zl_f1_8_), .B(Zl_f1_9_), .ZN(
        Inst_f1_phpplmul_lowmul_n308) );
  INV_X1 Inst_f1_phpplmul_lowmul_U18 ( .A(Zh_f1[5]), .ZN(
        Inst_f1_phpplmul_lowmul_n326) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U17 ( .A(Inst_f1_phpplmul_lowmul_n269), .B(
        Inst_f1_phpplmul_lowmul_n256), .ZN(Inst_f1_phpplmul_lowmul_n340) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U16 ( .A1(Zh_f1[4]), .A2(Zl_f1_4_), .ZN(
        Inst_f1_phpplmul_lowmul_n256) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U15 ( .A1(Zl_f1_5_), .A2(Zh_f1[5]), .ZN(
        Inst_f1_phpplmul_lowmul_n269) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U14 ( .A(Inst_f1_phpplmul_lowmul_n340), .B(
        Inst_f1_phpplmul_lowmul_n255), .Z(Inst_f1_phpplmul_Orig_pl[5]) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U13 ( .A(Inst_f1_phpplmul_lowmul_n254), .B(
        Inst_f1_phpplmul_lowmul_n252), .ZN(Inst_f1_phpplmul_lowmul_n255) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U12 ( .A1(Inst_f1_phpplmul_lowmul_n253), 
        .A2(Inst_f1_phpplmul_lowmul_n249), .ZN(Inst_f1_phpplmul_lowmul_n254)
         );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U11 ( .A1(Inst_f1_phpplmul_lowmul_n243), 
        .A2(Zl_f1_1_), .ZN(Inst_f1_phpplmul_lowmul_n253) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U10 ( .A(Inst_f1_phpplmul_lowmul_n339), .B(
        Inst_f1_phpplmul_lowmul_n251), .Z(Inst_f1_phpplmul_lowmul_n252) );
  NOR2_X1 Inst_f1_phpplmul_lowmul_U9 ( .A1(Inst_f1_phpplmul_lowmul_n338), .A2(
        Inst_f1_phpplmul_lowmul_n250), .ZN(Inst_f1_phpplmul_lowmul_n251) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U8 ( .A(Zl_f1_4_), .B(Zl_f1_5_), .ZN(
        Inst_f1_phpplmul_lowmul_n250) );
  XOR2_X1 Inst_f1_phpplmul_lowmul_U7 ( .A(Inst_f1_phpplmul_lowmul_n246), .B(
        Inst_f1_phpplmul_lowmul_n248), .Z(Inst_f1_phpplmul_lowmul_n249) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U6 ( .A1(Inst_f1_phpplmul_lowmul_n247), 
        .A2(Zh_f1[1]), .ZN(Inst_f1_phpplmul_lowmul_n248) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U5 ( .A1(Zl_f1_0_), .A2(
        Inst_f1_phpplmul_lowmul_n337), .ZN(Inst_f1_phpplmul_lowmul_n247) );
  NAND2_X1 Inst_f1_phpplmul_lowmul_U4 ( .A1(Zl_f1_0_), .A2(
        Inst_f1_phpplmul_lowmul_n245), .ZN(Inst_f1_phpplmul_lowmul_n246) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U3 ( .A(Inst_f1_phpplmul_lowmul_n244), .B(
        Zh_f1[5]), .ZN(Inst_f1_phpplmul_lowmul_n245) );
  XNOR2_X1 Inst_f1_phpplmul_lowmul_U2 ( .A(Zh_f1[0]), .B(Zh_f1[4]), .ZN(
        Inst_f1_phpplmul_lowmul_n244) );
  INV_X1 Inst_f1_phpplmul_lowmul_U1 ( .A(Zl_f1_0_), .ZN(
        Inst_f1_phpplmul_lowmul_n243) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_MaskXORInst_U2 ( .A(PRNGQ[8]), .B(
        PRNGQ[10]), .Z(Inst_f1_phpplmul_AddNewMaskpl_MaskXOR[0]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_MaskXORInst_U1 ( .A(PRNGQ[9]), .B(
        PRNGQ[11]), .Z(Inst_f1_phpplmul_AddNewMaskpl_MaskXOR[1]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_XORInst1_U2 ( .A(
        Inst_f1_phpplmul_Orig_pl[4]), .B(
        Inst_f1_phpplmul_AddNewMaskpl_MaskXOR[0]), .Z(pl[4]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_XORInst1_U1 ( .A(
        Inst_f1_phpplmul_Orig_pl[5]), .B(
        Inst_f1_phpplmul_AddNewMaskpl_MaskXOR[1]), .Z(pl[5]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_XORInst2_U4 ( .A(
        Inst_f1_phpplmul_Orig_pl[3]), .B(PRNGQ[11]), .Z(pl[3]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_XORInst2_U3 ( .A(
        Inst_f1_phpplmul_Orig_pl[2]), .B(PRNGQ[10]), .Z(pl[2]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_XORInst2_U2 ( .A(
        Inst_f1_phpplmul_Orig_pl[1]), .B(PRNGQ[9]), .Z(pl[1]) );
  XOR2_X1 Inst_f1_phpplmul_AddNewMaskpl_XORInst2_U1 ( .A(
        Inst_f1_phpplmul_Orig_pl[0]), .B(PRNGQ[8]), .Z(pl[0]) );
  DFF_X1 PL_1_s_current_state_reg_0_ ( .D(pl[0]), .CK(clk), .Q(FF1_out[0]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_1_ ( .D(pl[1]), .CK(clk), .Q(FF1_out[1]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_2_ ( .D(pl[2]), .CK(clk), .Q(FF1_out[2]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_3_ ( .D(pl[3]), .CK(clk), .Q(FF1_out[3]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_4_ ( .D(pl[4]), .CK(clk), .Q(FF1_out[4]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_5_ ( .D(pl[5]), .CK(clk), .Q(FF1_out[5]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_6_ ( .D(p[0]), .CK(clk), .Q(
        Inst_f2_abmul_pw2_1_), .QN() );
  DFF_X1 PL_1_s_current_state_reg_7_ ( .D(p[1]), .CK(clk), .Q(FF1_out[7]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_8_ ( .D(p[2]), .CK(clk), .Q(
        Inst_f2_abmul_pw2_3_), .QN() );
  DFF_X1 PL_1_s_current_state_reg_9_ ( .D(p[3]), .CK(clk), .Q(FF1_out[9]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_10_ ( .D(p[4]), .CK(clk), .Q(
        Inst_f2_abmul_pw2_5_), .QN() );
  DFF_X1 PL_1_s_current_state_reg_11_ ( .D(p[5]), .CK(clk), .Q(FF1_out[11]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_12_ ( .D(ph[0]), .CK(clk), .Q(FF1_out[12]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_13_ ( .D(ph[1]), .CK(clk), .Q(FF1_out[13]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_14_ ( .D(ph[2]), .CK(clk), .Q(FF1_out[14]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_15_ ( .D(ph[3]), .CK(clk), .Q(FF1_out[15]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_16_ ( .D(ph[4]), .CK(clk), .Q(FF1_out[16]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_17_ ( .D(ph[5]), .CK(clk), .Q(FF1_out[17]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_18_ ( .D(ab2[0]), .CK(clk), .Q(FF1_out[18]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_19_ ( .D(ab2[1]), .CK(clk), .Q(FF1_out[19]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_20_ ( .D(ab2[2]), .CK(clk), .Q(FF1_out[20]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_21_ ( .D(ab2[3]), .CK(clk), .Q(FF1_out[21]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_22_ ( .D(ab2[4]), .CK(clk), .Q(FF1_out[22]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_23_ ( .D(ab2[5]), .CK(clk), .Q(FF1_out[23]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_24_ ( .D(ab2[6]), .CK(clk), .Q(FF1_out[24]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_25_ ( .D(ab2[7]), .CK(clk), .Q(FF1_out[25]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_26_ ( .D(ab2[8]), .CK(clk), .Q(FF1_out[26]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_27_ ( .D(ab2[9]), .CK(clk), .Q(FF1_out[27]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_28_ ( .D(ab2[10]), .CK(clk), .Q(FF1_out[28]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_29_ ( .D(ab2[11]), .CK(clk), .Q(FF1_out[29]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_30_ ( .D(Zl_f1_0_), .CK(clk), .Q(Zl_f2[0]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_31_ ( .D(Zl_f1_1_), .CK(clk), .Q(Zl_f2[1]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_32_ ( .D(A[0]), .CK(clk), .Q(Zl_f2[2]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_33_ ( .D(Zl_f1_3_), .CK(clk), .Q(Zl_f2[3]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_34_ ( .D(Zl_f1_4_), .CK(clk), .Q(Zl_f2[4]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_35_ ( .D(Zl_f1_5_), .CK(clk), .Q(Zl_f2[5]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_36_ ( .D(A[8]), .CK(clk), .Q(Zl_f2[6]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_37_ ( .D(Zl_f1_7_), .CK(clk), .Q(Zl_f2[7]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_38_ ( .D(Zl_f1_8_), .CK(clk), .Q(Zl_f2[8]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_39_ ( .D(Zl_f1_9_), .CK(clk), .Q(Zl_f2[9]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_40_ ( .D(A[16]), .CK(clk), .Q(Zl_f2[10]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_41_ ( .D(Zl_f1_11_), .CK(clk), .Q(Zl_f2[11]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_42_ ( .D(Zh_f1[0]), .CK(clk), .Q(Zh_f2[0]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_43_ ( .D(Zh_f1[1]), .CK(clk), .Q(Zh_f2[1]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_44_ ( .D(Zh_f1[2]), .CK(clk), .Q(Zh_f2[2]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_45_ ( .D(Zh_f1[3]), .CK(clk), .Q(Zh_f2[3]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_46_ ( .D(Zh_f1[4]), .CK(clk), .Q(Zh_f2[4]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_47_ ( .D(Zh_f1[5]), .CK(clk), .Q(Zh_f2[5]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_48_ ( .D(Zh_f1[6]), .CK(clk), .Q(Zh_f2[6]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_49_ ( .D(Zh_f1[7]), .CK(clk), .Q(Zh_f2[7]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_50_ ( .D(Zh_f1[8]), .CK(clk), .Q(Zh_f2[8]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_51_ ( .D(Zh_f1[9]), .CK(clk), .Q(Zh_f2[9]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_52_ ( .D(Zh_f1[10]), .CK(clk), .Q(Zh_f2[10]), 
        .QN() );
  DFF_X1 PL_1_s_current_state_reg_53_ ( .D(Zh_f1[11]), .CK(clk), .Q(Zh_f2[11]), 
        .QN() );
  XOR2_X1 Inst_f2_U12 ( .A(FF1_out[27]), .B(Inst_f2_abin[9]), .Z(gamma0[5]) );
  XOR2_X1 Inst_f2_U11 ( .A(FF1_out[26]), .B(Inst_f2_abin[8]), .Z(gamma0[4]) );
  XOR2_X1 Inst_f2_U10 ( .A(FF1_out[25]), .B(Inst_f2_abin[7]), .Z(gamma1[3]) );
  XOR2_X1 Inst_f2_U9 ( .A(FF1_out[24]), .B(Inst_f2_abin[6]), .Z(gamma1[2]) );
  XOR2_X1 Inst_f2_U8 ( .A(FF1_out[23]), .B(Inst_f2_abin[5]), .Z(gamma0[3]) );
  XOR2_X1 Inst_f2_U7 ( .A(FF1_out[22]), .B(Inst_f2_abin[4]), .Z(gamma0[2]) );
  XOR2_X1 Inst_f2_U6 ( .A(FF1_out[21]), .B(Inst_f2_abin[3]), .Z(gamma1[1]) );
  XOR2_X1 Inst_f2_U5 ( .A(FF1_out[20]), .B(Inst_f2_abin[2]), .Z(gamma1[0]) );
  XOR2_X1 Inst_f2_U4 ( .A(FF1_out[19]), .B(Inst_f2_abin[1]), .Z(gamma0[1]) );
  XOR2_X1 Inst_f2_U3 ( .A(FF1_out[29]), .B(Inst_f2_abin[11]), .Z(gamma1[5]) );
  XOR2_X1 Inst_f2_U2 ( .A(FF1_out[18]), .B(Inst_f2_abin[0]), .Z(gamma0[0]) );
  XOR2_X2 Inst_f2_U1 ( .A(FF1_out[28]), .B(Inst_f2_abin[10]), .Z(gamma1[4]) );
  XOR2_X1 Inst_f2_abmul_U12 ( .A(Inst_f2_abmul_pw2_5_), .B(FF1_out[5]), .Z(
        Inst_f2_abin[9]) );
  XOR2_X1 Inst_f2_abmul_U11 ( .A(Inst_f2_abmul_pw2_4_), .B(FF1_out[4]), .Z(
        Inst_f2_abin[8]) );
  XOR2_X1 Inst_f2_abmul_U10 ( .A(Inst_f2_abmul_pw2_3_), .B(FF1_out[15]), .Z(
        Inst_f2_abin[7]) );
  XOR2_X1 Inst_f2_abmul_U9 ( .A(Inst_f2_abmul_pw2_2_), .B(FF1_out[14]), .Z(
        Inst_f2_abin[6]) );
  XOR2_X1 Inst_f2_abmul_U8 ( .A(Inst_f2_abmul_pw2_3_), .B(FF1_out[3]), .Z(
        Inst_f2_abin[5]) );
  XOR2_X1 Inst_f2_abmul_U7 ( .A(Inst_f2_abmul_pw2_2_), .B(FF1_out[2]), .Z(
        Inst_f2_abin[4]) );
  XOR2_X1 Inst_f2_abmul_U6 ( .A(Inst_f2_abmul_pw2_1_), .B(FF1_out[13]), .Z(
        Inst_f2_abin[3]) );
  XOR2_X1 Inst_f2_abmul_U5 ( .A(Inst_f2_abmul_pw2_0_), .B(FF1_out[12]), .Z(
        Inst_f2_abin[2]) );
  XOR2_X1 Inst_f2_abmul_U4 ( .A(Inst_f2_abmul_pw2_1_), .B(FF1_out[1]), .Z(
        Inst_f2_abin[1]) );
  XOR2_X1 Inst_f2_abmul_U3 ( .A(Inst_f2_abmul_pw2_5_), .B(FF1_out[17]), .Z(
        Inst_f2_abin[11]) );
  XOR2_X1 Inst_f2_abmul_U2 ( .A(Inst_f2_abmul_pw2_4_), .B(FF1_out[16]), .Z(
        Inst_f2_abin[10]) );
  XOR2_X1 Inst_f2_abmul_U1 ( .A(Inst_f2_abmul_pw2_0_), .B(FF1_out[0]), .Z(
        Inst_f2_abin[0]) );
  XOR2_X1 Inst_f2_abmul_NxGAMMA_U3 ( .A(Inst_f2_abmul_pw2_5_), .B(FF1_out[11]), 
        .Z(Inst_f2_abmul_pw2_4_) );
  XOR2_X1 Inst_f2_abmul_NxGAMMA_U2 ( .A(Inst_f2_abmul_pw2_3_), .B(FF1_out[9]), 
        .Z(Inst_f2_abmul_pw2_2_) );
  XOR2_X1 Inst_f2_abmul_NxGAMMA_U1 ( .A(Inst_f2_abmul_pw2_1_), .B(FF1_out[7]), 
        .Z(Inst_f2_abmul_pw2_0_) );
  XOR2_X1 Inst_f2_dinv_1_U6 ( .A(gamma1[5]), .B(gamma0[5]), .Z(
        Inst_f2_dinv_1_Orig_sA2N[5]) );
  XOR2_X1 Inst_f2_dinv_1_U5 ( .A(gamma1[4]), .B(gamma0[4]), .Z(
        Inst_f2_dinv_1_sA2[5]) );
  XOR2_X1 Inst_f2_dinv_1_U4 ( .A(gamma0[3]), .B(gamma1[3]), .Z(
        Inst_f2_dinv_1_Orig_sA2N[3]) );
  XOR2_X1 Inst_f2_dinv_1_U3 ( .A(gamma0[2]), .B(gamma1[2]), .Z(
        Inst_f2_dinv_1_sA2[3]) );
  XOR2_X1 Inst_f2_dinv_1_U2 ( .A(gamma0[1]), .B(gamma1[1]), .Z(
        Inst_f2_dinv_1_Orig_sA2N[1]) );
  XOR2_X1 Inst_f2_dinv_1_U1 ( .A(gamma0[0]), .B(gamma1[0]), .Z(
        Inst_f2_dinv_1_sA2[1]) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U104 ( .A(Inst_f2_dinv_1_mul_n340), .B(
        Inst_f2_dinv_1_mul_n339), .ZN(Inst_f2_dinv_1_Orig_ab[5]) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U103 ( .A(Inst_f2_dinv_1_mul_n338), .B(
        Inst_f2_dinv_1_mul_n337), .ZN(Inst_f2_dinv_1_mul_n340) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U102 ( .A(Inst_f2_dinv_1_mul_n336), .B(
        Inst_f2_dinv_1_mul_n335), .ZN(Inst_f2_dinv_1_mul_n337) );
  NOR2_X1 Inst_f2_dinv_1_mul_U101 ( .A1(Inst_f2_dinv_1_mul_n334), .A2(
        Inst_f2_dinv_1_mul_n333), .ZN(Inst_f2_dinv_1_mul_n336) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U100 ( .A(gamma0[2]), .B(gamma0[3]), .ZN(
        Inst_f2_dinv_1_mul_n334) );
  NAND2_X1 Inst_f2_dinv_1_mul_U99 ( .A1(Inst_f2_dinv_1_mul_n332), .A2(
        Inst_f2_dinv_1_mul_n331), .ZN(Inst_f2_dinv_1_mul_n338) );
  NAND2_X1 Inst_f2_dinv_1_mul_U98 ( .A1(Inst_f2_dinv_1_mul_n330), .A2(
        gamma0[1]), .ZN(Inst_f2_dinv_1_mul_n331) );
  NOR2_X1 Inst_f2_dinv_1_mul_U97 ( .A1(Inst_f2_dinv_1_mul_n329), .A2(gamma0[0]), .ZN(Inst_f2_dinv_1_mul_n330) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U96 ( .A(Inst_f2_dinv_1_mul_n329), .B(
        Inst_f2_dinv_1_mul_n328), .ZN(Inst_f2_dinv_1_mul_n332) );
  NAND2_X1 Inst_f2_dinv_1_mul_U95 ( .A1(gamma1[1]), .A2(
        Inst_f2_dinv_1_mul_n327), .ZN(Inst_f2_dinv_1_mul_n328) );
  NAND2_X1 Inst_f2_dinv_1_mul_U94 ( .A1(gamma0[0]), .A2(
        Inst_f2_dinv_1_mul_n326), .ZN(Inst_f2_dinv_1_mul_n327) );
  XOR2_X1 Inst_f2_dinv_1_mul_U93 ( .A(gamma1[2]), .B(gamma1[0]), .Z(
        Inst_f2_dinv_1_mul_n325) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U92 ( .A(Inst_f2_dinv_1_mul_n324), .B(
        Inst_f2_dinv_1_mul_n323), .ZN(Inst_f2_dinv_1_Orig_ab[4]) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U91 ( .A(Inst_f2_dinv_1_mul_n322), .B(
        Inst_f2_dinv_1_mul_n321), .ZN(Inst_f2_dinv_1_mul_n323) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U90 ( .A(Inst_f2_dinv_1_mul_n320), .B(
        Inst_f2_dinv_1_mul_n319), .ZN(Inst_f2_dinv_1_mul_n321) );
  NAND2_X1 Inst_f2_dinv_1_mul_U89 ( .A1(Inst_f2_dinv_1_mul_n318), .A2(
        gamma1[2]), .ZN(Inst_f2_dinv_1_mul_n320) );
  NAND2_X1 Inst_f2_dinv_1_mul_U88 ( .A1(Inst_f2_dinv_1_mul_n317), .A2(
        Inst_f2_dinv_1_mul_n316), .ZN(Inst_f2_dinv_1_mul_n322) );
  NAND2_X1 Inst_f2_dinv_1_mul_U87 ( .A1(gamma0[0]), .A2(
        Inst_f2_dinv_1_mul_n315), .ZN(Inst_f2_dinv_1_mul_n316) );
  OR2_X1 Inst_f2_dinv_1_mul_U86 ( .A1(Inst_f2_dinv_1_mul_n315), .A2(
        Inst_f2_dinv_1_mul_n326), .ZN(Inst_f2_dinv_1_mul_n317) );
  XOR2_X1 Inst_f2_dinv_1_mul_U85 ( .A(gamma1[1]), .B(Inst_f2_dinv_1_mul_n314), 
        .Z(Inst_f2_dinv_1_mul_n315) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U84 ( .A(Inst_f2_dinv_1_mul_n313), .B(
        Inst_f2_dinv_1_mul_n335), .ZN(Inst_f2_dinv_1_mul_n324) );
  XOR2_X1 Inst_f2_dinv_1_mul_U83 ( .A(Inst_f2_dinv_1_mul_n312), .B(
        Inst_f2_dinv_1_mul_n311), .Z(Inst_f2_dinv_1_mul_n335) );
  NAND2_X1 Inst_f2_dinv_1_mul_U82 ( .A1(gamma0[2]), .A2(gamma1[1]), .ZN(
        Inst_f2_dinv_1_mul_n311) );
  NOR2_X1 Inst_f2_dinv_1_mul_U81 ( .A1(Inst_f2_dinv_1_mul_n310), .A2(
        Inst_f2_dinv_1_mul_n326), .ZN(Inst_f2_dinv_1_mul_n312) );
  INV_X1 Inst_f2_dinv_1_mul_U80 ( .A(gamma0[1]), .ZN(Inst_f2_dinv_1_mul_n326)
         );
  XNOR2_X1 Inst_f2_dinv_1_mul_U79 ( .A(gamma1[0]), .B(gamma1[2]), .ZN(
        Inst_f2_dinv_1_mul_n310) );
  NAND2_X1 Inst_f2_dinv_1_mul_U78 ( .A1(Inst_f2_dinv_1_mul_n309), .A2(
        Inst_f2_dinv_1_mul_n308), .ZN(Inst_f2_dinv_1_mul_n313) );
  NAND2_X1 Inst_f2_dinv_1_mul_U77 ( .A1(gamma1[1]), .A2(
        Inst_f2_dinv_1_mul_n307), .ZN(Inst_f2_dinv_1_mul_n308) );
  NAND2_X1 Inst_f2_dinv_1_mul_U76 ( .A1(gamma1[0]), .A2(gamma0[3]), .ZN(
        Inst_f2_dinv_1_mul_n309) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U75 ( .A(Inst_f2_dinv_1_mul_n306), .B(
        Inst_f2_dinv_1_mul_n305), .ZN(Inst_f2_dinv_1_Orig_ab[3]) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U74 ( .A(Inst_f2_dinv_1_mul_n304), .B(
        Inst_f2_dinv_1_mul_n303), .ZN(Inst_f2_dinv_1_mul_n305) );
  XOR2_X1 Inst_f2_dinv_1_mul_U73 ( .A(Inst_f2_dinv_1_mul_n302), .B(
        Inst_f2_dinv_1_mul_n301), .Z(Inst_f2_dinv_1_mul_n304) );
  NAND2_X1 Inst_f2_dinv_1_mul_U72 ( .A1(gamma1[4]), .A2(gamma0[4]), .ZN(
        Inst_f2_dinv_1_mul_n301) );
  NAND2_X1 Inst_f2_dinv_1_mul_U71 ( .A1(gamma1[5]), .A2(gamma0[5]), .ZN(
        Inst_f2_dinv_1_mul_n302) );
  XOR2_X1 Inst_f2_dinv_1_mul_U70 ( .A(Inst_f2_dinv_1_mul_n300), .B(
        Inst_f2_dinv_1_mul_n299), .Z(Inst_f2_dinv_1_mul_n306) );
  XOR2_X1 Inst_f2_dinv_1_mul_U69 ( .A(Inst_f2_dinv_1_mul_n298), .B(
        Inst_f2_dinv_1_mul_n297), .Z(Inst_f2_dinv_1_mul_n299) );
  NAND2_X1 Inst_f2_dinv_1_mul_U68 ( .A1(gamma1[4]), .A2(
        Inst_f2_dinv_1_mul_n296), .ZN(Inst_f2_dinv_1_mul_n297) );
  NAND2_X1 Inst_f2_dinv_1_mul_U67 ( .A1(gamma1[0]), .A2(gamma0[5]), .ZN(
        Inst_f2_dinv_1_mul_n298) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U66 ( .A(Inst_f2_dinv_1_mul_n295), .B(
        Inst_f2_dinv_1_mul_n294), .ZN(Inst_f2_dinv_1_mul_n300) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U65 ( .A(gamma1[5]), .B(Inst_f2_dinv_1_mul_n293), 
        .ZN(Inst_f2_dinv_1_mul_n294) );
  XOR2_X1 Inst_f2_dinv_1_mul_U64 ( .A(Inst_f2_dinv_1_mul_n292), .B(
        Inst_f2_dinv_1_mul_n291), .Z(Inst_f2_dinv_1_mul_n293) );
  NAND2_X1 Inst_f2_dinv_1_mul_U63 ( .A1(gamma0[0]), .A2(gamma1[4]), .ZN(
        Inst_f2_dinv_1_mul_n291) );
  NOR2_X1 Inst_f2_dinv_1_mul_U62 ( .A1(Inst_f2_dinv_1_mul_n290), .A2(gamma0[1]), .ZN(Inst_f2_dinv_1_mul_n292) );
  NAND2_X1 Inst_f2_dinv_1_mul_U61 ( .A1(Inst_f2_dinv_1_mul_n289), .A2(
        gamma0[4]), .ZN(Inst_f2_dinv_1_mul_n295) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U60 ( .A(Inst_f2_dinv_1_mul_n333), .B(
        Inst_f2_dinv_1_mul_n288), .ZN(Inst_f2_dinv_1_mul_n289) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U59 ( .A(gamma1[1]), .B(Inst_f2_dinv_1_mul_n287), 
        .ZN(Inst_f2_dinv_1_mul_n288) );
  INV_X1 Inst_f2_dinv_1_mul_U58 ( .A(gamma1[0]), .ZN(Inst_f2_dinv_1_mul_n333)
         );
  XOR2_X1 Inst_f2_dinv_1_mul_U57 ( .A(Inst_f2_dinv_1_mul_n286), .B(
        Inst_f2_dinv_1_mul_n285), .Z(Inst_f2_dinv_1_Orig_ab[2]) );
  NAND2_X1 Inst_f2_dinv_1_mul_U56 ( .A1(Inst_f2_dinv_1_mul_n284), .A2(
        Inst_f2_dinv_1_mul_n283), .ZN(Inst_f2_dinv_1_mul_n285) );
  OR2_X1 Inst_f2_dinv_1_mul_U55 ( .A1(gamma0[5]), .A2(Inst_f2_dinv_1_mul_n290), 
        .ZN(Inst_f2_dinv_1_mul_n283) );
  NAND2_X1 Inst_f2_dinv_1_mul_U54 ( .A1(Inst_f2_dinv_1_mul_n282), .A2(
        gamma0[5]), .ZN(Inst_f2_dinv_1_mul_n284) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U53 ( .A(Inst_f2_dinv_1_mul_n281), .B(gamma1[0]), 
        .ZN(Inst_f2_dinv_1_mul_n282) );
  XOR2_X1 Inst_f2_dinv_1_mul_U52 ( .A(Inst_f2_dinv_1_mul_n280), .B(
        Inst_f2_dinv_1_mul_n279), .Z(Inst_f2_dinv_1_mul_n286) );
  NOR2_X1 Inst_f2_dinv_1_mul_U51 ( .A1(Inst_f2_dinv_1_mul_n287), .A2(
        Inst_f2_dinv_1_mul_n278), .ZN(Inst_f2_dinv_1_mul_n279) );
  XOR2_X1 Inst_f2_dinv_1_mul_U50 ( .A(Inst_f2_dinv_1_mul_n296), .B(gamma0[1]), 
        .Z(Inst_f2_dinv_1_mul_n278) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U49 ( .A(Inst_f2_dinv_1_mul_n277), .B(
        Inst_f2_dinv_1_mul_n276), .ZN(Inst_f2_dinv_1_mul_n280) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U48 ( .A(gamma0[0]), .B(Inst_f2_dinv_1_mul_n319), 
        .ZN(Inst_f2_dinv_1_mul_n276) );
  XOR2_X1 Inst_f2_dinv_1_mul_U47 ( .A(Inst_f2_dinv_1_mul_n275), .B(
        Inst_f2_dinv_1_mul_n274), .Z(Inst_f2_dinv_1_mul_n319) );
  NAND2_X1 Inst_f2_dinv_1_mul_U46 ( .A1(gamma1[1]), .A2(gamma0[0]), .ZN(
        Inst_f2_dinv_1_mul_n274) );
  NAND2_X1 Inst_f2_dinv_1_mul_U45 ( .A1(gamma1[0]), .A2(gamma0[1]), .ZN(
        Inst_f2_dinv_1_mul_n275) );
  XOR2_X1 Inst_f2_dinv_1_mul_U44 ( .A(Inst_f2_dinv_1_mul_n273), .B(
        Inst_f2_dinv_1_mul_n303), .Z(Inst_f2_dinv_1_mul_n277) );
  XOR2_X1 Inst_f2_dinv_1_mul_U43 ( .A(Inst_f2_dinv_1_mul_n272), .B(
        Inst_f2_dinv_1_mul_n271), .Z(Inst_f2_dinv_1_mul_n303) );
  NAND2_X1 Inst_f2_dinv_1_mul_U42 ( .A1(gamma1[4]), .A2(gamma0[1]), .ZN(
        Inst_f2_dinv_1_mul_n271) );
  NAND2_X1 Inst_f2_dinv_1_mul_U41 ( .A1(gamma1[5]), .A2(gamma0[0]), .ZN(
        Inst_f2_dinv_1_mul_n272) );
  XOR2_X1 Inst_f2_dinv_1_mul_U40 ( .A(Inst_f2_dinv_1_mul_n270), .B(
        Inst_f2_dinv_1_mul_n269), .Z(Inst_f2_dinv_1_mul_n273) );
  NAND2_X1 Inst_f2_dinv_1_mul_U39 ( .A1(gamma0[4]), .A2(
        Inst_f2_dinv_1_mul_n290), .ZN(Inst_f2_dinv_1_mul_n269) );
  INV_X1 Inst_f2_dinv_1_mul_U38 ( .A(gamma1[1]), .ZN(Inst_f2_dinv_1_mul_n290)
         );
  XNOR2_X1 Inst_f2_dinv_1_mul_U37 ( .A(Inst_f2_dinv_1_mul_n268), .B(
        Inst_f2_dinv_1_mul_n267), .ZN(Inst_f2_dinv_1_Orig_ab[1]) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U36 ( .A(Inst_f2_dinv_1_mul_n266), .B(
        Inst_f2_dinv_1_mul_n265), .ZN(Inst_f2_dinv_1_mul_n268) );
  NAND2_X1 Inst_f2_dinv_1_mul_U35 ( .A1(Inst_f2_dinv_1_mul_n264), .A2(
        gamma1[2]), .ZN(Inst_f2_dinv_1_mul_n265) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U34 ( .A(gamma0[2]), .B(Inst_f2_dinv_1_mul_n296), 
        .ZN(Inst_f2_dinv_1_mul_n264) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U33 ( .A(Inst_f2_dinv_1_mul_n263), .B(
        Inst_f2_dinv_1_mul_n262), .ZN(Inst_f2_dinv_1_mul_n266) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U32 ( .A(Inst_f2_dinv_1_mul_n261), .B(
        Inst_f2_dinv_1_mul_n260), .ZN(Inst_f2_dinv_1_mul_n262) );
  NAND2_X1 Inst_f2_dinv_1_mul_U31 ( .A1(Inst_f2_dinv_1_mul_n259), .A2(
        Inst_f2_dinv_1_mul_n318), .ZN(Inst_f2_dinv_1_mul_n260) );
  XOR2_X1 Inst_f2_dinv_1_mul_U30 ( .A(gamma0[2]), .B(gamma0[3]), .Z(
        Inst_f2_dinv_1_mul_n318) );
  XOR2_X1 Inst_f2_dinv_1_mul_U29 ( .A(gamma1[2]), .B(gamma1[4]), .Z(
        Inst_f2_dinv_1_mul_n259) );
  NAND2_X1 Inst_f2_dinv_1_mul_U28 ( .A1(gamma1[3]), .A2(gamma0[4]), .ZN(
        Inst_f2_dinv_1_mul_n261) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U27 ( .A(Inst_f2_dinv_1_mul_n258), .B(
        Inst_f2_dinv_1_mul_n257), .ZN(Inst_f2_dinv_1_mul_n263) );
  XOR2_X1 Inst_f2_dinv_1_mul_U26 ( .A(Inst_f2_dinv_1_mul_n256), .B(
        Inst_f2_dinv_1_mul_n255), .Z(Inst_f2_dinv_1_mul_n258) );
  NOR2_X1 Inst_f2_dinv_1_mul_U25 ( .A1(Inst_f2_dinv_1_mul_n281), .A2(gamma0[4]), .ZN(Inst_f2_dinv_1_mul_n255) );
  INV_X1 Inst_f2_dinv_1_mul_U24 ( .A(gamma1[4]), .ZN(Inst_f2_dinv_1_mul_n281)
         );
  NOR2_X1 Inst_f2_dinv_1_mul_U23 ( .A1(Inst_f2_dinv_1_mul_n287), .A2(gamma0[5]), .ZN(Inst_f2_dinv_1_mul_n256) );
  INV_X1 Inst_f2_dinv_1_mul_U22 ( .A(gamma1[5]), .ZN(Inst_f2_dinv_1_mul_n287)
         );
  XNOR2_X1 Inst_f2_dinv_1_mul_U21 ( .A(Inst_f2_dinv_1_mul_n254), .B(
        Inst_f2_dinv_1_mul_n253), .ZN(Inst_f2_dinv_1_Orig_ab[0]) );
  NAND2_X1 Inst_f2_dinv_1_mul_U20 ( .A1(gamma1[2]), .A2(gamma0[5]), .ZN(
        Inst_f2_dinv_1_mul_n253) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U19 ( .A(Inst_f2_dinv_1_mul_n339), .B(
        Inst_f2_dinv_1_mul_n252), .ZN(Inst_f2_dinv_1_mul_n254) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U18 ( .A(Inst_f2_dinv_1_mul_n251), .B(
        Inst_f2_dinv_1_mul_n250), .ZN(Inst_f2_dinv_1_mul_n252) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U17 ( .A(Inst_f2_dinv_1_mul_n249), .B(
        Inst_f2_dinv_1_mul_n248), .ZN(Inst_f2_dinv_1_mul_n250) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U16 ( .A(Inst_f2_dinv_1_mul_n247), .B(
        Inst_f2_dinv_1_mul_n267), .ZN(Inst_f2_dinv_1_mul_n248) );
  NAND2_X1 Inst_f2_dinv_1_mul_U15 ( .A1(gamma0[2]), .A2(
        Inst_f2_dinv_1_mul_n246), .ZN(Inst_f2_dinv_1_mul_n267) );
  XOR2_X1 Inst_f2_dinv_1_mul_U14 ( .A(gamma1[3]), .B(gamma1[5]), .Z(
        Inst_f2_dinv_1_mul_n246) );
  NOR2_X1 Inst_f2_dinv_1_mul_U13 ( .A1(Inst_f2_dinv_1_mul_n245), .A2(
        Inst_f2_dinv_1_mul_n307), .ZN(Inst_f2_dinv_1_mul_n247) );
  INV_X1 Inst_f2_dinv_1_mul_U12 ( .A(gamma0[3]), .ZN(Inst_f2_dinv_1_mul_n307)
         );
  XNOR2_X1 Inst_f2_dinv_1_mul_U11 ( .A(gamma1[5]), .B(gamma1[4]), .ZN(
        Inst_f2_dinv_1_mul_n245) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U10 ( .A(Inst_f2_dinv_1_mul_n270), .B(gamma0[4]), 
        .ZN(Inst_f2_dinv_1_mul_n249) );
  NAND2_X1 Inst_f2_dinv_1_mul_U9 ( .A1(gamma1[4]), .A2(gamma0[5]), .ZN(
        Inst_f2_dinv_1_mul_n270) );
  NOR2_X1 Inst_f2_dinv_1_mul_U8 ( .A1(Inst_f2_dinv_1_mul_n314), .A2(
        Inst_f2_dinv_1_mul_n296), .ZN(Inst_f2_dinv_1_mul_n251) );
  XNOR2_X1 Inst_f2_dinv_1_mul_U7 ( .A(gamma0[4]), .B(gamma0[5]), .ZN(
        Inst_f2_dinv_1_mul_n296) );
  INV_X1 Inst_f2_dinv_1_mul_U6 ( .A(gamma1[3]), .ZN(Inst_f2_dinv_1_mul_n314)
         );
  XNOR2_X1 Inst_f2_dinv_1_mul_U5 ( .A(Inst_f2_dinv_1_mul_n257), .B(
        Inst_f2_dinv_1_mul_n244), .ZN(Inst_f2_dinv_1_mul_n339) );
  NAND2_X1 Inst_f2_dinv_1_mul_U4 ( .A1(gamma1[2]), .A2(gamma0[2]), .ZN(
        Inst_f2_dinv_1_mul_n244) );
  NAND2_X1 Inst_f2_dinv_1_mul_U3 ( .A1(gamma0[3]), .A2(gamma1[3]), .ZN(
        Inst_f2_dinv_1_mul_n257) );
  AND2_X1 Inst_f2_dinv_1_mul_U2 ( .A1(gamma0[0]), .A2(Inst_f2_dinv_1_mul_n243), 
        .ZN(Inst_f2_dinv_1_mul_n329) );
  XOR2_X1 Inst_f2_dinv_1_mul_U1 ( .A(Inst_f2_dinv_1_mul_n325), .B(gamma1[3]), 
        .Z(Inst_f2_dinv_1_mul_n243) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_MaskXORInst_U2 ( .A(PRNGQ[13]), .B(
        PRNGQ[15]), .Z(Inst_f2_dinv_1_AddNewMaskab_MaskXOR[1]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_MaskXORInst_U1 ( .A(PRNGQ[12]), .B(
        PRNGQ[14]), .Z(Inst_f2_dinv_1_AddNewMaskab_MaskXOR[0]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_XORInst1_U2 ( .A(
        Inst_f2_dinv_1_Orig_ab[5]), .B(Inst_f2_dinv_1_AddNewMaskab_MaskXOR[1]), 
        .Z(ab[5]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_XORInst1_U1 ( .A(
        Inst_f2_dinv_1_Orig_ab[4]), .B(Inst_f2_dinv_1_AddNewMaskab_MaskXOR[0]), 
        .Z(ab[4]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_XORInst2_U4 ( .A(
        Inst_f2_dinv_1_Orig_ab[3]), .B(PRNGQ[15]), .Z(ab[3]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_XORInst2_U3 ( .A(
        Inst_f2_dinv_1_Orig_ab[2]), .B(PRNGQ[14]), .Z(ab[2]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_XORInst2_U2 ( .A(
        Inst_f2_dinv_1_Orig_ab[1]), .B(PRNGQ[13]), .Z(ab[1]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMaskab_XORInst2_U1 ( .A(
        Inst_f2_dinv_1_Orig_ab[0]), .B(PRNGQ[12]), .Z(ab[0]) );
  XOR2_X1 Inst_f2_dinv_1_NxGAMMA_U3 ( .A(Inst_f2_dinv_1_Orig_sA2N[5]), .B(
        Inst_f2_dinv_1_sA2[5]), .Z(Inst_f2_dinv_1_Orig_sA2N[4]) );
  XOR2_X1 Inst_f2_dinv_1_NxGAMMA_U2 ( .A(Inst_f2_dinv_1_Orig_sA2N[3]), .B(
        Inst_f2_dinv_1_sA2[3]), .Z(Inst_f2_dinv_1_Orig_sA2N[2]) );
  XOR2_X1 Inst_f2_dinv_1_NxGAMMA_U1 ( .A(Inst_f2_dinv_1_Orig_sA2N[1]), .B(
        Inst_f2_dinv_1_sA2[1]), .Z(Inst_f2_dinv_1_Orig_sA2N[0]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_MaskXORInst_U2 ( .A(PRNGQ[17]), .B(
        PRNGQ[19]), .Z(Inst_f2_dinv_1_AddNewMasksA2N_MaskXOR[1]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_MaskXORInst_U1 ( .A(PRNGQ[16]), .B(
        PRNGQ[18]), .Z(Inst_f2_dinv_1_AddNewMasksA2N_MaskXOR[0]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_XORInst1_U2 ( .A(
        Inst_f2_dinv_1_Orig_sA2N[5]), .B(
        Inst_f2_dinv_1_AddNewMasksA2N_MaskXOR[1]), .Z(sA2N[5]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_XORInst1_U1 ( .A(
        Inst_f2_dinv_1_Orig_sA2N[4]), .B(
        Inst_f2_dinv_1_AddNewMasksA2N_MaskXOR[0]), .Z(sA2N[4]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_XORInst2_U4 ( .A(
        Inst_f2_dinv_1_Orig_sA2N[3]), .B(PRNGQ[19]), .Z(sA2N[3]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_XORInst2_U3 ( .A(
        Inst_f2_dinv_1_Orig_sA2N[2]), .B(PRNGQ[18]), .Z(sA2N[2]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_XORInst2_U2 ( .A(
        Inst_f2_dinv_1_Orig_sA2N[1]), .B(PRNGQ[17]), .Z(sA2N[1]) );
  XOR2_X1 Inst_f2_dinv_1_AddNewMasksA2N_XORInst2_U1 ( .A(
        Inst_f2_dinv_1_Orig_sA2N[0]), .B(PRNGQ[16]), .Z(sA2N[0]) );
  DFF_X1 PL_2_s_current_state_reg_0_ ( .D(gamma0[0]), .CK(clk), .Q(FF2_out[0]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_1_ ( .D(gamma0[1]), .CK(clk), .Q(FF2_out[1]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_2_ ( .D(gamma0[2]), .CK(clk), .Q(FF2_out[2]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_3_ ( .D(gamma0[3]), .CK(clk), .Q(FF2_out[3]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_4_ ( .D(gamma0[4]), .CK(clk), .Q(FF2_out[4]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_5_ ( .D(gamma0[5]), .CK(clk), .Q(FF2_out[5]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_6_ ( .D(ab[0]), .CK(clk), .Q(FF2_out[6]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_7_ ( .D(ab[1]), .CK(clk), .Q(FF2_out[7]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_8_ ( .D(ab[2]), .CK(clk), .Q(FF2_out[8]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_9_ ( .D(ab[3]), .CK(clk), .Q(FF2_out[9]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_10_ ( .D(ab[4]), .CK(clk), .Q(FF2_out[10]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_11_ ( .D(ab[5]), .CK(clk), .Q(FF2_out[11]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_12_ ( .D(sA2N[0]), .CK(clk), .Q(FF2_out[12]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_13_ ( .D(sA2N[1]), .CK(clk), .Q(FF2_out[13]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_14_ ( .D(sA2N[2]), .CK(clk), .Q(FF2_out[14]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_15_ ( .D(sA2N[3]), .CK(clk), .Q(FF2_out[15]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_16_ ( .D(sA2N[4]), .CK(clk), .Q(FF2_out[16]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_17_ ( .D(sA2N[5]), .CK(clk), .Q(FF2_out[17]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_18_ ( .D(gamma1[0]), .CK(clk), .Q(
        FF2_out[18]), .QN() );
  DFF_X1 PL_2_s_current_state_reg_19_ ( .D(gamma1[1]), .CK(clk), .Q(
        FF2_out[19]), .QN() );
  DFF_X1 PL_2_s_current_state_reg_20_ ( .D(gamma1[2]), .CK(clk), .Q(
        FF2_out[20]), .QN() );
  DFF_X1 PL_2_s_current_state_reg_21_ ( .D(gamma1[3]), .CK(clk), .Q(
        FF2_out[21]), .QN() );
  DFF_X1 PL_2_s_current_state_reg_22_ ( .D(gamma1[4]), .CK(clk), .Q(
        FF2_out[22]), .QN() );
  DFF_X1 PL_2_s_current_state_reg_23_ ( .D(gamma1[5]), .CK(clk), .Q(
        FF2_out[23]), .QN() );
  DFF_X1 PL_2_s_current_state_reg_24_ ( .D(Zl_f2[0]), .CK(clk), .Q(Zl_f3[0]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_25_ ( .D(Zl_f2[1]), .CK(clk), .Q(Zl_f3[1]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_26_ ( .D(Zl_f2[2]), .CK(clk), .Q(Zl_f3[2]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_27_ ( .D(Zl_f2[3]), .CK(clk), .Q(Zl_f3[3]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_28_ ( .D(Zl_f2[4]), .CK(clk), .Q(Zl_f3[4]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_29_ ( .D(Zl_f2[5]), .CK(clk), .Q(Zl_f3[5]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_30_ ( .D(Zl_f2[6]), .CK(clk), .Q(Zl_f3[6]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_31_ ( .D(Zl_f2[7]), .CK(clk), .Q(Zl_f3[7]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_32_ ( .D(Zl_f2[8]), .CK(clk), .Q(Zl_f3[8]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_33_ ( .D(Zl_f2[9]), .CK(clk), .Q(Zl_f3[9]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_34_ ( .D(Zl_f2[10]), .CK(clk), .Q(Zl_f3[10]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_35_ ( .D(Zl_f2[11]), .CK(clk), .Q(Zl_f3[11]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_36_ ( .D(Zh_f2[0]), .CK(clk), .Q(Zh_f3[0]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_37_ ( .D(Zh_f2[1]), .CK(clk), .Q(Zh_f3[1]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_38_ ( .D(Zh_f2[2]), .CK(clk), .Q(Zh_f3[2]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_39_ ( .D(Zh_f2[3]), .CK(clk), .Q(Zh_f3[3]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_40_ ( .D(Zh_f2[4]), .CK(clk), .Q(Zh_f3[4]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_41_ ( .D(Zh_f2[5]), .CK(clk), .Q(Zh_f3[5]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_42_ ( .D(Zh_f2[6]), .CK(clk), .Q(Zh_f3[6]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_43_ ( .D(Zh_f2[7]), .CK(clk), .Q(Zh_f3[7]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_44_ ( .D(Zh_f2[8]), .CK(clk), .Q(Zh_f3[8]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_45_ ( .D(Zh_f2[9]), .CK(clk), .Q(Zh_f3[9]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_46_ ( .D(Zh_f2[10]), .CK(clk), .Q(Zh_f3[10]), 
        .QN() );
  DFF_X1 PL_2_s_current_state_reg_47_ ( .D(Zh_f2[11]), .CK(clk), .Q(Zh_f3[11]), 
        .QN() );
  XOR2_X2 Inst_f3_dinv_2_U6 ( .A(FF2_out[11]), .B(FF2_out[17]), .Z(
        Inst_f3_dinv_2_d_4_) );
  XOR2_X2 Inst_f3_dinv_2_U5 ( .A(FF2_out[7]), .B(FF2_out[13]), .Z(
        Inst_f3_dinv_2_d_0_) );
  XOR2_X2 Inst_f3_dinv_2_U4 ( .A(FF2_out[6]), .B(FF2_out[12]), .Z(
        Inst_f3_dinv_2_d_1_) );
  XOR2_X2 Inst_f3_dinv_2_U3 ( .A(FF2_out[10]), .B(FF2_out[16]), .Z(
        Inst_f3_dinv_2_d_5_) );
  XOR2_X2 Inst_f3_dinv_2_U2 ( .A(FF2_out[9]), .B(FF2_out[15]), .Z(
        Inst_f3_dinv_2_d_2_) );
  XOR2_X2 Inst_f3_dinv_2_U1 ( .A(FF2_out[8]), .B(FF2_out[14]), .Z(
        Inst_f3_dinv_2_d_3_) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U104 ( .A(Inst_f3_dinv_2_himul_n337), .B(
        Inst_f3_dinv_2_himul_n336), .ZN(Inst_f3_dinv_2_pl[4]) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U103 ( .A(Inst_f3_dinv_2_himul_n335), .B(
        Inst_f3_dinv_2_himul_n334), .ZN(Inst_f3_dinv_2_himul_n336) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U102 ( .A(Inst_f3_dinv_2_himul_n333), .B(
        Inst_f3_dinv_2_himul_n332), .ZN(Inst_f3_dinv_2_himul_n334) );
  NAND2_X1 Inst_f3_dinv_2_himul_U101 ( .A1(Inst_f3_dinv_2_himul_n331), .A2(
        FF2_out[20]), .ZN(Inst_f3_dinv_2_himul_n333) );
  NAND2_X1 Inst_f3_dinv_2_himul_U100 ( .A1(Inst_f3_dinv_2_himul_n330), .A2(
        Inst_f3_dinv_2_himul_n329), .ZN(Inst_f3_dinv_2_himul_n335) );
  NAND2_X1 Inst_f3_dinv_2_himul_U99 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        Inst_f3_dinv_2_himul_n328), .ZN(Inst_f3_dinv_2_himul_n329) );
  OR2_X1 Inst_f3_dinv_2_himul_U98 ( .A1(Inst_f3_dinv_2_himul_n328), .A2(
        Inst_f3_dinv_2_himul_n338), .ZN(Inst_f3_dinv_2_himul_n330) );
  XOR2_X1 Inst_f3_dinv_2_himul_U97 ( .A(FF2_out[19]), .B(
        Inst_f3_dinv_2_himul_n327), .Z(Inst_f3_dinv_2_himul_n328) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U96 ( .A(Inst_f3_dinv_2_himul_n326), .B(
        Inst_f3_dinv_2_himul_n340), .ZN(Inst_f3_dinv_2_himul_n337) );
  XOR2_X1 Inst_f3_dinv_2_himul_U95 ( .A(Inst_f3_dinv_2_himul_n325), .B(
        Inst_f3_dinv_2_himul_n324), .Z(Inst_f3_dinv_2_himul_n340) );
  NAND2_X1 Inst_f3_dinv_2_himul_U94 ( .A1(Inst_f3_dinv_2_d_2_), .A2(
        FF2_out[19]), .ZN(Inst_f3_dinv_2_himul_n324) );
  NOR2_X1 Inst_f3_dinv_2_himul_U93 ( .A1(Inst_f3_dinv_2_himul_n323), .A2(
        Inst_f3_dinv_2_himul_n338), .ZN(Inst_f3_dinv_2_himul_n325) );
  INV_X1 Inst_f3_dinv_2_himul_U92 ( .A(Inst_f3_dinv_2_d_1_), .ZN(
        Inst_f3_dinv_2_himul_n338) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U91 ( .A(FF2_out[18]), .B(FF2_out[20]), .ZN(
        Inst_f3_dinv_2_himul_n323) );
  NAND2_X1 Inst_f3_dinv_2_himul_U90 ( .A1(Inst_f3_dinv_2_himul_n322), .A2(
        Inst_f3_dinv_2_himul_n321), .ZN(Inst_f3_dinv_2_himul_n326) );
  NAND2_X1 Inst_f3_dinv_2_himul_U89 ( .A1(FF2_out[19]), .A2(
        Inst_f3_dinv_2_himul_n320), .ZN(Inst_f3_dinv_2_himul_n321) );
  NAND2_X1 Inst_f3_dinv_2_himul_U88 ( .A1(FF2_out[18]), .A2(
        Inst_f3_dinv_2_d_3_), .ZN(Inst_f3_dinv_2_himul_n322) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U87 ( .A(Inst_f3_dinv_2_himul_n319), .B(
        Inst_f3_dinv_2_himul_n318), .ZN(Inst_f3_dinv_2_pl[3]) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U86 ( .A(Inst_f3_dinv_2_himul_n317), .B(
        Inst_f3_dinv_2_himul_n316), .ZN(Inst_f3_dinv_2_himul_n318) );
  XOR2_X1 Inst_f3_dinv_2_himul_U85 ( .A(Inst_f3_dinv_2_himul_n315), .B(
        Inst_f3_dinv_2_himul_n314), .Z(Inst_f3_dinv_2_himul_n317) );
  NAND2_X1 Inst_f3_dinv_2_himul_U84 ( .A1(FF2_out[22]), .A2(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_himul_n314) );
  NAND2_X1 Inst_f3_dinv_2_himul_U83 ( .A1(FF2_out[23]), .A2(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n315) );
  XOR2_X1 Inst_f3_dinv_2_himul_U82 ( .A(Inst_f3_dinv_2_himul_n313), .B(
        Inst_f3_dinv_2_himul_n312), .Z(Inst_f3_dinv_2_himul_n319) );
  XOR2_X1 Inst_f3_dinv_2_himul_U81 ( .A(Inst_f3_dinv_2_himul_n311), .B(
        Inst_f3_dinv_2_himul_n310), .Z(Inst_f3_dinv_2_himul_n312) );
  NAND2_X1 Inst_f3_dinv_2_himul_U80 ( .A1(FF2_out[22]), .A2(
        Inst_f3_dinv_2_himul_n309), .ZN(Inst_f3_dinv_2_himul_n310) );
  NAND2_X1 Inst_f3_dinv_2_himul_U79 ( .A1(FF2_out[18]), .A2(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n311) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U78 ( .A(Inst_f3_dinv_2_himul_n308), .B(
        Inst_f3_dinv_2_himul_n307), .ZN(Inst_f3_dinv_2_himul_n313) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U77 ( .A(FF2_out[23]), .B(
        Inst_f3_dinv_2_himul_n306), .ZN(Inst_f3_dinv_2_himul_n307) );
  XOR2_X1 Inst_f3_dinv_2_himul_U76 ( .A(Inst_f3_dinv_2_himul_n305), .B(
        Inst_f3_dinv_2_himul_n304), .Z(Inst_f3_dinv_2_himul_n306) );
  NAND2_X1 Inst_f3_dinv_2_himul_U75 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        FF2_out[22]), .ZN(Inst_f3_dinv_2_himul_n304) );
  NOR2_X1 Inst_f3_dinv_2_himul_U74 ( .A1(Inst_f3_dinv_2_himul_n303), .A2(
        Inst_f3_dinv_2_d_1_), .ZN(Inst_f3_dinv_2_himul_n305) );
  NAND2_X1 Inst_f3_dinv_2_himul_U73 ( .A1(Inst_f3_dinv_2_himul_n302), .A2(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_himul_n308) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U72 ( .A(Inst_f3_dinv_2_himul_n339), .B(
        Inst_f3_dinv_2_himul_n301), .ZN(Inst_f3_dinv_2_himul_n302) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U71 ( .A(FF2_out[19]), .B(
        Inst_f3_dinv_2_himul_n300), .ZN(Inst_f3_dinv_2_himul_n301) );
  INV_X1 Inst_f3_dinv_2_himul_U70 ( .A(FF2_out[18]), .ZN(
        Inst_f3_dinv_2_himul_n339) );
  XOR2_X1 Inst_f3_dinv_2_himul_U69 ( .A(Inst_f3_dinv_2_himul_n299), .B(
        Inst_f3_dinv_2_himul_n298), .Z(Inst_f3_dinv_2_pl[2]) );
  NAND2_X1 Inst_f3_dinv_2_himul_U68 ( .A1(Inst_f3_dinv_2_himul_n297), .A2(
        Inst_f3_dinv_2_himul_n296), .ZN(Inst_f3_dinv_2_himul_n298) );
  OR2_X1 Inst_f3_dinv_2_himul_U67 ( .A1(Inst_f3_dinv_2_d_5_), .A2(
        Inst_f3_dinv_2_himul_n303), .ZN(Inst_f3_dinv_2_himul_n296) );
  NAND2_X1 Inst_f3_dinv_2_himul_U66 ( .A1(Inst_f3_dinv_2_himul_n295), .A2(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n297) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U65 ( .A(Inst_f3_dinv_2_himul_n294), .B(
        FF2_out[18]), .ZN(Inst_f3_dinv_2_himul_n295) );
  XOR2_X1 Inst_f3_dinv_2_himul_U64 ( .A(Inst_f3_dinv_2_himul_n293), .B(
        Inst_f3_dinv_2_himul_n292), .Z(Inst_f3_dinv_2_himul_n299) );
  NOR2_X1 Inst_f3_dinv_2_himul_U63 ( .A1(Inst_f3_dinv_2_himul_n300), .A2(
        Inst_f3_dinv_2_himul_n291), .ZN(Inst_f3_dinv_2_himul_n292) );
  XOR2_X1 Inst_f3_dinv_2_himul_U62 ( .A(Inst_f3_dinv_2_himul_n309), .B(
        Inst_f3_dinv_2_d_1_), .Z(Inst_f3_dinv_2_himul_n291) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U61 ( .A(Inst_f3_dinv_2_himul_n290), .B(
        Inst_f3_dinv_2_himul_n289), .ZN(Inst_f3_dinv_2_himul_n293) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U60 ( .A(Inst_f3_dinv_2_d_0_), .B(
        Inst_f3_dinv_2_himul_n332), .ZN(Inst_f3_dinv_2_himul_n289) );
  XOR2_X1 Inst_f3_dinv_2_himul_U59 ( .A(Inst_f3_dinv_2_himul_n288), .B(
        Inst_f3_dinv_2_himul_n287), .Z(Inst_f3_dinv_2_himul_n332) );
  NAND2_X1 Inst_f3_dinv_2_himul_U58 ( .A1(FF2_out[19]), .A2(
        Inst_f3_dinv_2_d_0_), .ZN(Inst_f3_dinv_2_himul_n287) );
  NAND2_X1 Inst_f3_dinv_2_himul_U57 ( .A1(FF2_out[18]), .A2(
        Inst_f3_dinv_2_d_1_), .ZN(Inst_f3_dinv_2_himul_n288) );
  XOR2_X1 Inst_f3_dinv_2_himul_U56 ( .A(Inst_f3_dinv_2_himul_n286), .B(
        Inst_f3_dinv_2_himul_n316), .Z(Inst_f3_dinv_2_himul_n290) );
  XOR2_X1 Inst_f3_dinv_2_himul_U55 ( .A(Inst_f3_dinv_2_himul_n285), .B(
        Inst_f3_dinv_2_himul_n284), .Z(Inst_f3_dinv_2_himul_n316) );
  NAND2_X1 Inst_f3_dinv_2_himul_U54 ( .A1(FF2_out[22]), .A2(
        Inst_f3_dinv_2_d_1_), .ZN(Inst_f3_dinv_2_himul_n284) );
  NAND2_X1 Inst_f3_dinv_2_himul_U53 ( .A1(FF2_out[23]), .A2(
        Inst_f3_dinv_2_d_0_), .ZN(Inst_f3_dinv_2_himul_n285) );
  XOR2_X1 Inst_f3_dinv_2_himul_U52 ( .A(Inst_f3_dinv_2_himul_n283), .B(
        Inst_f3_dinv_2_himul_n282), .Z(Inst_f3_dinv_2_himul_n286) );
  NAND2_X1 Inst_f3_dinv_2_himul_U51 ( .A1(Inst_f3_dinv_2_d_4_), .A2(
        Inst_f3_dinv_2_himul_n303), .ZN(Inst_f3_dinv_2_himul_n282) );
  INV_X1 Inst_f3_dinv_2_himul_U50 ( .A(FF2_out[19]), .ZN(
        Inst_f3_dinv_2_himul_n303) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U49 ( .A(Inst_f3_dinv_2_himul_n281), .B(
        Inst_f3_dinv_2_himul_n280), .ZN(Inst_f3_dinv_2_pl[1]) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U48 ( .A(Inst_f3_dinv_2_himul_n279), .B(
        Inst_f3_dinv_2_himul_n278), .ZN(Inst_f3_dinv_2_himul_n281) );
  NAND2_X1 Inst_f3_dinv_2_himul_U47 ( .A1(Inst_f3_dinv_2_himul_n277), .A2(
        FF2_out[20]), .ZN(Inst_f3_dinv_2_himul_n278) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U46 ( .A(Inst_f3_dinv_2_d_2_), .B(
        Inst_f3_dinv_2_himul_n309), .ZN(Inst_f3_dinv_2_himul_n277) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U45 ( .A(Inst_f3_dinv_2_himul_n276), .B(
        Inst_f3_dinv_2_himul_n275), .ZN(Inst_f3_dinv_2_himul_n279) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U44 ( .A(Inst_f3_dinv_2_himul_n274), .B(
        Inst_f3_dinv_2_himul_n273), .ZN(Inst_f3_dinv_2_himul_n275) );
  NAND2_X1 Inst_f3_dinv_2_himul_U43 ( .A1(Inst_f3_dinv_2_himul_n272), .A2(
        Inst_f3_dinv_2_himul_n331), .ZN(Inst_f3_dinv_2_himul_n273) );
  XOR2_X1 Inst_f3_dinv_2_himul_U42 ( .A(Inst_f3_dinv_2_d_2_), .B(
        Inst_f3_dinv_2_d_3_), .Z(Inst_f3_dinv_2_himul_n331) );
  XOR2_X1 Inst_f3_dinv_2_himul_U41 ( .A(FF2_out[20]), .B(FF2_out[22]), .Z(
        Inst_f3_dinv_2_himul_n272) );
  NAND2_X1 Inst_f3_dinv_2_himul_U40 ( .A1(FF2_out[21]), .A2(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_himul_n274) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U39 ( .A(Inst_f3_dinv_2_himul_n271), .B(
        Inst_f3_dinv_2_himul_n270), .ZN(Inst_f3_dinv_2_himul_n276) );
  XOR2_X1 Inst_f3_dinv_2_himul_U38 ( .A(Inst_f3_dinv_2_himul_n269), .B(
        Inst_f3_dinv_2_himul_n268), .Z(Inst_f3_dinv_2_himul_n271) );
  NOR2_X1 Inst_f3_dinv_2_himul_U37 ( .A1(Inst_f3_dinv_2_himul_n294), .A2(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_himul_n268) );
  INV_X1 Inst_f3_dinv_2_himul_U36 ( .A(FF2_out[22]), .ZN(
        Inst_f3_dinv_2_himul_n294) );
  NOR2_X1 Inst_f3_dinv_2_himul_U35 ( .A1(Inst_f3_dinv_2_himul_n300), .A2(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n269) );
  INV_X1 Inst_f3_dinv_2_himul_U34 ( .A(FF2_out[23]), .ZN(
        Inst_f3_dinv_2_himul_n300) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U33 ( .A(Inst_f3_dinv_2_himul_n267), .B(
        Inst_f3_dinv_2_himul_n266), .ZN(Inst_f3_dinv_2_pl[0]) );
  NAND2_X1 Inst_f3_dinv_2_himul_U32 ( .A1(FF2_out[20]), .A2(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n266) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U31 ( .A(Inst_f3_dinv_2_himul_n341), .B(
        Inst_f3_dinv_2_himul_n265), .ZN(Inst_f3_dinv_2_himul_n267) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U30 ( .A(Inst_f3_dinv_2_himul_n264), .B(
        Inst_f3_dinv_2_himul_n263), .ZN(Inst_f3_dinv_2_himul_n265) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U29 ( .A(Inst_f3_dinv_2_himul_n262), .B(
        Inst_f3_dinv_2_himul_n261), .ZN(Inst_f3_dinv_2_himul_n263) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U28 ( .A(Inst_f3_dinv_2_himul_n260), .B(
        Inst_f3_dinv_2_himul_n280), .ZN(Inst_f3_dinv_2_himul_n261) );
  NAND2_X1 Inst_f3_dinv_2_himul_U27 ( .A1(Inst_f3_dinv_2_d_2_), .A2(
        Inst_f3_dinv_2_himul_n259), .ZN(Inst_f3_dinv_2_himul_n280) );
  XOR2_X1 Inst_f3_dinv_2_himul_U26 ( .A(FF2_out[21]), .B(FF2_out[23]), .Z(
        Inst_f3_dinv_2_himul_n259) );
  NOR2_X1 Inst_f3_dinv_2_himul_U25 ( .A1(Inst_f3_dinv_2_himul_n258), .A2(
        Inst_f3_dinv_2_himul_n320), .ZN(Inst_f3_dinv_2_himul_n260) );
  INV_X1 Inst_f3_dinv_2_himul_U24 ( .A(Inst_f3_dinv_2_d_3_), .ZN(
        Inst_f3_dinv_2_himul_n320) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U23 ( .A(FF2_out[23]), .B(FF2_out[22]), .ZN(
        Inst_f3_dinv_2_himul_n258) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U22 ( .A(Inst_f3_dinv_2_himul_n283), .B(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_himul_n262) );
  NAND2_X1 Inst_f3_dinv_2_himul_U21 ( .A1(FF2_out[22]), .A2(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n283) );
  NOR2_X1 Inst_f3_dinv_2_himul_U20 ( .A1(Inst_f3_dinv_2_himul_n327), .A2(
        Inst_f3_dinv_2_himul_n309), .ZN(Inst_f3_dinv_2_himul_n264) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U19 ( .A(Inst_f3_dinv_2_d_4_), .B(
        Inst_f3_dinv_2_d_5_), .ZN(Inst_f3_dinv_2_himul_n309) );
  INV_X1 Inst_f3_dinv_2_himul_U18 ( .A(FF2_out[21]), .ZN(
        Inst_f3_dinv_2_himul_n327) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U17 ( .A(Inst_f3_dinv_2_himul_n270), .B(
        Inst_f3_dinv_2_himul_n257), .ZN(Inst_f3_dinv_2_himul_n341) );
  NAND2_X1 Inst_f3_dinv_2_himul_U16 ( .A1(FF2_out[20]), .A2(
        Inst_f3_dinv_2_d_2_), .ZN(Inst_f3_dinv_2_himul_n257) );
  NAND2_X1 Inst_f3_dinv_2_himul_U15 ( .A1(Inst_f3_dinv_2_d_3_), .A2(
        FF2_out[21]), .ZN(Inst_f3_dinv_2_himul_n270) );
  XOR2_X1 Inst_f3_dinv_2_himul_U14 ( .A(Inst_f3_dinv_2_himul_n256), .B(
        Inst_f3_dinv_2_himul_n341), .Z(Inst_f3_dinv_2_pl[5]) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U13 ( .A(Inst_f3_dinv_2_himul_n255), .B(
        Inst_f3_dinv_2_himul_n253), .ZN(Inst_f3_dinv_2_himul_n256) );
  NAND2_X1 Inst_f3_dinv_2_himul_U12 ( .A1(Inst_f3_dinv_2_himul_n254), .A2(
        Inst_f3_dinv_2_himul_n250), .ZN(Inst_f3_dinv_2_himul_n255) );
  NAND2_X1 Inst_f3_dinv_2_himul_U11 ( .A1(Inst_f3_dinv_2_himul_n244), .A2(
        Inst_f3_dinv_2_d_1_), .ZN(Inst_f3_dinv_2_himul_n254) );
  XOR2_X1 Inst_f3_dinv_2_himul_U10 ( .A(Inst_f3_dinv_2_himul_n252), .B(
        Inst_f3_dinv_2_himul_n340), .Z(Inst_f3_dinv_2_himul_n253) );
  NOR2_X1 Inst_f3_dinv_2_himul_U9 ( .A1(Inst_f3_dinv_2_himul_n339), .A2(
        Inst_f3_dinv_2_himul_n251), .ZN(Inst_f3_dinv_2_himul_n252) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U8 ( .A(Inst_f3_dinv_2_d_3_), .B(
        Inst_f3_dinv_2_d_2_), .ZN(Inst_f3_dinv_2_himul_n251) );
  XOR2_X1 Inst_f3_dinv_2_himul_U7 ( .A(Inst_f3_dinv_2_himul_n247), .B(
        Inst_f3_dinv_2_himul_n249), .Z(Inst_f3_dinv_2_himul_n250) );
  NAND2_X1 Inst_f3_dinv_2_himul_U6 ( .A1(Inst_f3_dinv_2_himul_n248), .A2(
        FF2_out[19]), .ZN(Inst_f3_dinv_2_himul_n249) );
  NAND2_X1 Inst_f3_dinv_2_himul_U5 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        Inst_f3_dinv_2_himul_n338), .ZN(Inst_f3_dinv_2_himul_n248) );
  NAND2_X1 Inst_f3_dinv_2_himul_U4 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        Inst_f3_dinv_2_himul_n246), .ZN(Inst_f3_dinv_2_himul_n247) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U3 ( .A(Inst_f3_dinv_2_himul_n245), .B(
        FF2_out[20]), .ZN(Inst_f3_dinv_2_himul_n246) );
  XNOR2_X1 Inst_f3_dinv_2_himul_U2 ( .A(FF2_out[18]), .B(FF2_out[21]), .ZN(
        Inst_f3_dinv_2_himul_n245) );
  INV_X1 Inst_f3_dinv_2_himul_U1 ( .A(Inst_f3_dinv_2_d_0_), .ZN(
        Inst_f3_dinv_2_himul_n244) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U104 ( .A(Inst_f3_dinv_2_lowmul_n336), .B(
        Inst_f3_dinv_2_lowmul_n335), .ZN(Inst_f3_dinv_2_ph[4]) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U103 ( .A(Inst_f3_dinv_2_lowmul_n334), .B(
        Inst_f3_dinv_2_lowmul_n333), .ZN(Inst_f3_dinv_2_lowmul_n335) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U102 ( .A(Inst_f3_dinv_2_lowmul_n332), .B(
        Inst_f3_dinv_2_lowmul_n331), .ZN(Inst_f3_dinv_2_lowmul_n333) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U101 ( .A1(Inst_f3_dinv_2_lowmul_n330), .A2(
        Inst_f3_dinv_2_d_2_), .ZN(Inst_f3_dinv_2_lowmul_n332) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U100 ( .A1(Inst_f3_dinv_2_lowmul_n329), .A2(
        Inst_f3_dinv_2_lowmul_n328), .ZN(Inst_f3_dinv_2_lowmul_n334) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U99 ( .A1(FF2_out[0]), .A2(
        Inst_f3_dinv_2_lowmul_n327), .ZN(Inst_f3_dinv_2_lowmul_n328) );
  OR2_X1 Inst_f3_dinv_2_lowmul_U98 ( .A1(Inst_f3_dinv_2_lowmul_n327), .A2(
        Inst_f3_dinv_2_lowmul_n337), .ZN(Inst_f3_dinv_2_lowmul_n329) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U97 ( .A(Inst_f3_dinv_2_d_1_), .B(
        Inst_f3_dinv_2_lowmul_n326), .Z(Inst_f3_dinv_2_lowmul_n327) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U96 ( .A(Inst_f3_dinv_2_lowmul_n325), .B(
        Inst_f3_dinv_2_lowmul_n339), .ZN(Inst_f3_dinv_2_lowmul_n336) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U95 ( .A(Inst_f3_dinv_2_lowmul_n324), .B(
        Inst_f3_dinv_2_lowmul_n323), .Z(Inst_f3_dinv_2_lowmul_n339) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U94 ( .A1(FF2_out[2]), .A2(
        Inst_f3_dinv_2_d_1_), .ZN(Inst_f3_dinv_2_lowmul_n323) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U93 ( .A1(Inst_f3_dinv_2_lowmul_n322), .A2(
        Inst_f3_dinv_2_lowmul_n337), .ZN(Inst_f3_dinv_2_lowmul_n324) );
  INV_X1 Inst_f3_dinv_2_lowmul_U92 ( .A(FF2_out[1]), .ZN(
        Inst_f3_dinv_2_lowmul_n337) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U91 ( .A(Inst_f3_dinv_2_d_0_), .B(
        Inst_f3_dinv_2_d_2_), .ZN(Inst_f3_dinv_2_lowmul_n322) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U90 ( .A1(Inst_f3_dinv_2_lowmul_n321), .A2(
        Inst_f3_dinv_2_lowmul_n320), .ZN(Inst_f3_dinv_2_lowmul_n325) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U89 ( .A1(Inst_f3_dinv_2_d_1_), .A2(
        Inst_f3_dinv_2_lowmul_n319), .ZN(Inst_f3_dinv_2_lowmul_n320) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U88 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        FF2_out[3]), .ZN(Inst_f3_dinv_2_lowmul_n321) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U87 ( .A(Inst_f3_dinv_2_lowmul_n318), .B(
        Inst_f3_dinv_2_lowmul_n317), .ZN(Inst_f3_dinv_2_ph[3]) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U86 ( .A(Inst_f3_dinv_2_lowmul_n316), .B(
        Inst_f3_dinv_2_lowmul_n315), .ZN(Inst_f3_dinv_2_lowmul_n317) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U85 ( .A(Inst_f3_dinv_2_lowmul_n314), .B(
        Inst_f3_dinv_2_lowmul_n313), .Z(Inst_f3_dinv_2_lowmul_n316) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U84 ( .A1(Inst_f3_dinv_2_d_4_), .A2(
        FF2_out[4]), .ZN(Inst_f3_dinv_2_lowmul_n313) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U83 ( .A1(Inst_f3_dinv_2_d_5_), .A2(
        FF2_out[5]), .ZN(Inst_f3_dinv_2_lowmul_n314) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U82 ( .A(Inst_f3_dinv_2_lowmul_n312), .B(
        Inst_f3_dinv_2_lowmul_n311), .Z(Inst_f3_dinv_2_lowmul_n318) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U81 ( .A(Inst_f3_dinv_2_lowmul_n310), .B(
        Inst_f3_dinv_2_lowmul_n309), .Z(Inst_f3_dinv_2_lowmul_n311) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U80 ( .A1(Inst_f3_dinv_2_d_4_), .A2(
        Inst_f3_dinv_2_lowmul_n308), .ZN(Inst_f3_dinv_2_lowmul_n309) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U79 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        FF2_out[5]), .ZN(Inst_f3_dinv_2_lowmul_n310) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U78 ( .A(Inst_f3_dinv_2_lowmul_n307), .B(
        Inst_f3_dinv_2_lowmul_n306), .ZN(Inst_f3_dinv_2_lowmul_n312) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U77 ( .A(Inst_f3_dinv_2_d_5_), .B(
        Inst_f3_dinv_2_lowmul_n305), .ZN(Inst_f3_dinv_2_lowmul_n306) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U76 ( .A(Inst_f3_dinv_2_lowmul_n304), .B(
        Inst_f3_dinv_2_lowmul_n303), .Z(Inst_f3_dinv_2_lowmul_n305) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U75 ( .A1(FF2_out[0]), .A2(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_lowmul_n303) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U74 ( .A1(Inst_f3_dinv_2_lowmul_n302), .A2(
        FF2_out[1]), .ZN(Inst_f3_dinv_2_lowmul_n304) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U73 ( .A1(Inst_f3_dinv_2_lowmul_n301), .A2(
        FF2_out[4]), .ZN(Inst_f3_dinv_2_lowmul_n307) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U72 ( .A(Inst_f3_dinv_2_lowmul_n338), .B(
        Inst_f3_dinv_2_lowmul_n300), .ZN(Inst_f3_dinv_2_lowmul_n301) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U71 ( .A(Inst_f3_dinv_2_d_1_), .B(
        Inst_f3_dinv_2_lowmul_n299), .ZN(Inst_f3_dinv_2_lowmul_n300) );
  INV_X1 Inst_f3_dinv_2_lowmul_U70 ( .A(Inst_f3_dinv_2_d_0_), .ZN(
        Inst_f3_dinv_2_lowmul_n338) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U69 ( .A(Inst_f3_dinv_2_lowmul_n298), .B(
        Inst_f3_dinv_2_lowmul_n297), .Z(Inst_f3_dinv_2_ph[2]) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U68 ( .A1(Inst_f3_dinv_2_lowmul_n296), .A2(
        Inst_f3_dinv_2_lowmul_n295), .ZN(Inst_f3_dinv_2_lowmul_n297) );
  OR2_X1 Inst_f3_dinv_2_lowmul_U67 ( .A1(FF2_out[5]), .A2(
        Inst_f3_dinv_2_lowmul_n302), .ZN(Inst_f3_dinv_2_lowmul_n295) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U66 ( .A1(Inst_f3_dinv_2_lowmul_n294), .A2(
        FF2_out[5]), .ZN(Inst_f3_dinv_2_lowmul_n296) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U65 ( .A(Inst_f3_dinv_2_lowmul_n293), .B(
        Inst_f3_dinv_2_d_0_), .ZN(Inst_f3_dinv_2_lowmul_n294) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U64 ( .A(Inst_f3_dinv_2_lowmul_n292), .B(
        Inst_f3_dinv_2_lowmul_n291), .Z(Inst_f3_dinv_2_lowmul_n298) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U63 ( .A1(Inst_f3_dinv_2_lowmul_n299), .A2(
        Inst_f3_dinv_2_lowmul_n290), .ZN(Inst_f3_dinv_2_lowmul_n291) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U62 ( .A(Inst_f3_dinv_2_lowmul_n308), .B(
        FF2_out[1]), .Z(Inst_f3_dinv_2_lowmul_n290) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U61 ( .A(Inst_f3_dinv_2_lowmul_n289), .B(
        Inst_f3_dinv_2_lowmul_n288), .ZN(Inst_f3_dinv_2_lowmul_n292) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U60 ( .A(FF2_out[0]), .B(
        Inst_f3_dinv_2_lowmul_n331), .ZN(Inst_f3_dinv_2_lowmul_n288) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U59 ( .A(Inst_f3_dinv_2_lowmul_n287), .B(
        Inst_f3_dinv_2_lowmul_n286), .Z(Inst_f3_dinv_2_lowmul_n331) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U58 ( .A1(Inst_f3_dinv_2_d_1_), .A2(
        FF2_out[0]), .ZN(Inst_f3_dinv_2_lowmul_n286) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U57 ( .A1(Inst_f3_dinv_2_d_0_), .A2(
        FF2_out[1]), .ZN(Inst_f3_dinv_2_lowmul_n287) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U56 ( .A(Inst_f3_dinv_2_lowmul_n285), .B(
        Inst_f3_dinv_2_lowmul_n315), .Z(Inst_f3_dinv_2_lowmul_n289) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U55 ( .A(Inst_f3_dinv_2_lowmul_n284), .B(
        Inst_f3_dinv_2_lowmul_n283), .Z(Inst_f3_dinv_2_lowmul_n315) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U54 ( .A1(Inst_f3_dinv_2_d_4_), .A2(
        FF2_out[1]), .ZN(Inst_f3_dinv_2_lowmul_n283) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U53 ( .A1(Inst_f3_dinv_2_d_5_), .A2(
        FF2_out[0]), .ZN(Inst_f3_dinv_2_lowmul_n284) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U52 ( .A(Inst_f3_dinv_2_lowmul_n282), .B(
        Inst_f3_dinv_2_lowmul_n281), .Z(Inst_f3_dinv_2_lowmul_n285) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U51 ( .A1(FF2_out[4]), .A2(
        Inst_f3_dinv_2_lowmul_n302), .ZN(Inst_f3_dinv_2_lowmul_n281) );
  INV_X1 Inst_f3_dinv_2_lowmul_U50 ( .A(Inst_f3_dinv_2_d_1_), .ZN(
        Inst_f3_dinv_2_lowmul_n302) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U49 ( .A(Inst_f3_dinv_2_lowmul_n280), .B(
        Inst_f3_dinv_2_lowmul_n279), .ZN(Inst_f3_dinv_2_ph[1]) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U48 ( .A(Inst_f3_dinv_2_lowmul_n278), .B(
        Inst_f3_dinv_2_lowmul_n277), .ZN(Inst_f3_dinv_2_lowmul_n280) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U47 ( .A1(Inst_f3_dinv_2_lowmul_n276), .A2(
        Inst_f3_dinv_2_d_2_), .ZN(Inst_f3_dinv_2_lowmul_n277) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U46 ( .A(FF2_out[2]), .B(
        Inst_f3_dinv_2_lowmul_n308), .ZN(Inst_f3_dinv_2_lowmul_n276) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U45 ( .A(Inst_f3_dinv_2_lowmul_n275), .B(
        Inst_f3_dinv_2_lowmul_n274), .ZN(Inst_f3_dinv_2_lowmul_n278) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U44 ( .A(Inst_f3_dinv_2_lowmul_n273), .B(
        Inst_f3_dinv_2_lowmul_n272), .ZN(Inst_f3_dinv_2_lowmul_n274) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U43 ( .A1(Inst_f3_dinv_2_lowmul_n271), .A2(
        Inst_f3_dinv_2_lowmul_n330), .ZN(Inst_f3_dinv_2_lowmul_n272) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U42 ( .A(FF2_out[2]), .B(FF2_out[3]), .Z(
        Inst_f3_dinv_2_lowmul_n330) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U41 ( .A(Inst_f3_dinv_2_d_2_), .B(
        Inst_f3_dinv_2_d_4_), .Z(Inst_f3_dinv_2_lowmul_n271) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U40 ( .A1(Inst_f3_dinv_2_d_3_), .A2(
        FF2_out[4]), .ZN(Inst_f3_dinv_2_lowmul_n273) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U39 ( .A(Inst_f3_dinv_2_lowmul_n270), .B(
        Inst_f3_dinv_2_lowmul_n269), .ZN(Inst_f3_dinv_2_lowmul_n275) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U38 ( .A(Inst_f3_dinv_2_lowmul_n268), .B(
        Inst_f3_dinv_2_lowmul_n267), .Z(Inst_f3_dinv_2_lowmul_n270) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U37 ( .A1(Inst_f3_dinv_2_lowmul_n293), .A2(
        FF2_out[4]), .ZN(Inst_f3_dinv_2_lowmul_n267) );
  INV_X1 Inst_f3_dinv_2_lowmul_U36 ( .A(Inst_f3_dinv_2_d_4_), .ZN(
        Inst_f3_dinv_2_lowmul_n293) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U35 ( .A1(Inst_f3_dinv_2_lowmul_n299), .A2(
        FF2_out[5]), .ZN(Inst_f3_dinv_2_lowmul_n268) );
  INV_X1 Inst_f3_dinv_2_lowmul_U34 ( .A(Inst_f3_dinv_2_d_5_), .ZN(
        Inst_f3_dinv_2_lowmul_n299) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U33 ( .A(Inst_f3_dinv_2_lowmul_n266), .B(
        Inst_f3_dinv_2_lowmul_n265), .ZN(Inst_f3_dinv_2_ph[0]) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U32 ( .A1(Inst_f3_dinv_2_d_2_), .A2(
        FF2_out[5]), .ZN(Inst_f3_dinv_2_lowmul_n265) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U31 ( .A(Inst_f3_dinv_2_lowmul_n340), .B(
        Inst_f3_dinv_2_lowmul_n264), .ZN(Inst_f3_dinv_2_lowmul_n266) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U30 ( .A(Inst_f3_dinv_2_lowmul_n263), .B(
        Inst_f3_dinv_2_lowmul_n262), .ZN(Inst_f3_dinv_2_lowmul_n264) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U29 ( .A(Inst_f3_dinv_2_lowmul_n261), .B(
        Inst_f3_dinv_2_lowmul_n260), .ZN(Inst_f3_dinv_2_lowmul_n262) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U28 ( .A(Inst_f3_dinv_2_lowmul_n259), .B(
        Inst_f3_dinv_2_lowmul_n279), .ZN(Inst_f3_dinv_2_lowmul_n260) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U27 ( .A1(FF2_out[2]), .A2(
        Inst_f3_dinv_2_lowmul_n258), .ZN(Inst_f3_dinv_2_lowmul_n279) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U26 ( .A(Inst_f3_dinv_2_d_3_), .B(
        Inst_f3_dinv_2_d_5_), .Z(Inst_f3_dinv_2_lowmul_n258) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U25 ( .A1(Inst_f3_dinv_2_lowmul_n257), .A2(
        Inst_f3_dinv_2_lowmul_n319), .ZN(Inst_f3_dinv_2_lowmul_n259) );
  INV_X1 Inst_f3_dinv_2_lowmul_U24 ( .A(FF2_out[3]), .ZN(
        Inst_f3_dinv_2_lowmul_n319) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U23 ( .A(Inst_f3_dinv_2_d_5_), .B(
        Inst_f3_dinv_2_d_4_), .ZN(Inst_f3_dinv_2_lowmul_n257) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U22 ( .A(Inst_f3_dinv_2_lowmul_n282), .B(
        FF2_out[4]), .ZN(Inst_f3_dinv_2_lowmul_n261) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U21 ( .A1(Inst_f3_dinv_2_d_4_), .A2(
        FF2_out[5]), .ZN(Inst_f3_dinv_2_lowmul_n282) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U20 ( .A1(Inst_f3_dinv_2_lowmul_n326), .A2(
        Inst_f3_dinv_2_lowmul_n308), .ZN(Inst_f3_dinv_2_lowmul_n263) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U19 ( .A(FF2_out[4]), .B(FF2_out[5]), .ZN(
        Inst_f3_dinv_2_lowmul_n308) );
  INV_X1 Inst_f3_dinv_2_lowmul_U18 ( .A(Inst_f3_dinv_2_d_3_), .ZN(
        Inst_f3_dinv_2_lowmul_n326) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U17 ( .A(Inst_f3_dinv_2_lowmul_n269), .B(
        Inst_f3_dinv_2_lowmul_n256), .ZN(Inst_f3_dinv_2_lowmul_n340) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U16 ( .A1(Inst_f3_dinv_2_d_2_), .A2(
        FF2_out[2]), .ZN(Inst_f3_dinv_2_lowmul_n256) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U15 ( .A1(FF2_out[3]), .A2(
        Inst_f3_dinv_2_d_3_), .ZN(Inst_f3_dinv_2_lowmul_n269) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U14 ( .A(Inst_f3_dinv_2_lowmul_n255), .B(
        Inst_f3_dinv_2_lowmul_n340), .Z(Inst_f3_dinv_2_ph[5]) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U13 ( .A(Inst_f3_dinv_2_lowmul_n254), .B(
        Inst_f3_dinv_2_lowmul_n252), .ZN(Inst_f3_dinv_2_lowmul_n255) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U12 ( .A1(Inst_f3_dinv_2_lowmul_n253), .A2(
        Inst_f3_dinv_2_lowmul_n249), .ZN(Inst_f3_dinv_2_lowmul_n254) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U11 ( .A1(Inst_f3_dinv_2_lowmul_n243), .A2(
        FF2_out[1]), .ZN(Inst_f3_dinv_2_lowmul_n253) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U10 ( .A(Inst_f3_dinv_2_lowmul_n251), .B(
        Inst_f3_dinv_2_lowmul_n339), .Z(Inst_f3_dinv_2_lowmul_n252) );
  NOR2_X1 Inst_f3_dinv_2_lowmul_U9 ( .A1(Inst_f3_dinv_2_lowmul_n338), .A2(
        Inst_f3_dinv_2_lowmul_n250), .ZN(Inst_f3_dinv_2_lowmul_n251) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U8 ( .A(FF2_out[2]), .B(FF2_out[3]), .ZN(
        Inst_f3_dinv_2_lowmul_n250) );
  XOR2_X1 Inst_f3_dinv_2_lowmul_U7 ( .A(Inst_f3_dinv_2_lowmul_n246), .B(
        Inst_f3_dinv_2_lowmul_n248), .Z(Inst_f3_dinv_2_lowmul_n249) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U6 ( .A1(Inst_f3_dinv_2_lowmul_n247), .A2(
        Inst_f3_dinv_2_d_1_), .ZN(Inst_f3_dinv_2_lowmul_n248) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U5 ( .A1(FF2_out[0]), .A2(
        Inst_f3_dinv_2_lowmul_n337), .ZN(Inst_f3_dinv_2_lowmul_n247) );
  NAND2_X1 Inst_f3_dinv_2_lowmul_U4 ( .A1(FF2_out[0]), .A2(
        Inst_f3_dinv_2_lowmul_n245), .ZN(Inst_f3_dinv_2_lowmul_n246) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U3 ( .A(Inst_f3_dinv_2_lowmul_n244), .B(
        Inst_f3_dinv_2_d_2_), .ZN(Inst_f3_dinv_2_lowmul_n245) );
  XNOR2_X1 Inst_f3_dinv_2_lowmul_U2 ( .A(Inst_f3_dinv_2_d_0_), .B(
        Inst_f3_dinv_2_d_3_), .ZN(Inst_f3_dinv_2_lowmul_n244) );
  INV_X1 Inst_f3_dinv_2_lowmul_U1 ( .A(FF2_out[0]), .ZN(
        Inst_f3_dinv_2_lowmul_n243) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_MaskXORInst_U4 ( .A(PRNGQ[24]), .B(
        PRNGQ[26]), .Z(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[2]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_MaskXORInst_U3 ( .A(PRNGQ[20]), .B(
        PRNGQ[22]), .Z(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[0]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_MaskXORInst_U2 ( .A(PRNGQ[25]), .B(
        PRNGQ[27]), .Z(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[3]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_MaskXORInst_U1 ( .A(PRNGQ[21]), .B(
        PRNGQ[23]), .Z(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[1]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst1_U4 ( .A(Inst_f3_dinv_2_ph[4]), 
        .B(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[2]), .Z(muld[10]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst1_U3 ( .A(Inst_f3_dinv_2_pl[4]), 
        .B(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[0]), .Z(muld[8]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst1_U2 ( .A(Inst_f3_dinv_2_ph[5]), 
        .B(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[3]), .Z(muld[11]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst1_U1 ( .A(Inst_f3_dinv_2_pl[5]), 
        .B(Inst_f3_dinv_2_AddNewMaskQ_MaskXOR[1]), .Z(muld[9]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U8 ( .A(Inst_f3_dinv_2_ph[3]), 
        .B(PRNGQ[27]), .Z(muld[7]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U7 ( .A(Inst_f3_dinv_2_ph[2]), 
        .B(PRNGQ[26]), .Z(muld[6]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U6 ( .A(Inst_f3_dinv_2_pl[3]), 
        .B(PRNGQ[23]), .Z(muld[5]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U5 ( .A(Inst_f3_dinv_2_pl[2]), 
        .B(PRNGQ[22]), .Z(muld[4]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U4 ( .A(Inst_f3_dinv_2_ph[1]), 
        .B(PRNGQ[25]), .Z(muld[3]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U3 ( .A(Inst_f3_dinv_2_ph[0]), 
        .B(PRNGQ[24]), .Z(muld[2]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U2 ( .A(Inst_f3_dinv_2_pl[1]), 
        .B(PRNGQ[21]), .Z(muld[1]) );
  XOR2_X1 Inst_f3_dinv_2_AddNewMaskQ_XORInst2_U1 ( .A(Inst_f3_dinv_2_pl[0]), 
        .B(PRNGQ[20]), .Z(muld[0]) );
  DFF_X1 PL_3_s_current_state_reg_0_ ( .D(muld[0]), .CK(clk), .Q(FF3_out[0]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_1_ ( .D(muld[1]), .CK(clk), .Q(FF3_out[1]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_2_ ( .D(muld[2]), .CK(clk), .Q(FF3_out[2]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_3_ ( .D(muld[3]), .CK(clk), .Q(FF3_out[3]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_4_ ( .D(muld[4]), .CK(clk), .Q(FF3_out[4]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_5_ ( .D(muld[5]), .CK(clk), .Q(FF3_out[5]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_6_ ( .D(muld[6]), .CK(clk), .Q(FF3_out[6]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_7_ ( .D(muld[7]), .CK(clk), .Q(FF3_out[7]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_8_ ( .D(muld[8]), .CK(clk), .Q(FF3_out[8]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_9_ ( .D(muld[9]), .CK(clk), .Q(FF3_out[9]), 
        .QN() );
  DFF_X1 PL_3_s_current_state_reg_10_ ( .D(muld[10]), .CK(clk), .Q(FF3_out[10]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_11_ ( .D(muld[11]), .CK(clk), .Q(FF3_out[11]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_12_ ( .D(Zl_f3[0]), .CK(clk), .Q(FF3_out[12]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_13_ ( .D(Zl_f3[1]), .CK(clk), .Q(FF3_out[13]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_14_ ( .D(Zl_f3[2]), .CK(clk), .Q(FF3_out[14]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_15_ ( .D(Zl_f3[3]), .CK(clk), .Q(FF3_out[15]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_16_ ( .D(Zl_f3[4]), .CK(clk), .Q(FF3_out[16]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_17_ ( .D(Zl_f3[5]), .CK(clk), .Q(FF3_out[17]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_18_ ( .D(Zl_f3[6]), .CK(clk), .Q(FF3_out[18]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_19_ ( .D(Zl_f3[7]), .CK(clk), .Q(FF3_out[19]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_20_ ( .D(Zl_f3[8]), .CK(clk), .Q(FF3_out[20]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_21_ ( .D(Zl_f3[9]), .CK(clk), .Q(FF3_out[21]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_22_ ( .D(Zl_f3[10]), .CK(clk), .Q(
        FF3_out[22]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_23_ ( .D(Zl_f3[11]), .CK(clk), .Q(
        FF3_out[23]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_24_ ( .D(Zh_f3[0]), .CK(clk), .Q(FF3_out[24]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_25_ ( .D(Zh_f3[1]), .CK(clk), .Q(FF3_out[25]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_26_ ( .D(Zh_f3[2]), .CK(clk), .Q(FF3_out[26]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_27_ ( .D(Zh_f3[3]), .CK(clk), .Q(FF3_out[27]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_28_ ( .D(Zh_f3[4]), .CK(clk), .Q(FF3_out[28]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_29_ ( .D(Zh_f3[5]), .CK(clk), .Q(FF3_out[29]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_30_ ( .D(Zh_f3[6]), .CK(clk), .Q(FF3_out[30]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_31_ ( .D(Zh_f3[7]), .CK(clk), .Q(FF3_out[31]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_32_ ( .D(Zh_f3[8]), .CK(clk), .Q(FF3_out[32]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_33_ ( .D(Zh_f3[9]), .CK(clk), .Q(FF3_out[33]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_34_ ( .D(Zh_f3[10]), .CK(clk), .Q(
        FF3_out[34]), .QN() );
  DFF_X1 PL_3_s_current_state_reg_35_ ( .D(Zh_f3[11]), .CK(clk), .Q(
        FF3_out[35]), .QN() );
  XOR2_X1 Inst_f4_multd_L_U12 ( .A(FF3_out[11]), .B(FF3_out[9]), .Z(
        Inst_f4_multd_L_sB[5]) );
  XOR2_X1 Inst_f4_multd_L_U11 ( .A(FF3_out[10]), .B(FF3_out[8]), .Z(
        Inst_f4_multd_L_sB[4]) );
  XOR2_X1 Inst_f4_multd_L_U10 ( .A(FF3_out[5]), .B(FF3_out[7]), .Z(
        Inst_f4_multd_L_sB[3]) );
  XOR2_X1 Inst_f4_multd_L_U9 ( .A(FF3_out[4]), .B(FF3_out[6]), .Z(
        Inst_f4_multd_L_sB[2]) );
  XOR2_X1 Inst_f4_multd_L_U8 ( .A(FF3_out[1]), .B(FF3_out[3]), .Z(
        Inst_f4_multd_L_sB[1]) );
  XOR2_X1 Inst_f4_multd_L_U7 ( .A(FF3_out[0]), .B(FF3_out[2]), .Z(
        Inst_f4_multd_L_sB[0]) );
  XOR2_X1 Inst_f4_multd_L_U6 ( .A(FF3_out[35]), .B(FF3_out[33]), .Z(
        Inst_f4_multd_L_sA[5]) );
  XOR2_X1 Inst_f4_multd_L_U5 ( .A(FF3_out[34]), .B(FF3_out[32]), .Z(
        Inst_f4_multd_L_sA[4]) );
  XOR2_X1 Inst_f4_multd_L_U4 ( .A(FF3_out[29]), .B(FF3_out[31]), .Z(
        Inst_f4_multd_L_sA[3]) );
  XOR2_X1 Inst_f4_multd_L_U3 ( .A(FF3_out[28]), .B(FF3_out[30]), .Z(
        Inst_f4_multd_L_sA[2]) );
  XOR2_X1 Inst_f4_multd_L_U2 ( .A(FF3_out[25]), .B(FF3_out[27]), .Z(
        Inst_f4_multd_L_sA[1]) );
  XOR2_X1 Inst_f4_multd_L_U1 ( .A(FF3_out[24]), .B(FF3_out[26]), .Z(
        Inst_f4_multd_L_sA[0]) );
  XNOR2_X1 Inst_f4_multd_L_himul_U104 ( .A(Inst_f4_multd_L_himul_n336), .B(
        Inst_f4_multd_L_himul_n335), .ZN(Inst_f4_multd_L_Orig_ph[4]) );
  XNOR2_X1 Inst_f4_multd_L_himul_U103 ( .A(Inst_f4_multd_L_himul_n334), .B(
        Inst_f4_multd_L_himul_n333), .ZN(Inst_f4_multd_L_himul_n335) );
  XNOR2_X1 Inst_f4_multd_L_himul_U102 ( .A(Inst_f4_multd_L_himul_n332), .B(
        Inst_f4_multd_L_himul_n331), .ZN(Inst_f4_multd_L_himul_n333) );
  NAND2_X1 Inst_f4_multd_L_himul_U101 ( .A1(Inst_f4_multd_L_himul_n330), .A2(
        FF3_out[30]), .ZN(Inst_f4_multd_L_himul_n332) );
  NAND2_X1 Inst_f4_multd_L_himul_U100 ( .A1(Inst_f4_multd_L_himul_n329), .A2(
        Inst_f4_multd_L_himul_n328), .ZN(Inst_f4_multd_L_himul_n334) );
  NAND2_X1 Inst_f4_multd_L_himul_U99 ( .A1(FF3_out[2]), .A2(
        Inst_f4_multd_L_himul_n327), .ZN(Inst_f4_multd_L_himul_n328) );
  OR2_X1 Inst_f4_multd_L_himul_U98 ( .A1(Inst_f4_multd_L_himul_n327), .A2(
        Inst_f4_multd_L_himul_n337), .ZN(Inst_f4_multd_L_himul_n329) );
  XOR2_X1 Inst_f4_multd_L_himul_U97 ( .A(FF3_out[27]), .B(
        Inst_f4_multd_L_himul_n326), .Z(Inst_f4_multd_L_himul_n327) );
  XNOR2_X1 Inst_f4_multd_L_himul_U96 ( .A(Inst_f4_multd_L_himul_n325), .B(
        Inst_f4_multd_L_himul_n339), .ZN(Inst_f4_multd_L_himul_n336) );
  XOR2_X1 Inst_f4_multd_L_himul_U95 ( .A(Inst_f4_multd_L_himul_n324), .B(
        Inst_f4_multd_L_himul_n323), .Z(Inst_f4_multd_L_himul_n339) );
  NAND2_X1 Inst_f4_multd_L_himul_U94 ( .A1(FF3_out[6]), .A2(FF3_out[27]), .ZN(
        Inst_f4_multd_L_himul_n323) );
  NOR2_X1 Inst_f4_multd_L_himul_U93 ( .A1(Inst_f4_multd_L_himul_n322), .A2(
        Inst_f4_multd_L_himul_n337), .ZN(Inst_f4_multd_L_himul_n324) );
  INV_X1 Inst_f4_multd_L_himul_U92 ( .A(FF3_out[3]), .ZN(
        Inst_f4_multd_L_himul_n337) );
  XNOR2_X1 Inst_f4_multd_L_himul_U91 ( .A(FF3_out[26]), .B(FF3_out[30]), .ZN(
        Inst_f4_multd_L_himul_n322) );
  NAND2_X1 Inst_f4_multd_L_himul_U90 ( .A1(Inst_f4_multd_L_himul_n321), .A2(
        Inst_f4_multd_L_himul_n320), .ZN(Inst_f4_multd_L_himul_n325) );
  NAND2_X1 Inst_f4_multd_L_himul_U89 ( .A1(FF3_out[27]), .A2(
        Inst_f4_multd_L_himul_n319), .ZN(Inst_f4_multd_L_himul_n320) );
  NAND2_X1 Inst_f4_multd_L_himul_U88 ( .A1(FF3_out[26]), .A2(FF3_out[7]), .ZN(
        Inst_f4_multd_L_himul_n321) );
  XNOR2_X1 Inst_f4_multd_L_himul_U87 ( .A(Inst_f4_multd_L_himul_n318), .B(
        Inst_f4_multd_L_himul_n317), .ZN(Inst_f4_multd_L_Orig_ph[3]) );
  XNOR2_X1 Inst_f4_multd_L_himul_U86 ( .A(Inst_f4_multd_L_himul_n316), .B(
        Inst_f4_multd_L_himul_n315), .ZN(Inst_f4_multd_L_himul_n317) );
  XOR2_X1 Inst_f4_multd_L_himul_U85 ( .A(Inst_f4_multd_L_himul_n314), .B(
        Inst_f4_multd_L_himul_n313), .Z(Inst_f4_multd_L_himul_n316) );
  NAND2_X1 Inst_f4_multd_L_himul_U84 ( .A1(FF3_out[34]), .A2(FF3_out[10]), 
        .ZN(Inst_f4_multd_L_himul_n313) );
  NAND2_X1 Inst_f4_multd_L_himul_U83 ( .A1(FF3_out[35]), .A2(FF3_out[11]), 
        .ZN(Inst_f4_multd_L_himul_n314) );
  XOR2_X1 Inst_f4_multd_L_himul_U82 ( .A(Inst_f4_multd_L_himul_n312), .B(
        Inst_f4_multd_L_himul_n311), .Z(Inst_f4_multd_L_himul_n318) );
  XOR2_X1 Inst_f4_multd_L_himul_U81 ( .A(Inst_f4_multd_L_himul_n310), .B(
        Inst_f4_multd_L_himul_n309), .Z(Inst_f4_multd_L_himul_n311) );
  NAND2_X1 Inst_f4_multd_L_himul_U80 ( .A1(FF3_out[34]), .A2(
        Inst_f4_multd_L_himul_n308), .ZN(Inst_f4_multd_L_himul_n309) );
  NAND2_X1 Inst_f4_multd_L_himul_U79 ( .A1(FF3_out[26]), .A2(FF3_out[11]), 
        .ZN(Inst_f4_multd_L_himul_n310) );
  XNOR2_X1 Inst_f4_multd_L_himul_U78 ( .A(Inst_f4_multd_L_himul_n307), .B(
        Inst_f4_multd_L_himul_n306), .ZN(Inst_f4_multd_L_himul_n312) );
  XNOR2_X1 Inst_f4_multd_L_himul_U77 ( .A(FF3_out[35]), .B(
        Inst_f4_multd_L_himul_n305), .ZN(Inst_f4_multd_L_himul_n306) );
  XOR2_X1 Inst_f4_multd_L_himul_U76 ( .A(Inst_f4_multd_L_himul_n304), .B(
        Inst_f4_multd_L_himul_n303), .Z(Inst_f4_multd_L_himul_n305) );
  NAND2_X1 Inst_f4_multd_L_himul_U75 ( .A1(FF3_out[2]), .A2(FF3_out[34]), .ZN(
        Inst_f4_multd_L_himul_n303) );
  NOR2_X1 Inst_f4_multd_L_himul_U74 ( .A1(Inst_f4_multd_L_himul_n302), .A2(
        FF3_out[3]), .ZN(Inst_f4_multd_L_himul_n304) );
  NAND2_X1 Inst_f4_multd_L_himul_U73 ( .A1(Inst_f4_multd_L_himul_n301), .A2(
        FF3_out[10]), .ZN(Inst_f4_multd_L_himul_n307) );
  XNOR2_X1 Inst_f4_multd_L_himul_U72 ( .A(Inst_f4_multd_L_himul_n338), .B(
        Inst_f4_multd_L_himul_n300), .ZN(Inst_f4_multd_L_himul_n301) );
  XNOR2_X1 Inst_f4_multd_L_himul_U71 ( .A(FF3_out[27]), .B(
        Inst_f4_multd_L_himul_n299), .ZN(Inst_f4_multd_L_himul_n300) );
  INV_X1 Inst_f4_multd_L_himul_U70 ( .A(FF3_out[26]), .ZN(
        Inst_f4_multd_L_himul_n338) );
  XOR2_X1 Inst_f4_multd_L_himul_U69 ( .A(Inst_f4_multd_L_himul_n298), .B(
        Inst_f4_multd_L_himul_n297), .Z(Inst_f4_multd_L_Orig_ph[2]) );
  NAND2_X1 Inst_f4_multd_L_himul_U68 ( .A1(Inst_f4_multd_L_himul_n296), .A2(
        Inst_f4_multd_L_himul_n295), .ZN(Inst_f4_multd_L_himul_n297) );
  OR2_X1 Inst_f4_multd_L_himul_U67 ( .A1(FF3_out[11]), .A2(
        Inst_f4_multd_L_himul_n302), .ZN(Inst_f4_multd_L_himul_n295) );
  NAND2_X1 Inst_f4_multd_L_himul_U66 ( .A1(Inst_f4_multd_L_himul_n294), .A2(
        FF3_out[11]), .ZN(Inst_f4_multd_L_himul_n296) );
  XNOR2_X1 Inst_f4_multd_L_himul_U65 ( .A(Inst_f4_multd_L_himul_n293), .B(
        FF3_out[26]), .ZN(Inst_f4_multd_L_himul_n294) );
  XOR2_X1 Inst_f4_multd_L_himul_U64 ( .A(Inst_f4_multd_L_himul_n292), .B(
        Inst_f4_multd_L_himul_n291), .Z(Inst_f4_multd_L_himul_n298) );
  NOR2_X1 Inst_f4_multd_L_himul_U63 ( .A1(Inst_f4_multd_L_himul_n299), .A2(
        Inst_f4_multd_L_himul_n290), .ZN(Inst_f4_multd_L_himul_n291) );
  XOR2_X1 Inst_f4_multd_L_himul_U62 ( .A(Inst_f4_multd_L_himul_n308), .B(
        FF3_out[3]), .Z(Inst_f4_multd_L_himul_n290) );
  XNOR2_X1 Inst_f4_multd_L_himul_U61 ( .A(Inst_f4_multd_L_himul_n289), .B(
        Inst_f4_multd_L_himul_n288), .ZN(Inst_f4_multd_L_himul_n292) );
  XNOR2_X1 Inst_f4_multd_L_himul_U60 ( .A(FF3_out[2]), .B(
        Inst_f4_multd_L_himul_n331), .ZN(Inst_f4_multd_L_himul_n288) );
  XOR2_X1 Inst_f4_multd_L_himul_U59 ( .A(Inst_f4_multd_L_himul_n287), .B(
        Inst_f4_multd_L_himul_n286), .Z(Inst_f4_multd_L_himul_n331) );
  NAND2_X1 Inst_f4_multd_L_himul_U58 ( .A1(FF3_out[27]), .A2(FF3_out[2]), .ZN(
        Inst_f4_multd_L_himul_n286) );
  NAND2_X1 Inst_f4_multd_L_himul_U57 ( .A1(FF3_out[26]), .A2(FF3_out[3]), .ZN(
        Inst_f4_multd_L_himul_n287) );
  XOR2_X1 Inst_f4_multd_L_himul_U56 ( .A(Inst_f4_multd_L_himul_n285), .B(
        Inst_f4_multd_L_himul_n315), .Z(Inst_f4_multd_L_himul_n289) );
  XOR2_X1 Inst_f4_multd_L_himul_U55 ( .A(Inst_f4_multd_L_himul_n284), .B(
        Inst_f4_multd_L_himul_n283), .Z(Inst_f4_multd_L_himul_n315) );
  NAND2_X1 Inst_f4_multd_L_himul_U54 ( .A1(FF3_out[34]), .A2(FF3_out[3]), .ZN(
        Inst_f4_multd_L_himul_n283) );
  NAND2_X1 Inst_f4_multd_L_himul_U53 ( .A1(FF3_out[35]), .A2(FF3_out[2]), .ZN(
        Inst_f4_multd_L_himul_n284) );
  XOR2_X1 Inst_f4_multd_L_himul_U52 ( .A(Inst_f4_multd_L_himul_n282), .B(
        Inst_f4_multd_L_himul_n281), .Z(Inst_f4_multd_L_himul_n285) );
  NAND2_X1 Inst_f4_multd_L_himul_U51 ( .A1(FF3_out[10]), .A2(
        Inst_f4_multd_L_himul_n302), .ZN(Inst_f4_multd_L_himul_n281) );
  INV_X1 Inst_f4_multd_L_himul_U50 ( .A(FF3_out[27]), .ZN(
        Inst_f4_multd_L_himul_n302) );
  XNOR2_X1 Inst_f4_multd_L_himul_U49 ( .A(Inst_f4_multd_L_himul_n280), .B(
        Inst_f4_multd_L_himul_n279), .ZN(Inst_f4_multd_L_Orig_ph[1]) );
  XNOR2_X1 Inst_f4_multd_L_himul_U48 ( .A(Inst_f4_multd_L_himul_n278), .B(
        Inst_f4_multd_L_himul_n277), .ZN(Inst_f4_multd_L_himul_n280) );
  NAND2_X1 Inst_f4_multd_L_himul_U47 ( .A1(Inst_f4_multd_L_himul_n276), .A2(
        FF3_out[30]), .ZN(Inst_f4_multd_L_himul_n277) );
  XNOR2_X1 Inst_f4_multd_L_himul_U46 ( .A(FF3_out[6]), .B(
        Inst_f4_multd_L_himul_n308), .ZN(Inst_f4_multd_L_himul_n276) );
  XNOR2_X1 Inst_f4_multd_L_himul_U45 ( .A(Inst_f4_multd_L_himul_n275), .B(
        Inst_f4_multd_L_himul_n274), .ZN(Inst_f4_multd_L_himul_n278) );
  XNOR2_X1 Inst_f4_multd_L_himul_U44 ( .A(Inst_f4_multd_L_himul_n273), .B(
        Inst_f4_multd_L_himul_n272), .ZN(Inst_f4_multd_L_himul_n274) );
  NAND2_X1 Inst_f4_multd_L_himul_U43 ( .A1(Inst_f4_multd_L_himul_n271), .A2(
        Inst_f4_multd_L_himul_n330), .ZN(Inst_f4_multd_L_himul_n272) );
  XOR2_X1 Inst_f4_multd_L_himul_U42 ( .A(FF3_out[6]), .B(FF3_out[7]), .Z(
        Inst_f4_multd_L_himul_n330) );
  XOR2_X1 Inst_f4_multd_L_himul_U41 ( .A(FF3_out[30]), .B(FF3_out[34]), .Z(
        Inst_f4_multd_L_himul_n271) );
  NAND2_X1 Inst_f4_multd_L_himul_U40 ( .A1(FF3_out[31]), .A2(FF3_out[10]), 
        .ZN(Inst_f4_multd_L_himul_n273) );
  XNOR2_X1 Inst_f4_multd_L_himul_U39 ( .A(Inst_f4_multd_L_himul_n270), .B(
        Inst_f4_multd_L_himul_n269), .ZN(Inst_f4_multd_L_himul_n275) );
  XOR2_X1 Inst_f4_multd_L_himul_U38 ( .A(Inst_f4_multd_L_himul_n268), .B(
        Inst_f4_multd_L_himul_n267), .Z(Inst_f4_multd_L_himul_n270) );
  NOR2_X1 Inst_f4_multd_L_himul_U37 ( .A1(Inst_f4_multd_L_himul_n293), .A2(
        FF3_out[10]), .ZN(Inst_f4_multd_L_himul_n267) );
  INV_X1 Inst_f4_multd_L_himul_U36 ( .A(FF3_out[34]), .ZN(
        Inst_f4_multd_L_himul_n293) );
  NOR2_X1 Inst_f4_multd_L_himul_U35 ( .A1(Inst_f4_multd_L_himul_n299), .A2(
        FF3_out[11]), .ZN(Inst_f4_multd_L_himul_n268) );
  INV_X1 Inst_f4_multd_L_himul_U34 ( .A(FF3_out[35]), .ZN(
        Inst_f4_multd_L_himul_n299) );
  XNOR2_X1 Inst_f4_multd_L_himul_U33 ( .A(Inst_f4_multd_L_himul_n266), .B(
        Inst_f4_multd_L_himul_n265), .ZN(Inst_f4_multd_L_Orig_ph[0]) );
  NAND2_X1 Inst_f4_multd_L_himul_U32 ( .A1(FF3_out[30]), .A2(FF3_out[11]), 
        .ZN(Inst_f4_multd_L_himul_n265) );
  XNOR2_X1 Inst_f4_multd_L_himul_U31 ( .A(Inst_f4_multd_L_himul_n340), .B(
        Inst_f4_multd_L_himul_n264), .ZN(Inst_f4_multd_L_himul_n266) );
  XNOR2_X1 Inst_f4_multd_L_himul_U30 ( .A(Inst_f4_multd_L_himul_n263), .B(
        Inst_f4_multd_L_himul_n262), .ZN(Inst_f4_multd_L_himul_n264) );
  XNOR2_X1 Inst_f4_multd_L_himul_U29 ( .A(Inst_f4_multd_L_himul_n261), .B(
        Inst_f4_multd_L_himul_n260), .ZN(Inst_f4_multd_L_himul_n262) );
  XNOR2_X1 Inst_f4_multd_L_himul_U28 ( .A(Inst_f4_multd_L_himul_n259), .B(
        Inst_f4_multd_L_himul_n279), .ZN(Inst_f4_multd_L_himul_n260) );
  NAND2_X1 Inst_f4_multd_L_himul_U27 ( .A1(FF3_out[6]), .A2(
        Inst_f4_multd_L_himul_n258), .ZN(Inst_f4_multd_L_himul_n279) );
  XOR2_X1 Inst_f4_multd_L_himul_U26 ( .A(FF3_out[31]), .B(FF3_out[35]), .Z(
        Inst_f4_multd_L_himul_n258) );
  NOR2_X1 Inst_f4_multd_L_himul_U25 ( .A1(Inst_f4_multd_L_himul_n257), .A2(
        Inst_f4_multd_L_himul_n319), .ZN(Inst_f4_multd_L_himul_n259) );
  INV_X1 Inst_f4_multd_L_himul_U24 ( .A(FF3_out[7]), .ZN(
        Inst_f4_multd_L_himul_n319) );
  XNOR2_X1 Inst_f4_multd_L_himul_U23 ( .A(FF3_out[35]), .B(FF3_out[34]), .ZN(
        Inst_f4_multd_L_himul_n257) );
  XNOR2_X1 Inst_f4_multd_L_himul_U22 ( .A(Inst_f4_multd_L_himul_n282), .B(
        FF3_out[10]), .ZN(Inst_f4_multd_L_himul_n261) );
  NAND2_X1 Inst_f4_multd_L_himul_U21 ( .A1(FF3_out[34]), .A2(FF3_out[11]), 
        .ZN(Inst_f4_multd_L_himul_n282) );
  NOR2_X1 Inst_f4_multd_L_himul_U20 ( .A1(Inst_f4_multd_L_himul_n326), .A2(
        Inst_f4_multd_L_himul_n308), .ZN(Inst_f4_multd_L_himul_n263) );
  XNOR2_X1 Inst_f4_multd_L_himul_U19 ( .A(FF3_out[10]), .B(FF3_out[11]), .ZN(
        Inst_f4_multd_L_himul_n308) );
  INV_X1 Inst_f4_multd_L_himul_U18 ( .A(FF3_out[31]), .ZN(
        Inst_f4_multd_L_himul_n326) );
  XNOR2_X1 Inst_f4_multd_L_himul_U17 ( .A(Inst_f4_multd_L_himul_n269), .B(
        Inst_f4_multd_L_himul_n256), .ZN(Inst_f4_multd_L_himul_n340) );
  NAND2_X1 Inst_f4_multd_L_himul_U16 ( .A1(FF3_out[30]), .A2(FF3_out[6]), .ZN(
        Inst_f4_multd_L_himul_n256) );
  NAND2_X1 Inst_f4_multd_L_himul_U15 ( .A1(FF3_out[7]), .A2(FF3_out[31]), .ZN(
        Inst_f4_multd_L_himul_n269) );
  XOR2_X1 Inst_f4_multd_L_himul_U14 ( .A(Inst_f4_multd_L_himul_n255), .B(
        Inst_f4_multd_L_himul_n340), .Z(Inst_f4_multd_L_Orig_ph[5]) );
  XNOR2_X1 Inst_f4_multd_L_himul_U13 ( .A(Inst_f4_multd_L_himul_n254), .B(
        Inst_f4_multd_L_himul_n252), .ZN(Inst_f4_multd_L_himul_n255) );
  NAND2_X1 Inst_f4_multd_L_himul_U12 ( .A1(Inst_f4_multd_L_himul_n253), .A2(
        Inst_f4_multd_L_himul_n249), .ZN(Inst_f4_multd_L_himul_n254) );
  NAND2_X1 Inst_f4_multd_L_himul_U11 ( .A1(Inst_f4_multd_L_himul_n243), .A2(
        FF3_out[3]), .ZN(Inst_f4_multd_L_himul_n253) );
  XOR2_X1 Inst_f4_multd_L_himul_U10 ( .A(Inst_f4_multd_L_himul_n251), .B(
        Inst_f4_multd_L_himul_n339), .Z(Inst_f4_multd_L_himul_n252) );
  NOR2_X1 Inst_f4_multd_L_himul_U9 ( .A1(Inst_f4_multd_L_himul_n338), .A2(
        Inst_f4_multd_L_himul_n250), .ZN(Inst_f4_multd_L_himul_n251) );
  XNOR2_X1 Inst_f4_multd_L_himul_U8 ( .A(FF3_out[6]), .B(FF3_out[7]), .ZN(
        Inst_f4_multd_L_himul_n250) );
  XOR2_X1 Inst_f4_multd_L_himul_U7 ( .A(Inst_f4_multd_L_himul_n246), .B(
        Inst_f4_multd_L_himul_n248), .Z(Inst_f4_multd_L_himul_n249) );
  NAND2_X1 Inst_f4_multd_L_himul_U6 ( .A1(Inst_f4_multd_L_himul_n247), .A2(
        FF3_out[27]), .ZN(Inst_f4_multd_L_himul_n248) );
  NAND2_X1 Inst_f4_multd_L_himul_U5 ( .A1(FF3_out[2]), .A2(
        Inst_f4_multd_L_himul_n337), .ZN(Inst_f4_multd_L_himul_n247) );
  NAND2_X1 Inst_f4_multd_L_himul_U4 ( .A1(FF3_out[2]), .A2(
        Inst_f4_multd_L_himul_n245), .ZN(Inst_f4_multd_L_himul_n246) );
  XNOR2_X1 Inst_f4_multd_L_himul_U3 ( .A(Inst_f4_multd_L_himul_n244), .B(
        FF3_out[30]), .ZN(Inst_f4_multd_L_himul_n245) );
  XNOR2_X1 Inst_f4_multd_L_himul_U2 ( .A(FF3_out[26]), .B(FF3_out[31]), .ZN(
        Inst_f4_multd_L_himul_n244) );
  INV_X1 Inst_f4_multd_L_himul_U1 ( .A(FF3_out[2]), .ZN(
        Inst_f4_multd_L_himul_n243) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_MaskXORInst_U2 ( .A(PRNGQ[40]), .B(
        PRNGQ[42]), .Z(Inst_f4_multd_L_AddNewMaskph_MaskXOR[0]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_MaskXORInst_U1 ( .A(PRNGQ[41]), .B(
        PRNGQ[43]), .Z(Inst_f4_multd_L_AddNewMaskph_MaskXOR[1]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_XORInst1_U2 ( .A(
        Inst_f4_multd_L_Orig_ph[4]), .B(
        Inst_f4_multd_L_AddNewMaskph_MaskXOR[0]), .Z(ph_L[4]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_XORInst1_U1 ( .A(
        Inst_f4_multd_L_Orig_ph[5]), .B(
        Inst_f4_multd_L_AddNewMaskph_MaskXOR[1]), .Z(ph_L[5]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_XORInst2_U4 ( .A(
        Inst_f4_multd_L_Orig_ph[3]), .B(PRNGQ[43]), .Z(ph_L[3]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_XORInst2_U3 ( .A(
        Inst_f4_multd_L_Orig_ph[2]), .B(PRNGQ[42]), .Z(ph_L[2]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_XORInst2_U2 ( .A(
        Inst_f4_multd_L_Orig_ph[1]), .B(PRNGQ[41]), .Z(ph_L[1]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskph_XORInst2_U1 ( .A(
        Inst_f4_multd_L_Orig_ph[0]), .B(PRNGQ[40]), .Z(ph_L[0]) );
  XOR2_X1 Inst_f4_multd_L_summul_U104 ( .A(Inst_f4_multd_L_sA[2]), .B(
        Inst_f4_multd_L_sA[0]), .Z(Inst_f4_multd_L_summul_n336) );
  XNOR2_X1 Inst_f4_multd_L_summul_U103 ( .A(Inst_f4_multd_L_summul_n335), .B(
        Inst_f4_multd_L_summul_n334), .ZN(Inst_f4_multd_L_Orig_p[4]) );
  XNOR2_X1 Inst_f4_multd_L_summul_U102 ( .A(Inst_f4_multd_L_summul_n333), .B(
        Inst_f4_multd_L_summul_n332), .ZN(Inst_f4_multd_L_summul_n334) );
  XNOR2_X1 Inst_f4_multd_L_summul_U101 ( .A(Inst_f4_multd_L_summul_n331), .B(
        Inst_f4_multd_L_summul_n330), .ZN(Inst_f4_multd_L_summul_n332) );
  NAND2_X1 Inst_f4_multd_L_summul_U100 ( .A1(Inst_f4_multd_L_summul_n329), 
        .A2(Inst_f4_multd_L_sA[2]), .ZN(Inst_f4_multd_L_summul_n331) );
  NAND2_X1 Inst_f4_multd_L_summul_U99 ( .A1(Inst_f4_multd_L_summul_n328), .A2(
        Inst_f4_multd_L_summul_n327), .ZN(Inst_f4_multd_L_summul_n333) );
  NAND2_X1 Inst_f4_multd_L_summul_U98 ( .A1(Inst_f4_multd_L_sB[0]), .A2(
        Inst_f4_multd_L_summul_n326), .ZN(Inst_f4_multd_L_summul_n327) );
  OR2_X1 Inst_f4_multd_L_summul_U97 ( .A1(Inst_f4_multd_L_summul_n326), .A2(
        Inst_f4_multd_L_summul_n337), .ZN(Inst_f4_multd_L_summul_n328) );
  XOR2_X1 Inst_f4_multd_L_summul_U96 ( .A(Inst_f4_multd_L_sA[1]), .B(
        Inst_f4_multd_L_summul_n325), .Z(Inst_f4_multd_L_summul_n326) );
  XNOR2_X1 Inst_f4_multd_L_summul_U95 ( .A(Inst_f4_multd_L_summul_n324), .B(
        Inst_f4_multd_L_summul_n339), .ZN(Inst_f4_multd_L_summul_n335) );
  XOR2_X1 Inst_f4_multd_L_summul_U94 ( .A(Inst_f4_multd_L_summul_n323), .B(
        Inst_f4_multd_L_summul_n322), .Z(Inst_f4_multd_L_summul_n339) );
  NAND2_X1 Inst_f4_multd_L_summul_U93 ( .A1(Inst_f4_multd_L_sB[2]), .A2(
        Inst_f4_multd_L_sA[1]), .ZN(Inst_f4_multd_L_summul_n322) );
  NOR2_X1 Inst_f4_multd_L_summul_U92 ( .A1(Inst_f4_multd_L_summul_n321), .A2(
        Inst_f4_multd_L_summul_n337), .ZN(Inst_f4_multd_L_summul_n323) );
  INV_X1 Inst_f4_multd_L_summul_U91 ( .A(Inst_f4_multd_L_sB[1]), .ZN(
        Inst_f4_multd_L_summul_n337) );
  XNOR2_X1 Inst_f4_multd_L_summul_U90 ( .A(Inst_f4_multd_L_sA[0]), .B(
        Inst_f4_multd_L_sA[2]), .ZN(Inst_f4_multd_L_summul_n321) );
  NAND2_X1 Inst_f4_multd_L_summul_U89 ( .A1(Inst_f4_multd_L_summul_n320), .A2(
        Inst_f4_multd_L_summul_n319), .ZN(Inst_f4_multd_L_summul_n324) );
  NAND2_X1 Inst_f4_multd_L_summul_U88 ( .A1(Inst_f4_multd_L_sA[1]), .A2(
        Inst_f4_multd_L_summul_n318), .ZN(Inst_f4_multd_L_summul_n319) );
  NAND2_X1 Inst_f4_multd_L_summul_U87 ( .A1(Inst_f4_multd_L_sA[0]), .A2(
        Inst_f4_multd_L_sB[3]), .ZN(Inst_f4_multd_L_summul_n320) );
  XNOR2_X1 Inst_f4_multd_L_summul_U86 ( .A(Inst_f4_multd_L_summul_n317), .B(
        Inst_f4_multd_L_summul_n316), .ZN(Inst_f4_multd_L_Orig_p[3]) );
  XNOR2_X1 Inst_f4_multd_L_summul_U85 ( .A(Inst_f4_multd_L_summul_n315), .B(
        Inst_f4_multd_L_summul_n314), .ZN(Inst_f4_multd_L_summul_n316) );
  XOR2_X1 Inst_f4_multd_L_summul_U84 ( .A(Inst_f4_multd_L_summul_n313), .B(
        Inst_f4_multd_L_summul_n312), .Z(Inst_f4_multd_L_summul_n315) );
  NAND2_X1 Inst_f4_multd_L_summul_U83 ( .A1(Inst_f4_multd_L_sA[4]), .A2(
        Inst_f4_multd_L_sB[4]), .ZN(Inst_f4_multd_L_summul_n312) );
  NAND2_X1 Inst_f4_multd_L_summul_U82 ( .A1(Inst_f4_multd_L_sA[5]), .A2(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n313) );
  XOR2_X1 Inst_f4_multd_L_summul_U81 ( .A(Inst_f4_multd_L_summul_n311), .B(
        Inst_f4_multd_L_summul_n310), .Z(Inst_f4_multd_L_summul_n317) );
  XOR2_X1 Inst_f4_multd_L_summul_U80 ( .A(Inst_f4_multd_L_summul_n309), .B(
        Inst_f4_multd_L_summul_n308), .Z(Inst_f4_multd_L_summul_n310) );
  NAND2_X1 Inst_f4_multd_L_summul_U79 ( .A1(Inst_f4_multd_L_sA[4]), .A2(
        Inst_f4_multd_L_summul_n307), .ZN(Inst_f4_multd_L_summul_n308) );
  NAND2_X1 Inst_f4_multd_L_summul_U78 ( .A1(Inst_f4_multd_L_sA[0]), .A2(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n309) );
  XNOR2_X1 Inst_f4_multd_L_summul_U77 ( .A(Inst_f4_multd_L_summul_n306), .B(
        Inst_f4_multd_L_summul_n305), .ZN(Inst_f4_multd_L_summul_n311) );
  XNOR2_X1 Inst_f4_multd_L_summul_U76 ( .A(Inst_f4_multd_L_sA[5]), .B(
        Inst_f4_multd_L_summul_n304), .ZN(Inst_f4_multd_L_summul_n305) );
  XOR2_X1 Inst_f4_multd_L_summul_U75 ( .A(Inst_f4_multd_L_summul_n303), .B(
        Inst_f4_multd_L_summul_n302), .Z(Inst_f4_multd_L_summul_n304) );
  NAND2_X1 Inst_f4_multd_L_summul_U74 ( .A1(Inst_f4_multd_L_sB[0]), .A2(
        Inst_f4_multd_L_sA[4]), .ZN(Inst_f4_multd_L_summul_n302) );
  NOR2_X1 Inst_f4_multd_L_summul_U73 ( .A1(Inst_f4_multd_L_summul_n301), .A2(
        Inst_f4_multd_L_sB[1]), .ZN(Inst_f4_multd_L_summul_n303) );
  NAND2_X1 Inst_f4_multd_L_summul_U72 ( .A1(Inst_f4_multd_L_summul_n300), .A2(
        Inst_f4_multd_L_sB[4]), .ZN(Inst_f4_multd_L_summul_n306) );
  XNOR2_X1 Inst_f4_multd_L_summul_U71 ( .A(Inst_f4_multd_L_summul_n338), .B(
        Inst_f4_multd_L_summul_n299), .ZN(Inst_f4_multd_L_summul_n300) );
  XNOR2_X1 Inst_f4_multd_L_summul_U70 ( .A(Inst_f4_multd_L_sA[1]), .B(
        Inst_f4_multd_L_summul_n298), .ZN(Inst_f4_multd_L_summul_n299) );
  INV_X1 Inst_f4_multd_L_summul_U69 ( .A(Inst_f4_multd_L_sA[0]), .ZN(
        Inst_f4_multd_L_summul_n338) );
  XOR2_X1 Inst_f4_multd_L_summul_U68 ( .A(Inst_f4_multd_L_summul_n297), .B(
        Inst_f4_multd_L_summul_n296), .Z(Inst_f4_multd_L_Orig_p[2]) );
  NAND2_X1 Inst_f4_multd_L_summul_U67 ( .A1(Inst_f4_multd_L_summul_n295), .A2(
        Inst_f4_multd_L_summul_n294), .ZN(Inst_f4_multd_L_summul_n296) );
  OR2_X1 Inst_f4_multd_L_summul_U66 ( .A1(Inst_f4_multd_L_sB[5]), .A2(
        Inst_f4_multd_L_summul_n301), .ZN(Inst_f4_multd_L_summul_n294) );
  NAND2_X1 Inst_f4_multd_L_summul_U65 ( .A1(Inst_f4_multd_L_summul_n293), .A2(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n295) );
  XNOR2_X1 Inst_f4_multd_L_summul_U64 ( .A(Inst_f4_multd_L_summul_n292), .B(
        Inst_f4_multd_L_sA[0]), .ZN(Inst_f4_multd_L_summul_n293) );
  XOR2_X1 Inst_f4_multd_L_summul_U63 ( .A(Inst_f4_multd_L_summul_n291), .B(
        Inst_f4_multd_L_summul_n290), .Z(Inst_f4_multd_L_summul_n297) );
  NOR2_X1 Inst_f4_multd_L_summul_U62 ( .A1(Inst_f4_multd_L_summul_n298), .A2(
        Inst_f4_multd_L_summul_n289), .ZN(Inst_f4_multd_L_summul_n290) );
  XOR2_X1 Inst_f4_multd_L_summul_U61 ( .A(Inst_f4_multd_L_summul_n307), .B(
        Inst_f4_multd_L_sB[1]), .Z(Inst_f4_multd_L_summul_n289) );
  XNOR2_X1 Inst_f4_multd_L_summul_U60 ( .A(Inst_f4_multd_L_summul_n288), .B(
        Inst_f4_multd_L_summul_n287), .ZN(Inst_f4_multd_L_summul_n291) );
  XNOR2_X1 Inst_f4_multd_L_summul_U59 ( .A(Inst_f4_multd_L_sB[0]), .B(
        Inst_f4_multd_L_summul_n330), .ZN(Inst_f4_multd_L_summul_n287) );
  XOR2_X1 Inst_f4_multd_L_summul_U58 ( .A(Inst_f4_multd_L_summul_n286), .B(
        Inst_f4_multd_L_summul_n285), .Z(Inst_f4_multd_L_summul_n330) );
  NAND2_X1 Inst_f4_multd_L_summul_U57 ( .A1(Inst_f4_multd_L_sA[1]), .A2(
        Inst_f4_multd_L_sB[0]), .ZN(Inst_f4_multd_L_summul_n285) );
  NAND2_X1 Inst_f4_multd_L_summul_U56 ( .A1(Inst_f4_multd_L_sA[0]), .A2(
        Inst_f4_multd_L_sB[1]), .ZN(Inst_f4_multd_L_summul_n286) );
  XOR2_X1 Inst_f4_multd_L_summul_U55 ( .A(Inst_f4_multd_L_summul_n284), .B(
        Inst_f4_multd_L_summul_n314), .Z(Inst_f4_multd_L_summul_n288) );
  XOR2_X1 Inst_f4_multd_L_summul_U54 ( .A(Inst_f4_multd_L_summul_n283), .B(
        Inst_f4_multd_L_summul_n282), .Z(Inst_f4_multd_L_summul_n314) );
  NAND2_X1 Inst_f4_multd_L_summul_U53 ( .A1(Inst_f4_multd_L_sA[4]), .A2(
        Inst_f4_multd_L_sB[1]), .ZN(Inst_f4_multd_L_summul_n282) );
  NAND2_X1 Inst_f4_multd_L_summul_U52 ( .A1(Inst_f4_multd_L_sA[5]), .A2(
        Inst_f4_multd_L_sB[0]), .ZN(Inst_f4_multd_L_summul_n283) );
  XOR2_X1 Inst_f4_multd_L_summul_U51 ( .A(Inst_f4_multd_L_summul_n281), .B(
        Inst_f4_multd_L_summul_n280), .Z(Inst_f4_multd_L_summul_n284) );
  NAND2_X1 Inst_f4_multd_L_summul_U50 ( .A1(Inst_f4_multd_L_sB[4]), .A2(
        Inst_f4_multd_L_summul_n301), .ZN(Inst_f4_multd_L_summul_n280) );
  INV_X1 Inst_f4_multd_L_summul_U49 ( .A(Inst_f4_multd_L_sA[1]), .ZN(
        Inst_f4_multd_L_summul_n301) );
  XNOR2_X1 Inst_f4_multd_L_summul_U48 ( .A(Inst_f4_multd_L_summul_n279), .B(
        Inst_f4_multd_L_summul_n278), .ZN(Inst_f4_multd_L_Orig_p[1]) );
  XNOR2_X1 Inst_f4_multd_L_summul_U47 ( .A(Inst_f4_multd_L_summul_n277), .B(
        Inst_f4_multd_L_summul_n276), .ZN(Inst_f4_multd_L_summul_n279) );
  NAND2_X1 Inst_f4_multd_L_summul_U46 ( .A1(Inst_f4_multd_L_summul_n275), .A2(
        Inst_f4_multd_L_sA[2]), .ZN(Inst_f4_multd_L_summul_n276) );
  XNOR2_X1 Inst_f4_multd_L_summul_U45 ( .A(Inst_f4_multd_L_sB[2]), .B(
        Inst_f4_multd_L_summul_n307), .ZN(Inst_f4_multd_L_summul_n275) );
  XNOR2_X1 Inst_f4_multd_L_summul_U44 ( .A(Inst_f4_multd_L_summul_n274), .B(
        Inst_f4_multd_L_summul_n273), .ZN(Inst_f4_multd_L_summul_n277) );
  XNOR2_X1 Inst_f4_multd_L_summul_U43 ( .A(Inst_f4_multd_L_summul_n272), .B(
        Inst_f4_multd_L_summul_n271), .ZN(Inst_f4_multd_L_summul_n273) );
  NAND2_X1 Inst_f4_multd_L_summul_U42 ( .A1(Inst_f4_multd_L_summul_n270), .A2(
        Inst_f4_multd_L_summul_n329), .ZN(Inst_f4_multd_L_summul_n271) );
  XOR2_X1 Inst_f4_multd_L_summul_U41 ( .A(Inst_f4_multd_L_sB[2]), .B(
        Inst_f4_multd_L_sB[3]), .Z(Inst_f4_multd_L_summul_n329) );
  XOR2_X1 Inst_f4_multd_L_summul_U40 ( .A(Inst_f4_multd_L_sA[2]), .B(
        Inst_f4_multd_L_sA[4]), .Z(Inst_f4_multd_L_summul_n270) );
  NAND2_X1 Inst_f4_multd_L_summul_U39 ( .A1(Inst_f4_multd_L_sA[3]), .A2(
        Inst_f4_multd_L_sB[4]), .ZN(Inst_f4_multd_L_summul_n272) );
  XNOR2_X1 Inst_f4_multd_L_summul_U38 ( .A(Inst_f4_multd_L_summul_n269), .B(
        Inst_f4_multd_L_summul_n268), .ZN(Inst_f4_multd_L_summul_n274) );
  XOR2_X1 Inst_f4_multd_L_summul_U37 ( .A(Inst_f4_multd_L_summul_n267), .B(
        Inst_f4_multd_L_summul_n266), .Z(Inst_f4_multd_L_summul_n269) );
  NOR2_X1 Inst_f4_multd_L_summul_U36 ( .A1(Inst_f4_multd_L_summul_n292), .A2(
        Inst_f4_multd_L_sB[4]), .ZN(Inst_f4_multd_L_summul_n266) );
  INV_X1 Inst_f4_multd_L_summul_U35 ( .A(Inst_f4_multd_L_sA[4]), .ZN(
        Inst_f4_multd_L_summul_n292) );
  NOR2_X1 Inst_f4_multd_L_summul_U34 ( .A1(Inst_f4_multd_L_summul_n298), .A2(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n267) );
  INV_X1 Inst_f4_multd_L_summul_U33 ( .A(Inst_f4_multd_L_sA[5]), .ZN(
        Inst_f4_multd_L_summul_n298) );
  XNOR2_X1 Inst_f4_multd_L_summul_U32 ( .A(Inst_f4_multd_L_summul_n265), .B(
        Inst_f4_multd_L_summul_n264), .ZN(Inst_f4_multd_L_Orig_p[0]) );
  NAND2_X1 Inst_f4_multd_L_summul_U31 ( .A1(Inst_f4_multd_L_sA[2]), .A2(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n264) );
  XNOR2_X1 Inst_f4_multd_L_summul_U30 ( .A(Inst_f4_multd_L_summul_n340), .B(
        Inst_f4_multd_L_summul_n263), .ZN(Inst_f4_multd_L_summul_n265) );
  XNOR2_X1 Inst_f4_multd_L_summul_U29 ( .A(Inst_f4_multd_L_summul_n262), .B(
        Inst_f4_multd_L_summul_n261), .ZN(Inst_f4_multd_L_summul_n263) );
  XNOR2_X1 Inst_f4_multd_L_summul_U28 ( .A(Inst_f4_multd_L_summul_n260), .B(
        Inst_f4_multd_L_summul_n259), .ZN(Inst_f4_multd_L_summul_n261) );
  XNOR2_X1 Inst_f4_multd_L_summul_U27 ( .A(Inst_f4_multd_L_summul_n258), .B(
        Inst_f4_multd_L_summul_n278), .ZN(Inst_f4_multd_L_summul_n259) );
  NAND2_X1 Inst_f4_multd_L_summul_U26 ( .A1(Inst_f4_multd_L_sB[2]), .A2(
        Inst_f4_multd_L_summul_n257), .ZN(Inst_f4_multd_L_summul_n278) );
  XOR2_X1 Inst_f4_multd_L_summul_U25 ( .A(Inst_f4_multd_L_sA[3]), .B(
        Inst_f4_multd_L_sA[5]), .Z(Inst_f4_multd_L_summul_n257) );
  NOR2_X1 Inst_f4_multd_L_summul_U24 ( .A1(Inst_f4_multd_L_summul_n256), .A2(
        Inst_f4_multd_L_summul_n318), .ZN(Inst_f4_multd_L_summul_n258) );
  INV_X1 Inst_f4_multd_L_summul_U23 ( .A(Inst_f4_multd_L_sB[3]), .ZN(
        Inst_f4_multd_L_summul_n318) );
  XNOR2_X1 Inst_f4_multd_L_summul_U22 ( .A(Inst_f4_multd_L_sA[5]), .B(
        Inst_f4_multd_L_sA[4]), .ZN(Inst_f4_multd_L_summul_n256) );
  XNOR2_X1 Inst_f4_multd_L_summul_U21 ( .A(Inst_f4_multd_L_summul_n281), .B(
        Inst_f4_multd_L_sB[4]), .ZN(Inst_f4_multd_L_summul_n260) );
  NAND2_X1 Inst_f4_multd_L_summul_U20 ( .A1(Inst_f4_multd_L_sA[4]), .A2(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n281) );
  NOR2_X1 Inst_f4_multd_L_summul_U19 ( .A1(Inst_f4_multd_L_summul_n325), .A2(
        Inst_f4_multd_L_summul_n307), .ZN(Inst_f4_multd_L_summul_n262) );
  XNOR2_X1 Inst_f4_multd_L_summul_U18 ( .A(Inst_f4_multd_L_sB[4]), .B(
        Inst_f4_multd_L_sB[5]), .ZN(Inst_f4_multd_L_summul_n307) );
  INV_X1 Inst_f4_multd_L_summul_U17 ( .A(Inst_f4_multd_L_sA[3]), .ZN(
        Inst_f4_multd_L_summul_n325) );
  XNOR2_X1 Inst_f4_multd_L_summul_U16 ( .A(Inst_f4_multd_L_summul_n268), .B(
        Inst_f4_multd_L_summul_n255), .ZN(Inst_f4_multd_L_summul_n340) );
  NAND2_X1 Inst_f4_multd_L_summul_U15 ( .A1(Inst_f4_multd_L_sA[2]), .A2(
        Inst_f4_multd_L_sB[2]), .ZN(Inst_f4_multd_L_summul_n255) );
  NAND2_X1 Inst_f4_multd_L_summul_U14 ( .A1(Inst_f4_multd_L_sB[3]), .A2(
        Inst_f4_multd_L_sA[3]), .ZN(Inst_f4_multd_L_summul_n268) );
  XNOR2_X1 Inst_f4_multd_L_summul_U13 ( .A(Inst_f4_multd_L_summul_n340), .B(
        Inst_f4_multd_L_summul_n254), .ZN(Inst_f4_multd_L_Orig_p[5]) );
  XNOR2_X1 Inst_f4_multd_L_summul_U12 ( .A(Inst_f4_multd_L_summul_n253), .B(
        Inst_f4_multd_L_summul_n339), .ZN(Inst_f4_multd_L_summul_n254) );
  XNOR2_X1 Inst_f4_multd_L_summul_U11 ( .A(Inst_f4_multd_L_summul_n250), .B(
        Inst_f4_multd_L_summul_n252), .ZN(Inst_f4_multd_L_summul_n253) );
  NOR2_X1 Inst_f4_multd_L_summul_U10 ( .A1(Inst_f4_multd_L_summul_n338), .A2(
        Inst_f4_multd_L_summul_n251), .ZN(Inst_f4_multd_L_summul_n252) );
  XNOR2_X1 Inst_f4_multd_L_summul_U9 ( .A(Inst_f4_multd_L_sB[2]), .B(
        Inst_f4_multd_L_sB[3]), .ZN(Inst_f4_multd_L_summul_n251) );
  NAND2_X1 Inst_f4_multd_L_summul_U8 ( .A1(Inst_f4_multd_L_summul_n244), .A2(
        Inst_f4_multd_L_summul_n249), .ZN(Inst_f4_multd_L_summul_n250) );
  XOR2_X1 Inst_f4_multd_L_summul_U7 ( .A(Inst_f4_multd_L_summul_n247), .B(
        Inst_f4_multd_L_summul_n248), .Z(Inst_f4_multd_L_summul_n249) );
  NAND2_X1 Inst_f4_multd_L_summul_U6 ( .A1(Inst_f4_multd_L_summul_n245), .A2(
        Inst_f4_multd_L_sA[1]), .ZN(Inst_f4_multd_L_summul_n248) );
  NAND2_X1 Inst_f4_multd_L_summul_U5 ( .A1(Inst_f4_multd_L_sB[0]), .A2(
        Inst_f4_multd_L_summul_n246), .ZN(Inst_f4_multd_L_summul_n247) );
  XOR2_X1 Inst_f4_multd_L_summul_U4 ( .A(Inst_f4_multd_L_sA[3]), .B(
        Inst_f4_multd_L_summul_n336), .Z(Inst_f4_multd_L_summul_n246) );
  NAND2_X1 Inst_f4_multd_L_summul_U3 ( .A1(Inst_f4_multd_L_sB[0]), .A2(
        Inst_f4_multd_L_summul_n337), .ZN(Inst_f4_multd_L_summul_n245) );
  NAND2_X1 Inst_f4_multd_L_summul_U2 ( .A1(Inst_f4_multd_L_sB[1]), .A2(
        Inst_f4_multd_L_summul_n243), .ZN(Inst_f4_multd_L_summul_n244) );
  INV_X1 Inst_f4_multd_L_summul_U1 ( .A(Inst_f4_multd_L_sB[0]), .ZN(
        Inst_f4_multd_L_summul_n243) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_MaskXORInst_U2 ( .A(PRNGQ[44]), .B(
        PRNGQ[46]), .Z(Inst_f4_multd_L_AddNewMaskp_MaskXOR[0]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_MaskXORInst_U1 ( .A(PRNGQ[45]), .B(
        PRNGQ[47]), .Z(Inst_f4_multd_L_AddNewMaskp_MaskXOR[1]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_XORInst1_U2 ( .A(
        Inst_f4_multd_L_Orig_p[4]), .B(Inst_f4_multd_L_AddNewMaskp_MaskXOR[0]), 
        .Z(p_L[4]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_XORInst1_U1 ( .A(
        Inst_f4_multd_L_Orig_p[5]), .B(Inst_f4_multd_L_AddNewMaskp_MaskXOR[1]), 
        .Z(p_L[5]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_XORInst2_U4 ( .A(
        Inst_f4_multd_L_Orig_p[3]), .B(PRNGQ[47]), .Z(p_L[3]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_XORInst2_U3 ( .A(
        Inst_f4_multd_L_Orig_p[2]), .B(PRNGQ[46]), .Z(p_L[2]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_XORInst2_U2 ( .A(
        Inst_f4_multd_L_Orig_p[1]), .B(PRNGQ[45]), .Z(p_L[1]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskp_XORInst2_U1 ( .A(
        Inst_f4_multd_L_Orig_p[0]), .B(PRNGQ[44]), .Z(p_L[0]) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U104 ( .A(Inst_f4_multd_L_lowmul_n336), .B(
        Inst_f4_multd_L_lowmul_n335), .ZN(Inst_f4_multd_L_Orig_pl[4]) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U103 ( .A(Inst_f4_multd_L_lowmul_n334), .B(
        Inst_f4_multd_L_lowmul_n333), .ZN(Inst_f4_multd_L_lowmul_n335) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U102 ( .A(Inst_f4_multd_L_lowmul_n332), .B(
        Inst_f4_multd_L_lowmul_n331), .ZN(Inst_f4_multd_L_lowmul_n333) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U101 ( .A1(Inst_f4_multd_L_lowmul_n330), 
        .A2(FF3_out[28]), .ZN(Inst_f4_multd_L_lowmul_n332) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U100 ( .A1(Inst_f4_multd_L_lowmul_n329), 
        .A2(Inst_f4_multd_L_lowmul_n328), .ZN(Inst_f4_multd_L_lowmul_n334) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U99 ( .A1(FF3_out[0]), .A2(
        Inst_f4_multd_L_lowmul_n327), .ZN(Inst_f4_multd_L_lowmul_n328) );
  OR2_X1 Inst_f4_multd_L_lowmul_U98 ( .A1(Inst_f4_multd_L_lowmul_n327), .A2(
        Inst_f4_multd_L_lowmul_n337), .ZN(Inst_f4_multd_L_lowmul_n329) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U97 ( .A(FF3_out[25]), .B(
        Inst_f4_multd_L_lowmul_n326), .Z(Inst_f4_multd_L_lowmul_n327) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U96 ( .A(Inst_f4_multd_L_lowmul_n325), .B(
        Inst_f4_multd_L_lowmul_n339), .ZN(Inst_f4_multd_L_lowmul_n336) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U95 ( .A(Inst_f4_multd_L_lowmul_n324), .B(
        Inst_f4_multd_L_lowmul_n323), .Z(Inst_f4_multd_L_lowmul_n339) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U94 ( .A1(FF3_out[4]), .A2(FF3_out[25]), 
        .ZN(Inst_f4_multd_L_lowmul_n323) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U93 ( .A1(Inst_f4_multd_L_lowmul_n322), .A2(
        Inst_f4_multd_L_lowmul_n337), .ZN(Inst_f4_multd_L_lowmul_n324) );
  INV_X1 Inst_f4_multd_L_lowmul_U92 ( .A(FF3_out[1]), .ZN(
        Inst_f4_multd_L_lowmul_n337) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U91 ( .A(FF3_out[24]), .B(FF3_out[28]), .ZN(
        Inst_f4_multd_L_lowmul_n322) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U90 ( .A1(Inst_f4_multd_L_lowmul_n321), .A2(
        Inst_f4_multd_L_lowmul_n320), .ZN(Inst_f4_multd_L_lowmul_n325) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U89 ( .A1(FF3_out[25]), .A2(
        Inst_f4_multd_L_lowmul_n319), .ZN(Inst_f4_multd_L_lowmul_n320) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U88 ( .A1(FF3_out[24]), .A2(FF3_out[5]), 
        .ZN(Inst_f4_multd_L_lowmul_n321) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U87 ( .A(Inst_f4_multd_L_lowmul_n318), .B(
        Inst_f4_multd_L_lowmul_n317), .ZN(Inst_f4_multd_L_Orig_pl[3]) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U86 ( .A(Inst_f4_multd_L_lowmul_n316), .B(
        Inst_f4_multd_L_lowmul_n315), .ZN(Inst_f4_multd_L_lowmul_n317) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U85 ( .A(Inst_f4_multd_L_lowmul_n314), .B(
        Inst_f4_multd_L_lowmul_n313), .Z(Inst_f4_multd_L_lowmul_n316) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U84 ( .A1(FF3_out[32]), .A2(FF3_out[8]), 
        .ZN(Inst_f4_multd_L_lowmul_n313) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U83 ( .A1(FF3_out[33]), .A2(FF3_out[9]), 
        .ZN(Inst_f4_multd_L_lowmul_n314) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U82 ( .A(Inst_f4_multd_L_lowmul_n312), .B(
        Inst_f4_multd_L_lowmul_n311), .Z(Inst_f4_multd_L_lowmul_n318) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U81 ( .A(Inst_f4_multd_L_lowmul_n310), .B(
        Inst_f4_multd_L_lowmul_n309), .Z(Inst_f4_multd_L_lowmul_n311) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U80 ( .A1(FF3_out[32]), .A2(
        Inst_f4_multd_L_lowmul_n308), .ZN(Inst_f4_multd_L_lowmul_n309) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U79 ( .A1(FF3_out[24]), .A2(FF3_out[9]), 
        .ZN(Inst_f4_multd_L_lowmul_n310) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U78 ( .A(Inst_f4_multd_L_lowmul_n307), .B(
        Inst_f4_multd_L_lowmul_n306), .ZN(Inst_f4_multd_L_lowmul_n312) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U77 ( .A(FF3_out[33]), .B(
        Inst_f4_multd_L_lowmul_n305), .ZN(Inst_f4_multd_L_lowmul_n306) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U76 ( .A(Inst_f4_multd_L_lowmul_n304), .B(
        Inst_f4_multd_L_lowmul_n303), .Z(Inst_f4_multd_L_lowmul_n305) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U75 ( .A1(FF3_out[0]), .A2(FF3_out[32]), 
        .ZN(Inst_f4_multd_L_lowmul_n303) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U74 ( .A1(Inst_f4_multd_L_lowmul_n302), .A2(
        FF3_out[1]), .ZN(Inst_f4_multd_L_lowmul_n304) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U73 ( .A1(Inst_f4_multd_L_lowmul_n301), .A2(
        FF3_out[8]), .ZN(Inst_f4_multd_L_lowmul_n307) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U72 ( .A(Inst_f4_multd_L_lowmul_n338), .B(
        Inst_f4_multd_L_lowmul_n300), .ZN(Inst_f4_multd_L_lowmul_n301) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U71 ( .A(FF3_out[25]), .B(
        Inst_f4_multd_L_lowmul_n299), .ZN(Inst_f4_multd_L_lowmul_n300) );
  INV_X1 Inst_f4_multd_L_lowmul_U70 ( .A(FF3_out[24]), .ZN(
        Inst_f4_multd_L_lowmul_n338) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U69 ( .A(Inst_f4_multd_L_lowmul_n298), .B(
        Inst_f4_multd_L_lowmul_n297), .Z(Inst_f4_multd_L_Orig_pl[2]) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U68 ( .A1(Inst_f4_multd_L_lowmul_n296), .A2(
        Inst_f4_multd_L_lowmul_n295), .ZN(Inst_f4_multd_L_lowmul_n297) );
  OR2_X1 Inst_f4_multd_L_lowmul_U67 ( .A1(FF3_out[9]), .A2(
        Inst_f4_multd_L_lowmul_n302), .ZN(Inst_f4_multd_L_lowmul_n295) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U66 ( .A1(Inst_f4_multd_L_lowmul_n294), .A2(
        FF3_out[9]), .ZN(Inst_f4_multd_L_lowmul_n296) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U65 ( .A(Inst_f4_multd_L_lowmul_n293), .B(
        FF3_out[24]), .ZN(Inst_f4_multd_L_lowmul_n294) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U64 ( .A(Inst_f4_multd_L_lowmul_n292), .B(
        Inst_f4_multd_L_lowmul_n291), .Z(Inst_f4_multd_L_lowmul_n298) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U63 ( .A1(Inst_f4_multd_L_lowmul_n299), .A2(
        Inst_f4_multd_L_lowmul_n290), .ZN(Inst_f4_multd_L_lowmul_n291) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U62 ( .A(Inst_f4_multd_L_lowmul_n308), .B(
        FF3_out[1]), .Z(Inst_f4_multd_L_lowmul_n290) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U61 ( .A(Inst_f4_multd_L_lowmul_n289), .B(
        Inst_f4_multd_L_lowmul_n288), .ZN(Inst_f4_multd_L_lowmul_n292) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U60 ( .A(FF3_out[0]), .B(
        Inst_f4_multd_L_lowmul_n331), .ZN(Inst_f4_multd_L_lowmul_n288) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U59 ( .A(Inst_f4_multd_L_lowmul_n287), .B(
        Inst_f4_multd_L_lowmul_n286), .Z(Inst_f4_multd_L_lowmul_n331) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U58 ( .A1(FF3_out[25]), .A2(FF3_out[0]), 
        .ZN(Inst_f4_multd_L_lowmul_n286) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U57 ( .A1(FF3_out[24]), .A2(FF3_out[1]), 
        .ZN(Inst_f4_multd_L_lowmul_n287) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U56 ( .A(Inst_f4_multd_L_lowmul_n285), .B(
        Inst_f4_multd_L_lowmul_n315), .Z(Inst_f4_multd_L_lowmul_n289) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U55 ( .A(Inst_f4_multd_L_lowmul_n284), .B(
        Inst_f4_multd_L_lowmul_n283), .Z(Inst_f4_multd_L_lowmul_n315) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U54 ( .A1(FF3_out[32]), .A2(FF3_out[1]), 
        .ZN(Inst_f4_multd_L_lowmul_n283) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U53 ( .A1(FF3_out[33]), .A2(FF3_out[0]), 
        .ZN(Inst_f4_multd_L_lowmul_n284) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U52 ( .A(Inst_f4_multd_L_lowmul_n282), .B(
        Inst_f4_multd_L_lowmul_n281), .Z(Inst_f4_multd_L_lowmul_n285) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U51 ( .A1(FF3_out[8]), .A2(
        Inst_f4_multd_L_lowmul_n302), .ZN(Inst_f4_multd_L_lowmul_n281) );
  INV_X1 Inst_f4_multd_L_lowmul_U50 ( .A(FF3_out[25]), .ZN(
        Inst_f4_multd_L_lowmul_n302) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U49 ( .A(Inst_f4_multd_L_lowmul_n280), .B(
        Inst_f4_multd_L_lowmul_n279), .ZN(Inst_f4_multd_L_Orig_pl[1]) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U48 ( .A(Inst_f4_multd_L_lowmul_n278), .B(
        Inst_f4_multd_L_lowmul_n277), .ZN(Inst_f4_multd_L_lowmul_n280) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U47 ( .A1(Inst_f4_multd_L_lowmul_n276), .A2(
        FF3_out[28]), .ZN(Inst_f4_multd_L_lowmul_n277) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U46 ( .A(FF3_out[4]), .B(
        Inst_f4_multd_L_lowmul_n308), .ZN(Inst_f4_multd_L_lowmul_n276) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U45 ( .A(Inst_f4_multd_L_lowmul_n275), .B(
        Inst_f4_multd_L_lowmul_n274), .ZN(Inst_f4_multd_L_lowmul_n278) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U44 ( .A(Inst_f4_multd_L_lowmul_n273), .B(
        Inst_f4_multd_L_lowmul_n272), .ZN(Inst_f4_multd_L_lowmul_n274) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U43 ( .A1(Inst_f4_multd_L_lowmul_n271), .A2(
        Inst_f4_multd_L_lowmul_n330), .ZN(Inst_f4_multd_L_lowmul_n272) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U42 ( .A(FF3_out[4]), .B(FF3_out[5]), .Z(
        Inst_f4_multd_L_lowmul_n330) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U41 ( .A(FF3_out[28]), .B(FF3_out[32]), .Z(
        Inst_f4_multd_L_lowmul_n271) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U40 ( .A1(FF3_out[29]), .A2(FF3_out[8]), 
        .ZN(Inst_f4_multd_L_lowmul_n273) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U39 ( .A(Inst_f4_multd_L_lowmul_n270), .B(
        Inst_f4_multd_L_lowmul_n269), .ZN(Inst_f4_multd_L_lowmul_n275) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U38 ( .A(Inst_f4_multd_L_lowmul_n268), .B(
        Inst_f4_multd_L_lowmul_n267), .Z(Inst_f4_multd_L_lowmul_n270) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U37 ( .A1(Inst_f4_multd_L_lowmul_n293), .A2(
        FF3_out[8]), .ZN(Inst_f4_multd_L_lowmul_n267) );
  INV_X1 Inst_f4_multd_L_lowmul_U36 ( .A(FF3_out[32]), .ZN(
        Inst_f4_multd_L_lowmul_n293) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U35 ( .A1(Inst_f4_multd_L_lowmul_n299), .A2(
        FF3_out[9]), .ZN(Inst_f4_multd_L_lowmul_n268) );
  INV_X1 Inst_f4_multd_L_lowmul_U34 ( .A(FF3_out[33]), .ZN(
        Inst_f4_multd_L_lowmul_n299) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U33 ( .A(Inst_f4_multd_L_lowmul_n266), .B(
        Inst_f4_multd_L_lowmul_n265), .ZN(Inst_f4_multd_L_Orig_pl[0]) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U32 ( .A1(FF3_out[28]), .A2(FF3_out[9]), 
        .ZN(Inst_f4_multd_L_lowmul_n265) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U31 ( .A(Inst_f4_multd_L_lowmul_n340), .B(
        Inst_f4_multd_L_lowmul_n264), .ZN(Inst_f4_multd_L_lowmul_n266) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U30 ( .A(Inst_f4_multd_L_lowmul_n263), .B(
        Inst_f4_multd_L_lowmul_n262), .ZN(Inst_f4_multd_L_lowmul_n264) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U29 ( .A(Inst_f4_multd_L_lowmul_n261), .B(
        Inst_f4_multd_L_lowmul_n260), .ZN(Inst_f4_multd_L_lowmul_n262) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U28 ( .A(Inst_f4_multd_L_lowmul_n259), .B(
        Inst_f4_multd_L_lowmul_n279), .ZN(Inst_f4_multd_L_lowmul_n260) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U27 ( .A1(FF3_out[4]), .A2(
        Inst_f4_multd_L_lowmul_n258), .ZN(Inst_f4_multd_L_lowmul_n279) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U26 ( .A(FF3_out[29]), .B(FF3_out[33]), .Z(
        Inst_f4_multd_L_lowmul_n258) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U25 ( .A1(Inst_f4_multd_L_lowmul_n257), .A2(
        Inst_f4_multd_L_lowmul_n319), .ZN(Inst_f4_multd_L_lowmul_n259) );
  INV_X1 Inst_f4_multd_L_lowmul_U24 ( .A(FF3_out[5]), .ZN(
        Inst_f4_multd_L_lowmul_n319) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U23 ( .A(FF3_out[33]), .B(FF3_out[32]), .ZN(
        Inst_f4_multd_L_lowmul_n257) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U22 ( .A(Inst_f4_multd_L_lowmul_n282), .B(
        FF3_out[8]), .ZN(Inst_f4_multd_L_lowmul_n261) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U21 ( .A1(FF3_out[32]), .A2(FF3_out[9]), 
        .ZN(Inst_f4_multd_L_lowmul_n282) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U20 ( .A1(Inst_f4_multd_L_lowmul_n326), .A2(
        Inst_f4_multd_L_lowmul_n308), .ZN(Inst_f4_multd_L_lowmul_n263) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U19 ( .A(FF3_out[8]), .B(FF3_out[9]), .ZN(
        Inst_f4_multd_L_lowmul_n308) );
  INV_X1 Inst_f4_multd_L_lowmul_U18 ( .A(FF3_out[29]), .ZN(
        Inst_f4_multd_L_lowmul_n326) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U17 ( .A(Inst_f4_multd_L_lowmul_n269), .B(
        Inst_f4_multd_L_lowmul_n256), .ZN(Inst_f4_multd_L_lowmul_n340) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U16 ( .A1(FF3_out[28]), .A2(FF3_out[4]), 
        .ZN(Inst_f4_multd_L_lowmul_n256) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U15 ( .A1(FF3_out[5]), .A2(FF3_out[29]), 
        .ZN(Inst_f4_multd_L_lowmul_n269) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U14 ( .A(Inst_f4_multd_L_lowmul_n255), .B(
        Inst_f4_multd_L_lowmul_n340), .Z(Inst_f4_multd_L_Orig_pl[5]) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U13 ( .A(Inst_f4_multd_L_lowmul_n254), .B(
        Inst_f4_multd_L_lowmul_n252), .ZN(Inst_f4_multd_L_lowmul_n255) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U12 ( .A1(Inst_f4_multd_L_lowmul_n253), .A2(
        Inst_f4_multd_L_lowmul_n249), .ZN(Inst_f4_multd_L_lowmul_n254) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U11 ( .A1(Inst_f4_multd_L_lowmul_n243), .A2(
        FF3_out[1]), .ZN(Inst_f4_multd_L_lowmul_n253) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U10 ( .A(Inst_f4_multd_L_lowmul_n251), .B(
        Inst_f4_multd_L_lowmul_n339), .Z(Inst_f4_multd_L_lowmul_n252) );
  NOR2_X1 Inst_f4_multd_L_lowmul_U9 ( .A1(Inst_f4_multd_L_lowmul_n338), .A2(
        Inst_f4_multd_L_lowmul_n250), .ZN(Inst_f4_multd_L_lowmul_n251) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U8 ( .A(FF3_out[4]), .B(FF3_out[5]), .ZN(
        Inst_f4_multd_L_lowmul_n250) );
  XOR2_X1 Inst_f4_multd_L_lowmul_U7 ( .A(Inst_f4_multd_L_lowmul_n246), .B(
        Inst_f4_multd_L_lowmul_n248), .Z(Inst_f4_multd_L_lowmul_n249) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U6 ( .A1(Inst_f4_multd_L_lowmul_n247), .A2(
        FF3_out[25]), .ZN(Inst_f4_multd_L_lowmul_n248) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U5 ( .A1(FF3_out[0]), .A2(
        Inst_f4_multd_L_lowmul_n337), .ZN(Inst_f4_multd_L_lowmul_n247) );
  NAND2_X1 Inst_f4_multd_L_lowmul_U4 ( .A1(FF3_out[0]), .A2(
        Inst_f4_multd_L_lowmul_n245), .ZN(Inst_f4_multd_L_lowmul_n246) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U3 ( .A(Inst_f4_multd_L_lowmul_n244), .B(
        FF3_out[28]), .ZN(Inst_f4_multd_L_lowmul_n245) );
  XNOR2_X1 Inst_f4_multd_L_lowmul_U2 ( .A(FF3_out[24]), .B(FF3_out[29]), .ZN(
        Inst_f4_multd_L_lowmul_n244) );
  INV_X1 Inst_f4_multd_L_lowmul_U1 ( .A(FF3_out[0]), .ZN(
        Inst_f4_multd_L_lowmul_n243) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_MaskXORInst_U2 ( .A(PRNGQ[48]), .B(
        PRNGQ[50]), .Z(Inst_f4_multd_L_AddNewMaskpl_MaskXOR[0]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_MaskXORInst_U1 ( .A(PRNGQ[49]), .B(
        PRNGQ[51]), .Z(Inst_f4_multd_L_AddNewMaskpl_MaskXOR[1]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_XORInst1_U2 ( .A(
        Inst_f4_multd_L_Orig_pl[4]), .B(
        Inst_f4_multd_L_AddNewMaskpl_MaskXOR[0]), .Z(pl_L[4]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_XORInst1_U1 ( .A(
        Inst_f4_multd_L_Orig_pl[5]), .B(
        Inst_f4_multd_L_AddNewMaskpl_MaskXOR[1]), .Z(pl_L[5]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_XORInst2_U4 ( .A(
        Inst_f4_multd_L_Orig_pl[3]), .B(PRNGQ[51]), .Z(pl_L[3]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_XORInst2_U3 ( .A(
        Inst_f4_multd_L_Orig_pl[2]), .B(PRNGQ[50]), .Z(pl_L[2]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_XORInst2_U2 ( .A(
        Inst_f4_multd_L_Orig_pl[1]), .B(PRNGQ[49]), .Z(pl_L[1]) );
  XOR2_X1 Inst_f4_multd_L_AddNewMaskpl_XORInst2_U1 ( .A(
        Inst_f4_multd_L_Orig_pl[0]), .B(PRNGQ[48]), .Z(pl_L[0]) );
  XOR2_X1 Inst_f4_multd_H_U12 ( .A(FF3_out[23]), .B(FF3_out[21]), .Z(
        Inst_f4_multd_H_sB[5]) );
  XOR2_X1 Inst_f4_multd_H_U11 ( .A(FF3_out[22]), .B(FF3_out[20]), .Z(
        Inst_f4_multd_H_sB[4]) );
  XOR2_X1 Inst_f4_multd_H_U10 ( .A(FF3_out[17]), .B(FF3_out[19]), .Z(
        Inst_f4_multd_H_sB[3]) );
  XOR2_X1 Inst_f4_multd_H_U9 ( .A(FF3_out[16]), .B(FF3_out[18]), .Z(
        Inst_f4_multd_H_sB[2]) );
  XOR2_X1 Inst_f4_multd_H_U8 ( .A(FF3_out[13]), .B(FF3_out[15]), .Z(
        Inst_f4_multd_H_sB[1]) );
  XOR2_X1 Inst_f4_multd_H_U7 ( .A(FF3_out[12]), .B(FF3_out[14]), .Z(
        Inst_f4_multd_H_sB[0]) );
  XOR2_X1 Inst_f4_multd_H_U6 ( .A(FF3_out[11]), .B(FF3_out[9]), .Z(
        Inst_f4_multd_H_sA[5]) );
  XOR2_X1 Inst_f4_multd_H_U5 ( .A(FF3_out[10]), .B(FF3_out[8]), .Z(
        Inst_f4_multd_H_sA[4]) );
  XOR2_X1 Inst_f4_multd_H_U4 ( .A(FF3_out[5]), .B(FF3_out[7]), .Z(
        Inst_f4_multd_H_sA[3]) );
  XOR2_X1 Inst_f4_multd_H_U3 ( .A(FF3_out[4]), .B(FF3_out[6]), .Z(
        Inst_f4_multd_H_sA[2]) );
  XOR2_X1 Inst_f4_multd_H_U2 ( .A(FF3_out[1]), .B(FF3_out[3]), .Z(
        Inst_f4_multd_H_sA[1]) );
  XOR2_X1 Inst_f4_multd_H_U1 ( .A(FF3_out[0]), .B(FF3_out[2]), .Z(
        Inst_f4_multd_H_sA[0]) );
  XNOR2_X1 Inst_f4_multd_H_himul_U104 ( .A(Inst_f4_multd_H_himul_n336), .B(
        Inst_f4_multd_H_himul_n335), .ZN(Inst_f4_multd_H_Orig_ph[4]) );
  XNOR2_X1 Inst_f4_multd_H_himul_U103 ( .A(Inst_f4_multd_H_himul_n334), .B(
        Inst_f4_multd_H_himul_n333), .ZN(Inst_f4_multd_H_himul_n335) );
  XNOR2_X1 Inst_f4_multd_H_himul_U102 ( .A(Inst_f4_multd_H_himul_n332), .B(
        Inst_f4_multd_H_himul_n331), .ZN(Inst_f4_multd_H_himul_n333) );
  NAND2_X1 Inst_f4_multd_H_himul_U101 ( .A1(Inst_f4_multd_H_himul_n330), .A2(
        FF3_out[6]), .ZN(Inst_f4_multd_H_himul_n332) );
  NAND2_X1 Inst_f4_multd_H_himul_U100 ( .A1(Inst_f4_multd_H_himul_n329), .A2(
        Inst_f4_multd_H_himul_n328), .ZN(Inst_f4_multd_H_himul_n334) );
  NAND2_X1 Inst_f4_multd_H_himul_U99 ( .A1(FF3_out[14]), .A2(
        Inst_f4_multd_H_himul_n327), .ZN(Inst_f4_multd_H_himul_n328) );
  OR2_X1 Inst_f4_multd_H_himul_U98 ( .A1(Inst_f4_multd_H_himul_n327), .A2(
        Inst_f4_multd_H_himul_n337), .ZN(Inst_f4_multd_H_himul_n329) );
  XOR2_X1 Inst_f4_multd_H_himul_U97 ( .A(FF3_out[3]), .B(
        Inst_f4_multd_H_himul_n326), .Z(Inst_f4_multd_H_himul_n327) );
  XNOR2_X1 Inst_f4_multd_H_himul_U96 ( .A(Inst_f4_multd_H_himul_n325), .B(
        Inst_f4_multd_H_himul_n339), .ZN(Inst_f4_multd_H_himul_n336) );
  XOR2_X1 Inst_f4_multd_H_himul_U95 ( .A(Inst_f4_multd_H_himul_n324), .B(
        Inst_f4_multd_H_himul_n323), .Z(Inst_f4_multd_H_himul_n339) );
  NAND2_X1 Inst_f4_multd_H_himul_U94 ( .A1(FF3_out[18]), .A2(FF3_out[3]), .ZN(
        Inst_f4_multd_H_himul_n323) );
  NOR2_X1 Inst_f4_multd_H_himul_U93 ( .A1(Inst_f4_multd_H_himul_n322), .A2(
        Inst_f4_multd_H_himul_n337), .ZN(Inst_f4_multd_H_himul_n324) );
  INV_X1 Inst_f4_multd_H_himul_U92 ( .A(FF3_out[15]), .ZN(
        Inst_f4_multd_H_himul_n337) );
  XNOR2_X1 Inst_f4_multd_H_himul_U91 ( .A(FF3_out[2]), .B(FF3_out[6]), .ZN(
        Inst_f4_multd_H_himul_n322) );
  NAND2_X1 Inst_f4_multd_H_himul_U90 ( .A1(Inst_f4_multd_H_himul_n321), .A2(
        Inst_f4_multd_H_himul_n320), .ZN(Inst_f4_multd_H_himul_n325) );
  NAND2_X1 Inst_f4_multd_H_himul_U89 ( .A1(FF3_out[3]), .A2(
        Inst_f4_multd_H_himul_n319), .ZN(Inst_f4_multd_H_himul_n320) );
  NAND2_X1 Inst_f4_multd_H_himul_U88 ( .A1(FF3_out[2]), .A2(FF3_out[19]), .ZN(
        Inst_f4_multd_H_himul_n321) );
  XNOR2_X1 Inst_f4_multd_H_himul_U87 ( .A(Inst_f4_multd_H_himul_n318), .B(
        Inst_f4_multd_H_himul_n317), .ZN(Inst_f4_multd_H_Orig_ph[3]) );
  XNOR2_X1 Inst_f4_multd_H_himul_U86 ( .A(Inst_f4_multd_H_himul_n316), .B(
        Inst_f4_multd_H_himul_n315), .ZN(Inst_f4_multd_H_himul_n317) );
  XOR2_X1 Inst_f4_multd_H_himul_U85 ( .A(Inst_f4_multd_H_himul_n314), .B(
        Inst_f4_multd_H_himul_n313), .Z(Inst_f4_multd_H_himul_n316) );
  NAND2_X1 Inst_f4_multd_H_himul_U84 ( .A1(FF3_out[10]), .A2(FF3_out[22]), 
        .ZN(Inst_f4_multd_H_himul_n313) );
  NAND2_X1 Inst_f4_multd_H_himul_U83 ( .A1(FF3_out[11]), .A2(FF3_out[23]), 
        .ZN(Inst_f4_multd_H_himul_n314) );
  XOR2_X1 Inst_f4_multd_H_himul_U82 ( .A(Inst_f4_multd_H_himul_n312), .B(
        Inst_f4_multd_H_himul_n311), .Z(Inst_f4_multd_H_himul_n318) );
  XOR2_X1 Inst_f4_multd_H_himul_U81 ( .A(Inst_f4_multd_H_himul_n310), .B(
        Inst_f4_multd_H_himul_n309), .Z(Inst_f4_multd_H_himul_n311) );
  NAND2_X1 Inst_f4_multd_H_himul_U80 ( .A1(FF3_out[10]), .A2(
        Inst_f4_multd_H_himul_n308), .ZN(Inst_f4_multd_H_himul_n309) );
  NAND2_X1 Inst_f4_multd_H_himul_U79 ( .A1(FF3_out[2]), .A2(FF3_out[23]), .ZN(
        Inst_f4_multd_H_himul_n310) );
  XNOR2_X1 Inst_f4_multd_H_himul_U78 ( .A(Inst_f4_multd_H_himul_n307), .B(
        Inst_f4_multd_H_himul_n306), .ZN(Inst_f4_multd_H_himul_n312) );
  XNOR2_X1 Inst_f4_multd_H_himul_U77 ( .A(FF3_out[11]), .B(
        Inst_f4_multd_H_himul_n305), .ZN(Inst_f4_multd_H_himul_n306) );
  XOR2_X1 Inst_f4_multd_H_himul_U76 ( .A(Inst_f4_multd_H_himul_n304), .B(
        Inst_f4_multd_H_himul_n303), .Z(Inst_f4_multd_H_himul_n305) );
  NAND2_X1 Inst_f4_multd_H_himul_U75 ( .A1(FF3_out[14]), .A2(FF3_out[10]), 
        .ZN(Inst_f4_multd_H_himul_n303) );
  NOR2_X1 Inst_f4_multd_H_himul_U74 ( .A1(Inst_f4_multd_H_himul_n302), .A2(
        FF3_out[15]), .ZN(Inst_f4_multd_H_himul_n304) );
  NAND2_X1 Inst_f4_multd_H_himul_U73 ( .A1(Inst_f4_multd_H_himul_n301), .A2(
        FF3_out[22]), .ZN(Inst_f4_multd_H_himul_n307) );
  XNOR2_X1 Inst_f4_multd_H_himul_U72 ( .A(Inst_f4_multd_H_himul_n338), .B(
        Inst_f4_multd_H_himul_n300), .ZN(Inst_f4_multd_H_himul_n301) );
  XNOR2_X1 Inst_f4_multd_H_himul_U71 ( .A(FF3_out[3]), .B(
        Inst_f4_multd_H_himul_n299), .ZN(Inst_f4_multd_H_himul_n300) );
  INV_X1 Inst_f4_multd_H_himul_U70 ( .A(FF3_out[2]), .ZN(
        Inst_f4_multd_H_himul_n338) );
  XOR2_X1 Inst_f4_multd_H_himul_U69 ( .A(Inst_f4_multd_H_himul_n298), .B(
        Inst_f4_multd_H_himul_n297), .Z(Inst_f4_multd_H_Orig_ph[2]) );
  NAND2_X1 Inst_f4_multd_H_himul_U68 ( .A1(Inst_f4_multd_H_himul_n296), .A2(
        Inst_f4_multd_H_himul_n295), .ZN(Inst_f4_multd_H_himul_n297) );
  OR2_X1 Inst_f4_multd_H_himul_U67 ( .A1(FF3_out[23]), .A2(
        Inst_f4_multd_H_himul_n302), .ZN(Inst_f4_multd_H_himul_n295) );
  NAND2_X1 Inst_f4_multd_H_himul_U66 ( .A1(Inst_f4_multd_H_himul_n294), .A2(
        FF3_out[23]), .ZN(Inst_f4_multd_H_himul_n296) );
  XNOR2_X1 Inst_f4_multd_H_himul_U65 ( .A(Inst_f4_multd_H_himul_n293), .B(
        FF3_out[2]), .ZN(Inst_f4_multd_H_himul_n294) );
  XOR2_X1 Inst_f4_multd_H_himul_U64 ( .A(Inst_f4_multd_H_himul_n292), .B(
        Inst_f4_multd_H_himul_n291), .Z(Inst_f4_multd_H_himul_n298) );
  NOR2_X1 Inst_f4_multd_H_himul_U63 ( .A1(Inst_f4_multd_H_himul_n299), .A2(
        Inst_f4_multd_H_himul_n290), .ZN(Inst_f4_multd_H_himul_n291) );
  XOR2_X1 Inst_f4_multd_H_himul_U62 ( .A(Inst_f4_multd_H_himul_n308), .B(
        FF3_out[15]), .Z(Inst_f4_multd_H_himul_n290) );
  XNOR2_X1 Inst_f4_multd_H_himul_U61 ( .A(Inst_f4_multd_H_himul_n289), .B(
        Inst_f4_multd_H_himul_n288), .ZN(Inst_f4_multd_H_himul_n292) );
  XNOR2_X1 Inst_f4_multd_H_himul_U60 ( .A(FF3_out[14]), .B(
        Inst_f4_multd_H_himul_n331), .ZN(Inst_f4_multd_H_himul_n288) );
  XOR2_X1 Inst_f4_multd_H_himul_U59 ( .A(Inst_f4_multd_H_himul_n287), .B(
        Inst_f4_multd_H_himul_n286), .Z(Inst_f4_multd_H_himul_n331) );
  NAND2_X1 Inst_f4_multd_H_himul_U58 ( .A1(FF3_out[3]), .A2(FF3_out[14]), .ZN(
        Inst_f4_multd_H_himul_n286) );
  NAND2_X1 Inst_f4_multd_H_himul_U57 ( .A1(FF3_out[2]), .A2(FF3_out[15]), .ZN(
        Inst_f4_multd_H_himul_n287) );
  XOR2_X1 Inst_f4_multd_H_himul_U56 ( .A(Inst_f4_multd_H_himul_n285), .B(
        Inst_f4_multd_H_himul_n315), .Z(Inst_f4_multd_H_himul_n289) );
  XOR2_X1 Inst_f4_multd_H_himul_U55 ( .A(Inst_f4_multd_H_himul_n284), .B(
        Inst_f4_multd_H_himul_n283), .Z(Inst_f4_multd_H_himul_n315) );
  NAND2_X1 Inst_f4_multd_H_himul_U54 ( .A1(FF3_out[10]), .A2(FF3_out[15]), 
        .ZN(Inst_f4_multd_H_himul_n283) );
  NAND2_X1 Inst_f4_multd_H_himul_U53 ( .A1(FF3_out[11]), .A2(FF3_out[14]), 
        .ZN(Inst_f4_multd_H_himul_n284) );
  XOR2_X1 Inst_f4_multd_H_himul_U52 ( .A(Inst_f4_multd_H_himul_n282), .B(
        Inst_f4_multd_H_himul_n281), .Z(Inst_f4_multd_H_himul_n285) );
  NAND2_X1 Inst_f4_multd_H_himul_U51 ( .A1(FF3_out[22]), .A2(
        Inst_f4_multd_H_himul_n302), .ZN(Inst_f4_multd_H_himul_n281) );
  INV_X1 Inst_f4_multd_H_himul_U50 ( .A(FF3_out[3]), .ZN(
        Inst_f4_multd_H_himul_n302) );
  XNOR2_X1 Inst_f4_multd_H_himul_U49 ( .A(Inst_f4_multd_H_himul_n280), .B(
        Inst_f4_multd_H_himul_n279), .ZN(Inst_f4_multd_H_Orig_ph[1]) );
  XNOR2_X1 Inst_f4_multd_H_himul_U48 ( .A(Inst_f4_multd_H_himul_n278), .B(
        Inst_f4_multd_H_himul_n277), .ZN(Inst_f4_multd_H_himul_n280) );
  NAND2_X1 Inst_f4_multd_H_himul_U47 ( .A1(Inst_f4_multd_H_himul_n276), .A2(
        FF3_out[6]), .ZN(Inst_f4_multd_H_himul_n277) );
  XNOR2_X1 Inst_f4_multd_H_himul_U46 ( .A(FF3_out[18]), .B(
        Inst_f4_multd_H_himul_n308), .ZN(Inst_f4_multd_H_himul_n276) );
  XNOR2_X1 Inst_f4_multd_H_himul_U45 ( .A(Inst_f4_multd_H_himul_n275), .B(
        Inst_f4_multd_H_himul_n274), .ZN(Inst_f4_multd_H_himul_n278) );
  XNOR2_X1 Inst_f4_multd_H_himul_U44 ( .A(Inst_f4_multd_H_himul_n273), .B(
        Inst_f4_multd_H_himul_n272), .ZN(Inst_f4_multd_H_himul_n274) );
  NAND2_X1 Inst_f4_multd_H_himul_U43 ( .A1(Inst_f4_multd_H_himul_n271), .A2(
        Inst_f4_multd_H_himul_n330), .ZN(Inst_f4_multd_H_himul_n272) );
  XOR2_X1 Inst_f4_multd_H_himul_U42 ( .A(FF3_out[18]), .B(FF3_out[19]), .Z(
        Inst_f4_multd_H_himul_n330) );
  XOR2_X1 Inst_f4_multd_H_himul_U41 ( .A(FF3_out[6]), .B(FF3_out[10]), .Z(
        Inst_f4_multd_H_himul_n271) );
  NAND2_X1 Inst_f4_multd_H_himul_U40 ( .A1(FF3_out[7]), .A2(FF3_out[22]), .ZN(
        Inst_f4_multd_H_himul_n273) );
  XNOR2_X1 Inst_f4_multd_H_himul_U39 ( .A(Inst_f4_multd_H_himul_n270), .B(
        Inst_f4_multd_H_himul_n269), .ZN(Inst_f4_multd_H_himul_n275) );
  XOR2_X1 Inst_f4_multd_H_himul_U38 ( .A(Inst_f4_multd_H_himul_n268), .B(
        Inst_f4_multd_H_himul_n267), .Z(Inst_f4_multd_H_himul_n270) );
  NOR2_X1 Inst_f4_multd_H_himul_U37 ( .A1(Inst_f4_multd_H_himul_n293), .A2(
        FF3_out[22]), .ZN(Inst_f4_multd_H_himul_n267) );
  INV_X1 Inst_f4_multd_H_himul_U36 ( .A(FF3_out[10]), .ZN(
        Inst_f4_multd_H_himul_n293) );
  NOR2_X1 Inst_f4_multd_H_himul_U35 ( .A1(Inst_f4_multd_H_himul_n299), .A2(
        FF3_out[23]), .ZN(Inst_f4_multd_H_himul_n268) );
  INV_X1 Inst_f4_multd_H_himul_U34 ( .A(FF3_out[11]), .ZN(
        Inst_f4_multd_H_himul_n299) );
  XNOR2_X1 Inst_f4_multd_H_himul_U33 ( .A(Inst_f4_multd_H_himul_n266), .B(
        Inst_f4_multd_H_himul_n265), .ZN(Inst_f4_multd_H_Orig_ph[0]) );
  NAND2_X1 Inst_f4_multd_H_himul_U32 ( .A1(FF3_out[6]), .A2(FF3_out[23]), .ZN(
        Inst_f4_multd_H_himul_n265) );
  XNOR2_X1 Inst_f4_multd_H_himul_U31 ( .A(Inst_f4_multd_H_himul_n340), .B(
        Inst_f4_multd_H_himul_n264), .ZN(Inst_f4_multd_H_himul_n266) );
  XNOR2_X1 Inst_f4_multd_H_himul_U30 ( .A(Inst_f4_multd_H_himul_n263), .B(
        Inst_f4_multd_H_himul_n262), .ZN(Inst_f4_multd_H_himul_n264) );
  XNOR2_X1 Inst_f4_multd_H_himul_U29 ( .A(Inst_f4_multd_H_himul_n261), .B(
        Inst_f4_multd_H_himul_n260), .ZN(Inst_f4_multd_H_himul_n262) );
  XNOR2_X1 Inst_f4_multd_H_himul_U28 ( .A(Inst_f4_multd_H_himul_n259), .B(
        Inst_f4_multd_H_himul_n279), .ZN(Inst_f4_multd_H_himul_n260) );
  NAND2_X1 Inst_f4_multd_H_himul_U27 ( .A1(FF3_out[18]), .A2(
        Inst_f4_multd_H_himul_n258), .ZN(Inst_f4_multd_H_himul_n279) );
  XOR2_X1 Inst_f4_multd_H_himul_U26 ( .A(FF3_out[7]), .B(FF3_out[11]), .Z(
        Inst_f4_multd_H_himul_n258) );
  NOR2_X1 Inst_f4_multd_H_himul_U25 ( .A1(Inst_f4_multd_H_himul_n257), .A2(
        Inst_f4_multd_H_himul_n319), .ZN(Inst_f4_multd_H_himul_n259) );
  INV_X1 Inst_f4_multd_H_himul_U24 ( .A(FF3_out[19]), .ZN(
        Inst_f4_multd_H_himul_n319) );
  XNOR2_X1 Inst_f4_multd_H_himul_U23 ( .A(FF3_out[11]), .B(FF3_out[10]), .ZN(
        Inst_f4_multd_H_himul_n257) );
  XNOR2_X1 Inst_f4_multd_H_himul_U22 ( .A(Inst_f4_multd_H_himul_n282), .B(
        FF3_out[22]), .ZN(Inst_f4_multd_H_himul_n261) );
  NAND2_X1 Inst_f4_multd_H_himul_U21 ( .A1(FF3_out[10]), .A2(FF3_out[23]), 
        .ZN(Inst_f4_multd_H_himul_n282) );
  NOR2_X1 Inst_f4_multd_H_himul_U20 ( .A1(Inst_f4_multd_H_himul_n326), .A2(
        Inst_f4_multd_H_himul_n308), .ZN(Inst_f4_multd_H_himul_n263) );
  XNOR2_X1 Inst_f4_multd_H_himul_U19 ( .A(FF3_out[22]), .B(FF3_out[23]), .ZN(
        Inst_f4_multd_H_himul_n308) );
  INV_X1 Inst_f4_multd_H_himul_U18 ( .A(FF3_out[7]), .ZN(
        Inst_f4_multd_H_himul_n326) );
  XNOR2_X1 Inst_f4_multd_H_himul_U17 ( .A(Inst_f4_multd_H_himul_n269), .B(
        Inst_f4_multd_H_himul_n256), .ZN(Inst_f4_multd_H_himul_n340) );
  NAND2_X1 Inst_f4_multd_H_himul_U16 ( .A1(FF3_out[6]), .A2(FF3_out[18]), .ZN(
        Inst_f4_multd_H_himul_n256) );
  NAND2_X1 Inst_f4_multd_H_himul_U15 ( .A1(FF3_out[19]), .A2(FF3_out[7]), .ZN(
        Inst_f4_multd_H_himul_n269) );
  XOR2_X1 Inst_f4_multd_H_himul_U14 ( .A(Inst_f4_multd_H_himul_n255), .B(
        Inst_f4_multd_H_himul_n340), .Z(Inst_f4_multd_H_Orig_ph[5]) );
  XNOR2_X1 Inst_f4_multd_H_himul_U13 ( .A(Inst_f4_multd_H_himul_n254), .B(
        Inst_f4_multd_H_himul_n252), .ZN(Inst_f4_multd_H_himul_n255) );
  NAND2_X1 Inst_f4_multd_H_himul_U12 ( .A1(Inst_f4_multd_H_himul_n253), .A2(
        Inst_f4_multd_H_himul_n249), .ZN(Inst_f4_multd_H_himul_n254) );
  NAND2_X1 Inst_f4_multd_H_himul_U11 ( .A1(Inst_f4_multd_H_himul_n243), .A2(
        FF3_out[15]), .ZN(Inst_f4_multd_H_himul_n253) );
  XOR2_X1 Inst_f4_multd_H_himul_U10 ( .A(Inst_f4_multd_H_himul_n251), .B(
        Inst_f4_multd_H_himul_n339), .Z(Inst_f4_multd_H_himul_n252) );
  NOR2_X1 Inst_f4_multd_H_himul_U9 ( .A1(Inst_f4_multd_H_himul_n338), .A2(
        Inst_f4_multd_H_himul_n250), .ZN(Inst_f4_multd_H_himul_n251) );
  XNOR2_X1 Inst_f4_multd_H_himul_U8 ( .A(FF3_out[18]), .B(FF3_out[19]), .ZN(
        Inst_f4_multd_H_himul_n250) );
  XOR2_X1 Inst_f4_multd_H_himul_U7 ( .A(Inst_f4_multd_H_himul_n246), .B(
        Inst_f4_multd_H_himul_n248), .Z(Inst_f4_multd_H_himul_n249) );
  NAND2_X1 Inst_f4_multd_H_himul_U6 ( .A1(Inst_f4_multd_H_himul_n247), .A2(
        FF3_out[3]), .ZN(Inst_f4_multd_H_himul_n248) );
  NAND2_X1 Inst_f4_multd_H_himul_U5 ( .A1(FF3_out[14]), .A2(
        Inst_f4_multd_H_himul_n337), .ZN(Inst_f4_multd_H_himul_n247) );
  NAND2_X1 Inst_f4_multd_H_himul_U4 ( .A1(FF3_out[14]), .A2(
        Inst_f4_multd_H_himul_n245), .ZN(Inst_f4_multd_H_himul_n246) );
  XNOR2_X1 Inst_f4_multd_H_himul_U3 ( .A(Inst_f4_multd_H_himul_n244), .B(
        FF3_out[6]), .ZN(Inst_f4_multd_H_himul_n245) );
  XNOR2_X1 Inst_f4_multd_H_himul_U2 ( .A(FF3_out[2]), .B(FF3_out[7]), .ZN(
        Inst_f4_multd_H_himul_n244) );
  INV_X1 Inst_f4_multd_H_himul_U1 ( .A(FF3_out[14]), .ZN(
        Inst_f4_multd_H_himul_n243) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_MaskXORInst_U2 ( .A(PRNGQ[28]), .B(
        PRNGQ[30]), .Z(Inst_f4_multd_H_AddNewMaskph_MaskXOR[0]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_MaskXORInst_U1 ( .A(PRNGQ[29]), .B(
        PRNGQ[31]), .Z(Inst_f4_multd_H_AddNewMaskph_MaskXOR[1]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_XORInst1_U2 ( .A(
        Inst_f4_multd_H_Orig_ph[4]), .B(
        Inst_f4_multd_H_AddNewMaskph_MaskXOR[0]), .Z(ph_H[4]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_XORInst1_U1 ( .A(
        Inst_f4_multd_H_Orig_ph[5]), .B(
        Inst_f4_multd_H_AddNewMaskph_MaskXOR[1]), .Z(ph_H[5]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_XORInst2_U4 ( .A(
        Inst_f4_multd_H_Orig_ph[3]), .B(PRNGQ[31]), .Z(ph_H[3]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_XORInst2_U3 ( .A(
        Inst_f4_multd_H_Orig_ph[2]), .B(PRNGQ[30]), .Z(ph_H[2]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_XORInst2_U2 ( .A(
        Inst_f4_multd_H_Orig_ph[1]), .B(PRNGQ[29]), .Z(ph_H[1]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskph_XORInst2_U1 ( .A(
        Inst_f4_multd_H_Orig_ph[0]), .B(PRNGQ[28]), .Z(ph_H[0]) );
  XNOR2_X1 Inst_f4_multd_H_summul_U104 ( .A(Inst_f4_multd_H_summul_n340), .B(
        Inst_f4_multd_H_summul_n339), .ZN(Inst_f4_multd_H_Orig_p[5]) );
  XNOR2_X1 Inst_f4_multd_H_summul_U103 ( .A(Inst_f4_multd_H_summul_n338), .B(
        Inst_f4_multd_H_summul_n337), .ZN(Inst_f4_multd_H_summul_n340) );
  XNOR2_X1 Inst_f4_multd_H_summul_U102 ( .A(Inst_f4_multd_H_summul_n336), .B(
        Inst_f4_multd_H_summul_n335), .ZN(Inst_f4_multd_H_summul_n337) );
  NOR2_X1 Inst_f4_multd_H_summul_U101 ( .A1(Inst_f4_multd_H_summul_n334), .A2(
        Inst_f4_multd_H_summul_n333), .ZN(Inst_f4_multd_H_summul_n336) );
  XNOR2_X1 Inst_f4_multd_H_summul_U100 ( .A(Inst_f4_multd_H_sB[2]), .B(
        Inst_f4_multd_H_sB[3]), .ZN(Inst_f4_multd_H_summul_n334) );
  NAND2_X1 Inst_f4_multd_H_summul_U99 ( .A1(Inst_f4_multd_H_summul_n332), .A2(
        Inst_f4_multd_H_summul_n331), .ZN(Inst_f4_multd_H_summul_n338) );
  NAND2_X1 Inst_f4_multd_H_summul_U98 ( .A1(Inst_f4_multd_H_summul_n330), .A2(
        Inst_f4_multd_H_sB[1]), .ZN(Inst_f4_multd_H_summul_n331) );
  NOR2_X1 Inst_f4_multd_H_summul_U97 ( .A1(Inst_f4_multd_H_summul_n329), .A2(
        Inst_f4_multd_H_sB[0]), .ZN(Inst_f4_multd_H_summul_n330) );
  XNOR2_X1 Inst_f4_multd_H_summul_U96 ( .A(Inst_f4_multd_H_summul_n329), .B(
        Inst_f4_multd_H_summul_n328), .ZN(Inst_f4_multd_H_summul_n332) );
  NAND2_X1 Inst_f4_multd_H_summul_U95 ( .A1(Inst_f4_multd_H_sA[1]), .A2(
        Inst_f4_multd_H_summul_n327), .ZN(Inst_f4_multd_H_summul_n328) );
  NAND2_X1 Inst_f4_multd_H_summul_U94 ( .A1(Inst_f4_multd_H_sB[0]), .A2(
        Inst_f4_multd_H_summul_n326), .ZN(Inst_f4_multd_H_summul_n327) );
  XNOR2_X1 Inst_f4_multd_H_summul_U93 ( .A(Inst_f4_multd_H_summul_n325), .B(
        Inst_f4_multd_H_summul_n324), .ZN(Inst_f4_multd_H_Orig_p[4]) );
  XNOR2_X1 Inst_f4_multd_H_summul_U92 ( .A(Inst_f4_multd_H_summul_n323), .B(
        Inst_f4_multd_H_summul_n322), .ZN(Inst_f4_multd_H_summul_n324) );
  XNOR2_X1 Inst_f4_multd_H_summul_U91 ( .A(Inst_f4_multd_H_summul_n321), .B(
        Inst_f4_multd_H_summul_n320), .ZN(Inst_f4_multd_H_summul_n322) );
  NAND2_X1 Inst_f4_multd_H_summul_U90 ( .A1(Inst_f4_multd_H_summul_n319), .A2(
        Inst_f4_multd_H_sA[2]), .ZN(Inst_f4_multd_H_summul_n321) );
  NAND2_X1 Inst_f4_multd_H_summul_U89 ( .A1(Inst_f4_multd_H_summul_n318), .A2(
        Inst_f4_multd_H_summul_n317), .ZN(Inst_f4_multd_H_summul_n323) );
  NAND2_X1 Inst_f4_multd_H_summul_U88 ( .A1(Inst_f4_multd_H_sB[0]), .A2(
        Inst_f4_multd_H_summul_n316), .ZN(Inst_f4_multd_H_summul_n317) );
  OR2_X1 Inst_f4_multd_H_summul_U87 ( .A1(Inst_f4_multd_H_summul_n316), .A2(
        Inst_f4_multd_H_summul_n326), .ZN(Inst_f4_multd_H_summul_n318) );
  XOR2_X1 Inst_f4_multd_H_summul_U86 ( .A(Inst_f4_multd_H_sA[1]), .B(
        Inst_f4_multd_H_summul_n315), .Z(Inst_f4_multd_H_summul_n316) );
  XNOR2_X1 Inst_f4_multd_H_summul_U85 ( .A(Inst_f4_multd_H_summul_n314), .B(
        Inst_f4_multd_H_summul_n335), .ZN(Inst_f4_multd_H_summul_n325) );
  XOR2_X1 Inst_f4_multd_H_summul_U84 ( .A(Inst_f4_multd_H_summul_n313), .B(
        Inst_f4_multd_H_summul_n312), .Z(Inst_f4_multd_H_summul_n335) );
  NAND2_X1 Inst_f4_multd_H_summul_U83 ( .A1(Inst_f4_multd_H_sB[2]), .A2(
        Inst_f4_multd_H_sA[1]), .ZN(Inst_f4_multd_H_summul_n312) );
  NOR2_X1 Inst_f4_multd_H_summul_U82 ( .A1(Inst_f4_multd_H_summul_n311), .A2(
        Inst_f4_multd_H_summul_n326), .ZN(Inst_f4_multd_H_summul_n313) );
  INV_X1 Inst_f4_multd_H_summul_U81 ( .A(Inst_f4_multd_H_sB[1]), .ZN(
        Inst_f4_multd_H_summul_n326) );
  XNOR2_X1 Inst_f4_multd_H_summul_U80 ( .A(Inst_f4_multd_H_sA[0]), .B(
        Inst_f4_multd_H_sA[2]), .ZN(Inst_f4_multd_H_summul_n311) );
  NAND2_X1 Inst_f4_multd_H_summul_U79 ( .A1(Inst_f4_multd_H_summul_n310), .A2(
        Inst_f4_multd_H_summul_n309), .ZN(Inst_f4_multd_H_summul_n314) );
  NAND2_X1 Inst_f4_multd_H_summul_U78 ( .A1(Inst_f4_multd_H_sA[1]), .A2(
        Inst_f4_multd_H_summul_n308), .ZN(Inst_f4_multd_H_summul_n309) );
  NAND2_X1 Inst_f4_multd_H_summul_U77 ( .A1(Inst_f4_multd_H_sA[0]), .A2(
        Inst_f4_multd_H_sB[3]), .ZN(Inst_f4_multd_H_summul_n310) );
  XNOR2_X1 Inst_f4_multd_H_summul_U76 ( .A(Inst_f4_multd_H_summul_n307), .B(
        Inst_f4_multd_H_summul_n306), .ZN(Inst_f4_multd_H_Orig_p[3]) );
  XNOR2_X1 Inst_f4_multd_H_summul_U75 ( .A(Inst_f4_multd_H_summul_n305), .B(
        Inst_f4_multd_H_summul_n304), .ZN(Inst_f4_multd_H_summul_n306) );
  XOR2_X1 Inst_f4_multd_H_summul_U74 ( .A(Inst_f4_multd_H_summul_n303), .B(
        Inst_f4_multd_H_summul_n302), .Z(Inst_f4_multd_H_summul_n305) );
  NAND2_X1 Inst_f4_multd_H_summul_U73 ( .A1(Inst_f4_multd_H_sA[4]), .A2(
        Inst_f4_multd_H_sB[4]), .ZN(Inst_f4_multd_H_summul_n302) );
  NAND2_X1 Inst_f4_multd_H_summul_U72 ( .A1(Inst_f4_multd_H_sA[5]), .A2(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n303) );
  XOR2_X1 Inst_f4_multd_H_summul_U71 ( .A(Inst_f4_multd_H_summul_n301), .B(
        Inst_f4_multd_H_summul_n300), .Z(Inst_f4_multd_H_summul_n307) );
  XOR2_X1 Inst_f4_multd_H_summul_U70 ( .A(Inst_f4_multd_H_summul_n299), .B(
        Inst_f4_multd_H_summul_n298), .Z(Inst_f4_multd_H_summul_n300) );
  NAND2_X1 Inst_f4_multd_H_summul_U69 ( .A1(Inst_f4_multd_H_sA[4]), .A2(
        Inst_f4_multd_H_summul_n297), .ZN(Inst_f4_multd_H_summul_n298) );
  NAND2_X1 Inst_f4_multd_H_summul_U68 ( .A1(Inst_f4_multd_H_sA[0]), .A2(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n299) );
  XNOR2_X1 Inst_f4_multd_H_summul_U67 ( .A(Inst_f4_multd_H_summul_n296), .B(
        Inst_f4_multd_H_summul_n295), .ZN(Inst_f4_multd_H_summul_n301) );
  XNOR2_X1 Inst_f4_multd_H_summul_U66 ( .A(Inst_f4_multd_H_sA[5]), .B(
        Inst_f4_multd_H_summul_n294), .ZN(Inst_f4_multd_H_summul_n295) );
  XOR2_X1 Inst_f4_multd_H_summul_U65 ( .A(Inst_f4_multd_H_summul_n293), .B(
        Inst_f4_multd_H_summul_n292), .Z(Inst_f4_multd_H_summul_n294) );
  NAND2_X1 Inst_f4_multd_H_summul_U64 ( .A1(Inst_f4_multd_H_sB[0]), .A2(
        Inst_f4_multd_H_sA[4]), .ZN(Inst_f4_multd_H_summul_n292) );
  NOR2_X1 Inst_f4_multd_H_summul_U63 ( .A1(Inst_f4_multd_H_summul_n291), .A2(
        Inst_f4_multd_H_sB[1]), .ZN(Inst_f4_multd_H_summul_n293) );
  NAND2_X1 Inst_f4_multd_H_summul_U62 ( .A1(Inst_f4_multd_H_summul_n290), .A2(
        Inst_f4_multd_H_sB[4]), .ZN(Inst_f4_multd_H_summul_n296) );
  XNOR2_X1 Inst_f4_multd_H_summul_U61 ( .A(Inst_f4_multd_H_summul_n333), .B(
        Inst_f4_multd_H_summul_n289), .ZN(Inst_f4_multd_H_summul_n290) );
  XNOR2_X1 Inst_f4_multd_H_summul_U60 ( .A(Inst_f4_multd_H_sA[1]), .B(
        Inst_f4_multd_H_summul_n288), .ZN(Inst_f4_multd_H_summul_n289) );
  INV_X1 Inst_f4_multd_H_summul_U59 ( .A(Inst_f4_multd_H_sA[0]), .ZN(
        Inst_f4_multd_H_summul_n333) );
  XOR2_X1 Inst_f4_multd_H_summul_U58 ( .A(Inst_f4_multd_H_summul_n287), .B(
        Inst_f4_multd_H_summul_n286), .Z(Inst_f4_multd_H_Orig_p[2]) );
  NAND2_X1 Inst_f4_multd_H_summul_U57 ( .A1(Inst_f4_multd_H_summul_n285), .A2(
        Inst_f4_multd_H_summul_n284), .ZN(Inst_f4_multd_H_summul_n286) );
  OR2_X1 Inst_f4_multd_H_summul_U56 ( .A1(Inst_f4_multd_H_sB[5]), .A2(
        Inst_f4_multd_H_summul_n291), .ZN(Inst_f4_multd_H_summul_n284) );
  NAND2_X1 Inst_f4_multd_H_summul_U55 ( .A1(Inst_f4_multd_H_summul_n283), .A2(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n285) );
  XNOR2_X1 Inst_f4_multd_H_summul_U54 ( .A(Inst_f4_multd_H_summul_n282), .B(
        Inst_f4_multd_H_sA[0]), .ZN(Inst_f4_multd_H_summul_n283) );
  XOR2_X1 Inst_f4_multd_H_summul_U53 ( .A(Inst_f4_multd_H_summul_n281), .B(
        Inst_f4_multd_H_summul_n280), .Z(Inst_f4_multd_H_summul_n287) );
  NOR2_X1 Inst_f4_multd_H_summul_U52 ( .A1(Inst_f4_multd_H_summul_n288), .A2(
        Inst_f4_multd_H_summul_n279), .ZN(Inst_f4_multd_H_summul_n280) );
  XOR2_X1 Inst_f4_multd_H_summul_U51 ( .A(Inst_f4_multd_H_summul_n297), .B(
        Inst_f4_multd_H_sB[1]), .Z(Inst_f4_multd_H_summul_n279) );
  XNOR2_X1 Inst_f4_multd_H_summul_U50 ( .A(Inst_f4_multd_H_summul_n278), .B(
        Inst_f4_multd_H_summul_n277), .ZN(Inst_f4_multd_H_summul_n281) );
  XNOR2_X1 Inst_f4_multd_H_summul_U49 ( .A(Inst_f4_multd_H_sB[0]), .B(
        Inst_f4_multd_H_summul_n320), .ZN(Inst_f4_multd_H_summul_n277) );
  XOR2_X1 Inst_f4_multd_H_summul_U48 ( .A(Inst_f4_multd_H_summul_n276), .B(
        Inst_f4_multd_H_summul_n275), .Z(Inst_f4_multd_H_summul_n320) );
  NAND2_X1 Inst_f4_multd_H_summul_U47 ( .A1(Inst_f4_multd_H_sA[1]), .A2(
        Inst_f4_multd_H_sB[0]), .ZN(Inst_f4_multd_H_summul_n275) );
  NAND2_X1 Inst_f4_multd_H_summul_U46 ( .A1(Inst_f4_multd_H_sA[0]), .A2(
        Inst_f4_multd_H_sB[1]), .ZN(Inst_f4_multd_H_summul_n276) );
  XOR2_X1 Inst_f4_multd_H_summul_U45 ( .A(Inst_f4_multd_H_summul_n274), .B(
        Inst_f4_multd_H_summul_n304), .Z(Inst_f4_multd_H_summul_n278) );
  XOR2_X1 Inst_f4_multd_H_summul_U44 ( .A(Inst_f4_multd_H_summul_n273), .B(
        Inst_f4_multd_H_summul_n272), .Z(Inst_f4_multd_H_summul_n304) );
  NAND2_X1 Inst_f4_multd_H_summul_U43 ( .A1(Inst_f4_multd_H_sA[4]), .A2(
        Inst_f4_multd_H_sB[1]), .ZN(Inst_f4_multd_H_summul_n272) );
  NAND2_X1 Inst_f4_multd_H_summul_U42 ( .A1(Inst_f4_multd_H_sA[5]), .A2(
        Inst_f4_multd_H_sB[0]), .ZN(Inst_f4_multd_H_summul_n273) );
  XOR2_X1 Inst_f4_multd_H_summul_U41 ( .A(Inst_f4_multd_H_summul_n271), .B(
        Inst_f4_multd_H_summul_n270), .Z(Inst_f4_multd_H_summul_n274) );
  NAND2_X1 Inst_f4_multd_H_summul_U40 ( .A1(Inst_f4_multd_H_sB[4]), .A2(
        Inst_f4_multd_H_summul_n291), .ZN(Inst_f4_multd_H_summul_n270) );
  INV_X1 Inst_f4_multd_H_summul_U39 ( .A(Inst_f4_multd_H_sA[1]), .ZN(
        Inst_f4_multd_H_summul_n291) );
  XNOR2_X1 Inst_f4_multd_H_summul_U38 ( .A(Inst_f4_multd_H_summul_n269), .B(
        Inst_f4_multd_H_summul_n268), .ZN(Inst_f4_multd_H_Orig_p[1]) );
  XNOR2_X1 Inst_f4_multd_H_summul_U37 ( .A(Inst_f4_multd_H_summul_n267), .B(
        Inst_f4_multd_H_summul_n266), .ZN(Inst_f4_multd_H_summul_n269) );
  NAND2_X1 Inst_f4_multd_H_summul_U36 ( .A1(Inst_f4_multd_H_summul_n265), .A2(
        Inst_f4_multd_H_sA[2]), .ZN(Inst_f4_multd_H_summul_n266) );
  XNOR2_X1 Inst_f4_multd_H_summul_U35 ( .A(Inst_f4_multd_H_sB[2]), .B(
        Inst_f4_multd_H_summul_n297), .ZN(Inst_f4_multd_H_summul_n265) );
  XNOR2_X1 Inst_f4_multd_H_summul_U34 ( .A(Inst_f4_multd_H_summul_n264), .B(
        Inst_f4_multd_H_summul_n263), .ZN(Inst_f4_multd_H_summul_n267) );
  XNOR2_X1 Inst_f4_multd_H_summul_U33 ( .A(Inst_f4_multd_H_summul_n262), .B(
        Inst_f4_multd_H_summul_n261), .ZN(Inst_f4_multd_H_summul_n263) );
  NAND2_X1 Inst_f4_multd_H_summul_U32 ( .A1(Inst_f4_multd_H_summul_n260), .A2(
        Inst_f4_multd_H_summul_n319), .ZN(Inst_f4_multd_H_summul_n261) );
  XOR2_X1 Inst_f4_multd_H_summul_U31 ( .A(Inst_f4_multd_H_sB[2]), .B(
        Inst_f4_multd_H_sB[3]), .Z(Inst_f4_multd_H_summul_n319) );
  XOR2_X1 Inst_f4_multd_H_summul_U30 ( .A(Inst_f4_multd_H_sA[2]), .B(
        Inst_f4_multd_H_sA[4]), .Z(Inst_f4_multd_H_summul_n260) );
  NAND2_X1 Inst_f4_multd_H_summul_U29 ( .A1(Inst_f4_multd_H_sA[3]), .A2(
        Inst_f4_multd_H_sB[4]), .ZN(Inst_f4_multd_H_summul_n262) );
  XNOR2_X1 Inst_f4_multd_H_summul_U28 ( .A(Inst_f4_multd_H_summul_n259), .B(
        Inst_f4_multd_H_summul_n258), .ZN(Inst_f4_multd_H_summul_n264) );
  XOR2_X1 Inst_f4_multd_H_summul_U27 ( .A(Inst_f4_multd_H_summul_n257), .B(
        Inst_f4_multd_H_summul_n256), .Z(Inst_f4_multd_H_summul_n259) );
  NOR2_X1 Inst_f4_multd_H_summul_U26 ( .A1(Inst_f4_multd_H_summul_n282), .A2(
        Inst_f4_multd_H_sB[4]), .ZN(Inst_f4_multd_H_summul_n256) );
  INV_X1 Inst_f4_multd_H_summul_U25 ( .A(Inst_f4_multd_H_sA[4]), .ZN(
        Inst_f4_multd_H_summul_n282) );
  NOR2_X1 Inst_f4_multd_H_summul_U24 ( .A1(Inst_f4_multd_H_summul_n288), .A2(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n257) );
  INV_X1 Inst_f4_multd_H_summul_U23 ( .A(Inst_f4_multd_H_sA[5]), .ZN(
        Inst_f4_multd_H_summul_n288) );
  XNOR2_X1 Inst_f4_multd_H_summul_U22 ( .A(Inst_f4_multd_H_summul_n255), .B(
        Inst_f4_multd_H_summul_n254), .ZN(Inst_f4_multd_H_Orig_p[0]) );
  NAND2_X1 Inst_f4_multd_H_summul_U21 ( .A1(Inst_f4_multd_H_sA[2]), .A2(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n254) );
  XNOR2_X1 Inst_f4_multd_H_summul_U20 ( .A(Inst_f4_multd_H_summul_n339), .B(
        Inst_f4_multd_H_summul_n253), .ZN(Inst_f4_multd_H_summul_n255) );
  XNOR2_X1 Inst_f4_multd_H_summul_U19 ( .A(Inst_f4_multd_H_summul_n252), .B(
        Inst_f4_multd_H_summul_n251), .ZN(Inst_f4_multd_H_summul_n253) );
  XNOR2_X1 Inst_f4_multd_H_summul_U18 ( .A(Inst_f4_multd_H_summul_n250), .B(
        Inst_f4_multd_H_summul_n249), .ZN(Inst_f4_multd_H_summul_n251) );
  XNOR2_X1 Inst_f4_multd_H_summul_U17 ( .A(Inst_f4_multd_H_summul_n248), .B(
        Inst_f4_multd_H_summul_n268), .ZN(Inst_f4_multd_H_summul_n249) );
  NAND2_X1 Inst_f4_multd_H_summul_U16 ( .A1(Inst_f4_multd_H_sB[2]), .A2(
        Inst_f4_multd_H_summul_n247), .ZN(Inst_f4_multd_H_summul_n268) );
  XOR2_X1 Inst_f4_multd_H_summul_U15 ( .A(Inst_f4_multd_H_sA[3]), .B(
        Inst_f4_multd_H_sA[5]), .Z(Inst_f4_multd_H_summul_n247) );
  NOR2_X1 Inst_f4_multd_H_summul_U14 ( .A1(Inst_f4_multd_H_summul_n246), .A2(
        Inst_f4_multd_H_summul_n308), .ZN(Inst_f4_multd_H_summul_n248) );
  INV_X1 Inst_f4_multd_H_summul_U13 ( .A(Inst_f4_multd_H_sB[3]), .ZN(
        Inst_f4_multd_H_summul_n308) );
  XNOR2_X1 Inst_f4_multd_H_summul_U12 ( .A(Inst_f4_multd_H_sA[5]), .B(
        Inst_f4_multd_H_sA[4]), .ZN(Inst_f4_multd_H_summul_n246) );
  XNOR2_X1 Inst_f4_multd_H_summul_U11 ( .A(Inst_f4_multd_H_summul_n271), .B(
        Inst_f4_multd_H_sB[4]), .ZN(Inst_f4_multd_H_summul_n250) );
  NAND2_X1 Inst_f4_multd_H_summul_U10 ( .A1(Inst_f4_multd_H_sA[4]), .A2(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n271) );
  NOR2_X1 Inst_f4_multd_H_summul_U9 ( .A1(Inst_f4_multd_H_summul_n315), .A2(
        Inst_f4_multd_H_summul_n297), .ZN(Inst_f4_multd_H_summul_n252) );
  XNOR2_X1 Inst_f4_multd_H_summul_U8 ( .A(Inst_f4_multd_H_sB[4]), .B(
        Inst_f4_multd_H_sB[5]), .ZN(Inst_f4_multd_H_summul_n297) );
  INV_X1 Inst_f4_multd_H_summul_U7 ( .A(Inst_f4_multd_H_sA[3]), .ZN(
        Inst_f4_multd_H_summul_n315) );
  XNOR2_X1 Inst_f4_multd_H_summul_U6 ( .A(Inst_f4_multd_H_summul_n258), .B(
        Inst_f4_multd_H_summul_n245), .ZN(Inst_f4_multd_H_summul_n339) );
  NAND2_X1 Inst_f4_multd_H_summul_U5 ( .A1(Inst_f4_multd_H_sA[2]), .A2(
        Inst_f4_multd_H_sB[2]), .ZN(Inst_f4_multd_H_summul_n245) );
  NAND2_X1 Inst_f4_multd_H_summul_U4 ( .A1(Inst_f4_multd_H_sB[3]), .A2(
        Inst_f4_multd_H_sA[3]), .ZN(Inst_f4_multd_H_summul_n258) );
  AND2_X1 Inst_f4_multd_H_summul_U3 ( .A1(Inst_f4_multd_H_summul_n244), .A2(
        Inst_f4_multd_H_sB[0]), .ZN(Inst_f4_multd_H_summul_n329) );
  XNOR2_X1 Inst_f4_multd_H_summul_U2 ( .A(Inst_f4_multd_H_summul_n243), .B(
        Inst_f4_multd_H_sA[0]), .ZN(Inst_f4_multd_H_summul_n244) );
  XNOR2_X1 Inst_f4_multd_H_summul_U1 ( .A(Inst_f4_multd_H_sA[3]), .B(
        Inst_f4_multd_H_sA[2]), .ZN(Inst_f4_multd_H_summul_n243) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_MaskXORInst_U2 ( .A(PRNGQ[33]), .B(
        PRNGQ[35]), .Z(Inst_f4_multd_H_AddNewMaskp_MaskXOR[1]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_MaskXORInst_U1 ( .A(PRNGQ[32]), .B(
        PRNGQ[34]), .Z(Inst_f4_multd_H_AddNewMaskp_MaskXOR[0]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_XORInst1_U2 ( .A(
        Inst_f4_multd_H_Orig_p[5]), .B(Inst_f4_multd_H_AddNewMaskp_MaskXOR[1]), 
        .Z(p_H[5]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_XORInst1_U1 ( .A(
        Inst_f4_multd_H_Orig_p[4]), .B(Inst_f4_multd_H_AddNewMaskp_MaskXOR[0]), 
        .Z(p_H[4]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_XORInst2_U4 ( .A(
        Inst_f4_multd_H_Orig_p[3]), .B(PRNGQ[35]), .Z(p_H[3]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_XORInst2_U3 ( .A(
        Inst_f4_multd_H_Orig_p[2]), .B(PRNGQ[34]), .Z(p_H[2]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_XORInst2_U2 ( .A(
        Inst_f4_multd_H_Orig_p[1]), .B(PRNGQ[33]), .Z(p_H[1]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskp_XORInst2_U1 ( .A(
        Inst_f4_multd_H_Orig_p[0]), .B(PRNGQ[32]), .Z(p_H[0]) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U104 ( .A(Inst_f4_multd_H_lowmul_n336), .B(
        Inst_f4_multd_H_lowmul_n335), .ZN(Inst_f4_multd_H_Orig_pl[4]) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U103 ( .A(Inst_f4_multd_H_lowmul_n334), .B(
        Inst_f4_multd_H_lowmul_n333), .ZN(Inst_f4_multd_H_lowmul_n335) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U102 ( .A(Inst_f4_multd_H_lowmul_n332), .B(
        Inst_f4_multd_H_lowmul_n331), .ZN(Inst_f4_multd_H_lowmul_n333) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U101 ( .A1(Inst_f4_multd_H_lowmul_n330), 
        .A2(FF3_out[4]), .ZN(Inst_f4_multd_H_lowmul_n332) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U100 ( .A1(Inst_f4_multd_H_lowmul_n329), 
        .A2(Inst_f4_multd_H_lowmul_n328), .ZN(Inst_f4_multd_H_lowmul_n334) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U99 ( .A1(FF3_out[12]), .A2(
        Inst_f4_multd_H_lowmul_n327), .ZN(Inst_f4_multd_H_lowmul_n328) );
  OR2_X1 Inst_f4_multd_H_lowmul_U98 ( .A1(Inst_f4_multd_H_lowmul_n327), .A2(
        Inst_f4_multd_H_lowmul_n337), .ZN(Inst_f4_multd_H_lowmul_n329) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U97 ( .A(FF3_out[1]), .B(
        Inst_f4_multd_H_lowmul_n326), .Z(Inst_f4_multd_H_lowmul_n327) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U96 ( .A(Inst_f4_multd_H_lowmul_n325), .B(
        Inst_f4_multd_H_lowmul_n339), .ZN(Inst_f4_multd_H_lowmul_n336) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U95 ( .A(Inst_f4_multd_H_lowmul_n324), .B(
        Inst_f4_multd_H_lowmul_n323), .Z(Inst_f4_multd_H_lowmul_n339) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U94 ( .A1(FF3_out[16]), .A2(FF3_out[1]), 
        .ZN(Inst_f4_multd_H_lowmul_n323) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U93 ( .A1(Inst_f4_multd_H_lowmul_n322), .A2(
        Inst_f4_multd_H_lowmul_n337), .ZN(Inst_f4_multd_H_lowmul_n324) );
  INV_X1 Inst_f4_multd_H_lowmul_U92 ( .A(FF3_out[13]), .ZN(
        Inst_f4_multd_H_lowmul_n337) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U91 ( .A(FF3_out[0]), .B(FF3_out[4]), .ZN(
        Inst_f4_multd_H_lowmul_n322) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U90 ( .A1(Inst_f4_multd_H_lowmul_n321), .A2(
        Inst_f4_multd_H_lowmul_n320), .ZN(Inst_f4_multd_H_lowmul_n325) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U89 ( .A1(FF3_out[1]), .A2(
        Inst_f4_multd_H_lowmul_n319), .ZN(Inst_f4_multd_H_lowmul_n320) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U88 ( .A1(FF3_out[0]), .A2(FF3_out[17]), 
        .ZN(Inst_f4_multd_H_lowmul_n321) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U87 ( .A(Inst_f4_multd_H_lowmul_n318), .B(
        Inst_f4_multd_H_lowmul_n317), .ZN(Inst_f4_multd_H_Orig_pl[3]) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U86 ( .A(Inst_f4_multd_H_lowmul_n316), .B(
        Inst_f4_multd_H_lowmul_n315), .ZN(Inst_f4_multd_H_lowmul_n317) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U85 ( .A(Inst_f4_multd_H_lowmul_n314), .B(
        Inst_f4_multd_H_lowmul_n313), .Z(Inst_f4_multd_H_lowmul_n316) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U84 ( .A1(FF3_out[8]), .A2(FF3_out[20]), 
        .ZN(Inst_f4_multd_H_lowmul_n313) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U83 ( .A1(FF3_out[9]), .A2(FF3_out[21]), 
        .ZN(Inst_f4_multd_H_lowmul_n314) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U82 ( .A(Inst_f4_multd_H_lowmul_n312), .B(
        Inst_f4_multd_H_lowmul_n311), .Z(Inst_f4_multd_H_lowmul_n318) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U81 ( .A(Inst_f4_multd_H_lowmul_n310), .B(
        Inst_f4_multd_H_lowmul_n309), .Z(Inst_f4_multd_H_lowmul_n311) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U80 ( .A1(FF3_out[8]), .A2(
        Inst_f4_multd_H_lowmul_n308), .ZN(Inst_f4_multd_H_lowmul_n309) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U79 ( .A1(FF3_out[0]), .A2(FF3_out[21]), 
        .ZN(Inst_f4_multd_H_lowmul_n310) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U78 ( .A(Inst_f4_multd_H_lowmul_n307), .B(
        Inst_f4_multd_H_lowmul_n306), .ZN(Inst_f4_multd_H_lowmul_n312) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U77 ( .A(FF3_out[9]), .B(
        Inst_f4_multd_H_lowmul_n305), .ZN(Inst_f4_multd_H_lowmul_n306) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U76 ( .A(Inst_f4_multd_H_lowmul_n304), .B(
        Inst_f4_multd_H_lowmul_n303), .Z(Inst_f4_multd_H_lowmul_n305) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U75 ( .A1(FF3_out[12]), .A2(FF3_out[8]), 
        .ZN(Inst_f4_multd_H_lowmul_n303) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U74 ( .A1(Inst_f4_multd_H_lowmul_n302), .A2(
        FF3_out[13]), .ZN(Inst_f4_multd_H_lowmul_n304) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U73 ( .A1(Inst_f4_multd_H_lowmul_n301), .A2(
        FF3_out[20]), .ZN(Inst_f4_multd_H_lowmul_n307) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U72 ( .A(Inst_f4_multd_H_lowmul_n338), .B(
        Inst_f4_multd_H_lowmul_n300), .ZN(Inst_f4_multd_H_lowmul_n301) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U71 ( .A(FF3_out[1]), .B(
        Inst_f4_multd_H_lowmul_n299), .ZN(Inst_f4_multd_H_lowmul_n300) );
  INV_X1 Inst_f4_multd_H_lowmul_U70 ( .A(FF3_out[0]), .ZN(
        Inst_f4_multd_H_lowmul_n338) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U69 ( .A(Inst_f4_multd_H_lowmul_n298), .B(
        Inst_f4_multd_H_lowmul_n297), .Z(Inst_f4_multd_H_Orig_pl[2]) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U68 ( .A1(Inst_f4_multd_H_lowmul_n296), .A2(
        Inst_f4_multd_H_lowmul_n295), .ZN(Inst_f4_multd_H_lowmul_n297) );
  OR2_X1 Inst_f4_multd_H_lowmul_U67 ( .A1(FF3_out[21]), .A2(
        Inst_f4_multd_H_lowmul_n302), .ZN(Inst_f4_multd_H_lowmul_n295) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U66 ( .A1(Inst_f4_multd_H_lowmul_n294), .A2(
        FF3_out[21]), .ZN(Inst_f4_multd_H_lowmul_n296) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U65 ( .A(Inst_f4_multd_H_lowmul_n293), .B(
        FF3_out[0]), .ZN(Inst_f4_multd_H_lowmul_n294) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U64 ( .A(Inst_f4_multd_H_lowmul_n292), .B(
        Inst_f4_multd_H_lowmul_n291), .Z(Inst_f4_multd_H_lowmul_n298) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U63 ( .A1(Inst_f4_multd_H_lowmul_n299), .A2(
        Inst_f4_multd_H_lowmul_n290), .ZN(Inst_f4_multd_H_lowmul_n291) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U62 ( .A(Inst_f4_multd_H_lowmul_n308), .B(
        FF3_out[13]), .Z(Inst_f4_multd_H_lowmul_n290) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U61 ( .A(Inst_f4_multd_H_lowmul_n289), .B(
        Inst_f4_multd_H_lowmul_n288), .ZN(Inst_f4_multd_H_lowmul_n292) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U60 ( .A(FF3_out[12]), .B(
        Inst_f4_multd_H_lowmul_n331), .ZN(Inst_f4_multd_H_lowmul_n288) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U59 ( .A(Inst_f4_multd_H_lowmul_n287), .B(
        Inst_f4_multd_H_lowmul_n286), .Z(Inst_f4_multd_H_lowmul_n331) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U58 ( .A1(FF3_out[1]), .A2(FF3_out[12]), 
        .ZN(Inst_f4_multd_H_lowmul_n286) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U57 ( .A1(FF3_out[0]), .A2(FF3_out[13]), 
        .ZN(Inst_f4_multd_H_lowmul_n287) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U56 ( .A(Inst_f4_multd_H_lowmul_n285), .B(
        Inst_f4_multd_H_lowmul_n315), .Z(Inst_f4_multd_H_lowmul_n289) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U55 ( .A(Inst_f4_multd_H_lowmul_n284), .B(
        Inst_f4_multd_H_lowmul_n283), .Z(Inst_f4_multd_H_lowmul_n315) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U54 ( .A1(FF3_out[8]), .A2(FF3_out[13]), 
        .ZN(Inst_f4_multd_H_lowmul_n283) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U53 ( .A1(FF3_out[9]), .A2(FF3_out[12]), 
        .ZN(Inst_f4_multd_H_lowmul_n284) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U52 ( .A(Inst_f4_multd_H_lowmul_n282), .B(
        Inst_f4_multd_H_lowmul_n281), .Z(Inst_f4_multd_H_lowmul_n285) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U51 ( .A1(FF3_out[20]), .A2(
        Inst_f4_multd_H_lowmul_n302), .ZN(Inst_f4_multd_H_lowmul_n281) );
  INV_X1 Inst_f4_multd_H_lowmul_U50 ( .A(FF3_out[1]), .ZN(
        Inst_f4_multd_H_lowmul_n302) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U49 ( .A(Inst_f4_multd_H_lowmul_n280), .B(
        Inst_f4_multd_H_lowmul_n279), .ZN(Inst_f4_multd_H_Orig_pl[1]) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U48 ( .A(Inst_f4_multd_H_lowmul_n278), .B(
        Inst_f4_multd_H_lowmul_n277), .ZN(Inst_f4_multd_H_lowmul_n280) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U47 ( .A1(Inst_f4_multd_H_lowmul_n276), .A2(
        FF3_out[4]), .ZN(Inst_f4_multd_H_lowmul_n277) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U46 ( .A(FF3_out[16]), .B(
        Inst_f4_multd_H_lowmul_n308), .ZN(Inst_f4_multd_H_lowmul_n276) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U45 ( .A(Inst_f4_multd_H_lowmul_n275), .B(
        Inst_f4_multd_H_lowmul_n274), .ZN(Inst_f4_multd_H_lowmul_n278) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U44 ( .A(Inst_f4_multd_H_lowmul_n273), .B(
        Inst_f4_multd_H_lowmul_n272), .ZN(Inst_f4_multd_H_lowmul_n274) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U43 ( .A1(Inst_f4_multd_H_lowmul_n271), .A2(
        Inst_f4_multd_H_lowmul_n330), .ZN(Inst_f4_multd_H_lowmul_n272) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U42 ( .A(FF3_out[16]), .B(FF3_out[17]), .Z(
        Inst_f4_multd_H_lowmul_n330) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U41 ( .A(FF3_out[4]), .B(FF3_out[8]), .Z(
        Inst_f4_multd_H_lowmul_n271) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U40 ( .A1(FF3_out[5]), .A2(FF3_out[20]), 
        .ZN(Inst_f4_multd_H_lowmul_n273) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U39 ( .A(Inst_f4_multd_H_lowmul_n270), .B(
        Inst_f4_multd_H_lowmul_n269), .ZN(Inst_f4_multd_H_lowmul_n275) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U38 ( .A(Inst_f4_multd_H_lowmul_n268), .B(
        Inst_f4_multd_H_lowmul_n267), .Z(Inst_f4_multd_H_lowmul_n270) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U37 ( .A1(Inst_f4_multd_H_lowmul_n293), .A2(
        FF3_out[20]), .ZN(Inst_f4_multd_H_lowmul_n267) );
  INV_X1 Inst_f4_multd_H_lowmul_U36 ( .A(FF3_out[8]), .ZN(
        Inst_f4_multd_H_lowmul_n293) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U35 ( .A1(Inst_f4_multd_H_lowmul_n299), .A2(
        FF3_out[21]), .ZN(Inst_f4_multd_H_lowmul_n268) );
  INV_X1 Inst_f4_multd_H_lowmul_U34 ( .A(FF3_out[9]), .ZN(
        Inst_f4_multd_H_lowmul_n299) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U33 ( .A(Inst_f4_multd_H_lowmul_n266), .B(
        Inst_f4_multd_H_lowmul_n265), .ZN(Inst_f4_multd_H_Orig_pl[0]) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U32 ( .A1(FF3_out[4]), .A2(FF3_out[21]), 
        .ZN(Inst_f4_multd_H_lowmul_n265) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U31 ( .A(Inst_f4_multd_H_lowmul_n340), .B(
        Inst_f4_multd_H_lowmul_n264), .ZN(Inst_f4_multd_H_lowmul_n266) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U30 ( .A(Inst_f4_multd_H_lowmul_n263), .B(
        Inst_f4_multd_H_lowmul_n262), .ZN(Inst_f4_multd_H_lowmul_n264) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U29 ( .A(Inst_f4_multd_H_lowmul_n261), .B(
        Inst_f4_multd_H_lowmul_n260), .ZN(Inst_f4_multd_H_lowmul_n262) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U28 ( .A(Inst_f4_multd_H_lowmul_n259), .B(
        Inst_f4_multd_H_lowmul_n279), .ZN(Inst_f4_multd_H_lowmul_n260) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U27 ( .A1(FF3_out[16]), .A2(
        Inst_f4_multd_H_lowmul_n258), .ZN(Inst_f4_multd_H_lowmul_n279) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U26 ( .A(FF3_out[5]), .B(FF3_out[9]), .Z(
        Inst_f4_multd_H_lowmul_n258) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U25 ( .A1(Inst_f4_multd_H_lowmul_n257), .A2(
        Inst_f4_multd_H_lowmul_n319), .ZN(Inst_f4_multd_H_lowmul_n259) );
  INV_X1 Inst_f4_multd_H_lowmul_U24 ( .A(FF3_out[17]), .ZN(
        Inst_f4_multd_H_lowmul_n319) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U23 ( .A(FF3_out[9]), .B(FF3_out[8]), .ZN(
        Inst_f4_multd_H_lowmul_n257) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U22 ( .A(Inst_f4_multd_H_lowmul_n282), .B(
        FF3_out[20]), .ZN(Inst_f4_multd_H_lowmul_n261) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U21 ( .A1(FF3_out[8]), .A2(FF3_out[21]), 
        .ZN(Inst_f4_multd_H_lowmul_n282) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U20 ( .A1(Inst_f4_multd_H_lowmul_n326), .A2(
        Inst_f4_multd_H_lowmul_n308), .ZN(Inst_f4_multd_H_lowmul_n263) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U19 ( .A(FF3_out[20]), .B(FF3_out[21]), .ZN(
        Inst_f4_multd_H_lowmul_n308) );
  INV_X1 Inst_f4_multd_H_lowmul_U18 ( .A(FF3_out[5]), .ZN(
        Inst_f4_multd_H_lowmul_n326) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U17 ( .A(Inst_f4_multd_H_lowmul_n269), .B(
        Inst_f4_multd_H_lowmul_n256), .ZN(Inst_f4_multd_H_lowmul_n340) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U16 ( .A1(FF3_out[4]), .A2(FF3_out[16]), 
        .ZN(Inst_f4_multd_H_lowmul_n256) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U15 ( .A1(FF3_out[17]), .A2(FF3_out[5]), 
        .ZN(Inst_f4_multd_H_lowmul_n269) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U14 ( .A(Inst_f4_multd_H_lowmul_n255), .B(
        Inst_f4_multd_H_lowmul_n340), .Z(Inst_f4_multd_H_Orig_pl[5]) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U13 ( .A(Inst_f4_multd_H_lowmul_n254), .B(
        Inst_f4_multd_H_lowmul_n252), .ZN(Inst_f4_multd_H_lowmul_n255) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U12 ( .A1(Inst_f4_multd_H_lowmul_n253), .A2(
        Inst_f4_multd_H_lowmul_n249), .ZN(Inst_f4_multd_H_lowmul_n254) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U11 ( .A1(Inst_f4_multd_H_lowmul_n243), .A2(
        FF3_out[13]), .ZN(Inst_f4_multd_H_lowmul_n253) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U10 ( .A(Inst_f4_multd_H_lowmul_n251), .B(
        Inst_f4_multd_H_lowmul_n339), .Z(Inst_f4_multd_H_lowmul_n252) );
  NOR2_X1 Inst_f4_multd_H_lowmul_U9 ( .A1(Inst_f4_multd_H_lowmul_n338), .A2(
        Inst_f4_multd_H_lowmul_n250), .ZN(Inst_f4_multd_H_lowmul_n251) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U8 ( .A(FF3_out[16]), .B(FF3_out[17]), .ZN(
        Inst_f4_multd_H_lowmul_n250) );
  XOR2_X1 Inst_f4_multd_H_lowmul_U7 ( .A(Inst_f4_multd_H_lowmul_n246), .B(
        Inst_f4_multd_H_lowmul_n248), .Z(Inst_f4_multd_H_lowmul_n249) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U6 ( .A1(Inst_f4_multd_H_lowmul_n247), .A2(
        FF3_out[1]), .ZN(Inst_f4_multd_H_lowmul_n248) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U5 ( .A1(FF3_out[12]), .A2(
        Inst_f4_multd_H_lowmul_n337), .ZN(Inst_f4_multd_H_lowmul_n247) );
  NAND2_X1 Inst_f4_multd_H_lowmul_U4 ( .A1(FF3_out[12]), .A2(
        Inst_f4_multd_H_lowmul_n245), .ZN(Inst_f4_multd_H_lowmul_n246) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U3 ( .A(Inst_f4_multd_H_lowmul_n244), .B(
        FF3_out[4]), .ZN(Inst_f4_multd_H_lowmul_n245) );
  XNOR2_X1 Inst_f4_multd_H_lowmul_U2 ( .A(FF3_out[0]), .B(FF3_out[5]), .ZN(
        Inst_f4_multd_H_lowmul_n244) );
  INV_X1 Inst_f4_multd_H_lowmul_U1 ( .A(FF3_out[12]), .ZN(
        Inst_f4_multd_H_lowmul_n243) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_MaskXORInst_U2 ( .A(PRNGQ[36]), .B(
        PRNGQ[38]), .Z(Inst_f4_multd_H_AddNewMaskpl_MaskXOR[0]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_MaskXORInst_U1 ( .A(PRNGQ[37]), .B(
        PRNGQ[39]), .Z(Inst_f4_multd_H_AddNewMaskpl_MaskXOR[1]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_XORInst1_U2 ( .A(
        Inst_f4_multd_H_Orig_pl[4]), .B(
        Inst_f4_multd_H_AddNewMaskpl_MaskXOR[0]), .Z(pl_H[4]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_XORInst1_U1 ( .A(
        Inst_f4_multd_H_Orig_pl[5]), .B(
        Inst_f4_multd_H_AddNewMaskpl_MaskXOR[1]), .Z(pl_H[5]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_XORInst2_U4 ( .A(
        Inst_f4_multd_H_Orig_pl[3]), .B(PRNGQ[39]), .Z(pl_H[3]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_XORInst2_U3 ( .A(
        Inst_f4_multd_H_Orig_pl[2]), .B(PRNGQ[38]), .Z(pl_H[2]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_XORInst2_U2 ( .A(
        Inst_f4_multd_H_Orig_pl[1]), .B(PRNGQ[37]), .Z(pl_H[1]) );
  XOR2_X1 Inst_f4_multd_H_AddNewMaskpl_XORInst2_U1 ( .A(
        Inst_f4_multd_H_Orig_pl[0]), .B(PRNGQ[36]), .Z(pl_H[0]) );
  DFF_X1 PL_4_s_current_state_reg_0_ ( .D(pl_L[0]), .CK(clk), .Q(FF4_out[0]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_1_ ( .D(pl_L[1]), .CK(clk), .Q(FF4_out[1]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_2_ ( .D(pl_L[2]), .CK(clk), .Q(FF4_out[2]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_3_ ( .D(pl_L[3]), .CK(clk), .Q(FF4_out[3]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_4_ ( .D(pl_L[4]), .CK(clk), .Q(FF4_out[4]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_5_ ( .D(pl_L[5]), .CK(clk), .Q(FF4_out[5]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_6_ ( .D(p_L[0]), .CK(clk), .Q(
        Inst_f5_plwillwin_pw2_1_), .QN() );
  DFF_X1 PL_4_s_current_state_reg_7_ ( .D(p_L[1]), .CK(clk), .Q(FF4_out[7]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_8_ ( .D(p_L[2]), .CK(clk), .Q(
        Inst_f5_plwillwin_pw2_3_), .QN() );
  DFF_X1 PL_4_s_current_state_reg_9_ ( .D(p_L[3]), .CK(clk), .Q(FF4_out[9]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_10_ ( .D(p_L[4]), .CK(clk), .Q(
        Inst_f5_plwillwin_pw2_5_), .QN() );
  DFF_X1 PL_4_s_current_state_reg_11_ ( .D(p_L[5]), .CK(clk), .Q(FF4_out[11]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_12_ ( .D(ph_L[0]), .CK(clk), .Q(FF4_out[12]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_13_ ( .D(ph_L[1]), .CK(clk), .Q(FF4_out[13]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_14_ ( .D(ph_L[2]), .CK(clk), .Q(FF4_out[14]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_15_ ( .D(ph_L[3]), .CK(clk), .Q(FF4_out[15]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_16_ ( .D(ph_L[4]), .CK(clk), .Q(FF4_out[16]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_17_ ( .D(ph_L[5]), .CK(clk), .Q(FF4_out[17]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_18_ ( .D(pl_H[0]), .CK(clk), .Q(FF4_out[18]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_19_ ( .D(pl_H[1]), .CK(clk), .Q(FF4_out[19]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_20_ ( .D(pl_H[2]), .CK(clk), .Q(FF4_out[20]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_21_ ( .D(pl_H[3]), .CK(clk), .Q(FF4_out[21]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_22_ ( .D(pl_H[4]), .CK(clk), .Q(FF4_out[22]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_23_ ( .D(pl_H[5]), .CK(clk), .Q(FF4_out[23]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_24_ ( .D(p_H[0]), .CK(clk), .Q(
        Inst_f5_phwillwin_pw2_1_), .QN() );
  DFF_X1 PL_4_s_current_state_reg_25_ ( .D(p_H[1]), .CK(clk), .Q(FF4_out[25]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_26_ ( .D(p_H[2]), .CK(clk), .Q(
        Inst_f5_phwillwin_pw2_3_), .QN() );
  DFF_X1 PL_4_s_current_state_reg_27_ ( .D(p_H[3]), .CK(clk), .Q(FF4_out[27]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_28_ ( .D(p_H[4]), .CK(clk), .Q(
        Inst_f5_phwillwin_pw2_5_), .QN() );
  DFF_X1 PL_4_s_current_state_reg_29_ ( .D(p_H[5]), .CK(clk), .Q(FF4_out[29]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_30_ ( .D(ph_H[0]), .CK(clk), .Q(FF4_out[30]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_31_ ( .D(ph_H[1]), .CK(clk), .Q(FF4_out[31]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_32_ ( .D(ph_H[2]), .CK(clk), .Q(FF4_out[32]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_33_ ( .D(ph_H[3]), .CK(clk), .Q(FF4_out[33]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_34_ ( .D(ph_H[4]), .CK(clk), .Q(FF4_out[34]), 
        .QN() );
  DFF_X1 PL_4_s_current_state_reg_35_ ( .D(ph_H[5]), .CK(clk), .Q(FF4_out[35]), 
        .QN() );
  XOR2_X1 Inst_f5_phwillwin_U12 ( .A(Inst_f5_phwillwin_pw2_5_), .B(FF4_out[23]), .Z(Inst_f5_ph[9]) );
  XOR2_X1 Inst_f5_phwillwin_U11 ( .A(Inst_f5_phwillwin_pw2_4_), .B(FF4_out[22]), .Z(Inst_f5_ph[8]) );
  XOR2_X1 Inst_f5_phwillwin_U10 ( .A(Inst_f5_phwillwin_pw2_3_), .B(FF4_out[33]), .Z(Inst_f5_ph[7]) );
  XOR2_X1 Inst_f5_phwillwin_U9 ( .A(Inst_f5_phwillwin_pw2_2_), .B(FF4_out[32]), 
        .Z(Inst_f5_ph[6]) );
  XOR2_X1 Inst_f5_phwillwin_U8 ( .A(Inst_f5_phwillwin_pw2_3_), .B(FF4_out[21]), 
        .Z(Inst_f5_ph[5]) );
  XOR2_X1 Inst_f5_phwillwin_U7 ( .A(Inst_f5_phwillwin_pw2_2_), .B(FF4_out[20]), 
        .Z(Inst_f5_ph[4]) );
  XOR2_X1 Inst_f5_phwillwin_U6 ( .A(Inst_f5_phwillwin_pw2_1_), .B(FF4_out[31]), 
        .Z(Inst_f5_ph[3]) );
  XOR2_X1 Inst_f5_phwillwin_U5 ( .A(Inst_f5_phwillwin_pw2_0_), .B(FF4_out[30]), 
        .Z(Inst_f5_ph[2]) );
  XOR2_X1 Inst_f5_phwillwin_U4 ( .A(Inst_f5_phwillwin_pw2_1_), .B(FF4_out[19]), 
        .Z(Inst_f5_ph[1]) );
  XOR2_X1 Inst_f5_phwillwin_U3 ( .A(Inst_f5_phwillwin_pw2_5_), .B(FF4_out[35]), 
        .Z(Inst_f5_ph[11]) );
  XOR2_X1 Inst_f5_phwillwin_U2 ( .A(Inst_f5_phwillwin_pw2_4_), .B(FF4_out[34]), 
        .Z(Inst_f5_ph[10]) );
  XOR2_X1 Inst_f5_phwillwin_U1 ( .A(Inst_f5_phwillwin_pw2_0_), .B(FF4_out[18]), 
        .Z(Inst_f5_ph[0]) );
  XOR2_X1 Inst_f5_phwillwin_NxGAMMA_U3 ( .A(Inst_f5_phwillwin_pw2_5_), .B(
        FF4_out[29]), .Z(Inst_f5_phwillwin_pw2_4_) );
  XOR2_X1 Inst_f5_phwillwin_NxGAMMA_U2 ( .A(Inst_f5_phwillwin_pw2_3_), .B(
        FF4_out[27]), .Z(Inst_f5_phwillwin_pw2_2_) );
  XOR2_X1 Inst_f5_phwillwin_NxGAMMA_U1 ( .A(Inst_f5_phwillwin_pw2_1_), .B(
        FF4_out[25]), .Z(Inst_f5_phwillwin_pw2_0_) );
  XOR2_X1 Inst_f5_plwillwin_U12 ( .A(Inst_f5_plwillwin_pw2_5_), .B(FF4_out[5]), 
        .Z(Inst_f5_pl[9]) );
  XOR2_X1 Inst_f5_plwillwin_U11 ( .A(Inst_f5_plwillwin_pw2_4_), .B(FF4_out[4]), 
        .Z(Inst_f5_pl[8]) );
  XOR2_X1 Inst_f5_plwillwin_U10 ( .A(Inst_f5_plwillwin_pw2_3_), .B(FF4_out[15]), .Z(Inst_f5_pl[7]) );
  XOR2_X1 Inst_f5_plwillwin_U9 ( .A(Inst_f5_plwillwin_pw2_2_), .B(FF4_out[14]), 
        .Z(Inst_f5_pl[6]) );
  XOR2_X1 Inst_f5_plwillwin_U8 ( .A(Inst_f5_plwillwin_pw2_3_), .B(FF4_out[3]), 
        .Z(Inst_f5_pl[5]) );
  XOR2_X1 Inst_f5_plwillwin_U7 ( .A(Inst_f5_plwillwin_pw2_2_), .B(FF4_out[2]), 
        .Z(Inst_f5_pl[4]) );
  XOR2_X1 Inst_f5_plwillwin_U6 ( .A(Inst_f5_plwillwin_pw2_1_), .B(FF4_out[13]), 
        .Z(Inst_f5_pl[3]) );
  XOR2_X1 Inst_f5_plwillwin_U5 ( .A(Inst_f5_plwillwin_pw2_0_), .B(FF4_out[12]), 
        .Z(Inst_f5_pl[2]) );
  XOR2_X1 Inst_f5_plwillwin_U4 ( .A(Inst_f5_plwillwin_pw2_1_), .B(FF4_out[1]), 
        .Z(Inst_f5_pl[1]) );
  XOR2_X1 Inst_f5_plwillwin_U3 ( .A(Inst_f5_plwillwin_pw2_5_), .B(FF4_out[17]), 
        .Z(Inst_f5_pl[11]) );
  XOR2_X1 Inst_f5_plwillwin_U2 ( .A(Inst_f5_plwillwin_pw2_4_), .B(FF4_out[16]), 
        .Z(Inst_f5_pl[10]) );
  XOR2_X1 Inst_f5_plwillwin_U1 ( .A(Inst_f5_plwillwin_pw2_0_), .B(FF4_out[0]), 
        .Z(Inst_f5_pl[0]) );
  XOR2_X1 Inst_f5_plwillwin_NxGAMMA_U3 ( .A(Inst_f5_plwillwin_pw2_5_), .B(
        FF4_out[11]), .Z(Inst_f5_plwillwin_pw2_4_) );
  XOR2_X1 Inst_f5_plwillwin_NxGAMMA_U2 ( .A(Inst_f5_plwillwin_pw2_3_), .B(
        FF4_out[9]), .Z(Inst_f5_plwillwin_pw2_2_) );
  XOR2_X1 Inst_f5_plwillwin_NxGAMMA_U1 ( .A(Inst_f5_plwillwin_pw2_1_), .B(
        FF4_out[7]), .Z(Inst_f5_plwillwin_pw2_0_) );
  XOR2_X1 Inst_f5_invlinearMapping_U33 ( .A(Inst_f5_pl[5]), .B(
        Inst_f5_invlinearMapping_n9), .Z(Q[8]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U32 ( .A(Q[4]), .B(
        Inst_f5_invlinearMapping_n8), .ZN(Q[3]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U31 ( .A(Q[5]), .B(
        Inst_f5_invlinearMapping_n7), .ZN(Q[2]) );
  XOR2_X1 Inst_f5_invlinearMapping_U30 ( .A(Q[7]), .B(Inst_f5_pl[2]), .Z(
        Inst_f5_invlinearMapping_n7) );
  XNOR2_X1 Inst_f5_invlinearMapping_U29 ( .A(Inst_f5_ph[2]), .B(Inst_f5_pl[0]), 
        .ZN(Q[5]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U28 ( .A(Q[20]), .B(
        Inst_f5_invlinearMapping_n6), .ZN(Q[19]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U27 ( .A(Q[21]), .B(
        Inst_f5_invlinearMapping_n5), .ZN(Q[18]) );
  XOR2_X1 Inst_f5_invlinearMapping_U26 ( .A(Q[23]), .B(Inst_f5_pl[10]), .Z(
        Inst_f5_invlinearMapping_n5) );
  XNOR2_X1 Inst_f5_invlinearMapping_U25 ( .A(Inst_f5_ph[10]), .B(Inst_f5_pl[8]), .ZN(Q[21]) );
  XOR2_X1 Inst_f5_invlinearMapping_U24 ( .A(Inst_f5_pl[9]), .B(
        Inst_f5_invlinearMapping_n6), .Z(Q[16]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U23 ( .A(Inst_f5_ph[10]), .B(Inst_f5_ph[8]), .ZN(Inst_f5_invlinearMapping_n6) );
  XNOR2_X1 Inst_f5_invlinearMapping_U22 ( .A(Q[12]), .B(
        Inst_f5_invlinearMapping_n9), .ZN(Q[11]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U21 ( .A(Inst_f5_ph[6]), .B(Inst_f5_ph[4]), 
        .ZN(Inst_f5_invlinearMapping_n9) );
  XNOR2_X1 Inst_f5_invlinearMapping_U20 ( .A(Q[13]), .B(
        Inst_f5_invlinearMapping_n4), .ZN(Q[10]) );
  XOR2_X1 Inst_f5_invlinearMapping_U19 ( .A(Q[15]), .B(Inst_f5_pl[6]), .Z(
        Inst_f5_invlinearMapping_n4) );
  XNOR2_X1 Inst_f5_invlinearMapping_U18 ( .A(Inst_f5_ph[6]), .B(Inst_f5_pl[4]), 
        .ZN(Q[13]) );
  XOR2_X1 Inst_f5_invlinearMapping_U17 ( .A(Inst_f5_pl[1]), .B(
        Inst_f5_invlinearMapping_n8), .Z(Q[0]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U16 ( .A(Inst_f5_ph[2]), .B(Inst_f5_ph[0]), 
        .ZN(Inst_f5_invlinearMapping_n8) );
  XNOR2_X1 Inst_f5_invlinearMapping_U15 ( .A(Inst_f5_ph[9]), .B(Q[22]), .ZN(
        Q[20]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U14 ( .A(Inst_f5_pl[11]), .B(
        Inst_f5_ph[11]), .ZN(Q[22]) );
  XOR2_X1 Inst_f5_invlinearMapping_U13 ( .A(Inst_f5_ph[9]), .B(Inst_f5_pl[11]), 
        .Z(Q[23]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U12 ( .A(Inst_f5_pl[5]), .B(
        Inst_f5_invlinearMapping_n3), .ZN(Q[9]) );
  XOR2_X1 Inst_f5_invlinearMapping_U11 ( .A(Inst_f5_ph[5]), .B(Inst_f5_ph[4]), 
        .Z(Inst_f5_invlinearMapping_n3) );
  XNOR2_X1 Inst_f5_invlinearMapping_U10 ( .A(Inst_f5_ph[5]), .B(Q[14]), .ZN(
        Q[12]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U9 ( .A(Inst_f5_pl[7]), .B(Inst_f5_ph[7]), 
        .ZN(Q[14]) );
  XOR2_X1 Inst_f5_invlinearMapping_U8 ( .A(Inst_f5_ph[5]), .B(Inst_f5_pl[7]), 
        .Z(Q[15]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U7 ( .A(Inst_f5_pl[1]), .B(
        Inst_f5_invlinearMapping_n2), .ZN(Q[1]) );
  XOR2_X1 Inst_f5_invlinearMapping_U6 ( .A(Inst_f5_ph[1]), .B(Inst_f5_ph[0]), 
        .Z(Inst_f5_invlinearMapping_n2) );
  XNOR2_X1 Inst_f5_invlinearMapping_U5 ( .A(Inst_f5_pl[9]), .B(
        Inst_f5_invlinearMapping_n1), .ZN(Q[17]) );
  XOR2_X1 Inst_f5_invlinearMapping_U4 ( .A(Inst_f5_ph[9]), .B(Inst_f5_ph[8]), 
        .Z(Inst_f5_invlinearMapping_n1) );
  XNOR2_X1 Inst_f5_invlinearMapping_U3 ( .A(Inst_f5_ph[1]), .B(Q[6]), .ZN(Q[4]) );
  XNOR2_X1 Inst_f5_invlinearMapping_U2 ( .A(Inst_f5_pl[3]), .B(Inst_f5_ph[3]), 
        .ZN(Q[6]) );
  XOR2_X1 Inst_f5_invlinearMapping_U1 ( .A(Inst_f5_ph[1]), .B(Inst_f5_pl[3]), 
        .Z(Q[7]) );
endmodule

