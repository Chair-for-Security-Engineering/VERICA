
module ICINI4 ( port_a_0, port_a_1, port_a_2, port_b_0, port_b_1, port_b_2, 
        port_c_0, port_c_1, port_c_2, port_rand_ref, port_rand_mul_0, 
        port_rand_mul_1, port_rand_mul_2, clk, reset );
  input [4:0] port_a_0;
  input [4:0] port_a_1;
  input [4:0] port_a_2;
  input [4:0] port_b_0;
  input [4:0] port_b_1;
  input [4:0] port_b_2;
  output [4:0] port_c_0;
  output [4:0] port_c_1;
  output [4:0] port_c_2;
  input [5:0] port_rand_ref;
  input [1:0] port_rand_mul_0;
  input [1:0] port_rand_mul_1;
  input [1:0] port_rand_mul_2;
  input clk, reset;
  wire   simpleXor_120_port_a0, simpleXor_120_port_z, simpleXor_121_port_z,
         simpleXor_122_port_a0, simpleXor_122_port_z, simpleXor_123_port_z,
         simpleXor_124_port_a0, simpleXor_124_port_z, simpleXor_125_port_z,
         simpleXor_126_port_a0, simpleXor_126_port_z, simpleXor_127_port_z,
         simpleXor_128_port_a0, simpleXor_128_port_z, simpleXor_129_port_z,
         simpleXor_130_port_a0, simpleXor_130_port_z, simpleXor_131_port_z,
         simpleXor_132_port_a0, simpleXor_132_port_z, simpleXor_133_port_z,
         simpleXor_134_port_a0, simpleXor_134_port_z, simpleXor_135_port_z,
         simpleXor_136_port_a0, simpleXor_136_port_z, simpleXor_137_port_z,
         simpleXor_138_port_a0, simpleXor_138_port_z, simpleXor_139_port_z,
         simpleXor_140_port_a0, simpleXor_140_port_z, simpleXor_141_port_z,
         simpleXor_142_port_a0, simpleXor_142_port_z, simpleXor_143_port_z,
         simpleXor_144_port_a0, simpleXor_144_port_z, simpleXor_145_port_z,
         simpleXor_146_port_a0, simpleXor_146_port_z, simpleXor_147_port_z,
         simpleXor_148_port_a0, simpleXor_148_port_z, simpleXor_149_port_z,
         simpleXor_150_port_a0, simpleXor_150_port_z, simpleXor_151_port_z,
         simpleXor_152_port_a0, simpleXor_152_port_z, simpleXor_153_port_z,
         simpleXor_154_port_a0, simpleXor_154_port_z, simpleXor_155_port_z,
         simpleXor_156_port_a0, simpleXor_156_port_z, simpleXor_157_port_z,
         simpleXor_158_port_a0, simpleXor_158_port_z, simpleXor_159_port_z,
         simpleXor_160_port_a0, simpleXor_160_port_z, simpleXor_161_port_z,
         simpleXor_162_port_a0, simpleXor_162_port_z, simpleXor_163_port_z,
         simpleXor_164_port_a0, simpleXor_164_port_z, simpleXor_165_port_z,
         simpleXor_166_port_a0, simpleXor_166_port_z, simpleXor_167_port_z,
         simpleXor_168_port_a0, simpleXor_168_port_z, simpleXor_169_port_z,
         simpleXor_170_port_a0, simpleXor_170_port_z, simpleXor_171_port_z,
         simpleXor_172_port_a0, simpleXor_172_port_z, simpleXor_173_port_z,
         simpleXor_174_port_a0, simpleXor_174_port_z, simpleXor_175_port_z,
         simpleXor_176_port_a0, simpleXor_176_port_z, simpleXor_177_port_z,
         simpleXor_178_port_a0, simpleXor_178_port_z, simpleXor_179_port_z, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, ref_1_n30,
         ref_1_n29, ref_1_n28, ref_1_n27, ref_1_n26, ref_1_n25, ref_1_n24,
         ref_1_n23, ref_1_n22, ref_1_n21, ref_1_n20, ref_1_n19, ref_1_n18,
         ref_1_n17, ref_1_n16, ref_1_n15, ref_1_n14, ref_1_n13, ref_1_n12,
         ref_1_n11, ref_1_n10, ref_1_n9, ref_1_n8, ref_1_n7, ref_1_n6,
         ref_1_n5, ref_1_n4, ref_1_n3, ref_1_n2, ref_1_n1, ref_1_maj_89_port_o,
         ref_1_maj_88_port_o, ref_1_maj_87_port_o, ref_1_maj_86_port_o,
         ref_1_maj_85_port_o, ref_1_maj_84_port_o, ref_1_maj_83_port_o,
         ref_1_maj_82_port_o, ref_1_maj_81_port_o, ref_1_maj_80_port_o,
         ref_1_maj_79_port_o, ref_1_maj_78_port_o, ref_1_maj_77_port_o,
         ref_1_maj_76_port_o, ref_1_maj_75_port_o, ref_1_maj_74_port_o,
         ref_1_maj_73_port_o, ref_1_maj_72_port_o, ref_1_maj_71_port_o,
         ref_1_maj_70_port_o, ref_1_maj_69_port_o, ref_1_maj_68_port_o,
         ref_1_maj_67_port_o, ref_1_maj_66_port_o, ref_1_maj_65_port_o,
         ref_1_maj_64_port_o, ref_1_maj_63_port_o, ref_1_maj_62_port_o,
         ref_1_maj_61_port_o, ref_1_maj_60_port_o, ref_1_maj_59_port_o,
         ref_1_maj_58_port_o, ref_1_maj_57_port_o, ref_1_maj_56_port_o,
         ref_1_maj_55_port_o, ref_1_maj_54_port_o, ref_1_maj_53_port_o,
         ref_1_maj_52_port_o, ref_1_maj_51_port_o, ref_1_refreshed_2_0_,
         ref_1_refreshed_2_1_, ref_1_refreshed_2_2_, ref_1_refreshed_2_3_,
         ref_1_refreshed_2_4_, ref_1_maj_50_port_o, ref_1_maj_49_port_o,
         ref_1_maj_48_port_o, ref_1_refreshed_1_0_, ref_1_refreshed_1_1_,
         ref_1_refreshed_1_2_, ref_1_refreshed_1_3_, ref_1_refreshed_1_4_,
         ref_1_maj_47_port_o, ref_1_maj_46_port_o, ref_1_maj_45_port_o,
         ref_1_refreshed_0_0_, ref_1_refreshed_0_1_, ref_1_refreshed_0_2_,
         ref_1_refreshed_0_3_, ref_1_refreshed_0_4_,
         ref_1_simpleXor_178_port_z, ref_1_simpleXor_177_port_z,
         ref_1_simpleXor_176_port_z, ref_1_simpleXor_174_port_z,
         ref_1_simpleXor_173_port_z, ref_1_simpleXor_172_port_z,
         ref_1_simpleXor_170_port_z, ref_1_simpleXor_169_port_z,
         ref_1_simpleXor_168_port_z, ref_1_simpleXor_166_port_z,
         ref_1_simpleXor_165_port_z, ref_1_simpleXor_164_port_z,
         ref_1_simpleXor_162_port_z, ref_1_simpleXor_161_port_z,
         ref_1_simpleXor_160_port_z, ref_1_simpleXor_158_port_z,
         ref_1_simpleXor_157_port_z, ref_1_simpleXor_156_port_z,
         ref_1_simpleXor_154_port_z, ref_1_simpleXor_153_port_z,
         ref_1_simpleXor_152_port_z, ref_1_simpleXor_150_port_z,
         ref_1_simpleXor_149_port_z, ref_1_simpleXor_148_port_z,
         ref_1_simpleXor_146_port_z, ref_1_simpleXor_145_port_z,
         ref_1_simpleXor_144_port_z, ref_1_simpleXor_142_port_z,
         ref_1_simpleXor_141_port_z, ref_1_simpleXor_140_port_z,
         ref_1_simpleXor_138_port_z, ref_1_simpleXor_137_port_z,
         ref_1_simpleXor_136_port_z, ref_1_simpleXor_134_port_z,
         ref_1_simpleXor_133_port_z, ref_1_simpleXor_132_port_z,
         ref_1_simpleXor_130_port_z, ref_1_simpleXor_129_port_z,
         ref_1_simpleXor_128_port_z, ref_1_simpleXor_126_port_z,
         ref_1_simpleXor_125_port_z, ref_1_simpleXor_124_port_z,
         ref_1_simpleXor_122_port_z, ref_1_simpleXor_121_port_z,
         ref_1_simpleXor_120_port_z, ref_1_maj_45_n13, ref_1_maj_45_n12,
         ref_1_maj_45_n11, ref_1_maj_45_n10, ref_1_maj_45_n9, ref_1_maj_45_n8,
         ref_1_maj_45_n7, ref_1_maj_45_n6, ref_1_maj_45_n5, ref_1_maj_45_n4,
         ref_1_maj_45_n3, ref_1_maj_45_n2, ref_1_maj_45_n1, ref_1_maj_46_n26,
         ref_1_maj_46_n25, ref_1_maj_46_n24, ref_1_maj_46_n23,
         ref_1_maj_46_n22, ref_1_maj_46_n21, ref_1_maj_46_n20,
         ref_1_maj_46_n19, ref_1_maj_46_n18, ref_1_maj_46_n17,
         ref_1_maj_46_n16, ref_1_maj_46_n15, ref_1_maj_46_n14,
         ref_1_maj_47_n26, ref_1_maj_47_n25, ref_1_maj_47_n24,
         ref_1_maj_47_n23, ref_1_maj_47_n22, ref_1_maj_47_n21,
         ref_1_maj_47_n20, ref_1_maj_47_n19, ref_1_maj_47_n18,
         ref_1_maj_47_n17, ref_1_maj_47_n16, ref_1_maj_47_n15,
         ref_1_maj_47_n14, ref_1_maj_48_n26, ref_1_maj_48_n25,
         ref_1_maj_48_n24, ref_1_maj_48_n23, ref_1_maj_48_n22,
         ref_1_maj_48_n21, ref_1_maj_48_n20, ref_1_maj_48_n19,
         ref_1_maj_48_n18, ref_1_maj_48_n17, ref_1_maj_48_n16,
         ref_1_maj_48_n15, ref_1_maj_48_n14, ref_1_maj_49_n26,
         ref_1_maj_49_n25, ref_1_maj_49_n24, ref_1_maj_49_n23,
         ref_1_maj_49_n22, ref_1_maj_49_n21, ref_1_maj_49_n20,
         ref_1_maj_49_n19, ref_1_maj_49_n18, ref_1_maj_49_n17,
         ref_1_maj_49_n16, ref_1_maj_49_n15, ref_1_maj_49_n14,
         ref_1_maj_50_n26, ref_1_maj_50_n25, ref_1_maj_50_n24,
         ref_1_maj_50_n23, ref_1_maj_50_n22, ref_1_maj_50_n21,
         ref_1_maj_50_n20, ref_1_maj_50_n19, ref_1_maj_50_n18,
         ref_1_maj_50_n17, ref_1_maj_50_n16, ref_1_maj_50_n15,
         ref_1_maj_50_n14, ref_1_maj_51_n26, ref_1_maj_51_n25,
         ref_1_maj_51_n24, ref_1_maj_51_n23, ref_1_maj_51_n22,
         ref_1_maj_51_n21, ref_1_maj_51_n20, ref_1_maj_51_n19,
         ref_1_maj_51_n18, ref_1_maj_51_n17, ref_1_maj_51_n16,
         ref_1_maj_51_n15, ref_1_maj_51_n14, ref_1_maj_52_n26,
         ref_1_maj_52_n25, ref_1_maj_52_n24, ref_1_maj_52_n23,
         ref_1_maj_52_n22, ref_1_maj_52_n21, ref_1_maj_52_n20,
         ref_1_maj_52_n19, ref_1_maj_52_n18, ref_1_maj_52_n17,
         ref_1_maj_52_n16, ref_1_maj_52_n15, ref_1_maj_52_n14,
         ref_1_maj_53_n26, ref_1_maj_53_n25, ref_1_maj_53_n24,
         ref_1_maj_53_n23, ref_1_maj_53_n22, ref_1_maj_53_n21,
         ref_1_maj_53_n20, ref_1_maj_53_n19, ref_1_maj_53_n18,
         ref_1_maj_53_n17, ref_1_maj_53_n16, ref_1_maj_53_n15,
         ref_1_maj_53_n14, ref_1_maj_54_n26, ref_1_maj_54_n25,
         ref_1_maj_54_n24, ref_1_maj_54_n23, ref_1_maj_54_n22,
         ref_1_maj_54_n21, ref_1_maj_54_n20, ref_1_maj_54_n19,
         ref_1_maj_54_n18, ref_1_maj_54_n17, ref_1_maj_54_n16,
         ref_1_maj_54_n15, ref_1_maj_54_n14, ref_1_maj_55_n26,
         ref_1_maj_55_n25, ref_1_maj_55_n24, ref_1_maj_55_n23,
         ref_1_maj_55_n22, ref_1_maj_55_n21, ref_1_maj_55_n20,
         ref_1_maj_55_n19, ref_1_maj_55_n18, ref_1_maj_55_n17,
         ref_1_maj_55_n16, ref_1_maj_55_n15, ref_1_maj_55_n14,
         ref_1_maj_56_n26, ref_1_maj_56_n25, ref_1_maj_56_n24,
         ref_1_maj_56_n23, ref_1_maj_56_n22, ref_1_maj_56_n21,
         ref_1_maj_56_n20, ref_1_maj_56_n19, ref_1_maj_56_n18,
         ref_1_maj_56_n17, ref_1_maj_56_n16, ref_1_maj_56_n15,
         ref_1_maj_56_n14, ref_1_maj_57_n26, ref_1_maj_57_n25,
         ref_1_maj_57_n24, ref_1_maj_57_n23, ref_1_maj_57_n22,
         ref_1_maj_57_n21, ref_1_maj_57_n20, ref_1_maj_57_n19,
         ref_1_maj_57_n18, ref_1_maj_57_n17, ref_1_maj_57_n16,
         ref_1_maj_57_n15, ref_1_maj_57_n14, ref_1_maj_58_n26,
         ref_1_maj_58_n25, ref_1_maj_58_n24, ref_1_maj_58_n23,
         ref_1_maj_58_n22, ref_1_maj_58_n21, ref_1_maj_58_n20,
         ref_1_maj_58_n19, ref_1_maj_58_n18, ref_1_maj_58_n17,
         ref_1_maj_58_n16, ref_1_maj_58_n15, ref_1_maj_58_n14,
         ref_1_maj_59_n26, ref_1_maj_59_n25, ref_1_maj_59_n24,
         ref_1_maj_59_n23, ref_1_maj_59_n22, ref_1_maj_59_n21,
         ref_1_maj_59_n20, ref_1_maj_59_n19, ref_1_maj_59_n18,
         ref_1_maj_59_n17, ref_1_maj_59_n16, ref_1_maj_59_n15,
         ref_1_maj_59_n14, ref_1_maj_60_n26, ref_1_maj_60_n25,
         ref_1_maj_60_n24, ref_1_maj_60_n23, ref_1_maj_60_n22,
         ref_1_maj_60_n21, ref_1_maj_60_n20, ref_1_maj_60_n19,
         ref_1_maj_60_n18, ref_1_maj_60_n17, ref_1_maj_60_n16,
         ref_1_maj_60_n15, ref_1_maj_60_n14, ref_1_maj_61_n26,
         ref_1_maj_61_n25, ref_1_maj_61_n24, ref_1_maj_61_n23,
         ref_1_maj_61_n22, ref_1_maj_61_n21, ref_1_maj_61_n20,
         ref_1_maj_61_n19, ref_1_maj_61_n18, ref_1_maj_61_n17,
         ref_1_maj_61_n16, ref_1_maj_61_n15, ref_1_maj_61_n14,
         ref_1_maj_62_n26, ref_1_maj_62_n25, ref_1_maj_62_n24,
         ref_1_maj_62_n23, ref_1_maj_62_n22, ref_1_maj_62_n21,
         ref_1_maj_62_n20, ref_1_maj_62_n19, ref_1_maj_62_n18,
         ref_1_maj_62_n17, ref_1_maj_62_n16, ref_1_maj_62_n15,
         ref_1_maj_62_n14, ref_1_maj_63_n26, ref_1_maj_63_n25,
         ref_1_maj_63_n24, ref_1_maj_63_n23, ref_1_maj_63_n22,
         ref_1_maj_63_n21, ref_1_maj_63_n20, ref_1_maj_63_n19,
         ref_1_maj_63_n18, ref_1_maj_63_n17, ref_1_maj_63_n16,
         ref_1_maj_63_n15, ref_1_maj_63_n14, ref_1_maj_64_n26,
         ref_1_maj_64_n25, ref_1_maj_64_n24, ref_1_maj_64_n23,
         ref_1_maj_64_n22, ref_1_maj_64_n21, ref_1_maj_64_n20,
         ref_1_maj_64_n19, ref_1_maj_64_n18, ref_1_maj_64_n17,
         ref_1_maj_64_n16, ref_1_maj_64_n15, ref_1_maj_64_n14,
         ref_1_maj_65_n26, ref_1_maj_65_n25, ref_1_maj_65_n24,
         ref_1_maj_65_n23, ref_1_maj_65_n22, ref_1_maj_65_n21,
         ref_1_maj_65_n20, ref_1_maj_65_n19, ref_1_maj_65_n18,
         ref_1_maj_65_n17, ref_1_maj_65_n16, ref_1_maj_65_n15,
         ref_1_maj_65_n14, ref_1_maj_66_n26, ref_1_maj_66_n25,
         ref_1_maj_66_n24, ref_1_maj_66_n23, ref_1_maj_66_n22,
         ref_1_maj_66_n21, ref_1_maj_66_n20, ref_1_maj_66_n19,
         ref_1_maj_66_n18, ref_1_maj_66_n17, ref_1_maj_66_n16,
         ref_1_maj_66_n15, ref_1_maj_66_n14, ref_1_maj_67_n26,
         ref_1_maj_67_n25, ref_1_maj_67_n24, ref_1_maj_67_n23,
         ref_1_maj_67_n22, ref_1_maj_67_n21, ref_1_maj_67_n20,
         ref_1_maj_67_n19, ref_1_maj_67_n18, ref_1_maj_67_n17,
         ref_1_maj_67_n16, ref_1_maj_67_n15, ref_1_maj_67_n14,
         ref_1_maj_68_n26, ref_1_maj_68_n25, ref_1_maj_68_n24,
         ref_1_maj_68_n23, ref_1_maj_68_n22, ref_1_maj_68_n21,
         ref_1_maj_68_n20, ref_1_maj_68_n19, ref_1_maj_68_n18,
         ref_1_maj_68_n17, ref_1_maj_68_n16, ref_1_maj_68_n15,
         ref_1_maj_68_n14, ref_1_maj_69_n26, ref_1_maj_69_n25,
         ref_1_maj_69_n24, ref_1_maj_69_n23, ref_1_maj_69_n22,
         ref_1_maj_69_n21, ref_1_maj_69_n20, ref_1_maj_69_n19,
         ref_1_maj_69_n18, ref_1_maj_69_n17, ref_1_maj_69_n16,
         ref_1_maj_69_n15, ref_1_maj_69_n14, ref_1_maj_70_n26,
         ref_1_maj_70_n25, ref_1_maj_70_n24, ref_1_maj_70_n23,
         ref_1_maj_70_n22, ref_1_maj_70_n21, ref_1_maj_70_n20,
         ref_1_maj_70_n19, ref_1_maj_70_n18, ref_1_maj_70_n17,
         ref_1_maj_70_n16, ref_1_maj_70_n15, ref_1_maj_70_n14,
         ref_1_maj_71_n26, ref_1_maj_71_n25, ref_1_maj_71_n24,
         ref_1_maj_71_n23, ref_1_maj_71_n22, ref_1_maj_71_n21,
         ref_1_maj_71_n20, ref_1_maj_71_n19, ref_1_maj_71_n18,
         ref_1_maj_71_n17, ref_1_maj_71_n16, ref_1_maj_71_n15,
         ref_1_maj_71_n14, ref_1_maj_72_n26, ref_1_maj_72_n25,
         ref_1_maj_72_n24, ref_1_maj_72_n23, ref_1_maj_72_n22,
         ref_1_maj_72_n21, ref_1_maj_72_n20, ref_1_maj_72_n19,
         ref_1_maj_72_n18, ref_1_maj_72_n17, ref_1_maj_72_n16,
         ref_1_maj_72_n15, ref_1_maj_72_n14, ref_1_maj_73_n26,
         ref_1_maj_73_n25, ref_1_maj_73_n24, ref_1_maj_73_n23,
         ref_1_maj_73_n22, ref_1_maj_73_n21, ref_1_maj_73_n20,
         ref_1_maj_73_n19, ref_1_maj_73_n18, ref_1_maj_73_n17,
         ref_1_maj_73_n16, ref_1_maj_73_n15, ref_1_maj_73_n14,
         ref_1_maj_74_n26, ref_1_maj_74_n25, ref_1_maj_74_n24,
         ref_1_maj_74_n23, ref_1_maj_74_n22, ref_1_maj_74_n21,
         ref_1_maj_74_n20, ref_1_maj_74_n19, ref_1_maj_74_n18,
         ref_1_maj_74_n17, ref_1_maj_74_n16, ref_1_maj_74_n15,
         ref_1_maj_74_n14, ref_1_maj_75_n26, ref_1_maj_75_n25,
         ref_1_maj_75_n24, ref_1_maj_75_n23, ref_1_maj_75_n22,
         ref_1_maj_75_n21, ref_1_maj_75_n20, ref_1_maj_75_n19,
         ref_1_maj_75_n18, ref_1_maj_75_n17, ref_1_maj_75_n16,
         ref_1_maj_75_n15, ref_1_maj_75_n14, ref_1_maj_76_n26,
         ref_1_maj_76_n25, ref_1_maj_76_n24, ref_1_maj_76_n23,
         ref_1_maj_76_n22, ref_1_maj_76_n21, ref_1_maj_76_n20,
         ref_1_maj_76_n19, ref_1_maj_76_n18, ref_1_maj_76_n17,
         ref_1_maj_76_n16, ref_1_maj_76_n15, ref_1_maj_76_n14,
         ref_1_maj_77_n26, ref_1_maj_77_n25, ref_1_maj_77_n24,
         ref_1_maj_77_n23, ref_1_maj_77_n22, ref_1_maj_77_n21,
         ref_1_maj_77_n20, ref_1_maj_77_n19, ref_1_maj_77_n18,
         ref_1_maj_77_n17, ref_1_maj_77_n16, ref_1_maj_77_n15,
         ref_1_maj_77_n14, ref_1_maj_78_n26, ref_1_maj_78_n25,
         ref_1_maj_78_n24, ref_1_maj_78_n23, ref_1_maj_78_n22,
         ref_1_maj_78_n21, ref_1_maj_78_n20, ref_1_maj_78_n19,
         ref_1_maj_78_n18, ref_1_maj_78_n17, ref_1_maj_78_n16,
         ref_1_maj_78_n15, ref_1_maj_78_n14, ref_1_maj_79_n26,
         ref_1_maj_79_n25, ref_1_maj_79_n24, ref_1_maj_79_n23,
         ref_1_maj_79_n22, ref_1_maj_79_n21, ref_1_maj_79_n20,
         ref_1_maj_79_n19, ref_1_maj_79_n18, ref_1_maj_79_n17,
         ref_1_maj_79_n16, ref_1_maj_79_n15, ref_1_maj_79_n14,
         ref_1_maj_80_n26, ref_1_maj_80_n25, ref_1_maj_80_n24,
         ref_1_maj_80_n23, ref_1_maj_80_n22, ref_1_maj_80_n21,
         ref_1_maj_80_n20, ref_1_maj_80_n19, ref_1_maj_80_n18,
         ref_1_maj_80_n17, ref_1_maj_80_n16, ref_1_maj_80_n15,
         ref_1_maj_80_n14, ref_1_maj_81_n26, ref_1_maj_81_n25,
         ref_1_maj_81_n24, ref_1_maj_81_n23, ref_1_maj_81_n22,
         ref_1_maj_81_n21, ref_1_maj_81_n20, ref_1_maj_81_n19,
         ref_1_maj_81_n18, ref_1_maj_81_n17, ref_1_maj_81_n16,
         ref_1_maj_81_n15, ref_1_maj_81_n14, ref_1_maj_82_n26,
         ref_1_maj_82_n25, ref_1_maj_82_n24, ref_1_maj_82_n23,
         ref_1_maj_82_n22, ref_1_maj_82_n21, ref_1_maj_82_n20,
         ref_1_maj_82_n19, ref_1_maj_82_n18, ref_1_maj_82_n17,
         ref_1_maj_82_n16, ref_1_maj_82_n15, ref_1_maj_82_n14,
         ref_1_maj_83_n26, ref_1_maj_83_n25, ref_1_maj_83_n24,
         ref_1_maj_83_n23, ref_1_maj_83_n22, ref_1_maj_83_n21,
         ref_1_maj_83_n20, ref_1_maj_83_n19, ref_1_maj_83_n18,
         ref_1_maj_83_n17, ref_1_maj_83_n16, ref_1_maj_83_n15,
         ref_1_maj_83_n14, ref_1_maj_84_n26, ref_1_maj_84_n25,
         ref_1_maj_84_n24, ref_1_maj_84_n23, ref_1_maj_84_n22,
         ref_1_maj_84_n21, ref_1_maj_84_n20, ref_1_maj_84_n19,
         ref_1_maj_84_n18, ref_1_maj_84_n17, ref_1_maj_84_n16,
         ref_1_maj_84_n15, ref_1_maj_84_n14, ref_1_maj_85_n26,
         ref_1_maj_85_n25, ref_1_maj_85_n24, ref_1_maj_85_n23,
         ref_1_maj_85_n22, ref_1_maj_85_n21, ref_1_maj_85_n20,
         ref_1_maj_85_n19, ref_1_maj_85_n18, ref_1_maj_85_n17,
         ref_1_maj_85_n16, ref_1_maj_85_n15, ref_1_maj_85_n14,
         ref_1_maj_86_n26, ref_1_maj_86_n25, ref_1_maj_86_n24,
         ref_1_maj_86_n23, ref_1_maj_86_n22, ref_1_maj_86_n21,
         ref_1_maj_86_n20, ref_1_maj_86_n19, ref_1_maj_86_n18,
         ref_1_maj_86_n17, ref_1_maj_86_n16, ref_1_maj_86_n15,
         ref_1_maj_86_n14, ref_1_maj_87_n26, ref_1_maj_87_n25,
         ref_1_maj_87_n24, ref_1_maj_87_n23, ref_1_maj_87_n22,
         ref_1_maj_87_n21, ref_1_maj_87_n20, ref_1_maj_87_n19,
         ref_1_maj_87_n18, ref_1_maj_87_n17, ref_1_maj_87_n16,
         ref_1_maj_87_n15, ref_1_maj_87_n14, ref_1_maj_88_n26,
         ref_1_maj_88_n25, ref_1_maj_88_n24, ref_1_maj_88_n23,
         ref_1_maj_88_n22, ref_1_maj_88_n21, ref_1_maj_88_n20,
         ref_1_maj_88_n19, ref_1_maj_88_n18, ref_1_maj_88_n17,
         ref_1_maj_88_n16, ref_1_maj_88_n15, ref_1_maj_88_n14,
         ref_1_maj_89_n26, ref_1_maj_89_n25, ref_1_maj_89_n24,
         ref_1_maj_89_n23, ref_1_maj_89_n22, ref_1_maj_89_n21,
         ref_1_maj_89_n20, ref_1_maj_89_n19, ref_1_maj_89_n18,
         ref_1_maj_89_n17, ref_1_maj_89_n16, ref_1_maj_89_n15,
         ref_1_maj_89_n14;
  wire   [4:0] ref_1_port_o_0_0;
  wire   [4:0] ref_1_port_o_0_1;
  wire   [4:0] ref_1_port_o_0_2;
  wire   [4:0] ref_1_port_o_1_0;
  wire   [4:0] ref_1_port_o_1_1;
  wire   [4:0] ref_1_port_o_1_2;
  wire   [4:0] ref_1_port_o_2_0;
  wire   [4:0] ref_1_port_o_2_1;
  wire   [4:0] ref_1_port_o_2_2;
  wire   [4:0] temp_0_0;
  wire   [4:0] mult_ab_0_1;
  wire   [4:0] mult_ab_0_2;
  wire   [4:0] temp_0_1;
  wire   [4:0] mult_ab_1_0;
  wire   [4:0] mult_ab_1_2;
  wire   [4:0] temp_0_2;
  wire   [4:0] mult_ab_2_0;
  wire   [4:0] mult_ab_2_1;

  DFF_X1 mult_ab_2_1_reg_4_ ( .D(simpleXor_179_port_z), .CK(clk), .Q(
        mult_ab_2_1[4]), .QN() );
  DFF_X1 mult_ab_2_1_reg_3_ ( .D(simpleXor_167_port_z), .CK(clk), .Q(
        mult_ab_2_1[3]), .QN() );
  DFF_X1 mult_ab_2_1_reg_2_ ( .D(simpleXor_155_port_z), .CK(clk), .Q(
        mult_ab_2_1[2]), .QN() );
  DFF_X1 mult_ab_2_1_reg_1_ ( .D(simpleXor_143_port_z), .CK(clk), .Q(
        mult_ab_2_1[1]), .QN() );
  DFF_X1 mult_ab_2_1_reg_0_ ( .D(simpleXor_131_port_z), .CK(clk), .Q(
        mult_ab_2_1[0]), .QN() );
  DFF_X1 mult_ab_2_2_reg_4_ ( .D(N14), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 mult_ab_2_2_reg_3_ ( .D(N11), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 mult_ab_2_2_reg_2_ ( .D(N8), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 mult_ab_2_2_reg_1_ ( .D(N5), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 mult_ab_2_2_reg_0_ ( .D(N2), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 mult_ab_1_2_reg_4_ ( .D(simpleXor_175_port_z), .CK(clk), .Q(
        mult_ab_1_2[4]), .QN() );
  DFF_X1 mult_ab_1_2_reg_3_ ( .D(simpleXor_163_port_z), .CK(clk), .Q(
        mult_ab_1_2[3]), .QN() );
  DFF_X1 mult_ab_1_2_reg_2_ ( .D(simpleXor_151_port_z), .CK(clk), .Q(
        mult_ab_1_2[2]), .QN() );
  DFF_X1 mult_ab_1_2_reg_1_ ( .D(simpleXor_139_port_z), .CK(clk), .Q(
        mult_ab_1_2[1]), .QN() );
  DFF_X1 mult_ab_1_2_reg_0_ ( .D(simpleXor_127_port_z), .CK(clk), .Q(
        mult_ab_1_2[0]), .QN() );
  DFF_X1 mult_ab_2_0_reg_4_ ( .D(simpleXor_177_port_z), .CK(clk), .Q(
        mult_ab_2_0[4]), .QN() );
  DFF_X1 mult_ab_2_0_reg_3_ ( .D(simpleXor_165_port_z), .CK(clk), .Q(
        mult_ab_2_0[3]), .QN() );
  DFF_X1 mult_ab_2_0_reg_2_ ( .D(simpleXor_153_port_z), .CK(clk), .Q(
        mult_ab_2_0[2]), .QN() );
  DFF_X1 mult_ab_2_0_reg_1_ ( .D(simpleXor_141_port_z), .CK(clk), .Q(
        mult_ab_2_0[1]), .QN() );
  DFF_X1 mult_ab_2_0_reg_0_ ( .D(simpleXor_129_port_z), .CK(clk), .Q(
        mult_ab_2_0[0]), .QN() );
  DFF_X1 mult_ab_1_0_reg_4_ ( .D(simpleXor_173_port_z), .CK(clk), .Q(
        mult_ab_1_0[4]), .QN() );
  DFF_X1 mult_ab_1_0_reg_3_ ( .D(simpleXor_161_port_z), .CK(clk), .Q(
        mult_ab_1_0[3]), .QN() );
  DFF_X1 mult_ab_1_0_reg_2_ ( .D(simpleXor_149_port_z), .CK(clk), .Q(
        mult_ab_1_0[2]), .QN() );
  DFF_X1 mult_ab_1_0_reg_1_ ( .D(simpleXor_137_port_z), .CK(clk), .Q(
        mult_ab_1_0[1]), .QN() );
  DFF_X1 mult_ab_1_0_reg_0_ ( .D(simpleXor_125_port_z), .CK(clk), .Q(
        mult_ab_1_0[0]), .QN() );
  DFF_X1 mult_ab_1_1_reg_4_ ( .D(N13), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 mult_ab_1_1_reg_3_ ( .D(N10), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 mult_ab_1_1_reg_2_ ( .D(N7), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 mult_ab_1_1_reg_1_ ( .D(N4), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 mult_ab_1_1_reg_0_ ( .D(N1), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 mult_ab_0_0_reg_4_ ( .D(N12), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 mult_ab_0_0_reg_3_ ( .D(N9), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 mult_ab_0_0_reg_2_ ( .D(N6), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 mult_ab_0_0_reg_1_ ( .D(N3), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 mult_ab_0_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 mult_ab_0_1_reg_4_ ( .D(simpleXor_169_port_z), .CK(clk), .Q(
        mult_ab_0_1[4]), .QN() );
  DFF_X1 mult_ab_0_1_reg_3_ ( .D(simpleXor_157_port_z), .CK(clk), .Q(
        mult_ab_0_1[3]), .QN() );
  DFF_X1 mult_ab_0_1_reg_2_ ( .D(simpleXor_145_port_z), .CK(clk), .Q(
        mult_ab_0_1[2]), .QN() );
  DFF_X1 mult_ab_0_1_reg_1_ ( .D(simpleXor_133_port_z), .CK(clk), .Q(
        mult_ab_0_1[1]), .QN() );
  DFF_X1 mult_ab_0_1_reg_0_ ( .D(simpleXor_121_port_z), .CK(clk), .Q(
        mult_ab_0_1[0]), .QN() );
  DFF_X1 mult_ab_0_2_reg_4_ ( .D(simpleXor_171_port_z), .CK(clk), .Q(
        mult_ab_0_2[4]), .QN() );
  DFF_X1 mult_ab_0_2_reg_3_ ( .D(simpleXor_159_port_z), .CK(clk), .Q(
        mult_ab_0_2[3]), .QN() );
  DFF_X1 mult_ab_0_2_reg_2_ ( .D(simpleXor_147_port_z), .CK(clk), .Q(
        mult_ab_0_2[2]), .QN() );
  DFF_X1 mult_ab_0_2_reg_1_ ( .D(simpleXor_135_port_z), .CK(clk), .Q(
        mult_ab_0_2[1]), .QN() );
  DFF_X1 mult_ab_0_2_reg_0_ ( .D(simpleXor_123_port_z), .CK(clk), .Q(
        mult_ab_0_2[0]), .QN() );
  AND2_X1 U78 ( .A1(ref_1_port_o_0_2[0]), .A2(port_a_0[0]), .ZN(
        simpleXor_122_port_a0) );
  AND2_X1 U79 ( .A1(ref_1_port_o_0_2[1]), .A2(port_a_0[1]), .ZN(
        simpleXor_134_port_a0) );
  AND2_X1 U80 ( .A1(ref_1_port_o_0_2[2]), .A2(port_a_0[2]), .ZN(
        simpleXor_146_port_a0) );
  AND2_X1 U81 ( .A1(ref_1_port_o_0_2[3]), .A2(port_a_0[3]), .ZN(
        simpleXor_158_port_a0) );
  AND2_X1 U82 ( .A1(ref_1_port_o_0_2[4]), .A2(port_a_0[4]), .ZN(
        simpleXor_170_port_a0) );
  AND2_X1 U83 ( .A1(ref_1_port_o_0_1[0]), .A2(port_a_0[0]), .ZN(
        simpleXor_120_port_a0) );
  AND2_X1 U84 ( .A1(ref_1_port_o_0_1[1]), .A2(port_a_0[1]), .ZN(
        simpleXor_132_port_a0) );
  AND2_X1 U85 ( .A1(ref_1_port_o_0_1[2]), .A2(port_a_0[2]), .ZN(
        simpleXor_144_port_a0) );
  AND2_X1 U86 ( .A1(ref_1_port_o_0_1[3]), .A2(port_a_0[3]), .ZN(
        simpleXor_156_port_a0) );
  AND2_X1 U87 ( .A1(ref_1_port_o_0_1[4]), .A2(port_a_0[4]), .ZN(
        simpleXor_168_port_a0) );
  AND2_X1 U88 ( .A1(ref_1_port_o_1_0[0]), .A2(port_a_1[0]), .ZN(
        simpleXor_124_port_a0) );
  AND2_X1 U89 ( .A1(ref_1_port_o_1_0[1]), .A2(port_a_1[1]), .ZN(
        simpleXor_136_port_a0) );
  AND2_X1 U90 ( .A1(ref_1_port_o_1_0[2]), .A2(port_a_1[2]), .ZN(
        simpleXor_148_port_a0) );
  AND2_X1 U91 ( .A1(ref_1_port_o_1_0[3]), .A2(port_a_1[3]), .ZN(
        simpleXor_160_port_a0) );
  AND2_X1 U92 ( .A1(ref_1_port_o_1_0[4]), .A2(port_a_1[4]), .ZN(
        simpleXor_172_port_a0) );
  AND2_X1 U93 ( .A1(ref_1_port_o_2_0[0]), .A2(port_a_2[0]), .ZN(
        simpleXor_128_port_a0) );
  AND2_X1 U94 ( .A1(ref_1_port_o_2_0[1]), .A2(port_a_2[1]), .ZN(
        simpleXor_140_port_a0) );
  AND2_X1 U95 ( .A1(ref_1_port_o_2_0[2]), .A2(port_a_2[2]), .ZN(
        simpleXor_152_port_a0) );
  AND2_X1 U96 ( .A1(ref_1_port_o_2_0[3]), .A2(port_a_2[3]), .ZN(
        simpleXor_164_port_a0) );
  AND2_X1 U97 ( .A1(ref_1_port_o_2_0[4]), .A2(port_a_2[4]), .ZN(
        simpleXor_176_port_a0) );
  AND2_X1 U98 ( .A1(ref_1_port_o_1_2[0]), .A2(port_a_1[0]), .ZN(
        simpleXor_126_port_a0) );
  AND2_X1 U99 ( .A1(ref_1_port_o_1_2[1]), .A2(port_a_1[1]), .ZN(
        simpleXor_138_port_a0) );
  AND2_X1 U100 ( .A1(ref_1_port_o_1_2[2]), .A2(port_a_1[2]), .ZN(
        simpleXor_150_port_a0) );
  AND2_X1 U101 ( .A1(ref_1_port_o_1_2[3]), .A2(port_a_1[3]), .ZN(
        simpleXor_162_port_a0) );
  AND2_X1 U102 ( .A1(ref_1_port_o_1_2[4]), .A2(port_a_1[4]), .ZN(
        simpleXor_174_port_a0) );
  AND2_X1 U103 ( .A1(ref_1_port_o_2_1[0]), .A2(port_a_2[0]), .ZN(
        simpleXor_130_port_a0) );
  AND2_X1 U104 ( .A1(ref_1_port_o_2_1[1]), .A2(port_a_2[1]), .ZN(
        simpleXor_142_port_a0) );
  AND2_X1 U105 ( .A1(ref_1_port_o_2_1[2]), .A2(port_a_2[2]), .ZN(
        simpleXor_154_port_a0) );
  AND2_X1 U106 ( .A1(ref_1_port_o_2_1[3]), .A2(port_a_2[3]), .ZN(
        simpleXor_166_port_a0) );
  AND2_X1 U107 ( .A1(ref_1_port_o_2_1[4]), .A2(port_a_2[4]), .ZN(
        simpleXor_178_port_a0) );
  AND2_X1 U108 ( .A1(ref_1_port_o_0_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U109 ( .A1(ref_1_port_o_0_0[1]), .A2(port_a_0[1]), .ZN(N3) );
  AND2_X1 U110 ( .A1(ref_1_port_o_0_0[2]), .A2(port_a_0[2]), .ZN(N6) );
  AND2_X1 U111 ( .A1(ref_1_port_o_0_0[3]), .A2(port_a_0[3]), .ZN(N9) );
  AND2_X1 U112 ( .A1(ref_1_port_o_0_0[4]), .A2(port_a_0[4]), .ZN(N12) );
  AND2_X1 U113 ( .A1(ref_1_port_o_1_1[0]), .A2(port_a_1[0]), .ZN(N1) );
  AND2_X1 U114 ( .A1(ref_1_port_o_1_1[1]), .A2(port_a_1[1]), .ZN(N4) );
  AND2_X1 U115 ( .A1(ref_1_port_o_1_1[2]), .A2(port_a_1[2]), .ZN(N7) );
  AND2_X1 U116 ( .A1(ref_1_port_o_1_1[3]), .A2(port_a_1[3]), .ZN(N10) );
  AND2_X1 U117 ( .A1(ref_1_port_o_1_1[4]), .A2(port_a_1[4]), .ZN(N13) );
  AND2_X1 U118 ( .A1(ref_1_port_o_2_2[0]), .A2(port_a_2[0]), .ZN(N2) );
  AND2_X1 U119 ( .A1(ref_1_port_o_2_2[1]), .A2(port_a_2[1]), .ZN(N5) );
  AND2_X1 U120 ( .A1(ref_1_port_o_2_2[2]), .A2(port_a_2[2]), .ZN(N8) );
  AND2_X1 U121 ( .A1(ref_1_port_o_2_2[3]), .A2(port_a_2[3]), .ZN(N11) );
  AND2_X1 U122 ( .A1(ref_1_port_o_2_2[4]), .A2(port_a_2[4]), .ZN(N14) );
  XOR2_X1 U123 ( .A(mult_ab_2_0[0]), .B(n5), .Z(port_c_2[0]) );
  XOR2_X1 U124 ( .A(temp_0_2[0]), .B(mult_ab_2_1[0]), .Z(n5) );
  XOR2_X1 U125 ( .A(mult_ab_2_0[1]), .B(n4), .Z(port_c_2[1]) );
  XOR2_X1 U126 ( .A(temp_0_2[1]), .B(mult_ab_2_1[1]), .Z(n4) );
  XOR2_X1 U127 ( .A(mult_ab_2_0[2]), .B(n3), .Z(port_c_2[2]) );
  XOR2_X1 U128 ( .A(temp_0_2[2]), .B(mult_ab_2_1[2]), .Z(n3) );
  XOR2_X1 U129 ( .A(mult_ab_2_0[3]), .B(n2), .Z(port_c_2[3]) );
  XOR2_X1 U130 ( .A(temp_0_2[3]), .B(mult_ab_2_1[3]), .Z(n2) );
  XOR2_X1 U131 ( .A(mult_ab_2_0[4]), .B(n1), .Z(port_c_2[4]) );
  XOR2_X1 U132 ( .A(temp_0_2[4]), .B(mult_ab_2_1[4]), .Z(n1) );
  XOR2_X1 U133 ( .A(mult_ab_1_0[0]), .B(n10), .Z(port_c_1[0]) );
  XOR2_X1 U134 ( .A(temp_0_1[0]), .B(mult_ab_1_2[0]), .Z(n10) );
  XOR2_X1 U135 ( .A(mult_ab_1_0[1]), .B(n9), .Z(port_c_1[1]) );
  XOR2_X1 U136 ( .A(temp_0_1[1]), .B(mult_ab_1_2[1]), .Z(n9) );
  XOR2_X1 U137 ( .A(mult_ab_1_0[2]), .B(n8), .Z(port_c_1[2]) );
  XOR2_X1 U138 ( .A(temp_0_1[2]), .B(mult_ab_1_2[2]), .Z(n8) );
  XOR2_X1 U139 ( .A(mult_ab_1_0[3]), .B(n7), .Z(port_c_1[3]) );
  XOR2_X1 U140 ( .A(temp_0_1[3]), .B(mult_ab_1_2[3]), .Z(n7) );
  XOR2_X1 U141 ( .A(mult_ab_1_0[4]), .B(n6), .Z(port_c_1[4]) );
  XOR2_X1 U142 ( .A(temp_0_1[4]), .B(mult_ab_1_2[4]), .Z(n6) );
  XOR2_X1 U143 ( .A(mult_ab_0_1[0]), .B(n15), .Z(port_c_0[0]) );
  XOR2_X1 U144 ( .A(temp_0_0[0]), .B(mult_ab_0_2[0]), .Z(n15) );
  XOR2_X1 U145 ( .A(mult_ab_0_1[1]), .B(n14), .Z(port_c_0[1]) );
  XOR2_X1 U146 ( .A(temp_0_0[1]), .B(mult_ab_0_2[1]), .Z(n14) );
  XOR2_X1 U147 ( .A(mult_ab_0_1[2]), .B(n13), .Z(port_c_0[2]) );
  XOR2_X1 U148 ( .A(temp_0_0[2]), .B(mult_ab_0_2[2]), .Z(n13) );
  XOR2_X1 U149 ( .A(mult_ab_0_1[3]), .B(n12), .Z(port_c_0[3]) );
  XOR2_X1 U150 ( .A(temp_0_0[3]), .B(mult_ab_0_2[3]), .Z(n12) );
  XOR2_X1 U151 ( .A(mult_ab_0_1[4]), .B(n11), .Z(port_c_0[4]) );
  XOR2_X1 U152 ( .A(temp_0_0[4]), .B(mult_ab_0_2[4]), .Z(n11) );
  BUF_X1 ref_1_U32 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n30) );
  BUF_X1 ref_1_U31 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n29) );
  BUF_X1 ref_1_U30 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n28) );
  BUF_X1 ref_1_U29 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n27) );
  BUF_X1 ref_1_U28 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n26) );
  BUF_X1 ref_1_U27 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n25) );
  BUF_X1 ref_1_U26 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n24) );
  BUF_X1 ref_1_U25 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n23) );
  BUF_X1 ref_1_U24 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n22) );
  BUF_X1 ref_1_U23 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n21) );
  BUF_X1 ref_1_U22 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n20) );
  BUF_X1 ref_1_U21 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n19) );
  BUF_X1 ref_1_U20 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n18) );
  BUF_X1 ref_1_U19 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n17) );
  BUF_X1 ref_1_U18 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n16) );
  BUF_X1 ref_1_U17 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n15) );
  BUF_X1 ref_1_U16 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n14) );
  BUF_X1 ref_1_U15 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n13) );
  BUF_X1 ref_1_U14 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n12) );
  BUF_X1 ref_1_U13 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n11) );
  BUF_X1 ref_1_U12 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n10) );
  BUF_X1 ref_1_U11 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n9) );
  BUF_X1 ref_1_U10 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n8) );
  BUF_X1 ref_1_U9 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n7) );
  BUF_X1 ref_1_U8 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n6) );
  BUF_X1 ref_1_U7 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n5) );
  BUF_X1 ref_1_U6 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n4) );
  BUF_X1 ref_1_U5 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n3) );
  BUF_X1 ref_1_U4 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n2) );
  BUF_X1 ref_1_U3 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n1) );
  DFF_X1 ref_1_reg_out_2_2_reg_0_ ( .D(ref_1_maj_53_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_1_ ( .D(ref_1_maj_62_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_2_ ( .D(ref_1_maj_71_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_3_ ( .D(ref_1_maj_80_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_4_ ( .D(ref_1_maj_89_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_0_ ( .D(ref_1_maj_52_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_1_ ( .D(ref_1_maj_61_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_2_ ( .D(ref_1_maj_70_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_3_ ( .D(ref_1_maj_79_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_4_ ( .D(ref_1_maj_88_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_0_ ( .D(ref_1_maj_51_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_1_ ( .D(ref_1_maj_60_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_2_ ( .D(ref_1_maj_69_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_3_ ( .D(ref_1_maj_78_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_4_ ( .D(ref_1_maj_87_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_0_ ( .D(ref_1_maj_50_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_1_ ( .D(ref_1_maj_59_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_2_ ( .D(ref_1_maj_68_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_3_ ( .D(ref_1_maj_77_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_4_ ( .D(ref_1_maj_86_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_0_ ( .D(ref_1_maj_49_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_1_ ( .D(ref_1_maj_58_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_2_ ( .D(ref_1_maj_67_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_3_ ( .D(ref_1_maj_76_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_4_ ( .D(ref_1_maj_85_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_0_ ( .D(ref_1_maj_48_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_1_ ( .D(ref_1_maj_57_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_2_ ( .D(ref_1_maj_66_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_3_ ( .D(ref_1_maj_75_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_4_ ( .D(ref_1_maj_84_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_0_ ( .D(ref_1_maj_47_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_1_ ( .D(ref_1_maj_56_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_2_ ( .D(ref_1_maj_65_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_3_ ( .D(ref_1_maj_74_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_4_ ( .D(ref_1_maj_83_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_0_ ( .D(ref_1_maj_46_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_1_ ( .D(ref_1_maj_55_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_2_ ( .D(ref_1_maj_64_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_3_ ( .D(ref_1_maj_73_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_4_ ( .D(ref_1_maj_82_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_0_ ( .D(ref_1_maj_45_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_1_ ( .D(ref_1_maj_54_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_2_ ( .D(ref_1_maj_63_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_3_ ( .D(ref_1_maj_72_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_4_ ( .D(ref_1_maj_81_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[4]), .QN() );
  XOR2_X1 ref_1_simpleXor_120_U1 ( .A(port_rand_ref[0]), .B(port_b_0[0]), .Z(
        ref_1_simpleXor_120_port_z) );
  XOR2_X1 ref_1_simpleXor_121_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_120_port_z), .Z(ref_1_simpleXor_121_port_z) );
  XOR2_X1 ref_1_simpleXor_122_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_121_port_z), .Z(ref_1_simpleXor_122_port_z) );
  XOR2_X1 ref_1_simpleXor_123_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_122_port_z), .Z(ref_1_refreshed_0_0_) );
  XOR2_X1 ref_1_simpleXor_124_U1 ( .A(port_rand_ref[0]), .B(port_b_1[0]), .Z(
        ref_1_simpleXor_124_port_z) );
  XOR2_X1 ref_1_simpleXor_125_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_124_port_z), .Z(ref_1_simpleXor_125_port_z) );
  XOR2_X1 ref_1_simpleXor_126_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_125_port_z), .Z(ref_1_simpleXor_126_port_z) );
  XOR2_X1 ref_1_simpleXor_127_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_126_port_z), .Z(ref_1_refreshed_1_0_) );
  XOR2_X1 ref_1_simpleXor_128_U1 ( .A(port_rand_ref[2]), .B(port_b_2[0]), .Z(
        ref_1_simpleXor_128_port_z) );
  XOR2_X1 ref_1_simpleXor_129_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_128_port_z), .Z(ref_1_simpleXor_129_port_z) );
  XOR2_X1 ref_1_simpleXor_130_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_129_port_z), .Z(ref_1_simpleXor_130_port_z) );
  XOR2_X1 ref_1_simpleXor_131_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_130_port_z), .Z(ref_1_refreshed_2_0_) );
  XOR2_X1 ref_1_simpleXor_132_U1 ( .A(port_rand_ref[0]), .B(port_b_0[1]), .Z(
        ref_1_simpleXor_132_port_z) );
  XOR2_X1 ref_1_simpleXor_133_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_132_port_z), .Z(ref_1_simpleXor_133_port_z) );
  XOR2_X1 ref_1_simpleXor_134_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_133_port_z), .Z(ref_1_simpleXor_134_port_z) );
  XOR2_X1 ref_1_simpleXor_135_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_134_port_z), .Z(ref_1_refreshed_0_1_) );
  XOR2_X1 ref_1_simpleXor_136_U1 ( .A(port_rand_ref[0]), .B(port_b_1[1]), .Z(
        ref_1_simpleXor_136_port_z) );
  XOR2_X1 ref_1_simpleXor_137_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_136_port_z), .Z(ref_1_simpleXor_137_port_z) );
  XOR2_X1 ref_1_simpleXor_138_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_137_port_z), .Z(ref_1_simpleXor_138_port_z) );
  XOR2_X1 ref_1_simpleXor_139_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_138_port_z), .Z(ref_1_refreshed_1_1_) );
  XOR2_X1 ref_1_simpleXor_140_U1 ( .A(port_rand_ref[2]), .B(port_b_2[1]), .Z(
        ref_1_simpleXor_140_port_z) );
  XOR2_X1 ref_1_simpleXor_141_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_140_port_z), .Z(ref_1_simpleXor_141_port_z) );
  XOR2_X1 ref_1_simpleXor_142_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_141_port_z), .Z(ref_1_simpleXor_142_port_z) );
  XOR2_X1 ref_1_simpleXor_143_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_142_port_z), .Z(ref_1_refreshed_2_1_) );
  XOR2_X1 ref_1_simpleXor_144_U1 ( .A(port_rand_ref[0]), .B(port_b_0[2]), .Z(
        ref_1_simpleXor_144_port_z) );
  XOR2_X1 ref_1_simpleXor_145_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_144_port_z), .Z(ref_1_simpleXor_145_port_z) );
  XOR2_X1 ref_1_simpleXor_146_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_145_port_z), .Z(ref_1_simpleXor_146_port_z) );
  XOR2_X1 ref_1_simpleXor_147_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_146_port_z), .Z(ref_1_refreshed_0_2_) );
  XOR2_X1 ref_1_simpleXor_148_U1 ( .A(port_rand_ref[0]), .B(port_b_1[2]), .Z(
        ref_1_simpleXor_148_port_z) );
  XOR2_X1 ref_1_simpleXor_149_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_148_port_z), .Z(ref_1_simpleXor_149_port_z) );
  XOR2_X1 ref_1_simpleXor_150_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_149_port_z), .Z(ref_1_simpleXor_150_port_z) );
  XOR2_X1 ref_1_simpleXor_151_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_150_port_z), .Z(ref_1_refreshed_1_2_) );
  XOR2_X1 ref_1_simpleXor_152_U1 ( .A(port_rand_ref[2]), .B(port_b_2[2]), .Z(
        ref_1_simpleXor_152_port_z) );
  XOR2_X1 ref_1_simpleXor_153_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_152_port_z), .Z(ref_1_simpleXor_153_port_z) );
  XOR2_X1 ref_1_simpleXor_154_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_153_port_z), .Z(ref_1_simpleXor_154_port_z) );
  XOR2_X1 ref_1_simpleXor_155_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_154_port_z), .Z(ref_1_refreshed_2_2_) );
  XOR2_X1 ref_1_simpleXor_156_U1 ( .A(port_rand_ref[0]), .B(port_b_0[3]), .Z(
        ref_1_simpleXor_156_port_z) );
  XOR2_X1 ref_1_simpleXor_157_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_156_port_z), .Z(ref_1_simpleXor_157_port_z) );
  XOR2_X1 ref_1_simpleXor_158_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_157_port_z), .Z(ref_1_simpleXor_158_port_z) );
  XOR2_X1 ref_1_simpleXor_159_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_158_port_z), .Z(ref_1_refreshed_0_3_) );
  XOR2_X1 ref_1_simpleXor_160_U1 ( .A(port_rand_ref[0]), .B(port_b_1[3]), .Z(
        ref_1_simpleXor_160_port_z) );
  XOR2_X1 ref_1_simpleXor_161_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_160_port_z), .Z(ref_1_simpleXor_161_port_z) );
  XOR2_X1 ref_1_simpleXor_162_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_161_port_z), .Z(ref_1_simpleXor_162_port_z) );
  XOR2_X1 ref_1_simpleXor_163_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_162_port_z), .Z(ref_1_refreshed_1_3_) );
  XOR2_X1 ref_1_simpleXor_164_U1 ( .A(port_rand_ref[2]), .B(port_b_2[3]), .Z(
        ref_1_simpleXor_164_port_z) );
  XOR2_X1 ref_1_simpleXor_165_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_164_port_z), .Z(ref_1_simpleXor_165_port_z) );
  XOR2_X1 ref_1_simpleXor_166_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_165_port_z), .Z(ref_1_simpleXor_166_port_z) );
  XOR2_X1 ref_1_simpleXor_167_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_166_port_z), .Z(ref_1_refreshed_2_3_) );
  XOR2_X1 ref_1_simpleXor_168_U1 ( .A(port_rand_ref[0]), .B(port_b_0[4]), .Z(
        ref_1_simpleXor_168_port_z) );
  XOR2_X1 ref_1_simpleXor_169_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_168_port_z), .Z(ref_1_simpleXor_169_port_z) );
  XOR2_X1 ref_1_simpleXor_170_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_169_port_z), .Z(ref_1_simpleXor_170_port_z) );
  XOR2_X1 ref_1_simpleXor_171_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_170_port_z), .Z(ref_1_refreshed_0_4_) );
  XOR2_X1 ref_1_simpleXor_172_U1 ( .A(port_rand_ref[0]), .B(port_b_1[4]), .Z(
        ref_1_simpleXor_172_port_z) );
  XOR2_X1 ref_1_simpleXor_173_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_172_port_z), .Z(ref_1_simpleXor_173_port_z) );
  XOR2_X1 ref_1_simpleXor_174_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_173_port_z), .Z(ref_1_simpleXor_174_port_z) );
  XOR2_X1 ref_1_simpleXor_175_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_174_port_z), .Z(ref_1_refreshed_1_4_) );
  XOR2_X1 ref_1_simpleXor_176_U1 ( .A(port_rand_ref[2]), .B(port_b_2[4]), .Z(
        ref_1_simpleXor_176_port_z) );
  XOR2_X1 ref_1_simpleXor_177_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_176_port_z), .Z(ref_1_simpleXor_177_port_z) );
  XOR2_X1 ref_1_simpleXor_178_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_177_port_z), .Z(ref_1_simpleXor_178_port_z) );
  XOR2_X1 ref_1_simpleXor_179_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_178_port_z), .Z(ref_1_refreshed_2_4_) );
  NAND2_X1 ref_1_maj_45_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_45_n9) );
  NAND2_X1 ref_1_maj_45_U14 ( .A1(ref_1_maj_45_n6), .A2(ref_1_maj_45_n5), .ZN(
        ref_1_maj_45_n10) );
  NAND2_X1 ref_1_maj_45_U13 ( .A1(ref_1_maj_45_n9), .A2(ref_1_maj_45_n10), 
        .ZN(ref_1_maj_45_n8) );
  NAND2_X1 ref_1_maj_45_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_45_n11), .ZN(
        ref_1_maj_45_n13) );
  NAND2_X1 ref_1_maj_45_U11 ( .A1(ref_1_n22), .A2(ref_1_n23), .ZN(
        ref_1_maj_45_n12) );
  NAND2_X1 ref_1_maj_45_U10 ( .A1(ref_1_maj_45_n12), .A2(ref_1_maj_45_n13), 
        .ZN(ref_1_maj_45_n7) );
  XOR2_X1 ref_1_maj_45_U9 ( .A(ref_1_n26), .B(ref_1_maj_45_n11), .Z(
        ref_1_maj_45_n6) );
  XOR2_X1 ref_1_maj_45_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_45_n5)
         );
  XOR2_X1 ref_1_maj_45_U7 ( .A(ref_1_n22), .B(ref_1_n23), .Z(ref_1_maj_45_n11)
         );
  OR2_X1 ref_1_maj_45_U6 ( .A1(ref_1_maj_45_n7), .A2(ref_1_maj_45_n8), .ZN(
        ref_1_maj_45_n3) );
  NAND2_X1 ref_1_maj_45_U5 ( .A1(ref_1_maj_45_n3), .A2(ref_1_maj_45_n4), .ZN(
        ref_1_maj_45_n2) );
  NAND2_X1 ref_1_maj_45_U4 ( .A1(ref_1_maj_45_n7), .A2(ref_1_maj_45_n8), .ZN(
        ref_1_maj_45_n1) );
  NAND2_X1 ref_1_maj_45_U3 ( .A1(ref_1_maj_45_n1), .A2(ref_1_maj_45_n2), .ZN(
        ref_1_maj_45_port_o) );
  XOR2_X1 ref_1_maj_45_U2 ( .A(ref_1_maj_45_n5), .B(ref_1_maj_45_n6), .Z(
        ref_1_maj_45_n4) );
  NAND2_X1 ref_1_maj_46_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_46_n18) );
  NAND2_X1 ref_1_maj_46_U14 ( .A1(ref_1_maj_46_n21), .A2(ref_1_maj_46_n22), 
        .ZN(ref_1_maj_46_n17) );
  NAND2_X1 ref_1_maj_46_U13 ( .A1(ref_1_maj_46_n18), .A2(ref_1_maj_46_n17), 
        .ZN(ref_1_maj_46_n19) );
  NAND2_X1 ref_1_maj_46_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_46_n16), .ZN(
        ref_1_maj_46_n14) );
  NAND2_X1 ref_1_maj_46_U11 ( .A1(ref_1_n22), .A2(ref_1_n23), .ZN(
        ref_1_maj_46_n15) );
  NAND2_X1 ref_1_maj_46_U10 ( .A1(ref_1_maj_46_n15), .A2(ref_1_maj_46_n14), 
        .ZN(ref_1_maj_46_n20) );
  XOR2_X1 ref_1_maj_46_U9 ( .A(ref_1_n26), .B(ref_1_maj_46_n16), .Z(
        ref_1_maj_46_n21) );
  XOR2_X1 ref_1_maj_46_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_46_n22)
         );
  XOR2_X1 ref_1_maj_46_U7 ( .A(ref_1_n22), .B(ref_1_n23), .Z(ref_1_maj_46_n16)
         );
  OR2_X1 ref_1_maj_46_U6 ( .A1(ref_1_maj_46_n20), .A2(ref_1_maj_46_n19), .ZN(
        ref_1_maj_46_n24) );
  NAND2_X1 ref_1_maj_46_U5 ( .A1(ref_1_maj_46_n24), .A2(ref_1_maj_46_n23), 
        .ZN(ref_1_maj_46_n25) );
  NAND2_X1 ref_1_maj_46_U4 ( .A1(ref_1_maj_46_n20), .A2(ref_1_maj_46_n19), 
        .ZN(ref_1_maj_46_n26) );
  NAND2_X1 ref_1_maj_46_U3 ( .A1(ref_1_maj_46_n26), .A2(ref_1_maj_46_n25), 
        .ZN(ref_1_maj_46_port_o) );
  XOR2_X1 ref_1_maj_46_U2 ( .A(ref_1_maj_46_n22), .B(ref_1_maj_46_n21), .Z(
        ref_1_maj_46_n23) );
  NAND2_X1 ref_1_maj_47_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_47_n18) );
  NAND2_X1 ref_1_maj_47_U14 ( .A1(ref_1_maj_47_n21), .A2(ref_1_maj_47_n22), 
        .ZN(ref_1_maj_47_n17) );
  NAND2_X1 ref_1_maj_47_U13 ( .A1(ref_1_maj_47_n18), .A2(ref_1_maj_47_n17), 
        .ZN(ref_1_maj_47_n19) );
  NAND2_X1 ref_1_maj_47_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_47_n16), 
        .ZN(ref_1_maj_47_n14) );
  NAND2_X1 ref_1_maj_47_U11 ( .A1(ref_1_refreshed_0_0_), .A2(ref_1_n23), .ZN(
        ref_1_maj_47_n15) );
  NAND2_X1 ref_1_maj_47_U10 ( .A1(ref_1_maj_47_n15), .A2(ref_1_maj_47_n14), 
        .ZN(ref_1_maj_47_n20) );
  XOR2_X1 ref_1_maj_47_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_47_n16), 
        .Z(ref_1_maj_47_n21) );
  XOR2_X1 ref_1_maj_47_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_47_n22) );
  XOR2_X1 ref_1_maj_47_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_n23), .Z(
        ref_1_maj_47_n16) );
  OR2_X1 ref_1_maj_47_U6 ( .A1(ref_1_maj_47_n20), .A2(ref_1_maj_47_n19), .ZN(
        ref_1_maj_47_n24) );
  NAND2_X1 ref_1_maj_47_U5 ( .A1(ref_1_maj_47_n24), .A2(ref_1_maj_47_n23), 
        .ZN(ref_1_maj_47_n25) );
  NAND2_X1 ref_1_maj_47_U4 ( .A1(ref_1_maj_47_n20), .A2(ref_1_maj_47_n19), 
        .ZN(ref_1_maj_47_n26) );
  NAND2_X1 ref_1_maj_47_U3 ( .A1(ref_1_maj_47_n26), .A2(ref_1_maj_47_n25), 
        .ZN(ref_1_maj_47_port_o) );
  XOR2_X1 ref_1_maj_47_U2 ( .A(ref_1_maj_47_n22), .B(ref_1_maj_47_n21), .Z(
        ref_1_maj_47_n23) );
  NAND2_X1 ref_1_maj_48_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_48_n18) );
  NAND2_X1 ref_1_maj_48_U14 ( .A1(ref_1_maj_48_n21), .A2(ref_1_maj_48_n22), 
        .ZN(ref_1_maj_48_n17) );
  NAND2_X1 ref_1_maj_48_U13 ( .A1(ref_1_maj_48_n18), .A2(ref_1_maj_48_n17), 
        .ZN(ref_1_maj_48_n19) );
  NAND2_X1 ref_1_maj_48_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_48_n16), .ZN(
        ref_1_maj_48_n14) );
  NAND2_X1 ref_1_maj_48_U11 ( .A1(ref_1_n12), .A2(ref_1_n13), .ZN(
        ref_1_maj_48_n15) );
  NAND2_X1 ref_1_maj_48_U10 ( .A1(ref_1_maj_48_n15), .A2(ref_1_maj_48_n14), 
        .ZN(ref_1_maj_48_n20) );
  XOR2_X1 ref_1_maj_48_U9 ( .A(ref_1_n16), .B(ref_1_maj_48_n16), .Z(
        ref_1_maj_48_n21) );
  XOR2_X1 ref_1_maj_48_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_48_n22)
         );
  XOR2_X1 ref_1_maj_48_U7 ( .A(ref_1_n12), .B(ref_1_n13), .Z(ref_1_maj_48_n16)
         );
  OR2_X1 ref_1_maj_48_U6 ( .A1(ref_1_maj_48_n20), .A2(ref_1_maj_48_n19), .ZN(
        ref_1_maj_48_n24) );
  NAND2_X1 ref_1_maj_48_U5 ( .A1(ref_1_maj_48_n24), .A2(ref_1_maj_48_n23), 
        .ZN(ref_1_maj_48_n25) );
  NAND2_X1 ref_1_maj_48_U4 ( .A1(ref_1_maj_48_n20), .A2(ref_1_maj_48_n19), 
        .ZN(ref_1_maj_48_n26) );
  NAND2_X1 ref_1_maj_48_U3 ( .A1(ref_1_maj_48_n26), .A2(ref_1_maj_48_n25), 
        .ZN(ref_1_maj_48_port_o) );
  XOR2_X1 ref_1_maj_48_U2 ( .A(ref_1_maj_48_n22), .B(ref_1_maj_48_n21), .Z(
        ref_1_maj_48_n23) );
  NAND2_X1 ref_1_maj_49_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_49_n18) );
  NAND2_X1 ref_1_maj_49_U14 ( .A1(ref_1_maj_49_n21), .A2(ref_1_maj_49_n22), 
        .ZN(ref_1_maj_49_n17) );
  NAND2_X1 ref_1_maj_49_U13 ( .A1(ref_1_maj_49_n18), .A2(ref_1_maj_49_n17), 
        .ZN(ref_1_maj_49_n19) );
  NAND2_X1 ref_1_maj_49_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_49_n16), 
        .ZN(ref_1_maj_49_n14) );
  NAND2_X1 ref_1_maj_49_U11 ( .A1(ref_1_refreshed_1_0_), .A2(ref_1_n13), .ZN(
        ref_1_maj_49_n15) );
  NAND2_X1 ref_1_maj_49_U10 ( .A1(ref_1_maj_49_n15), .A2(ref_1_maj_49_n14), 
        .ZN(ref_1_maj_49_n20) );
  XOR2_X1 ref_1_maj_49_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_49_n16), 
        .Z(ref_1_maj_49_n21) );
  XOR2_X1 ref_1_maj_49_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_49_n22) );
  XOR2_X1 ref_1_maj_49_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_n13), .Z(
        ref_1_maj_49_n16) );
  OR2_X1 ref_1_maj_49_U6 ( .A1(ref_1_maj_49_n20), .A2(ref_1_maj_49_n19), .ZN(
        ref_1_maj_49_n24) );
  NAND2_X1 ref_1_maj_49_U5 ( .A1(ref_1_maj_49_n24), .A2(ref_1_maj_49_n23), 
        .ZN(ref_1_maj_49_n25) );
  NAND2_X1 ref_1_maj_49_U4 ( .A1(ref_1_maj_49_n20), .A2(ref_1_maj_49_n19), 
        .ZN(ref_1_maj_49_n26) );
  NAND2_X1 ref_1_maj_49_U3 ( .A1(ref_1_maj_49_n26), .A2(ref_1_maj_49_n25), 
        .ZN(ref_1_maj_49_port_o) );
  XOR2_X1 ref_1_maj_49_U2 ( .A(ref_1_maj_49_n22), .B(ref_1_maj_49_n21), .Z(
        ref_1_maj_49_n23) );
  NAND2_X1 ref_1_maj_50_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_50_n18) );
  NAND2_X1 ref_1_maj_50_U14 ( .A1(ref_1_maj_50_n21), .A2(ref_1_maj_50_n22), 
        .ZN(ref_1_maj_50_n17) );
  NAND2_X1 ref_1_maj_50_U13 ( .A1(ref_1_maj_50_n18), .A2(ref_1_maj_50_n17), 
        .ZN(ref_1_maj_50_n19) );
  NAND2_X1 ref_1_maj_50_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_50_n16), 
        .ZN(ref_1_maj_50_n14) );
  NAND2_X1 ref_1_maj_50_U11 ( .A1(ref_1_refreshed_1_0_), .A2(ref_1_n13), .ZN(
        ref_1_maj_50_n15) );
  NAND2_X1 ref_1_maj_50_U10 ( .A1(ref_1_maj_50_n15), .A2(ref_1_maj_50_n14), 
        .ZN(ref_1_maj_50_n20) );
  XOR2_X1 ref_1_maj_50_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_50_n16), 
        .Z(ref_1_maj_50_n21) );
  XOR2_X1 ref_1_maj_50_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_50_n22) );
  XOR2_X1 ref_1_maj_50_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_n13), .Z(
        ref_1_maj_50_n16) );
  OR2_X1 ref_1_maj_50_U6 ( .A1(ref_1_maj_50_n20), .A2(ref_1_maj_50_n19), .ZN(
        ref_1_maj_50_n24) );
  NAND2_X1 ref_1_maj_50_U5 ( .A1(ref_1_maj_50_n24), .A2(ref_1_maj_50_n23), 
        .ZN(ref_1_maj_50_n25) );
  NAND2_X1 ref_1_maj_50_U4 ( .A1(ref_1_maj_50_n20), .A2(ref_1_maj_50_n19), 
        .ZN(ref_1_maj_50_n26) );
  NAND2_X1 ref_1_maj_50_U3 ( .A1(ref_1_maj_50_n26), .A2(ref_1_maj_50_n25), 
        .ZN(ref_1_maj_50_port_o) );
  XOR2_X1 ref_1_maj_50_U2 ( .A(ref_1_maj_50_n22), .B(ref_1_maj_50_n21), .Z(
        ref_1_maj_50_n23) );
  NAND2_X1 ref_1_maj_51_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_51_n18) );
  NAND2_X1 ref_1_maj_51_U14 ( .A1(ref_1_maj_51_n21), .A2(ref_1_maj_51_n22), 
        .ZN(ref_1_maj_51_n17) );
  NAND2_X1 ref_1_maj_51_U13 ( .A1(ref_1_maj_51_n18), .A2(ref_1_maj_51_n17), 
        .ZN(ref_1_maj_51_n19) );
  NAND2_X1 ref_1_maj_51_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_51_n16), .ZN(
        ref_1_maj_51_n14) );
  NAND2_X1 ref_1_maj_51_U11 ( .A1(ref_1_n2), .A2(ref_1_n3), .ZN(
        ref_1_maj_51_n15) );
  NAND2_X1 ref_1_maj_51_U10 ( .A1(ref_1_maj_51_n15), .A2(ref_1_maj_51_n14), 
        .ZN(ref_1_maj_51_n20) );
  XOR2_X1 ref_1_maj_51_U9 ( .A(ref_1_n6), .B(ref_1_maj_51_n16), .Z(
        ref_1_maj_51_n21) );
  XOR2_X1 ref_1_maj_51_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_51_n22)
         );
  XOR2_X1 ref_1_maj_51_U7 ( .A(ref_1_n2), .B(ref_1_n3), .Z(ref_1_maj_51_n16)
         );
  OR2_X1 ref_1_maj_51_U6 ( .A1(ref_1_maj_51_n20), .A2(ref_1_maj_51_n19), .ZN(
        ref_1_maj_51_n24) );
  NAND2_X1 ref_1_maj_51_U5 ( .A1(ref_1_maj_51_n24), .A2(ref_1_maj_51_n23), 
        .ZN(ref_1_maj_51_n25) );
  NAND2_X1 ref_1_maj_51_U4 ( .A1(ref_1_maj_51_n20), .A2(ref_1_maj_51_n19), 
        .ZN(ref_1_maj_51_n26) );
  NAND2_X1 ref_1_maj_51_U3 ( .A1(ref_1_maj_51_n26), .A2(ref_1_maj_51_n25), 
        .ZN(ref_1_maj_51_port_o) );
  XOR2_X1 ref_1_maj_51_U2 ( .A(ref_1_maj_51_n22), .B(ref_1_maj_51_n21), .Z(
        ref_1_maj_51_n23) );
  NAND2_X1 ref_1_maj_52_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_52_n18) );
  NAND2_X1 ref_1_maj_52_U14 ( .A1(ref_1_maj_52_n21), .A2(ref_1_maj_52_n22), 
        .ZN(ref_1_maj_52_n17) );
  NAND2_X1 ref_1_maj_52_U13 ( .A1(ref_1_maj_52_n18), .A2(ref_1_maj_52_n17), 
        .ZN(ref_1_maj_52_n19) );
  NAND2_X1 ref_1_maj_52_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_52_n16), 
        .ZN(ref_1_maj_52_n14) );
  NAND2_X1 ref_1_maj_52_U11 ( .A1(ref_1_refreshed_2_0_), .A2(ref_1_n3), .ZN(
        ref_1_maj_52_n15) );
  NAND2_X1 ref_1_maj_52_U10 ( .A1(ref_1_maj_52_n15), .A2(ref_1_maj_52_n14), 
        .ZN(ref_1_maj_52_n20) );
  XOR2_X1 ref_1_maj_52_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_52_n16), 
        .Z(ref_1_maj_52_n21) );
  XOR2_X1 ref_1_maj_52_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_52_n22) );
  XOR2_X1 ref_1_maj_52_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_n3), .Z(
        ref_1_maj_52_n16) );
  OR2_X1 ref_1_maj_52_U6 ( .A1(ref_1_maj_52_n20), .A2(ref_1_maj_52_n19), .ZN(
        ref_1_maj_52_n24) );
  NAND2_X1 ref_1_maj_52_U5 ( .A1(ref_1_maj_52_n24), .A2(ref_1_maj_52_n23), 
        .ZN(ref_1_maj_52_n25) );
  NAND2_X1 ref_1_maj_52_U4 ( .A1(ref_1_maj_52_n20), .A2(ref_1_maj_52_n19), 
        .ZN(ref_1_maj_52_n26) );
  NAND2_X1 ref_1_maj_52_U3 ( .A1(ref_1_maj_52_n26), .A2(ref_1_maj_52_n25), 
        .ZN(ref_1_maj_52_port_o) );
  XOR2_X1 ref_1_maj_52_U2 ( .A(ref_1_maj_52_n22), .B(ref_1_maj_52_n21), .Z(
        ref_1_maj_52_n23) );
  NAND2_X1 ref_1_maj_53_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_53_n18) );
  NAND2_X1 ref_1_maj_53_U14 ( .A1(ref_1_maj_53_n21), .A2(ref_1_maj_53_n22), 
        .ZN(ref_1_maj_53_n17) );
  NAND2_X1 ref_1_maj_53_U13 ( .A1(ref_1_maj_53_n18), .A2(ref_1_maj_53_n17), 
        .ZN(ref_1_maj_53_n19) );
  NAND2_X1 ref_1_maj_53_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_53_n16), 
        .ZN(ref_1_maj_53_n14) );
  NAND2_X1 ref_1_maj_53_U11 ( .A1(ref_1_refreshed_2_0_), .A2(ref_1_n3), .ZN(
        ref_1_maj_53_n15) );
  NAND2_X1 ref_1_maj_53_U10 ( .A1(ref_1_maj_53_n15), .A2(ref_1_maj_53_n14), 
        .ZN(ref_1_maj_53_n20) );
  XOR2_X1 ref_1_maj_53_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_53_n16), 
        .Z(ref_1_maj_53_n21) );
  XOR2_X1 ref_1_maj_53_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_53_n22) );
  XOR2_X1 ref_1_maj_53_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_n3), .Z(
        ref_1_maj_53_n16) );
  OR2_X1 ref_1_maj_53_U6 ( .A1(ref_1_maj_53_n20), .A2(ref_1_maj_53_n19), .ZN(
        ref_1_maj_53_n24) );
  NAND2_X1 ref_1_maj_53_U5 ( .A1(ref_1_maj_53_n24), .A2(ref_1_maj_53_n23), 
        .ZN(ref_1_maj_53_n25) );
  NAND2_X1 ref_1_maj_53_U4 ( .A1(ref_1_maj_53_n20), .A2(ref_1_maj_53_n19), 
        .ZN(ref_1_maj_53_n26) );
  NAND2_X1 ref_1_maj_53_U3 ( .A1(ref_1_maj_53_n26), .A2(ref_1_maj_53_n25), 
        .ZN(ref_1_maj_53_port_o) );
  XOR2_X1 ref_1_maj_53_U2 ( .A(ref_1_maj_53_n22), .B(ref_1_maj_53_n21), .Z(
        ref_1_maj_53_n23) );
  NAND2_X1 ref_1_maj_54_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_54_n18) );
  NAND2_X1 ref_1_maj_54_U14 ( .A1(ref_1_maj_54_n21), .A2(ref_1_maj_54_n22), 
        .ZN(ref_1_maj_54_n17) );
  NAND2_X1 ref_1_maj_54_U13 ( .A1(ref_1_maj_54_n18), .A2(ref_1_maj_54_n17), 
        .ZN(ref_1_maj_54_n19) );
  NAND2_X1 ref_1_maj_54_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_54_n16), 
        .ZN(ref_1_maj_54_n14) );
  NAND2_X1 ref_1_maj_54_U11 ( .A1(ref_1_refreshed_0_0_), .A2(ref_1_n23), .ZN(
        ref_1_maj_54_n15) );
  NAND2_X1 ref_1_maj_54_U10 ( .A1(ref_1_maj_54_n15), .A2(ref_1_maj_54_n14), 
        .ZN(ref_1_maj_54_n20) );
  XOR2_X1 ref_1_maj_54_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_54_n16), 
        .Z(ref_1_maj_54_n21) );
  XOR2_X1 ref_1_maj_54_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_54_n22) );
  XOR2_X1 ref_1_maj_54_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_n23), .Z(
        ref_1_maj_54_n16) );
  OR2_X1 ref_1_maj_54_U6 ( .A1(ref_1_maj_54_n20), .A2(ref_1_maj_54_n19), .ZN(
        ref_1_maj_54_n24) );
  NAND2_X1 ref_1_maj_54_U5 ( .A1(ref_1_maj_54_n24), .A2(ref_1_maj_54_n23), 
        .ZN(ref_1_maj_54_n25) );
  NAND2_X1 ref_1_maj_54_U4 ( .A1(ref_1_maj_54_n20), .A2(ref_1_maj_54_n19), 
        .ZN(ref_1_maj_54_n26) );
  NAND2_X1 ref_1_maj_54_U3 ( .A1(ref_1_maj_54_n26), .A2(ref_1_maj_54_n25), 
        .ZN(ref_1_maj_54_port_o) );
  XOR2_X1 ref_1_maj_54_U2 ( .A(ref_1_maj_54_n22), .B(ref_1_maj_54_n21), .Z(
        ref_1_maj_54_n23) );
  NAND2_X1 ref_1_maj_55_U15 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_55_n18) );
  NAND2_X1 ref_1_maj_55_U14 ( .A1(ref_1_maj_55_n21), .A2(ref_1_maj_55_n22), 
        .ZN(ref_1_maj_55_n17) );
  NAND2_X1 ref_1_maj_55_U13 ( .A1(ref_1_maj_55_n18), .A2(ref_1_maj_55_n17), 
        .ZN(ref_1_maj_55_n19) );
  NAND2_X1 ref_1_maj_55_U12 ( .A1(ref_1_refreshed_0_2_), .A2(ref_1_maj_55_n16), 
        .ZN(ref_1_maj_55_n14) );
  NAND2_X1 ref_1_maj_55_U11 ( .A1(ref_1_refreshed_0_0_), .A2(ref_1_n23), .ZN(
        ref_1_maj_55_n15) );
  NAND2_X1 ref_1_maj_55_U10 ( .A1(ref_1_maj_55_n15), .A2(ref_1_maj_55_n14), 
        .ZN(ref_1_maj_55_n20) );
  XOR2_X1 ref_1_maj_55_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_55_n16), 
        .Z(ref_1_maj_55_n21) );
  XOR2_X1 ref_1_maj_55_U8 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), 
        .Z(ref_1_maj_55_n22) );
  XOR2_X1 ref_1_maj_55_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_n23), .Z(
        ref_1_maj_55_n16) );
  OR2_X1 ref_1_maj_55_U6 ( .A1(ref_1_maj_55_n20), .A2(ref_1_maj_55_n19), .ZN(
        ref_1_maj_55_n24) );
  NAND2_X1 ref_1_maj_55_U5 ( .A1(ref_1_maj_55_n24), .A2(ref_1_maj_55_n23), 
        .ZN(ref_1_maj_55_n25) );
  NAND2_X1 ref_1_maj_55_U4 ( .A1(ref_1_maj_55_n20), .A2(ref_1_maj_55_n19), 
        .ZN(ref_1_maj_55_n26) );
  NAND2_X1 ref_1_maj_55_U3 ( .A1(ref_1_maj_55_n26), .A2(ref_1_maj_55_n25), 
        .ZN(ref_1_maj_55_port_o) );
  XOR2_X1 ref_1_maj_55_U2 ( .A(ref_1_maj_55_n22), .B(ref_1_maj_55_n21), .Z(
        ref_1_maj_55_n23) );
  NAND2_X1 ref_1_maj_56_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_56_n18) );
  NAND2_X1 ref_1_maj_56_U14 ( .A1(ref_1_maj_56_n21), .A2(ref_1_maj_56_n22), 
        .ZN(ref_1_maj_56_n17) );
  NAND2_X1 ref_1_maj_56_U13 ( .A1(ref_1_maj_56_n18), .A2(ref_1_maj_56_n17), 
        .ZN(ref_1_maj_56_n19) );
  NAND2_X1 ref_1_maj_56_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_56_n16), .ZN(
        ref_1_maj_56_n14) );
  NAND2_X1 ref_1_maj_56_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_56_n15) );
  NAND2_X1 ref_1_maj_56_U10 ( .A1(ref_1_maj_56_n15), .A2(ref_1_maj_56_n14), 
        .ZN(ref_1_maj_56_n20) );
  XOR2_X1 ref_1_maj_56_U9 ( .A(ref_1_n25), .B(ref_1_maj_56_n16), .Z(
        ref_1_maj_56_n21) );
  XOR2_X1 ref_1_maj_56_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(ref_1_maj_56_n22)
         );
  XOR2_X1 ref_1_maj_56_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(ref_1_maj_56_n16)
         );
  OR2_X1 ref_1_maj_56_U6 ( .A1(ref_1_maj_56_n20), .A2(ref_1_maj_56_n19), .ZN(
        ref_1_maj_56_n24) );
  NAND2_X1 ref_1_maj_56_U5 ( .A1(ref_1_maj_56_n24), .A2(ref_1_maj_56_n23), 
        .ZN(ref_1_maj_56_n25) );
  NAND2_X1 ref_1_maj_56_U4 ( .A1(ref_1_maj_56_n20), .A2(ref_1_maj_56_n19), 
        .ZN(ref_1_maj_56_n26) );
  NAND2_X1 ref_1_maj_56_U3 ( .A1(ref_1_maj_56_n26), .A2(ref_1_maj_56_n25), 
        .ZN(ref_1_maj_56_port_o) );
  XOR2_X1 ref_1_maj_56_U2 ( .A(ref_1_maj_56_n22), .B(ref_1_maj_56_n21), .Z(
        ref_1_maj_56_n23) );
  NAND2_X1 ref_1_maj_57_U15 ( .A1(ref_1_refreshed_1_3_), .A2(
        ref_1_refreshed_1_4_), .ZN(ref_1_maj_57_n18) );
  NAND2_X1 ref_1_maj_57_U14 ( .A1(ref_1_maj_57_n21), .A2(ref_1_maj_57_n22), 
        .ZN(ref_1_maj_57_n17) );
  NAND2_X1 ref_1_maj_57_U13 ( .A1(ref_1_maj_57_n18), .A2(ref_1_maj_57_n17), 
        .ZN(ref_1_maj_57_n19) );
  NAND2_X1 ref_1_maj_57_U12 ( .A1(ref_1_refreshed_1_2_), .A2(ref_1_maj_57_n16), 
        .ZN(ref_1_maj_57_n14) );
  NAND2_X1 ref_1_maj_57_U11 ( .A1(ref_1_refreshed_1_0_), .A2(ref_1_n13), .ZN(
        ref_1_maj_57_n15) );
  NAND2_X1 ref_1_maj_57_U10 ( .A1(ref_1_maj_57_n15), .A2(ref_1_maj_57_n14), 
        .ZN(ref_1_maj_57_n20) );
  XOR2_X1 ref_1_maj_57_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_57_n16), 
        .Z(ref_1_maj_57_n21) );
  XOR2_X1 ref_1_maj_57_U8 ( .A(ref_1_refreshed_1_3_), .B(ref_1_refreshed_1_4_), 
        .Z(ref_1_maj_57_n22) );
  XOR2_X1 ref_1_maj_57_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_n13), .Z(
        ref_1_maj_57_n16) );
  OR2_X1 ref_1_maj_57_U6 ( .A1(ref_1_maj_57_n20), .A2(ref_1_maj_57_n19), .ZN(
        ref_1_maj_57_n24) );
  NAND2_X1 ref_1_maj_57_U5 ( .A1(ref_1_maj_57_n24), .A2(ref_1_maj_57_n23), 
        .ZN(ref_1_maj_57_n25) );
  NAND2_X1 ref_1_maj_57_U4 ( .A1(ref_1_maj_57_n20), .A2(ref_1_maj_57_n19), 
        .ZN(ref_1_maj_57_n26) );
  NAND2_X1 ref_1_maj_57_U3 ( .A1(ref_1_maj_57_n26), .A2(ref_1_maj_57_n25), 
        .ZN(ref_1_maj_57_port_o) );
  XOR2_X1 ref_1_maj_57_U2 ( .A(ref_1_maj_57_n22), .B(ref_1_maj_57_n21), .Z(
        ref_1_maj_57_n23) );
  NAND2_X1 ref_1_maj_58_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_58_n18) );
  NAND2_X1 ref_1_maj_58_U14 ( .A1(ref_1_maj_58_n21), .A2(ref_1_maj_58_n22), 
        .ZN(ref_1_maj_58_n17) );
  NAND2_X1 ref_1_maj_58_U13 ( .A1(ref_1_maj_58_n18), .A2(ref_1_maj_58_n17), 
        .ZN(ref_1_maj_58_n19) );
  NAND2_X1 ref_1_maj_58_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_58_n16), .ZN(
        ref_1_maj_58_n14) );
  NAND2_X1 ref_1_maj_58_U11 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_58_n15) );
  NAND2_X1 ref_1_maj_58_U10 ( .A1(ref_1_maj_58_n15), .A2(ref_1_maj_58_n14), 
        .ZN(ref_1_maj_58_n20) );
  XOR2_X1 ref_1_maj_58_U9 ( .A(ref_1_n15), .B(ref_1_maj_58_n16), .Z(
        ref_1_maj_58_n21) );
  XOR2_X1 ref_1_maj_58_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(ref_1_maj_58_n22)
         );
  XOR2_X1 ref_1_maj_58_U7 ( .A(ref_1_n11), .B(ref_1_n14), .Z(ref_1_maj_58_n16)
         );
  OR2_X1 ref_1_maj_58_U6 ( .A1(ref_1_maj_58_n20), .A2(ref_1_maj_58_n19), .ZN(
        ref_1_maj_58_n24) );
  NAND2_X1 ref_1_maj_58_U5 ( .A1(ref_1_maj_58_n24), .A2(ref_1_maj_58_n23), 
        .ZN(ref_1_maj_58_n25) );
  NAND2_X1 ref_1_maj_58_U4 ( .A1(ref_1_maj_58_n20), .A2(ref_1_maj_58_n19), 
        .ZN(ref_1_maj_58_n26) );
  NAND2_X1 ref_1_maj_58_U3 ( .A1(ref_1_maj_58_n26), .A2(ref_1_maj_58_n25), 
        .ZN(ref_1_maj_58_port_o) );
  XOR2_X1 ref_1_maj_58_U2 ( .A(ref_1_maj_58_n22), .B(ref_1_maj_58_n21), .Z(
        ref_1_maj_58_n23) );
  NAND2_X1 ref_1_maj_59_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_59_n18) );
  NAND2_X1 ref_1_maj_59_U14 ( .A1(ref_1_maj_59_n21), .A2(ref_1_maj_59_n22), 
        .ZN(ref_1_maj_59_n17) );
  NAND2_X1 ref_1_maj_59_U13 ( .A1(ref_1_maj_59_n18), .A2(ref_1_maj_59_n17), 
        .ZN(ref_1_maj_59_n19) );
  NAND2_X1 ref_1_maj_59_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_59_n16), .ZN(
        ref_1_maj_59_n14) );
  NAND2_X1 ref_1_maj_59_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_59_n15) );
  NAND2_X1 ref_1_maj_59_U10 ( .A1(ref_1_maj_59_n15), .A2(ref_1_maj_59_n14), 
        .ZN(ref_1_maj_59_n20) );
  XOR2_X1 ref_1_maj_59_U9 ( .A(ref_1_n16), .B(ref_1_maj_59_n16), .Z(
        ref_1_maj_59_n21) );
  XOR2_X1 ref_1_maj_59_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_59_n22)
         );
  XOR2_X1 ref_1_maj_59_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(ref_1_maj_59_n16)
         );
  OR2_X1 ref_1_maj_59_U6 ( .A1(ref_1_maj_59_n20), .A2(ref_1_maj_59_n19), .ZN(
        ref_1_maj_59_n24) );
  NAND2_X1 ref_1_maj_59_U5 ( .A1(ref_1_maj_59_n24), .A2(ref_1_maj_59_n23), 
        .ZN(ref_1_maj_59_n25) );
  NAND2_X1 ref_1_maj_59_U4 ( .A1(ref_1_maj_59_n20), .A2(ref_1_maj_59_n19), 
        .ZN(ref_1_maj_59_n26) );
  NAND2_X1 ref_1_maj_59_U3 ( .A1(ref_1_maj_59_n26), .A2(ref_1_maj_59_n25), 
        .ZN(ref_1_maj_59_port_o) );
  XOR2_X1 ref_1_maj_59_U2 ( .A(ref_1_maj_59_n22), .B(ref_1_maj_59_n21), .Z(
        ref_1_maj_59_n23) );
  NAND2_X1 ref_1_maj_60_U15 ( .A1(ref_1_refreshed_2_3_), .A2(
        ref_1_refreshed_2_4_), .ZN(ref_1_maj_60_n18) );
  NAND2_X1 ref_1_maj_60_U14 ( .A1(ref_1_maj_60_n21), .A2(ref_1_maj_60_n22), 
        .ZN(ref_1_maj_60_n17) );
  NAND2_X1 ref_1_maj_60_U13 ( .A1(ref_1_maj_60_n18), .A2(ref_1_maj_60_n17), 
        .ZN(ref_1_maj_60_n19) );
  NAND2_X1 ref_1_maj_60_U12 ( .A1(ref_1_refreshed_2_2_), .A2(ref_1_maj_60_n16), 
        .ZN(ref_1_maj_60_n14) );
  NAND2_X1 ref_1_maj_60_U11 ( .A1(ref_1_refreshed_2_0_), .A2(ref_1_n3), .ZN(
        ref_1_maj_60_n15) );
  NAND2_X1 ref_1_maj_60_U10 ( .A1(ref_1_maj_60_n15), .A2(ref_1_maj_60_n14), 
        .ZN(ref_1_maj_60_n20) );
  XOR2_X1 ref_1_maj_60_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_60_n16), 
        .Z(ref_1_maj_60_n21) );
  XOR2_X1 ref_1_maj_60_U8 ( .A(ref_1_refreshed_2_3_), .B(ref_1_refreshed_2_4_), 
        .Z(ref_1_maj_60_n22) );
  XOR2_X1 ref_1_maj_60_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_n3), .Z(
        ref_1_maj_60_n16) );
  OR2_X1 ref_1_maj_60_U6 ( .A1(ref_1_maj_60_n20), .A2(ref_1_maj_60_n19), .ZN(
        ref_1_maj_60_n24) );
  NAND2_X1 ref_1_maj_60_U5 ( .A1(ref_1_maj_60_n24), .A2(ref_1_maj_60_n23), 
        .ZN(ref_1_maj_60_n25) );
  NAND2_X1 ref_1_maj_60_U4 ( .A1(ref_1_maj_60_n20), .A2(ref_1_maj_60_n19), 
        .ZN(ref_1_maj_60_n26) );
  NAND2_X1 ref_1_maj_60_U3 ( .A1(ref_1_maj_60_n26), .A2(ref_1_maj_60_n25), 
        .ZN(ref_1_maj_60_port_o) );
  XOR2_X1 ref_1_maj_60_U2 ( .A(ref_1_maj_60_n22), .B(ref_1_maj_60_n21), .Z(
        ref_1_maj_60_n23) );
  NAND2_X1 ref_1_maj_61_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_61_n18) );
  NAND2_X1 ref_1_maj_61_U14 ( .A1(ref_1_maj_61_n21), .A2(ref_1_maj_61_n22), 
        .ZN(ref_1_maj_61_n17) );
  NAND2_X1 ref_1_maj_61_U13 ( .A1(ref_1_maj_61_n18), .A2(ref_1_maj_61_n17), 
        .ZN(ref_1_maj_61_n19) );
  NAND2_X1 ref_1_maj_61_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_61_n16), .ZN(
        ref_1_maj_61_n14) );
  NAND2_X1 ref_1_maj_61_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_61_n15) );
  NAND2_X1 ref_1_maj_61_U10 ( .A1(ref_1_maj_61_n15), .A2(ref_1_maj_61_n14), 
        .ZN(ref_1_maj_61_n20) );
  XOR2_X1 ref_1_maj_61_U9 ( .A(ref_1_n5), .B(ref_1_maj_61_n16), .Z(
        ref_1_maj_61_n21) );
  XOR2_X1 ref_1_maj_61_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_61_n22)
         );
  XOR2_X1 ref_1_maj_61_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_61_n16)
         );
  OR2_X1 ref_1_maj_61_U6 ( .A1(ref_1_maj_61_n20), .A2(ref_1_maj_61_n19), .ZN(
        ref_1_maj_61_n24) );
  NAND2_X1 ref_1_maj_61_U5 ( .A1(ref_1_maj_61_n24), .A2(ref_1_maj_61_n23), 
        .ZN(ref_1_maj_61_n25) );
  NAND2_X1 ref_1_maj_61_U4 ( .A1(ref_1_maj_61_n20), .A2(ref_1_maj_61_n19), 
        .ZN(ref_1_maj_61_n26) );
  NAND2_X1 ref_1_maj_61_U3 ( .A1(ref_1_maj_61_n26), .A2(ref_1_maj_61_n25), 
        .ZN(ref_1_maj_61_port_o) );
  XOR2_X1 ref_1_maj_61_U2 ( .A(ref_1_maj_61_n22), .B(ref_1_maj_61_n21), .Z(
        ref_1_maj_61_n23) );
  NAND2_X1 ref_1_maj_62_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_62_n18) );
  NAND2_X1 ref_1_maj_62_U14 ( .A1(ref_1_maj_62_n21), .A2(ref_1_maj_62_n22), 
        .ZN(ref_1_maj_62_n17) );
  NAND2_X1 ref_1_maj_62_U13 ( .A1(ref_1_maj_62_n18), .A2(ref_1_maj_62_n17), 
        .ZN(ref_1_maj_62_n19) );
  NAND2_X1 ref_1_maj_62_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_62_n16), .ZN(
        ref_1_maj_62_n14) );
  NAND2_X1 ref_1_maj_62_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_62_n15) );
  NAND2_X1 ref_1_maj_62_U10 ( .A1(ref_1_maj_62_n15), .A2(ref_1_maj_62_n14), 
        .ZN(ref_1_maj_62_n20) );
  XOR2_X1 ref_1_maj_62_U9 ( .A(ref_1_n6), .B(ref_1_maj_62_n16), .Z(
        ref_1_maj_62_n21) );
  XOR2_X1 ref_1_maj_62_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_62_n22)
         );
  XOR2_X1 ref_1_maj_62_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_62_n16)
         );
  OR2_X1 ref_1_maj_62_U6 ( .A1(ref_1_maj_62_n20), .A2(ref_1_maj_62_n19), .ZN(
        ref_1_maj_62_n24) );
  NAND2_X1 ref_1_maj_62_U5 ( .A1(ref_1_maj_62_n24), .A2(ref_1_maj_62_n23), 
        .ZN(ref_1_maj_62_n25) );
  NAND2_X1 ref_1_maj_62_U4 ( .A1(ref_1_maj_62_n20), .A2(ref_1_maj_62_n19), 
        .ZN(ref_1_maj_62_n26) );
  NAND2_X1 ref_1_maj_62_U3 ( .A1(ref_1_maj_62_n26), .A2(ref_1_maj_62_n25), 
        .ZN(ref_1_maj_62_port_o) );
  XOR2_X1 ref_1_maj_62_U2 ( .A(ref_1_maj_62_n22), .B(ref_1_maj_62_n21), .Z(
        ref_1_maj_62_n23) );
  NAND2_X1 ref_1_maj_63_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_63_n18) );
  NAND2_X1 ref_1_maj_63_U14 ( .A1(ref_1_maj_63_n21), .A2(ref_1_maj_63_n22), 
        .ZN(ref_1_maj_63_n17) );
  NAND2_X1 ref_1_maj_63_U13 ( .A1(ref_1_maj_63_n18), .A2(ref_1_maj_63_n17), 
        .ZN(ref_1_maj_63_n19) );
  NAND2_X1 ref_1_maj_63_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_63_n16), .ZN(
        ref_1_maj_63_n14) );
  NAND2_X1 ref_1_maj_63_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_63_n15) );
  NAND2_X1 ref_1_maj_63_U10 ( .A1(ref_1_maj_63_n15), .A2(ref_1_maj_63_n14), 
        .ZN(ref_1_maj_63_n20) );
  XOR2_X1 ref_1_maj_63_U9 ( .A(ref_1_n26), .B(ref_1_maj_63_n16), .Z(
        ref_1_maj_63_n21) );
  XOR2_X1 ref_1_maj_63_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_63_n22)
         );
  XOR2_X1 ref_1_maj_63_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(ref_1_maj_63_n16)
         );
  OR2_X1 ref_1_maj_63_U6 ( .A1(ref_1_maj_63_n20), .A2(ref_1_maj_63_n19), .ZN(
        ref_1_maj_63_n24) );
  NAND2_X1 ref_1_maj_63_U5 ( .A1(ref_1_maj_63_n24), .A2(ref_1_maj_63_n23), 
        .ZN(ref_1_maj_63_n25) );
  NAND2_X1 ref_1_maj_63_U4 ( .A1(ref_1_maj_63_n20), .A2(ref_1_maj_63_n19), 
        .ZN(ref_1_maj_63_n26) );
  NAND2_X1 ref_1_maj_63_U3 ( .A1(ref_1_maj_63_n26), .A2(ref_1_maj_63_n25), 
        .ZN(ref_1_maj_63_port_o) );
  XOR2_X1 ref_1_maj_63_U2 ( .A(ref_1_maj_63_n22), .B(ref_1_maj_63_n21), .Z(
        ref_1_maj_63_n23) );
  NAND2_X1 ref_1_maj_64_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_64_n18) );
  NAND2_X1 ref_1_maj_64_U14 ( .A1(ref_1_maj_64_n21), .A2(ref_1_maj_64_n22), 
        .ZN(ref_1_maj_64_n17) );
  NAND2_X1 ref_1_maj_64_U13 ( .A1(ref_1_maj_64_n18), .A2(ref_1_maj_64_n17), 
        .ZN(ref_1_maj_64_n19) );
  NAND2_X1 ref_1_maj_64_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_64_n16), .ZN(
        ref_1_maj_64_n14) );
  NAND2_X1 ref_1_maj_64_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_64_n15) );
  NAND2_X1 ref_1_maj_64_U10 ( .A1(ref_1_maj_64_n15), .A2(ref_1_maj_64_n14), 
        .ZN(ref_1_maj_64_n20) );
  XOR2_X1 ref_1_maj_64_U9 ( .A(ref_1_n25), .B(ref_1_maj_64_n16), .Z(
        ref_1_maj_64_n21) );
  XOR2_X1 ref_1_maj_64_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(ref_1_maj_64_n22)
         );
  XOR2_X1 ref_1_maj_64_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(ref_1_maj_64_n16)
         );
  OR2_X1 ref_1_maj_64_U6 ( .A1(ref_1_maj_64_n20), .A2(ref_1_maj_64_n19), .ZN(
        ref_1_maj_64_n24) );
  NAND2_X1 ref_1_maj_64_U5 ( .A1(ref_1_maj_64_n24), .A2(ref_1_maj_64_n23), 
        .ZN(ref_1_maj_64_n25) );
  NAND2_X1 ref_1_maj_64_U4 ( .A1(ref_1_maj_64_n20), .A2(ref_1_maj_64_n19), 
        .ZN(ref_1_maj_64_n26) );
  NAND2_X1 ref_1_maj_64_U3 ( .A1(ref_1_maj_64_n26), .A2(ref_1_maj_64_n25), 
        .ZN(ref_1_maj_64_port_o) );
  XOR2_X1 ref_1_maj_64_U2 ( .A(ref_1_maj_64_n22), .B(ref_1_maj_64_n21), .Z(
        ref_1_maj_64_n23) );
  NAND2_X1 ref_1_maj_65_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_65_n18) );
  NAND2_X1 ref_1_maj_65_U14 ( .A1(ref_1_maj_65_n21), .A2(ref_1_maj_65_n22), 
        .ZN(ref_1_maj_65_n17) );
  NAND2_X1 ref_1_maj_65_U13 ( .A1(ref_1_maj_65_n18), .A2(ref_1_maj_65_n17), 
        .ZN(ref_1_maj_65_n19) );
  NAND2_X1 ref_1_maj_65_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_65_n16), .ZN(
        ref_1_maj_65_n14) );
  NAND2_X1 ref_1_maj_65_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_65_n15) );
  NAND2_X1 ref_1_maj_65_U10 ( .A1(ref_1_maj_65_n15), .A2(ref_1_maj_65_n14), 
        .ZN(ref_1_maj_65_n20) );
  XOR2_X1 ref_1_maj_65_U9 ( .A(ref_1_n26), .B(ref_1_maj_65_n16), .Z(
        ref_1_maj_65_n21) );
  XOR2_X1 ref_1_maj_65_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_65_n22)
         );
  XOR2_X1 ref_1_maj_65_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(ref_1_maj_65_n16)
         );
  OR2_X1 ref_1_maj_65_U6 ( .A1(ref_1_maj_65_n20), .A2(ref_1_maj_65_n19), .ZN(
        ref_1_maj_65_n24) );
  NAND2_X1 ref_1_maj_65_U5 ( .A1(ref_1_maj_65_n24), .A2(ref_1_maj_65_n23), 
        .ZN(ref_1_maj_65_n25) );
  NAND2_X1 ref_1_maj_65_U4 ( .A1(ref_1_maj_65_n20), .A2(ref_1_maj_65_n19), 
        .ZN(ref_1_maj_65_n26) );
  NAND2_X1 ref_1_maj_65_U3 ( .A1(ref_1_maj_65_n26), .A2(ref_1_maj_65_n25), 
        .ZN(ref_1_maj_65_port_o) );
  XOR2_X1 ref_1_maj_65_U2 ( .A(ref_1_maj_65_n22), .B(ref_1_maj_65_n21), .Z(
        ref_1_maj_65_n23) );
  NAND2_X1 ref_1_maj_66_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_66_n18) );
  NAND2_X1 ref_1_maj_66_U14 ( .A1(ref_1_maj_66_n21), .A2(ref_1_maj_66_n22), 
        .ZN(ref_1_maj_66_n17) );
  NAND2_X1 ref_1_maj_66_U13 ( .A1(ref_1_maj_66_n18), .A2(ref_1_maj_66_n17), 
        .ZN(ref_1_maj_66_n19) );
  NAND2_X1 ref_1_maj_66_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_66_n16), .ZN(
        ref_1_maj_66_n14) );
  NAND2_X1 ref_1_maj_66_U11 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_66_n15) );
  NAND2_X1 ref_1_maj_66_U10 ( .A1(ref_1_maj_66_n15), .A2(ref_1_maj_66_n14), 
        .ZN(ref_1_maj_66_n20) );
  XOR2_X1 ref_1_maj_66_U9 ( .A(ref_1_n15), .B(ref_1_maj_66_n16), .Z(
        ref_1_maj_66_n21) );
  XOR2_X1 ref_1_maj_66_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(ref_1_maj_66_n22)
         );
  XOR2_X1 ref_1_maj_66_U7 ( .A(ref_1_n11), .B(ref_1_n14), .Z(ref_1_maj_66_n16)
         );
  OR2_X1 ref_1_maj_66_U6 ( .A1(ref_1_maj_66_n20), .A2(ref_1_maj_66_n19), .ZN(
        ref_1_maj_66_n24) );
  NAND2_X1 ref_1_maj_66_U5 ( .A1(ref_1_maj_66_n24), .A2(ref_1_maj_66_n23), 
        .ZN(ref_1_maj_66_n25) );
  NAND2_X1 ref_1_maj_66_U4 ( .A1(ref_1_maj_66_n20), .A2(ref_1_maj_66_n19), 
        .ZN(ref_1_maj_66_n26) );
  NAND2_X1 ref_1_maj_66_U3 ( .A1(ref_1_maj_66_n26), .A2(ref_1_maj_66_n25), 
        .ZN(ref_1_maj_66_port_o) );
  XOR2_X1 ref_1_maj_66_U2 ( .A(ref_1_maj_66_n22), .B(ref_1_maj_66_n21), .Z(
        ref_1_maj_66_n23) );
  NAND2_X1 ref_1_maj_67_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_67_n18) );
  NAND2_X1 ref_1_maj_67_U14 ( .A1(ref_1_maj_67_n21), .A2(ref_1_maj_67_n22), 
        .ZN(ref_1_maj_67_n17) );
  NAND2_X1 ref_1_maj_67_U13 ( .A1(ref_1_maj_67_n18), .A2(ref_1_maj_67_n17), 
        .ZN(ref_1_maj_67_n19) );
  NAND2_X1 ref_1_maj_67_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_67_n16), .ZN(
        ref_1_maj_67_n14) );
  NAND2_X1 ref_1_maj_67_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_67_n15) );
  NAND2_X1 ref_1_maj_67_U10 ( .A1(ref_1_maj_67_n15), .A2(ref_1_maj_67_n14), 
        .ZN(ref_1_maj_67_n20) );
  XOR2_X1 ref_1_maj_67_U9 ( .A(ref_1_n16), .B(ref_1_maj_67_n16), .Z(
        ref_1_maj_67_n21) );
  XOR2_X1 ref_1_maj_67_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_67_n22)
         );
  XOR2_X1 ref_1_maj_67_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(ref_1_maj_67_n16)
         );
  OR2_X1 ref_1_maj_67_U6 ( .A1(ref_1_maj_67_n20), .A2(ref_1_maj_67_n19), .ZN(
        ref_1_maj_67_n24) );
  NAND2_X1 ref_1_maj_67_U5 ( .A1(ref_1_maj_67_n24), .A2(ref_1_maj_67_n23), 
        .ZN(ref_1_maj_67_n25) );
  NAND2_X1 ref_1_maj_67_U4 ( .A1(ref_1_maj_67_n20), .A2(ref_1_maj_67_n19), 
        .ZN(ref_1_maj_67_n26) );
  NAND2_X1 ref_1_maj_67_U3 ( .A1(ref_1_maj_67_n26), .A2(ref_1_maj_67_n25), 
        .ZN(ref_1_maj_67_port_o) );
  XOR2_X1 ref_1_maj_67_U2 ( .A(ref_1_maj_67_n22), .B(ref_1_maj_67_n21), .Z(
        ref_1_maj_67_n23) );
  NAND2_X1 ref_1_maj_68_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_68_n18) );
  NAND2_X1 ref_1_maj_68_U14 ( .A1(ref_1_maj_68_n21), .A2(ref_1_maj_68_n22), 
        .ZN(ref_1_maj_68_n17) );
  NAND2_X1 ref_1_maj_68_U13 ( .A1(ref_1_maj_68_n18), .A2(ref_1_maj_68_n17), 
        .ZN(ref_1_maj_68_n19) );
  NAND2_X1 ref_1_maj_68_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_68_n16), .ZN(
        ref_1_maj_68_n14) );
  NAND2_X1 ref_1_maj_68_U11 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_68_n15) );
  NAND2_X1 ref_1_maj_68_U10 ( .A1(ref_1_maj_68_n15), .A2(ref_1_maj_68_n14), 
        .ZN(ref_1_maj_68_n20) );
  XOR2_X1 ref_1_maj_68_U9 ( .A(ref_1_n15), .B(ref_1_maj_68_n16), .Z(
        ref_1_maj_68_n21) );
  XOR2_X1 ref_1_maj_68_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(ref_1_maj_68_n22)
         );
  XOR2_X1 ref_1_maj_68_U7 ( .A(ref_1_n11), .B(ref_1_n14), .Z(ref_1_maj_68_n16)
         );
  OR2_X1 ref_1_maj_68_U6 ( .A1(ref_1_maj_68_n20), .A2(ref_1_maj_68_n19), .ZN(
        ref_1_maj_68_n24) );
  NAND2_X1 ref_1_maj_68_U5 ( .A1(ref_1_maj_68_n24), .A2(ref_1_maj_68_n23), 
        .ZN(ref_1_maj_68_n25) );
  NAND2_X1 ref_1_maj_68_U4 ( .A1(ref_1_maj_68_n20), .A2(ref_1_maj_68_n19), 
        .ZN(ref_1_maj_68_n26) );
  NAND2_X1 ref_1_maj_68_U3 ( .A1(ref_1_maj_68_n26), .A2(ref_1_maj_68_n25), 
        .ZN(ref_1_maj_68_port_o) );
  XOR2_X1 ref_1_maj_68_U2 ( .A(ref_1_maj_68_n22), .B(ref_1_maj_68_n21), .Z(
        ref_1_maj_68_n23) );
  NAND2_X1 ref_1_maj_69_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_69_n18) );
  NAND2_X1 ref_1_maj_69_U14 ( .A1(ref_1_maj_69_n21), .A2(ref_1_maj_69_n22), 
        .ZN(ref_1_maj_69_n17) );
  NAND2_X1 ref_1_maj_69_U13 ( .A1(ref_1_maj_69_n18), .A2(ref_1_maj_69_n17), 
        .ZN(ref_1_maj_69_n19) );
  NAND2_X1 ref_1_maj_69_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_69_n16), .ZN(
        ref_1_maj_69_n14) );
  NAND2_X1 ref_1_maj_69_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_69_n15) );
  NAND2_X1 ref_1_maj_69_U10 ( .A1(ref_1_maj_69_n15), .A2(ref_1_maj_69_n14), 
        .ZN(ref_1_maj_69_n20) );
  XOR2_X1 ref_1_maj_69_U9 ( .A(ref_1_n5), .B(ref_1_maj_69_n16), .Z(
        ref_1_maj_69_n21) );
  XOR2_X1 ref_1_maj_69_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_69_n22)
         );
  XOR2_X1 ref_1_maj_69_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_69_n16)
         );
  OR2_X1 ref_1_maj_69_U6 ( .A1(ref_1_maj_69_n20), .A2(ref_1_maj_69_n19), .ZN(
        ref_1_maj_69_n24) );
  NAND2_X1 ref_1_maj_69_U5 ( .A1(ref_1_maj_69_n24), .A2(ref_1_maj_69_n23), 
        .ZN(ref_1_maj_69_n25) );
  NAND2_X1 ref_1_maj_69_U4 ( .A1(ref_1_maj_69_n20), .A2(ref_1_maj_69_n19), 
        .ZN(ref_1_maj_69_n26) );
  NAND2_X1 ref_1_maj_69_U3 ( .A1(ref_1_maj_69_n26), .A2(ref_1_maj_69_n25), 
        .ZN(ref_1_maj_69_port_o) );
  XOR2_X1 ref_1_maj_69_U2 ( .A(ref_1_maj_69_n22), .B(ref_1_maj_69_n21), .Z(
        ref_1_maj_69_n23) );
  NAND2_X1 ref_1_maj_70_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_70_n18) );
  NAND2_X1 ref_1_maj_70_U14 ( .A1(ref_1_maj_70_n21), .A2(ref_1_maj_70_n22), 
        .ZN(ref_1_maj_70_n17) );
  NAND2_X1 ref_1_maj_70_U13 ( .A1(ref_1_maj_70_n18), .A2(ref_1_maj_70_n17), 
        .ZN(ref_1_maj_70_n19) );
  NAND2_X1 ref_1_maj_70_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_70_n16), .ZN(
        ref_1_maj_70_n14) );
  NAND2_X1 ref_1_maj_70_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_70_n15) );
  NAND2_X1 ref_1_maj_70_U10 ( .A1(ref_1_maj_70_n15), .A2(ref_1_maj_70_n14), 
        .ZN(ref_1_maj_70_n20) );
  XOR2_X1 ref_1_maj_70_U9 ( .A(ref_1_n6), .B(ref_1_maj_70_n16), .Z(
        ref_1_maj_70_n21) );
  XOR2_X1 ref_1_maj_70_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_70_n22)
         );
  XOR2_X1 ref_1_maj_70_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_70_n16)
         );
  OR2_X1 ref_1_maj_70_U6 ( .A1(ref_1_maj_70_n20), .A2(ref_1_maj_70_n19), .ZN(
        ref_1_maj_70_n24) );
  NAND2_X1 ref_1_maj_70_U5 ( .A1(ref_1_maj_70_n24), .A2(ref_1_maj_70_n23), 
        .ZN(ref_1_maj_70_n25) );
  NAND2_X1 ref_1_maj_70_U4 ( .A1(ref_1_maj_70_n20), .A2(ref_1_maj_70_n19), 
        .ZN(ref_1_maj_70_n26) );
  NAND2_X1 ref_1_maj_70_U3 ( .A1(ref_1_maj_70_n26), .A2(ref_1_maj_70_n25), 
        .ZN(ref_1_maj_70_port_o) );
  XOR2_X1 ref_1_maj_70_U2 ( .A(ref_1_maj_70_n22), .B(ref_1_maj_70_n21), .Z(
        ref_1_maj_70_n23) );
  NAND2_X1 ref_1_maj_71_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_71_n18) );
  NAND2_X1 ref_1_maj_71_U14 ( .A1(ref_1_maj_71_n21), .A2(ref_1_maj_71_n22), 
        .ZN(ref_1_maj_71_n17) );
  NAND2_X1 ref_1_maj_71_U13 ( .A1(ref_1_maj_71_n18), .A2(ref_1_maj_71_n17), 
        .ZN(ref_1_maj_71_n19) );
  NAND2_X1 ref_1_maj_71_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_71_n16), .ZN(
        ref_1_maj_71_n14) );
  NAND2_X1 ref_1_maj_71_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_71_n15) );
  NAND2_X1 ref_1_maj_71_U10 ( .A1(ref_1_maj_71_n15), .A2(ref_1_maj_71_n14), 
        .ZN(ref_1_maj_71_n20) );
  XOR2_X1 ref_1_maj_71_U9 ( .A(ref_1_n5), .B(ref_1_maj_71_n16), .Z(
        ref_1_maj_71_n21) );
  XOR2_X1 ref_1_maj_71_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_71_n22)
         );
  XOR2_X1 ref_1_maj_71_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_71_n16)
         );
  OR2_X1 ref_1_maj_71_U6 ( .A1(ref_1_maj_71_n20), .A2(ref_1_maj_71_n19), .ZN(
        ref_1_maj_71_n24) );
  NAND2_X1 ref_1_maj_71_U5 ( .A1(ref_1_maj_71_n24), .A2(ref_1_maj_71_n23), 
        .ZN(ref_1_maj_71_n25) );
  NAND2_X1 ref_1_maj_71_U4 ( .A1(ref_1_maj_71_n20), .A2(ref_1_maj_71_n19), 
        .ZN(ref_1_maj_71_n26) );
  NAND2_X1 ref_1_maj_71_U3 ( .A1(ref_1_maj_71_n26), .A2(ref_1_maj_71_n25), 
        .ZN(ref_1_maj_71_port_o) );
  XOR2_X1 ref_1_maj_71_U2 ( .A(ref_1_maj_71_n22), .B(ref_1_maj_71_n21), .Z(
        ref_1_maj_71_n23) );
  NAND2_X1 ref_1_maj_72_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_72_n18) );
  NAND2_X1 ref_1_maj_72_U14 ( .A1(ref_1_maj_72_n21), .A2(ref_1_maj_72_n22), 
        .ZN(ref_1_maj_72_n17) );
  NAND2_X1 ref_1_maj_72_U13 ( .A1(ref_1_maj_72_n18), .A2(ref_1_maj_72_n17), 
        .ZN(ref_1_maj_72_n19) );
  NAND2_X1 ref_1_maj_72_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_72_n16), .ZN(
        ref_1_maj_72_n14) );
  NAND2_X1 ref_1_maj_72_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_72_n15) );
  NAND2_X1 ref_1_maj_72_U10 ( .A1(ref_1_maj_72_n15), .A2(ref_1_maj_72_n14), 
        .ZN(ref_1_maj_72_n20) );
  XOR2_X1 ref_1_maj_72_U9 ( .A(ref_1_n25), .B(ref_1_maj_72_n16), .Z(
        ref_1_maj_72_n21) );
  XOR2_X1 ref_1_maj_72_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(ref_1_maj_72_n22)
         );
  XOR2_X1 ref_1_maj_72_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(ref_1_maj_72_n16)
         );
  OR2_X1 ref_1_maj_72_U6 ( .A1(ref_1_maj_72_n20), .A2(ref_1_maj_72_n19), .ZN(
        ref_1_maj_72_n24) );
  NAND2_X1 ref_1_maj_72_U5 ( .A1(ref_1_maj_72_n24), .A2(ref_1_maj_72_n23), 
        .ZN(ref_1_maj_72_n25) );
  NAND2_X1 ref_1_maj_72_U4 ( .A1(ref_1_maj_72_n20), .A2(ref_1_maj_72_n19), 
        .ZN(ref_1_maj_72_n26) );
  NAND2_X1 ref_1_maj_72_U3 ( .A1(ref_1_maj_72_n26), .A2(ref_1_maj_72_n25), 
        .ZN(ref_1_maj_72_port_o) );
  XOR2_X1 ref_1_maj_72_U2 ( .A(ref_1_maj_72_n22), .B(ref_1_maj_72_n21), .Z(
        ref_1_maj_72_n23) );
  NAND2_X1 ref_1_maj_73_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_73_n18) );
  NAND2_X1 ref_1_maj_73_U14 ( .A1(ref_1_maj_73_n21), .A2(ref_1_maj_73_n22), 
        .ZN(ref_1_maj_73_n17) );
  NAND2_X1 ref_1_maj_73_U13 ( .A1(ref_1_maj_73_n18), .A2(ref_1_maj_73_n17), 
        .ZN(ref_1_maj_73_n19) );
  NAND2_X1 ref_1_maj_73_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_73_n16), .ZN(
        ref_1_maj_73_n14) );
  NAND2_X1 ref_1_maj_73_U11 ( .A1(ref_1_n21), .A2(ref_1_refreshed_0_1_), .ZN(
        ref_1_maj_73_n15) );
  NAND2_X1 ref_1_maj_73_U10 ( .A1(ref_1_maj_73_n15), .A2(ref_1_maj_73_n14), 
        .ZN(ref_1_maj_73_n20) );
  XOR2_X1 ref_1_maj_73_U9 ( .A(ref_1_n25), .B(ref_1_maj_73_n16), .Z(
        ref_1_maj_73_n21) );
  XOR2_X1 ref_1_maj_73_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(ref_1_maj_73_n22)
         );
  XOR2_X1 ref_1_maj_73_U7 ( .A(ref_1_n21), .B(ref_1_refreshed_0_1_), .Z(
        ref_1_maj_73_n16) );
  OR2_X1 ref_1_maj_73_U6 ( .A1(ref_1_maj_73_n20), .A2(ref_1_maj_73_n19), .ZN(
        ref_1_maj_73_n24) );
  NAND2_X1 ref_1_maj_73_U5 ( .A1(ref_1_maj_73_n24), .A2(ref_1_maj_73_n23), 
        .ZN(ref_1_maj_73_n25) );
  NAND2_X1 ref_1_maj_73_U4 ( .A1(ref_1_maj_73_n20), .A2(ref_1_maj_73_n19), 
        .ZN(ref_1_maj_73_n26) );
  NAND2_X1 ref_1_maj_73_U3 ( .A1(ref_1_maj_73_n26), .A2(ref_1_maj_73_n25), 
        .ZN(ref_1_maj_73_port_o) );
  XOR2_X1 ref_1_maj_73_U2 ( .A(ref_1_maj_73_n22), .B(ref_1_maj_73_n21), .Z(
        ref_1_maj_73_n23) );
  NAND2_X1 ref_1_maj_74_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_74_n18) );
  NAND2_X1 ref_1_maj_74_U14 ( .A1(ref_1_maj_74_n21), .A2(ref_1_maj_74_n22), 
        .ZN(ref_1_maj_74_n17) );
  NAND2_X1 ref_1_maj_74_U13 ( .A1(ref_1_maj_74_n18), .A2(ref_1_maj_74_n17), 
        .ZN(ref_1_maj_74_n19) );
  NAND2_X1 ref_1_maj_74_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_74_n16), .ZN(
        ref_1_maj_74_n14) );
  NAND2_X1 ref_1_maj_74_U11 ( .A1(ref_1_n21), .A2(ref_1_refreshed_0_1_), .ZN(
        ref_1_maj_74_n15) );
  NAND2_X1 ref_1_maj_74_U10 ( .A1(ref_1_maj_74_n15), .A2(ref_1_maj_74_n14), 
        .ZN(ref_1_maj_74_n20) );
  XOR2_X1 ref_1_maj_74_U9 ( .A(ref_1_n25), .B(ref_1_maj_74_n16), .Z(
        ref_1_maj_74_n21) );
  XOR2_X1 ref_1_maj_74_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(ref_1_maj_74_n22)
         );
  XOR2_X1 ref_1_maj_74_U7 ( .A(ref_1_n21), .B(ref_1_refreshed_0_1_), .Z(
        ref_1_maj_74_n16) );
  OR2_X1 ref_1_maj_74_U6 ( .A1(ref_1_maj_74_n20), .A2(ref_1_maj_74_n19), .ZN(
        ref_1_maj_74_n24) );
  NAND2_X1 ref_1_maj_74_U5 ( .A1(ref_1_maj_74_n24), .A2(ref_1_maj_74_n23), 
        .ZN(ref_1_maj_74_n25) );
  NAND2_X1 ref_1_maj_74_U4 ( .A1(ref_1_maj_74_n20), .A2(ref_1_maj_74_n19), 
        .ZN(ref_1_maj_74_n26) );
  NAND2_X1 ref_1_maj_74_U3 ( .A1(ref_1_maj_74_n26), .A2(ref_1_maj_74_n25), 
        .ZN(ref_1_maj_74_port_o) );
  XOR2_X1 ref_1_maj_74_U2 ( .A(ref_1_maj_74_n22), .B(ref_1_maj_74_n21), .Z(
        ref_1_maj_74_n23) );
  NAND2_X1 ref_1_maj_75_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_75_n18) );
  NAND2_X1 ref_1_maj_75_U14 ( .A1(ref_1_maj_75_n21), .A2(ref_1_maj_75_n22), 
        .ZN(ref_1_maj_75_n17) );
  NAND2_X1 ref_1_maj_75_U13 ( .A1(ref_1_maj_75_n18), .A2(ref_1_maj_75_n17), 
        .ZN(ref_1_maj_75_n19) );
  NAND2_X1 ref_1_maj_75_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_75_n16), .ZN(
        ref_1_maj_75_n14) );
  NAND2_X1 ref_1_maj_75_U11 ( .A1(ref_1_n11), .A2(ref_1_refreshed_1_1_), .ZN(
        ref_1_maj_75_n15) );
  NAND2_X1 ref_1_maj_75_U10 ( .A1(ref_1_maj_75_n15), .A2(ref_1_maj_75_n14), 
        .ZN(ref_1_maj_75_n20) );
  XOR2_X1 ref_1_maj_75_U9 ( .A(ref_1_n15), .B(ref_1_maj_75_n16), .Z(
        ref_1_maj_75_n21) );
  XOR2_X1 ref_1_maj_75_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(ref_1_maj_75_n22)
         );
  XOR2_X1 ref_1_maj_75_U7 ( .A(ref_1_n11), .B(ref_1_refreshed_1_1_), .Z(
        ref_1_maj_75_n16) );
  OR2_X1 ref_1_maj_75_U6 ( .A1(ref_1_maj_75_n20), .A2(ref_1_maj_75_n19), .ZN(
        ref_1_maj_75_n24) );
  NAND2_X1 ref_1_maj_75_U5 ( .A1(ref_1_maj_75_n24), .A2(ref_1_maj_75_n23), 
        .ZN(ref_1_maj_75_n25) );
  NAND2_X1 ref_1_maj_75_U4 ( .A1(ref_1_maj_75_n20), .A2(ref_1_maj_75_n19), 
        .ZN(ref_1_maj_75_n26) );
  NAND2_X1 ref_1_maj_75_U3 ( .A1(ref_1_maj_75_n26), .A2(ref_1_maj_75_n25), 
        .ZN(ref_1_maj_75_port_o) );
  XOR2_X1 ref_1_maj_75_U2 ( .A(ref_1_maj_75_n22), .B(ref_1_maj_75_n21), .Z(
        ref_1_maj_75_n23) );
  NAND2_X1 ref_1_maj_76_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_76_n18) );
  NAND2_X1 ref_1_maj_76_U14 ( .A1(ref_1_maj_76_n21), .A2(ref_1_maj_76_n22), 
        .ZN(ref_1_maj_76_n17) );
  NAND2_X1 ref_1_maj_76_U13 ( .A1(ref_1_maj_76_n18), .A2(ref_1_maj_76_n17), 
        .ZN(ref_1_maj_76_n19) );
  NAND2_X1 ref_1_maj_76_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_76_n16), .ZN(
        ref_1_maj_76_n14) );
  NAND2_X1 ref_1_maj_76_U11 ( .A1(ref_1_n11), .A2(ref_1_refreshed_1_1_), .ZN(
        ref_1_maj_76_n15) );
  NAND2_X1 ref_1_maj_76_U10 ( .A1(ref_1_maj_76_n15), .A2(ref_1_maj_76_n14), 
        .ZN(ref_1_maj_76_n20) );
  XOR2_X1 ref_1_maj_76_U9 ( .A(ref_1_n15), .B(ref_1_maj_76_n16), .Z(
        ref_1_maj_76_n21) );
  XOR2_X1 ref_1_maj_76_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(ref_1_maj_76_n22)
         );
  XOR2_X1 ref_1_maj_76_U7 ( .A(ref_1_n11), .B(ref_1_refreshed_1_1_), .Z(
        ref_1_maj_76_n16) );
  OR2_X1 ref_1_maj_76_U6 ( .A1(ref_1_maj_76_n20), .A2(ref_1_maj_76_n19), .ZN(
        ref_1_maj_76_n24) );
  NAND2_X1 ref_1_maj_76_U5 ( .A1(ref_1_maj_76_n24), .A2(ref_1_maj_76_n23), 
        .ZN(ref_1_maj_76_n25) );
  NAND2_X1 ref_1_maj_76_U4 ( .A1(ref_1_maj_76_n20), .A2(ref_1_maj_76_n19), 
        .ZN(ref_1_maj_76_n26) );
  NAND2_X1 ref_1_maj_76_U3 ( .A1(ref_1_maj_76_n26), .A2(ref_1_maj_76_n25), 
        .ZN(ref_1_maj_76_port_o) );
  XOR2_X1 ref_1_maj_76_U2 ( .A(ref_1_maj_76_n22), .B(ref_1_maj_76_n21), .Z(
        ref_1_maj_76_n23) );
  NAND2_X1 ref_1_maj_77_U15 ( .A1(ref_1_n17), .A2(ref_1_n19), .ZN(
        ref_1_maj_77_n18) );
  NAND2_X1 ref_1_maj_77_U14 ( .A1(ref_1_maj_77_n21), .A2(ref_1_maj_77_n22), 
        .ZN(ref_1_maj_77_n17) );
  NAND2_X1 ref_1_maj_77_U13 ( .A1(ref_1_maj_77_n18), .A2(ref_1_maj_77_n17), 
        .ZN(ref_1_maj_77_n19) );
  NAND2_X1 ref_1_maj_77_U12 ( .A1(ref_1_n15), .A2(ref_1_maj_77_n16), .ZN(
        ref_1_maj_77_n14) );
  NAND2_X1 ref_1_maj_77_U11 ( .A1(ref_1_n11), .A2(ref_1_refreshed_1_1_), .ZN(
        ref_1_maj_77_n15) );
  NAND2_X1 ref_1_maj_77_U10 ( .A1(ref_1_maj_77_n15), .A2(ref_1_maj_77_n14), 
        .ZN(ref_1_maj_77_n20) );
  XOR2_X1 ref_1_maj_77_U9 ( .A(ref_1_n15), .B(ref_1_maj_77_n16), .Z(
        ref_1_maj_77_n21) );
  XOR2_X1 ref_1_maj_77_U8 ( .A(ref_1_n17), .B(ref_1_n19), .Z(ref_1_maj_77_n22)
         );
  XOR2_X1 ref_1_maj_77_U7 ( .A(ref_1_n11), .B(ref_1_refreshed_1_1_), .Z(
        ref_1_maj_77_n16) );
  OR2_X1 ref_1_maj_77_U6 ( .A1(ref_1_maj_77_n20), .A2(ref_1_maj_77_n19), .ZN(
        ref_1_maj_77_n24) );
  NAND2_X1 ref_1_maj_77_U5 ( .A1(ref_1_maj_77_n24), .A2(ref_1_maj_77_n23), 
        .ZN(ref_1_maj_77_n25) );
  NAND2_X1 ref_1_maj_77_U4 ( .A1(ref_1_maj_77_n20), .A2(ref_1_maj_77_n19), 
        .ZN(ref_1_maj_77_n26) );
  NAND2_X1 ref_1_maj_77_U3 ( .A1(ref_1_maj_77_n26), .A2(ref_1_maj_77_n25), 
        .ZN(ref_1_maj_77_port_o) );
  XOR2_X1 ref_1_maj_77_U2 ( .A(ref_1_maj_77_n22), .B(ref_1_maj_77_n21), .Z(
        ref_1_maj_77_n23) );
  NAND2_X1 ref_1_maj_78_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_78_n18) );
  NAND2_X1 ref_1_maj_78_U14 ( .A1(ref_1_maj_78_n21), .A2(ref_1_maj_78_n22), 
        .ZN(ref_1_maj_78_n17) );
  NAND2_X1 ref_1_maj_78_U13 ( .A1(ref_1_maj_78_n18), .A2(ref_1_maj_78_n17), 
        .ZN(ref_1_maj_78_n19) );
  NAND2_X1 ref_1_maj_78_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_78_n16), .ZN(
        ref_1_maj_78_n14) );
  NAND2_X1 ref_1_maj_78_U11 ( .A1(ref_1_n1), .A2(ref_1_refreshed_2_1_), .ZN(
        ref_1_maj_78_n15) );
  NAND2_X1 ref_1_maj_78_U10 ( .A1(ref_1_maj_78_n15), .A2(ref_1_maj_78_n14), 
        .ZN(ref_1_maj_78_n20) );
  XOR2_X1 ref_1_maj_78_U9 ( .A(ref_1_n5), .B(ref_1_maj_78_n16), .Z(
        ref_1_maj_78_n21) );
  XOR2_X1 ref_1_maj_78_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_78_n22)
         );
  XOR2_X1 ref_1_maj_78_U7 ( .A(ref_1_n1), .B(ref_1_refreshed_2_1_), .Z(
        ref_1_maj_78_n16) );
  OR2_X1 ref_1_maj_78_U6 ( .A1(ref_1_maj_78_n20), .A2(ref_1_maj_78_n19), .ZN(
        ref_1_maj_78_n24) );
  NAND2_X1 ref_1_maj_78_U5 ( .A1(ref_1_maj_78_n24), .A2(ref_1_maj_78_n23), 
        .ZN(ref_1_maj_78_n25) );
  NAND2_X1 ref_1_maj_78_U4 ( .A1(ref_1_maj_78_n20), .A2(ref_1_maj_78_n19), 
        .ZN(ref_1_maj_78_n26) );
  NAND2_X1 ref_1_maj_78_U3 ( .A1(ref_1_maj_78_n26), .A2(ref_1_maj_78_n25), 
        .ZN(ref_1_maj_78_port_o) );
  XOR2_X1 ref_1_maj_78_U2 ( .A(ref_1_maj_78_n22), .B(ref_1_maj_78_n21), .Z(
        ref_1_maj_78_n23) );
  NAND2_X1 ref_1_maj_79_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_79_n18) );
  NAND2_X1 ref_1_maj_79_U14 ( .A1(ref_1_maj_79_n21), .A2(ref_1_maj_79_n22), 
        .ZN(ref_1_maj_79_n17) );
  NAND2_X1 ref_1_maj_79_U13 ( .A1(ref_1_maj_79_n18), .A2(ref_1_maj_79_n17), 
        .ZN(ref_1_maj_79_n19) );
  NAND2_X1 ref_1_maj_79_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_79_n16), .ZN(
        ref_1_maj_79_n14) );
  NAND2_X1 ref_1_maj_79_U11 ( .A1(ref_1_n1), .A2(ref_1_refreshed_2_1_), .ZN(
        ref_1_maj_79_n15) );
  NAND2_X1 ref_1_maj_79_U10 ( .A1(ref_1_maj_79_n15), .A2(ref_1_maj_79_n14), 
        .ZN(ref_1_maj_79_n20) );
  XOR2_X1 ref_1_maj_79_U9 ( .A(ref_1_n5), .B(ref_1_maj_79_n16), .Z(
        ref_1_maj_79_n21) );
  XOR2_X1 ref_1_maj_79_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_79_n22)
         );
  XOR2_X1 ref_1_maj_79_U7 ( .A(ref_1_n1), .B(ref_1_refreshed_2_1_), .Z(
        ref_1_maj_79_n16) );
  OR2_X1 ref_1_maj_79_U6 ( .A1(ref_1_maj_79_n20), .A2(ref_1_maj_79_n19), .ZN(
        ref_1_maj_79_n24) );
  NAND2_X1 ref_1_maj_79_U5 ( .A1(ref_1_maj_79_n24), .A2(ref_1_maj_79_n23), 
        .ZN(ref_1_maj_79_n25) );
  NAND2_X1 ref_1_maj_79_U4 ( .A1(ref_1_maj_79_n20), .A2(ref_1_maj_79_n19), 
        .ZN(ref_1_maj_79_n26) );
  NAND2_X1 ref_1_maj_79_U3 ( .A1(ref_1_maj_79_n26), .A2(ref_1_maj_79_n25), 
        .ZN(ref_1_maj_79_port_o) );
  XOR2_X1 ref_1_maj_79_U2 ( .A(ref_1_maj_79_n22), .B(ref_1_maj_79_n21), .Z(
        ref_1_maj_79_n23) );
  NAND2_X1 ref_1_maj_80_U15 ( .A1(ref_1_n7), .A2(ref_1_n9), .ZN(
        ref_1_maj_80_n18) );
  NAND2_X1 ref_1_maj_80_U14 ( .A1(ref_1_maj_80_n21), .A2(ref_1_maj_80_n22), 
        .ZN(ref_1_maj_80_n17) );
  NAND2_X1 ref_1_maj_80_U13 ( .A1(ref_1_maj_80_n18), .A2(ref_1_maj_80_n17), 
        .ZN(ref_1_maj_80_n19) );
  NAND2_X1 ref_1_maj_80_U12 ( .A1(ref_1_n5), .A2(ref_1_maj_80_n16), .ZN(
        ref_1_maj_80_n14) );
  NAND2_X1 ref_1_maj_80_U11 ( .A1(ref_1_n1), .A2(ref_1_refreshed_2_1_), .ZN(
        ref_1_maj_80_n15) );
  NAND2_X1 ref_1_maj_80_U10 ( .A1(ref_1_maj_80_n15), .A2(ref_1_maj_80_n14), 
        .ZN(ref_1_maj_80_n20) );
  XOR2_X1 ref_1_maj_80_U9 ( .A(ref_1_n5), .B(ref_1_maj_80_n16), .Z(
        ref_1_maj_80_n21) );
  XOR2_X1 ref_1_maj_80_U8 ( .A(ref_1_n7), .B(ref_1_n9), .Z(ref_1_maj_80_n22)
         );
  XOR2_X1 ref_1_maj_80_U7 ( .A(ref_1_n1), .B(ref_1_refreshed_2_1_), .Z(
        ref_1_maj_80_n16) );
  OR2_X1 ref_1_maj_80_U6 ( .A1(ref_1_maj_80_n20), .A2(ref_1_maj_80_n19), .ZN(
        ref_1_maj_80_n24) );
  NAND2_X1 ref_1_maj_80_U5 ( .A1(ref_1_maj_80_n24), .A2(ref_1_maj_80_n23), 
        .ZN(ref_1_maj_80_n25) );
  NAND2_X1 ref_1_maj_80_U4 ( .A1(ref_1_maj_80_n20), .A2(ref_1_maj_80_n19), 
        .ZN(ref_1_maj_80_n26) );
  NAND2_X1 ref_1_maj_80_U3 ( .A1(ref_1_maj_80_n26), .A2(ref_1_maj_80_n25), 
        .ZN(ref_1_maj_80_port_o) );
  XOR2_X1 ref_1_maj_80_U2 ( .A(ref_1_maj_80_n22), .B(ref_1_maj_80_n21), .Z(
        ref_1_maj_80_n23) );
  NAND2_X1 ref_1_maj_81_U15 ( .A1(ref_1_n27), .A2(ref_1_n29), .ZN(
        ref_1_maj_81_n18) );
  NAND2_X1 ref_1_maj_81_U14 ( .A1(ref_1_maj_81_n21), .A2(ref_1_maj_81_n22), 
        .ZN(ref_1_maj_81_n17) );
  NAND2_X1 ref_1_maj_81_U13 ( .A1(ref_1_maj_81_n18), .A2(ref_1_maj_81_n17), 
        .ZN(ref_1_maj_81_n19) );
  NAND2_X1 ref_1_maj_81_U12 ( .A1(ref_1_n25), .A2(ref_1_maj_81_n16), .ZN(
        ref_1_maj_81_n14) );
  NAND2_X1 ref_1_maj_81_U11 ( .A1(ref_1_n21), .A2(ref_1_refreshed_0_1_), .ZN(
        ref_1_maj_81_n15) );
  NAND2_X1 ref_1_maj_81_U10 ( .A1(ref_1_maj_81_n15), .A2(ref_1_maj_81_n14), 
        .ZN(ref_1_maj_81_n20) );
  XOR2_X1 ref_1_maj_81_U9 ( .A(ref_1_n25), .B(ref_1_maj_81_n16), .Z(
        ref_1_maj_81_n21) );
  XOR2_X1 ref_1_maj_81_U8 ( .A(ref_1_n27), .B(ref_1_n29), .Z(ref_1_maj_81_n22)
         );
  XOR2_X1 ref_1_maj_81_U7 ( .A(ref_1_n21), .B(ref_1_refreshed_0_1_), .Z(
        ref_1_maj_81_n16) );
  OR2_X1 ref_1_maj_81_U6 ( .A1(ref_1_maj_81_n20), .A2(ref_1_maj_81_n19), .ZN(
        ref_1_maj_81_n24) );
  NAND2_X1 ref_1_maj_81_U5 ( .A1(ref_1_maj_81_n24), .A2(ref_1_maj_81_n23), 
        .ZN(ref_1_maj_81_n25) );
  NAND2_X1 ref_1_maj_81_U4 ( .A1(ref_1_maj_81_n20), .A2(ref_1_maj_81_n19), 
        .ZN(ref_1_maj_81_n26) );
  NAND2_X1 ref_1_maj_81_U3 ( .A1(ref_1_maj_81_n26), .A2(ref_1_maj_81_n25), 
        .ZN(ref_1_maj_81_port_o) );
  XOR2_X1 ref_1_maj_81_U2 ( .A(ref_1_maj_81_n22), .B(ref_1_maj_81_n21), .Z(
        ref_1_maj_81_n23) );
  NAND2_X1 ref_1_maj_82_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_82_n18) );
  NAND2_X1 ref_1_maj_82_U14 ( .A1(ref_1_maj_82_n21), .A2(ref_1_maj_82_n22), 
        .ZN(ref_1_maj_82_n17) );
  NAND2_X1 ref_1_maj_82_U13 ( .A1(ref_1_maj_82_n18), .A2(ref_1_maj_82_n17), 
        .ZN(ref_1_maj_82_n19) );
  NAND2_X1 ref_1_maj_82_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_82_n16), .ZN(
        ref_1_maj_82_n14) );
  NAND2_X1 ref_1_maj_82_U11 ( .A1(ref_1_n22), .A2(ref_1_n23), .ZN(
        ref_1_maj_82_n15) );
  NAND2_X1 ref_1_maj_82_U10 ( .A1(ref_1_maj_82_n15), .A2(ref_1_maj_82_n14), 
        .ZN(ref_1_maj_82_n20) );
  XOR2_X1 ref_1_maj_82_U9 ( .A(ref_1_n26), .B(ref_1_maj_82_n16), .Z(
        ref_1_maj_82_n21) );
  XOR2_X1 ref_1_maj_82_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_82_n22)
         );
  XOR2_X1 ref_1_maj_82_U7 ( .A(ref_1_n22), .B(ref_1_n23), .Z(ref_1_maj_82_n16)
         );
  OR2_X1 ref_1_maj_82_U6 ( .A1(ref_1_maj_82_n20), .A2(ref_1_maj_82_n19), .ZN(
        ref_1_maj_82_n24) );
  NAND2_X1 ref_1_maj_82_U5 ( .A1(ref_1_maj_82_n24), .A2(ref_1_maj_82_n23), 
        .ZN(ref_1_maj_82_n25) );
  NAND2_X1 ref_1_maj_82_U4 ( .A1(ref_1_maj_82_n20), .A2(ref_1_maj_82_n19), 
        .ZN(ref_1_maj_82_n26) );
  NAND2_X1 ref_1_maj_82_U3 ( .A1(ref_1_maj_82_n26), .A2(ref_1_maj_82_n25), 
        .ZN(ref_1_maj_82_port_o) );
  XOR2_X1 ref_1_maj_82_U2 ( .A(ref_1_maj_82_n22), .B(ref_1_maj_82_n21), .Z(
        ref_1_maj_82_n23) );
  NAND2_X1 ref_1_maj_83_U15 ( .A1(ref_1_n28), .A2(ref_1_n30), .ZN(
        ref_1_maj_83_n18) );
  NAND2_X1 ref_1_maj_83_U14 ( .A1(ref_1_maj_83_n21), .A2(ref_1_maj_83_n22), 
        .ZN(ref_1_maj_83_n17) );
  NAND2_X1 ref_1_maj_83_U13 ( .A1(ref_1_maj_83_n18), .A2(ref_1_maj_83_n17), 
        .ZN(ref_1_maj_83_n19) );
  NAND2_X1 ref_1_maj_83_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_83_n16), .ZN(
        ref_1_maj_83_n14) );
  NAND2_X1 ref_1_maj_83_U11 ( .A1(ref_1_n22), .A2(ref_1_n24), .ZN(
        ref_1_maj_83_n15) );
  NAND2_X1 ref_1_maj_83_U10 ( .A1(ref_1_maj_83_n15), .A2(ref_1_maj_83_n14), 
        .ZN(ref_1_maj_83_n20) );
  XOR2_X1 ref_1_maj_83_U9 ( .A(ref_1_n26), .B(ref_1_maj_83_n16), .Z(
        ref_1_maj_83_n21) );
  XOR2_X1 ref_1_maj_83_U8 ( .A(ref_1_n28), .B(ref_1_n30), .Z(ref_1_maj_83_n22)
         );
  XOR2_X1 ref_1_maj_83_U7 ( .A(ref_1_n22), .B(ref_1_n24), .Z(ref_1_maj_83_n16)
         );
  OR2_X1 ref_1_maj_83_U6 ( .A1(ref_1_maj_83_n20), .A2(ref_1_maj_83_n19), .ZN(
        ref_1_maj_83_n24) );
  NAND2_X1 ref_1_maj_83_U5 ( .A1(ref_1_maj_83_n24), .A2(ref_1_maj_83_n23), 
        .ZN(ref_1_maj_83_n25) );
  NAND2_X1 ref_1_maj_83_U4 ( .A1(ref_1_maj_83_n20), .A2(ref_1_maj_83_n19), 
        .ZN(ref_1_maj_83_n26) );
  NAND2_X1 ref_1_maj_83_U3 ( .A1(ref_1_maj_83_n26), .A2(ref_1_maj_83_n25), 
        .ZN(ref_1_maj_83_port_o) );
  XOR2_X1 ref_1_maj_83_U2 ( .A(ref_1_maj_83_n22), .B(ref_1_maj_83_n21), .Z(
        ref_1_maj_83_n23) );
  NAND2_X1 ref_1_maj_84_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_84_n18) );
  NAND2_X1 ref_1_maj_84_U14 ( .A1(ref_1_maj_84_n21), .A2(ref_1_maj_84_n22), 
        .ZN(ref_1_maj_84_n17) );
  NAND2_X1 ref_1_maj_84_U13 ( .A1(ref_1_maj_84_n18), .A2(ref_1_maj_84_n17), 
        .ZN(ref_1_maj_84_n19) );
  NAND2_X1 ref_1_maj_84_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_84_n16), .ZN(
        ref_1_maj_84_n14) );
  NAND2_X1 ref_1_maj_84_U11 ( .A1(ref_1_n12), .A2(ref_1_n13), .ZN(
        ref_1_maj_84_n15) );
  NAND2_X1 ref_1_maj_84_U10 ( .A1(ref_1_maj_84_n15), .A2(ref_1_maj_84_n14), 
        .ZN(ref_1_maj_84_n20) );
  XOR2_X1 ref_1_maj_84_U9 ( .A(ref_1_n16), .B(ref_1_maj_84_n16), .Z(
        ref_1_maj_84_n21) );
  XOR2_X1 ref_1_maj_84_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_84_n22)
         );
  XOR2_X1 ref_1_maj_84_U7 ( .A(ref_1_n12), .B(ref_1_n13), .Z(ref_1_maj_84_n16)
         );
  OR2_X1 ref_1_maj_84_U6 ( .A1(ref_1_maj_84_n20), .A2(ref_1_maj_84_n19), .ZN(
        ref_1_maj_84_n24) );
  NAND2_X1 ref_1_maj_84_U5 ( .A1(ref_1_maj_84_n24), .A2(ref_1_maj_84_n23), 
        .ZN(ref_1_maj_84_n25) );
  NAND2_X1 ref_1_maj_84_U4 ( .A1(ref_1_maj_84_n20), .A2(ref_1_maj_84_n19), 
        .ZN(ref_1_maj_84_n26) );
  NAND2_X1 ref_1_maj_84_U3 ( .A1(ref_1_maj_84_n26), .A2(ref_1_maj_84_n25), 
        .ZN(ref_1_maj_84_port_o) );
  XOR2_X1 ref_1_maj_84_U2 ( .A(ref_1_maj_84_n22), .B(ref_1_maj_84_n21), .Z(
        ref_1_maj_84_n23) );
  NAND2_X1 ref_1_maj_85_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_85_n18) );
  NAND2_X1 ref_1_maj_85_U14 ( .A1(ref_1_maj_85_n21), .A2(ref_1_maj_85_n22), 
        .ZN(ref_1_maj_85_n17) );
  NAND2_X1 ref_1_maj_85_U13 ( .A1(ref_1_maj_85_n18), .A2(ref_1_maj_85_n17), 
        .ZN(ref_1_maj_85_n19) );
  NAND2_X1 ref_1_maj_85_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_85_n16), .ZN(
        ref_1_maj_85_n14) );
  NAND2_X1 ref_1_maj_85_U11 ( .A1(ref_1_n12), .A2(ref_1_n14), .ZN(
        ref_1_maj_85_n15) );
  NAND2_X1 ref_1_maj_85_U10 ( .A1(ref_1_maj_85_n15), .A2(ref_1_maj_85_n14), 
        .ZN(ref_1_maj_85_n20) );
  XOR2_X1 ref_1_maj_85_U9 ( .A(ref_1_n16), .B(ref_1_maj_85_n16), .Z(
        ref_1_maj_85_n21) );
  XOR2_X1 ref_1_maj_85_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_85_n22)
         );
  XOR2_X1 ref_1_maj_85_U7 ( .A(ref_1_n12), .B(ref_1_n14), .Z(ref_1_maj_85_n16)
         );
  OR2_X1 ref_1_maj_85_U6 ( .A1(ref_1_maj_85_n20), .A2(ref_1_maj_85_n19), .ZN(
        ref_1_maj_85_n24) );
  NAND2_X1 ref_1_maj_85_U5 ( .A1(ref_1_maj_85_n24), .A2(ref_1_maj_85_n23), 
        .ZN(ref_1_maj_85_n25) );
  NAND2_X1 ref_1_maj_85_U4 ( .A1(ref_1_maj_85_n20), .A2(ref_1_maj_85_n19), 
        .ZN(ref_1_maj_85_n26) );
  NAND2_X1 ref_1_maj_85_U3 ( .A1(ref_1_maj_85_n26), .A2(ref_1_maj_85_n25), 
        .ZN(ref_1_maj_85_port_o) );
  XOR2_X1 ref_1_maj_85_U2 ( .A(ref_1_maj_85_n22), .B(ref_1_maj_85_n21), .Z(
        ref_1_maj_85_n23) );
  NAND2_X1 ref_1_maj_86_U15 ( .A1(ref_1_n18), .A2(ref_1_n20), .ZN(
        ref_1_maj_86_n18) );
  NAND2_X1 ref_1_maj_86_U14 ( .A1(ref_1_maj_86_n21), .A2(ref_1_maj_86_n22), 
        .ZN(ref_1_maj_86_n17) );
  NAND2_X1 ref_1_maj_86_U13 ( .A1(ref_1_maj_86_n18), .A2(ref_1_maj_86_n17), 
        .ZN(ref_1_maj_86_n19) );
  NAND2_X1 ref_1_maj_86_U12 ( .A1(ref_1_n16), .A2(ref_1_maj_86_n16), .ZN(
        ref_1_maj_86_n14) );
  NAND2_X1 ref_1_maj_86_U11 ( .A1(ref_1_n12), .A2(ref_1_n13), .ZN(
        ref_1_maj_86_n15) );
  NAND2_X1 ref_1_maj_86_U10 ( .A1(ref_1_maj_86_n15), .A2(ref_1_maj_86_n14), 
        .ZN(ref_1_maj_86_n20) );
  XOR2_X1 ref_1_maj_86_U9 ( .A(ref_1_n16), .B(ref_1_maj_86_n16), .Z(
        ref_1_maj_86_n21) );
  XOR2_X1 ref_1_maj_86_U8 ( .A(ref_1_n18), .B(ref_1_n20), .Z(ref_1_maj_86_n22)
         );
  XOR2_X1 ref_1_maj_86_U7 ( .A(ref_1_n12), .B(ref_1_n13), .Z(ref_1_maj_86_n16)
         );
  OR2_X1 ref_1_maj_86_U6 ( .A1(ref_1_maj_86_n20), .A2(ref_1_maj_86_n19), .ZN(
        ref_1_maj_86_n24) );
  NAND2_X1 ref_1_maj_86_U5 ( .A1(ref_1_maj_86_n24), .A2(ref_1_maj_86_n23), 
        .ZN(ref_1_maj_86_n25) );
  NAND2_X1 ref_1_maj_86_U4 ( .A1(ref_1_maj_86_n20), .A2(ref_1_maj_86_n19), 
        .ZN(ref_1_maj_86_n26) );
  NAND2_X1 ref_1_maj_86_U3 ( .A1(ref_1_maj_86_n26), .A2(ref_1_maj_86_n25), 
        .ZN(ref_1_maj_86_port_o) );
  XOR2_X1 ref_1_maj_86_U2 ( .A(ref_1_maj_86_n22), .B(ref_1_maj_86_n21), .Z(
        ref_1_maj_86_n23) );
  NAND2_X1 ref_1_maj_87_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_87_n18) );
  NAND2_X1 ref_1_maj_87_U14 ( .A1(ref_1_maj_87_n21), .A2(ref_1_maj_87_n22), 
        .ZN(ref_1_maj_87_n17) );
  NAND2_X1 ref_1_maj_87_U13 ( .A1(ref_1_maj_87_n18), .A2(ref_1_maj_87_n17), 
        .ZN(ref_1_maj_87_n19) );
  NAND2_X1 ref_1_maj_87_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_87_n16), .ZN(
        ref_1_maj_87_n14) );
  NAND2_X1 ref_1_maj_87_U11 ( .A1(ref_1_n2), .A2(ref_1_n3), .ZN(
        ref_1_maj_87_n15) );
  NAND2_X1 ref_1_maj_87_U10 ( .A1(ref_1_maj_87_n15), .A2(ref_1_maj_87_n14), 
        .ZN(ref_1_maj_87_n20) );
  XOR2_X1 ref_1_maj_87_U9 ( .A(ref_1_n6), .B(ref_1_maj_87_n16), .Z(
        ref_1_maj_87_n21) );
  XOR2_X1 ref_1_maj_87_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_87_n22)
         );
  XOR2_X1 ref_1_maj_87_U7 ( .A(ref_1_n2), .B(ref_1_n3), .Z(ref_1_maj_87_n16)
         );
  OR2_X1 ref_1_maj_87_U6 ( .A1(ref_1_maj_87_n20), .A2(ref_1_maj_87_n19), .ZN(
        ref_1_maj_87_n24) );
  NAND2_X1 ref_1_maj_87_U5 ( .A1(ref_1_maj_87_n24), .A2(ref_1_maj_87_n23), 
        .ZN(ref_1_maj_87_n25) );
  NAND2_X1 ref_1_maj_87_U4 ( .A1(ref_1_maj_87_n20), .A2(ref_1_maj_87_n19), 
        .ZN(ref_1_maj_87_n26) );
  NAND2_X1 ref_1_maj_87_U3 ( .A1(ref_1_maj_87_n26), .A2(ref_1_maj_87_n25), 
        .ZN(ref_1_maj_87_port_o) );
  XOR2_X1 ref_1_maj_87_U2 ( .A(ref_1_maj_87_n22), .B(ref_1_maj_87_n21), .Z(
        ref_1_maj_87_n23) );
  NAND2_X1 ref_1_maj_88_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_88_n18) );
  NAND2_X1 ref_1_maj_88_U14 ( .A1(ref_1_maj_88_n21), .A2(ref_1_maj_88_n22), 
        .ZN(ref_1_maj_88_n17) );
  NAND2_X1 ref_1_maj_88_U13 ( .A1(ref_1_maj_88_n18), .A2(ref_1_maj_88_n17), 
        .ZN(ref_1_maj_88_n19) );
  NAND2_X1 ref_1_maj_88_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_88_n16), .ZN(
        ref_1_maj_88_n14) );
  NAND2_X1 ref_1_maj_88_U11 ( .A1(ref_1_n2), .A2(ref_1_n4), .ZN(
        ref_1_maj_88_n15) );
  NAND2_X1 ref_1_maj_88_U10 ( .A1(ref_1_maj_88_n15), .A2(ref_1_maj_88_n14), 
        .ZN(ref_1_maj_88_n20) );
  XOR2_X1 ref_1_maj_88_U9 ( .A(ref_1_n6), .B(ref_1_maj_88_n16), .Z(
        ref_1_maj_88_n21) );
  XOR2_X1 ref_1_maj_88_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_88_n22)
         );
  XOR2_X1 ref_1_maj_88_U7 ( .A(ref_1_n2), .B(ref_1_n4), .Z(ref_1_maj_88_n16)
         );
  OR2_X1 ref_1_maj_88_U6 ( .A1(ref_1_maj_88_n20), .A2(ref_1_maj_88_n19), .ZN(
        ref_1_maj_88_n24) );
  NAND2_X1 ref_1_maj_88_U5 ( .A1(ref_1_maj_88_n24), .A2(ref_1_maj_88_n23), 
        .ZN(ref_1_maj_88_n25) );
  NAND2_X1 ref_1_maj_88_U4 ( .A1(ref_1_maj_88_n20), .A2(ref_1_maj_88_n19), 
        .ZN(ref_1_maj_88_n26) );
  NAND2_X1 ref_1_maj_88_U3 ( .A1(ref_1_maj_88_n26), .A2(ref_1_maj_88_n25), 
        .ZN(ref_1_maj_88_port_o) );
  XOR2_X1 ref_1_maj_88_U2 ( .A(ref_1_maj_88_n22), .B(ref_1_maj_88_n21), .Z(
        ref_1_maj_88_n23) );
  NAND2_X1 ref_1_maj_89_U15 ( .A1(ref_1_n8), .A2(ref_1_n10), .ZN(
        ref_1_maj_89_n18) );
  NAND2_X1 ref_1_maj_89_U14 ( .A1(ref_1_maj_89_n21), .A2(ref_1_maj_89_n22), 
        .ZN(ref_1_maj_89_n17) );
  NAND2_X1 ref_1_maj_89_U13 ( .A1(ref_1_maj_89_n18), .A2(ref_1_maj_89_n17), 
        .ZN(ref_1_maj_89_n19) );
  NAND2_X1 ref_1_maj_89_U12 ( .A1(ref_1_n6), .A2(ref_1_maj_89_n16), .ZN(
        ref_1_maj_89_n14) );
  NAND2_X1 ref_1_maj_89_U11 ( .A1(ref_1_n2), .A2(ref_1_n3), .ZN(
        ref_1_maj_89_n15) );
  NAND2_X1 ref_1_maj_89_U10 ( .A1(ref_1_maj_89_n15), .A2(ref_1_maj_89_n14), 
        .ZN(ref_1_maj_89_n20) );
  XOR2_X1 ref_1_maj_89_U9 ( .A(ref_1_n6), .B(ref_1_maj_89_n16), .Z(
        ref_1_maj_89_n21) );
  XOR2_X1 ref_1_maj_89_U8 ( .A(ref_1_n8), .B(ref_1_n10), .Z(ref_1_maj_89_n22)
         );
  XOR2_X1 ref_1_maj_89_U7 ( .A(ref_1_n2), .B(ref_1_n3), .Z(ref_1_maj_89_n16)
         );
  OR2_X1 ref_1_maj_89_U6 ( .A1(ref_1_maj_89_n20), .A2(ref_1_maj_89_n19), .ZN(
        ref_1_maj_89_n24) );
  NAND2_X1 ref_1_maj_89_U5 ( .A1(ref_1_maj_89_n24), .A2(ref_1_maj_89_n23), 
        .ZN(ref_1_maj_89_n25) );
  NAND2_X1 ref_1_maj_89_U4 ( .A1(ref_1_maj_89_n20), .A2(ref_1_maj_89_n19), 
        .ZN(ref_1_maj_89_n26) );
  NAND2_X1 ref_1_maj_89_U3 ( .A1(ref_1_maj_89_n26), .A2(ref_1_maj_89_n25), 
        .ZN(ref_1_maj_89_port_o) );
  XOR2_X1 ref_1_maj_89_U2 ( .A(ref_1_maj_89_n22), .B(ref_1_maj_89_n21), .Z(
        ref_1_maj_89_n23) );
  XOR2_X1 simpleXor_120_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_120_port_a0), 
        .Z(simpleXor_120_port_z) );
  XOR2_X1 simpleXor_121_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_120_port_z), 
        .Z(simpleXor_121_port_z) );
  XOR2_X1 simpleXor_122_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_122_port_a0), 
        .Z(simpleXor_122_port_z) );
  XOR2_X1 simpleXor_123_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_122_port_z), 
        .Z(simpleXor_123_port_z) );
  XOR2_X1 simpleXor_124_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_124_port_a0), 
        .Z(simpleXor_124_port_z) );
  XOR2_X1 simpleXor_125_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_124_port_z), 
        .Z(simpleXor_125_port_z) );
  XOR2_X1 simpleXor_126_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_126_port_a0), 
        .Z(simpleXor_126_port_z) );
  XOR2_X1 simpleXor_127_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_126_port_z), 
        .Z(simpleXor_127_port_z) );
  XOR2_X1 simpleXor_128_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_128_port_a0), 
        .Z(simpleXor_128_port_z) );
  XOR2_X1 simpleXor_129_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_128_port_z), 
        .Z(simpleXor_129_port_z) );
  XOR2_X1 simpleXor_130_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_130_port_a0), 
        .Z(simpleXor_130_port_z) );
  XOR2_X1 simpleXor_131_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_130_port_z), 
        .Z(simpleXor_131_port_z) );
  XOR2_X1 simpleXor_132_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_132_port_a0), 
        .Z(simpleXor_132_port_z) );
  XOR2_X1 simpleXor_133_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_132_port_z), 
        .Z(simpleXor_133_port_z) );
  XOR2_X1 simpleXor_134_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_134_port_a0), 
        .Z(simpleXor_134_port_z) );
  XOR2_X1 simpleXor_135_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_134_port_z), 
        .Z(simpleXor_135_port_z) );
  XOR2_X1 simpleXor_136_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_136_port_a0), 
        .Z(simpleXor_136_port_z) );
  XOR2_X1 simpleXor_137_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_136_port_z), 
        .Z(simpleXor_137_port_z) );
  XOR2_X1 simpleXor_138_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_138_port_a0), 
        .Z(simpleXor_138_port_z) );
  XOR2_X1 simpleXor_139_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_138_port_z), 
        .Z(simpleXor_139_port_z) );
  XOR2_X1 simpleXor_140_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_140_port_a0), 
        .Z(simpleXor_140_port_z) );
  XOR2_X1 simpleXor_141_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_140_port_z), 
        .Z(simpleXor_141_port_z) );
  XOR2_X1 simpleXor_142_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_142_port_a0), 
        .Z(simpleXor_142_port_z) );
  XOR2_X1 simpleXor_143_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_142_port_z), 
        .Z(simpleXor_143_port_z) );
  XOR2_X1 simpleXor_144_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_144_port_a0), 
        .Z(simpleXor_144_port_z) );
  XOR2_X1 simpleXor_145_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_144_port_z), 
        .Z(simpleXor_145_port_z) );
  XOR2_X1 simpleXor_146_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_146_port_a0), 
        .Z(simpleXor_146_port_z) );
  XOR2_X1 simpleXor_147_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_146_port_z), 
        .Z(simpleXor_147_port_z) );
  XOR2_X1 simpleXor_148_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_148_port_a0), 
        .Z(simpleXor_148_port_z) );
  XOR2_X1 simpleXor_149_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_148_port_z), 
        .Z(simpleXor_149_port_z) );
  XOR2_X1 simpleXor_150_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_150_port_a0), 
        .Z(simpleXor_150_port_z) );
  XOR2_X1 simpleXor_151_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_150_port_z), 
        .Z(simpleXor_151_port_z) );
  XOR2_X1 simpleXor_152_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_152_port_a0), 
        .Z(simpleXor_152_port_z) );
  XOR2_X1 simpleXor_153_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_152_port_z), 
        .Z(simpleXor_153_port_z) );
  XOR2_X1 simpleXor_154_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_154_port_a0), 
        .Z(simpleXor_154_port_z) );
  XOR2_X1 simpleXor_155_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_154_port_z), 
        .Z(simpleXor_155_port_z) );
  XOR2_X1 simpleXor_156_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_156_port_a0), 
        .Z(simpleXor_156_port_z) );
  XOR2_X1 simpleXor_157_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_156_port_z), 
        .Z(simpleXor_157_port_z) );
  XOR2_X1 simpleXor_158_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_158_port_a0), 
        .Z(simpleXor_158_port_z) );
  XOR2_X1 simpleXor_159_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_158_port_z), 
        .Z(simpleXor_159_port_z) );
  XOR2_X1 simpleXor_160_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_160_port_a0), 
        .Z(simpleXor_160_port_z) );
  XOR2_X1 simpleXor_161_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_160_port_z), 
        .Z(simpleXor_161_port_z) );
  XOR2_X1 simpleXor_162_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_162_port_a0), 
        .Z(simpleXor_162_port_z) );
  XOR2_X1 simpleXor_163_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_162_port_z), 
        .Z(simpleXor_163_port_z) );
  XOR2_X1 simpleXor_164_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_164_port_a0), 
        .Z(simpleXor_164_port_z) );
  XOR2_X1 simpleXor_165_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_164_port_z), 
        .Z(simpleXor_165_port_z) );
  XOR2_X1 simpleXor_166_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_166_port_a0), 
        .Z(simpleXor_166_port_z) );
  XOR2_X1 simpleXor_167_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_166_port_z), 
        .Z(simpleXor_167_port_z) );
  XOR2_X1 simpleXor_168_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_168_port_a0), 
        .Z(simpleXor_168_port_z) );
  XOR2_X1 simpleXor_169_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_168_port_z), 
        .Z(simpleXor_169_port_z) );
  XOR2_X1 simpleXor_170_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_170_port_a0), 
        .Z(simpleXor_170_port_z) );
  XOR2_X1 simpleXor_171_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_170_port_z), 
        .Z(simpleXor_171_port_z) );
  XOR2_X1 simpleXor_172_U1 ( .A(port_rand_mul_0[0]), .B(simpleXor_172_port_a0), 
        .Z(simpleXor_172_port_z) );
  XOR2_X1 simpleXor_173_U1 ( .A(port_rand_mul_0[1]), .B(simpleXor_172_port_z), 
        .Z(simpleXor_173_port_z) );
  XOR2_X1 simpleXor_174_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_174_port_a0), 
        .Z(simpleXor_174_port_z) );
  XOR2_X1 simpleXor_175_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_174_port_z), 
        .Z(simpleXor_175_port_z) );
  XOR2_X1 simpleXor_176_U1 ( .A(port_rand_mul_1[0]), .B(simpleXor_176_port_a0), 
        .Z(simpleXor_176_port_z) );
  XOR2_X1 simpleXor_177_U1 ( .A(port_rand_mul_1[1]), .B(simpleXor_176_port_z), 
        .Z(simpleXor_177_port_z) );
  XOR2_X1 simpleXor_178_U1 ( .A(port_rand_mul_2[0]), .B(simpleXor_178_port_a0), 
        .Z(simpleXor_178_port_z) );
  XOR2_X1 simpleXor_179_U1 ( .A(port_rand_mul_2[1]), .B(simpleXor_178_port_z), 
        .Z(simpleXor_179_port_z) );
endmodule

