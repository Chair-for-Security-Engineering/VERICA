
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i0_s5, io_i0_s6, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, 
        io_i1_s4, io_i1_s5, io_i1_s6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, 
        p_rand_4, p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, 
        p_rand_11, p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16, 
        p_rand_17, p_rand_18, p_rand_19, p_rand_20, io_o0_s0, io_o0_s1, 
        io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5, io_o0_s6 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i0_s5, io_i0_s6, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4,
         io_i1_s5, io_i1_s6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4,
         p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10,
         p_rand_11, p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16,
         p_rand_17, p_rand_18, p_rand_19, p_rand_20;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5, io_o0_s6;
  wire   n_dom_0_n105, n_dom_0_n104, n_dom_0_n103, n_dom_0_n102, n_dom_0_n101,
         n_dom_0_n100, n_dom_0_n99, n_dom_0_n98, n_dom_0_n97, n_dom_0_n96,
         n_dom_0_n95, n_dom_0_n94, n_dom_0_n93, n_dom_0_n92, n_dom_0_n91,
         n_dom_0_n90, n_dom_0_n89, n_dom_0_n88, n_dom_0_n87, n_dom_0_n86,
         n_dom_0_n85, n_dom_0_n84, n_dom_0_n83, n_dom_0_n82, n_dom_0_n81,
         n_dom_0_n80, n_dom_0_n79, n_dom_0_n78, n_dom_0_n77, n_dom_0_n76,
         n_dom_0_n75, n_dom_0_n74, n_dom_0_n73, n_dom_0_n72, n_dom_0_n71,
         n_dom_0_n70, n_dom_0_n69, n_dom_0_n68, n_dom_0_n67, n_dom_0_n66,
         n_dom_0_n65, n_dom_0_n64, n_dom_0_n63, n_dom_0_n62, n_dom_0_n61,
         n_dom_0_n60, n_dom_0_n59, n_dom_0_n58, n_dom_0_n57, n_dom_0_n56,
         n_dom_0_n55, n_dom_0_n54, n_dom_0_n53, n_dom_0_n52, n_dom_0_n51,
         n_dom_0_n50, n_dom_0_n49, n_dom_0_n48, n_dom_0_n47, n_dom_0_n46,
         n_dom_0_n45, n_dom_0_n44, n_dom_0_n43, n_dom_0_n42, n_dom_0_n41,
         n_dom_0_n40, n_dom_0_n39, n_dom_0_n38, n_dom_0_n37, n_dom_0_n36,
         n_dom_0_n35, n_dom_0_n34, n_dom_0_n33, n_dom_0_n32, n_dom_0_n31,
         n_dom_0_n30, n_dom_0_n29, n_dom_0_n28, n_dom_0_n27, n_dom_0_n26,
         n_dom_0_n25, n_dom_0_n24, n_dom_0_n23, n_dom_0_n22, n_dom_0_n21,
         n_dom_0_n20, n_dom_0_n19, n_dom_0_n18, n_dom_0_n17, n_dom_0_n16,
         n_dom_0_n15, n_dom_0_n14, n_dom_0_n13, n_dom_0_n12, n_dom_0_n11,
         n_dom_0_n10, n_dom_0_n9, n_dom_0_n8, n_dom_0_n7, n_dom_0_n6,
         n_dom_0_n5, n_dom_0_n4, n_dom_0_n3, n_dom_0_n2, n_dom_0_n1,
         n_dom_0_N55, n_dom_0_N54, n_dom_0_N53, n_dom_0_N52, n_dom_0_N51,
         n_dom_0_N50, n_dom_0_N49, n_dom_0_N48, n_dom_0__dom_inter6_2,
         n_dom_0__dom_inter6_1, n_dom_0_reg_pipeline, n_dom_0_N47,
         n_dom_0__dom_inter5_7, n_dom_0__dom_inter5_6, n_dom_0_reg_pipeline_5,
         n_dom_0_N46, n_dom_0__dom_inter4_14, n_dom_0__dom_inter4_13,
         n_dom_0_reg_pipeline_11, n_dom_0_N45, n_dom_0__dom_inter3_20,
         n_dom_0__dom_inter3_19, n_dom_0_reg_pipeline_17, n_dom_0_N44,
         n_dom_0__dom_inter2_26, n_dom_0__dom_inter2_25,
         n_dom_0_reg_pipeline_23, n_dom_0_N43, n_dom_0__dom_inter1_32,
         n_dom_0__dom_inter1_31, n_dom_0_reg_pipeline_29, n_dom_0_N42,
         n_dom_0__dom_inter0_38, n_dom_0__dom_inter0_37,
         n_dom_0_reg_pipeline_35, n_dom_0_N41, n_dom_0_N40, n_dom_0_N39,
         n_dom_0_N38, n_dom_0_N37, n_dom_0_N36, n_dom_0_N35, n_dom_0_N34,
         n_dom_0_N33, n_dom_0_N32, n_dom_0_N31, n_dom_0_N30, n_dom_0_N29,
         n_dom_0_N28, n_dom_0_N27, n_dom_0_N26, n_dom_0_N25, n_dom_0_N24,
         n_dom_0_N23, n_dom_0_N22, n_dom_0_N21, n_dom_0_N20, n_dom_0_N19,
         n_dom_0_N18, n_dom_0_N17, n_dom_0_N16, n_dom_0_N15, n_dom_0_N14,
         n_dom_0_N13, n_dom_0_N12, n_dom_0_N11, n_dom_0_N10, n_dom_0_N9,
         n_dom_0_N8, n_dom_0_N7, n_dom_0_N6, n_dom_0_N5, n_dom_0_N4,
         n_dom_0_N3, n_dom_0_N2, n_dom_0_N1, n_dom_0_N0;

  NAND2_X1 u_dom_0_U135 ( .A1(io_i0_s0), .A2(io_i1_s6), .ZN(n_dom_0_n77) );
  XNOR2_X1 u_dom_0_U134 ( .A(p_rand_5), .B(n_dom_0_n77), .ZN(n_dom_0_N0) );
  NAND2_X1 u_dom_0_U133 ( .A1(io_i0_s0), .A2(io_i1_s5), .ZN(n_dom_0_n76) );
  XNOR2_X1 u_dom_0_U132 ( .A(p_rand_4), .B(n_dom_0_n76), .ZN(n_dom_0_N1) );
  NAND2_X1 u_dom_0_U131 ( .A1(io_i1_s2), .A2(io_i0_s1), .ZN(n_dom_0_n75) );
  XNOR2_X1 u_dom_0_U130 ( .A(p_rand_6), .B(n_dom_0_n75), .ZN(n_dom_0_N10) );
  NAND2_X1 u_dom_0_U129 ( .A1(io_i1_s0), .A2(io_i0_s1), .ZN(n_dom_0_n74) );
  XNOR2_X1 u_dom_0_U128 ( .A(p_rand_0), .B(n_dom_0_n74), .ZN(n_dom_0_N11) );
  NAND2_X1 u_dom_0_U127 ( .A1(io_i0_s2), .A2(io_i1_s6), .ZN(n_dom_0_n73) );
  XNOR2_X1 u_dom_0_U126 ( .A(p_rand_14), .B(n_dom_0_n73), .ZN(n_dom_0_N12) );
  NAND2_X1 u_dom_0_U125 ( .A1(io_i0_s2), .A2(io_i1_s5), .ZN(n_dom_0_n72) );
  XNOR2_X1 u_dom_0_U124 ( .A(p_rand_13), .B(n_dom_0_n72), .ZN(n_dom_0_N13) );
  NAND2_X1 u_dom_0_U123 ( .A1(io_i0_s2), .A2(io_i1_s4), .ZN(n_dom_0_n71) );
  XNOR2_X1 u_dom_0_U122 ( .A(p_rand_12), .B(n_dom_0_n71), .ZN(n_dom_0_N14) );
  NAND2_X1 u_dom_0_U121 ( .A1(io_i0_s2), .A2(io_i1_s3), .ZN(n_dom_0_n70) );
  XNOR2_X1 u_dom_0_U120 ( .A(p_rand_11), .B(n_dom_0_n70), .ZN(n_dom_0_N15) );
  NAND2_X1 u_dom_0_U119 ( .A1(io_i0_s2), .A2(io_i1_s1), .ZN(n_dom_0_n69) );
  XNOR2_X1 u_dom_0_U118 ( .A(p_rand_6), .B(n_dom_0_n69), .ZN(n_dom_0_N16) );
  NAND2_X1 u_dom_0_U117 ( .A1(io_i0_s2), .A2(io_i1_s0), .ZN(n_dom_0_n68) );
  XNOR2_X1 u_dom_0_U116 ( .A(p_rand_1), .B(n_dom_0_n68), .ZN(n_dom_0_N17) );
  NAND2_X1 u_dom_0_U115 ( .A1(io_i0_s3), .A2(io_i1_s6), .ZN(n_dom_0_n67) );
  XNOR2_X1 u_dom_0_U114 ( .A(p_rand_17), .B(n_dom_0_n67), .ZN(n_dom_0_N18) );
  NAND2_X1 u_dom_0_U113 ( .A1(io_i0_s3), .A2(io_i1_s5), .ZN(n_dom_0_n66) );
  XNOR2_X1 u_dom_0_U112 ( .A(p_rand_16), .B(n_dom_0_n66), .ZN(n_dom_0_N19) );
  NAND2_X1 u_dom_0_U111 ( .A1(io_i0_s0), .A2(io_i1_s4), .ZN(n_dom_0_n65) );
  XNOR2_X1 u_dom_0_U110 ( .A(p_rand_3), .B(n_dom_0_n65), .ZN(n_dom_0_N2) );
  NAND2_X1 u_dom_0_U109 ( .A1(io_i0_s3), .A2(io_i1_s4), .ZN(n_dom_0_n64) );
  XNOR2_X1 u_dom_0_U108 ( .A(p_rand_15), .B(n_dom_0_n64), .ZN(n_dom_0_N20) );
  NAND2_X1 u_dom_0_U107 ( .A1(io_i0_s3), .A2(io_i1_s2), .ZN(n_dom_0_n63) );
  XNOR2_X1 u_dom_0_U106 ( .A(p_rand_11), .B(n_dom_0_n63), .ZN(n_dom_0_N21) );
  NAND2_X1 u_dom_0_U105 ( .A1(io_i0_s3), .A2(io_i1_s1), .ZN(n_dom_0_n62) );
  XNOR2_X1 u_dom_0_U104 ( .A(p_rand_7), .B(n_dom_0_n62), .ZN(n_dom_0_N22) );
  NAND2_X1 u_dom_0_U103 ( .A1(io_i0_s3), .A2(io_i1_s0), .ZN(n_dom_0_n61) );
  XNOR2_X1 u_dom_0_U102 ( .A(p_rand_2), .B(n_dom_0_n61), .ZN(n_dom_0_N23) );
  NAND2_X1 u_dom_0_U101 ( .A1(io_i0_s4), .A2(io_i1_s6), .ZN(n_dom_0_n60) );
  XNOR2_X1 u_dom_0_U100 ( .A(p_rand_19), .B(n_dom_0_n60), .ZN(n_dom_0_N24) );
  NAND2_X1 u_dom_0_U99 ( .A1(io_i0_s4), .A2(io_i1_s5), .ZN(n_dom_0_n59) );
  XNOR2_X1 u_dom_0_U98 ( .A(p_rand_18), .B(n_dom_0_n59), .ZN(n_dom_0_N25) );
  NAND2_X1 u_dom_0_U97 ( .A1(io_i0_s4), .A2(io_i1_s3), .ZN(n_dom_0_n58) );
  XNOR2_X1 u_dom_0_U96 ( .A(p_rand_15), .B(n_dom_0_n58), .ZN(n_dom_0_N26) );
  NAND2_X1 u_dom_0_U95 ( .A1(io_i0_s4), .A2(io_i1_s2), .ZN(n_dom_0_n57) );
  XNOR2_X1 u_dom_0_U94 ( .A(p_rand_12), .B(n_dom_0_n57), .ZN(n_dom_0_N27) );
  NAND2_X1 u_dom_0_U93 ( .A1(io_i0_s4), .A2(io_i1_s1), .ZN(n_dom_0_n56) );
  XNOR2_X1 u_dom_0_U92 ( .A(p_rand_8), .B(n_dom_0_n56), .ZN(n_dom_0_N28) );
  NAND2_X1 u_dom_0_U91 ( .A1(io_i0_s4), .A2(io_i1_s0), .ZN(n_dom_0_n55) );
  XNOR2_X1 u_dom_0_U90 ( .A(p_rand_3), .B(n_dom_0_n55), .ZN(n_dom_0_N29) );
  NAND2_X1 u_dom_0_U89 ( .A1(io_i0_s0), .A2(io_i1_s3), .ZN(n_dom_0_n54) );
  XNOR2_X1 u_dom_0_U88 ( .A(p_rand_2), .B(n_dom_0_n54), .ZN(n_dom_0_N3) );
  NAND2_X1 u_dom_0_U87 ( .A1(io_i0_s5), .A2(io_i1_s6), .ZN(n_dom_0_n53) );
  XNOR2_X1 u_dom_0_U86 ( .A(p_rand_20), .B(n_dom_0_n53), .ZN(n_dom_0_N30) );
  NAND2_X1 u_dom_0_U85 ( .A1(io_i1_s0), .A2(io_i0_s5), .ZN(n_dom_0_n52) );
  XNOR2_X1 u_dom_0_U84 ( .A(p_rand_4), .B(n_dom_0_n52), .ZN(n_dom_0_N31) );
  NAND2_X1 u_dom_0_U83 ( .A1(io_i0_s5), .A2(io_i1_s4), .ZN(n_dom_0_n51) );
  XNOR2_X1 u_dom_0_U82 ( .A(p_rand_18), .B(n_dom_0_n51), .ZN(n_dom_0_N32) );
  NAND2_X1 u_dom_0_U81 ( .A1(io_i0_s5), .A2(io_i1_s3), .ZN(n_dom_0_n50) );
  XNOR2_X1 u_dom_0_U80 ( .A(p_rand_16), .B(n_dom_0_n50), .ZN(n_dom_0_N33) );
  NAND2_X1 u_dom_0_U79 ( .A1(io_i1_s2), .A2(io_i0_s5), .ZN(n_dom_0_n49) );
  XNOR2_X1 u_dom_0_U78 ( .A(p_rand_13), .B(n_dom_0_n49), .ZN(n_dom_0_N34) );
  NAND2_X1 u_dom_0_U77 ( .A1(io_i1_s1), .A2(io_i0_s5), .ZN(n_dom_0_n48) );
  XNOR2_X1 u_dom_0_U76 ( .A(p_rand_9), .B(n_dom_0_n48), .ZN(n_dom_0_N35) );
  NAND2_X1 u_dom_0_U75 ( .A1(io_i0_s6), .A2(io_i1_s5), .ZN(n_dom_0_n47) );
  XNOR2_X1 u_dom_0_U74 ( .A(p_rand_20), .B(n_dom_0_n47), .ZN(n_dom_0_N36) );
  NAND2_X1 u_dom_0_U73 ( .A1(io_i0_s6), .A2(io_i1_s4), .ZN(n_dom_0_n46) );
  XNOR2_X1 u_dom_0_U72 ( .A(p_rand_19), .B(n_dom_0_n46), .ZN(n_dom_0_N37) );
  NAND2_X1 u_dom_0_U71 ( .A1(io_i0_s6), .A2(io_i1_s3), .ZN(n_dom_0_n45) );
  XNOR2_X1 u_dom_0_U70 ( .A(p_rand_17), .B(n_dom_0_n45), .ZN(n_dom_0_N38) );
  NAND2_X1 u_dom_0_U69 ( .A1(io_i0_s6), .A2(io_i1_s2), .ZN(n_dom_0_n44) );
  XNOR2_X1 u_dom_0_U68 ( .A(p_rand_14), .B(n_dom_0_n44), .ZN(n_dom_0_N39) );
  NAND2_X1 u_dom_0_U67 ( .A1(io_i1_s2), .A2(io_i0_s0), .ZN(n_dom_0_n43) );
  XNOR2_X1 u_dom_0_U66 ( .A(p_rand_1), .B(n_dom_0_n43), .ZN(n_dom_0_N4) );
  NAND2_X1 u_dom_0_U65 ( .A1(io_i0_s6), .A2(io_i1_s1), .ZN(n_dom_0_n42) );
  XNOR2_X1 u_dom_0_U64 ( .A(p_rand_10), .B(n_dom_0_n42), .ZN(n_dom_0_N40) );
  NAND2_X1 u_dom_0_U63 ( .A1(io_i0_s6), .A2(io_i1_s0), .ZN(n_dom_0_n41) );
  XNOR2_X1 u_dom_0_U62 ( .A(p_rand_5), .B(n_dom_0_n41), .ZN(n_dom_0_N41) );
  XOR2_X1 u_dom_0_U61 ( .A(n_dom_0__dom_inter0_37), .B(n_dom_0_n103), .Z(
        n_dom_0_n39) );
  XOR2_X1 u_dom_0_U60 ( .A(n_dom_0_reg_pipeline_35), .B(n_dom_0_n102), .Z(
        n_dom_0_n40) );
  XOR2_X1 u_dom_0_U59 ( .A(n_dom_0_n39), .B(n_dom_0_n40), .Z(n_dom_0_n36) );
  XOR2_X1 u_dom_0_U58 ( .A(n_dom_0__dom_inter0_38), .B(n_dom_0_n104), .Z(
        n_dom_0_n38) );
  XOR2_X1 u_dom_0_U57 ( .A(n_dom_0_n38), .B(n_dom_0_n105), .Z(n_dom_0_n37) );
  XOR2_X1 u_dom_0_U56 ( .A(n_dom_0_n36), .B(n_dom_0_n37), .Z(n_dom_0_N42) );
  XOR2_X1 u_dom_0_U55 ( .A(n_dom_0__dom_inter1_31), .B(n_dom_0_n99), .Z(
        n_dom_0_n34) );
  XOR2_X1 u_dom_0_U54 ( .A(n_dom_0_reg_pipeline_29), .B(n_dom_0_n98), .Z(
        n_dom_0_n35) );
  XOR2_X1 u_dom_0_U53 ( .A(n_dom_0_n34), .B(n_dom_0_n35), .Z(n_dom_0_n31) );
  XOR2_X1 u_dom_0_U52 ( .A(n_dom_0__dom_inter1_32), .B(n_dom_0_n100), .Z(
        n_dom_0_n33) );
  XOR2_X1 u_dom_0_U51 ( .A(n_dom_0_n33), .B(n_dom_0_n101), .Z(n_dom_0_n32) );
  XOR2_X1 u_dom_0_U50 ( .A(n_dom_0_n31), .B(n_dom_0_n32), .Z(n_dom_0_N43) );
  XOR2_X1 u_dom_0_U49 ( .A(n_dom_0__dom_inter2_25), .B(n_dom_0_n95), .Z(
        n_dom_0_n29) );
  XOR2_X1 u_dom_0_U48 ( .A(n_dom_0_reg_pipeline_23), .B(n_dom_0_n94), .Z(
        n_dom_0_n30) );
  XOR2_X1 u_dom_0_U47 ( .A(n_dom_0_n29), .B(n_dom_0_n30), .Z(n_dom_0_n26) );
  XOR2_X1 u_dom_0_U46 ( .A(n_dom_0__dom_inter2_26), .B(n_dom_0_n96), .Z(
        n_dom_0_n28) );
  XOR2_X1 u_dom_0_U45 ( .A(n_dom_0_n28), .B(n_dom_0_n97), .Z(n_dom_0_n27) );
  XOR2_X1 u_dom_0_U44 ( .A(n_dom_0_n26), .B(n_dom_0_n27), .Z(n_dom_0_N44) );
  XOR2_X1 u_dom_0_U43 ( .A(n_dom_0__dom_inter3_19), .B(n_dom_0_n91), .Z(
        n_dom_0_n24) );
  XOR2_X1 u_dom_0_U42 ( .A(n_dom_0_reg_pipeline_17), .B(n_dom_0_n90), .Z(
        n_dom_0_n25) );
  XOR2_X1 u_dom_0_U41 ( .A(n_dom_0_n24), .B(n_dom_0_n25), .Z(n_dom_0_n21) );
  XOR2_X1 u_dom_0_U40 ( .A(n_dom_0__dom_inter3_20), .B(n_dom_0_n92), .Z(
        n_dom_0_n23) );
  XOR2_X1 u_dom_0_U39 ( .A(n_dom_0_n23), .B(n_dom_0_n93), .Z(n_dom_0_n22) );
  XOR2_X1 u_dom_0_U38 ( .A(n_dom_0_n21), .B(n_dom_0_n22), .Z(n_dom_0_N45) );
  XOR2_X1 u_dom_0_U37 ( .A(n_dom_0__dom_inter4_13), .B(n_dom_0_n87), .Z(
        n_dom_0_n19) );
  XOR2_X1 u_dom_0_U36 ( .A(n_dom_0_reg_pipeline_11), .B(n_dom_0_n86), .Z(
        n_dom_0_n20) );
  XOR2_X1 u_dom_0_U35 ( .A(n_dom_0_n19), .B(n_dom_0_n20), .Z(n_dom_0_n16) );
  XOR2_X1 u_dom_0_U34 ( .A(n_dom_0__dom_inter4_14), .B(n_dom_0_n88), .Z(
        n_dom_0_n18) );
  XOR2_X1 u_dom_0_U33 ( .A(n_dom_0_n18), .B(n_dom_0_n89), .Z(n_dom_0_n17) );
  XOR2_X1 u_dom_0_U32 ( .A(n_dom_0_n16), .B(n_dom_0_n17), .Z(n_dom_0_N46) );
  XOR2_X1 u_dom_0_U31 ( .A(n_dom_0__dom_inter5_6), .B(n_dom_0_n83), .Z(
        n_dom_0_n14) );
  XOR2_X1 u_dom_0_U30 ( .A(n_dom_0_reg_pipeline_5), .B(n_dom_0_n82), .Z(
        n_dom_0_n15) );
  XOR2_X1 u_dom_0_U29 ( .A(n_dom_0_n14), .B(n_dom_0_n15), .Z(n_dom_0_n11) );
  XOR2_X1 u_dom_0_U28 ( .A(n_dom_0__dom_inter5_7), .B(n_dom_0_n84), .Z(
        n_dom_0_n13) );
  XOR2_X1 u_dom_0_U27 ( .A(n_dom_0_n13), .B(n_dom_0_n85), .Z(n_dom_0_n12) );
  XOR2_X1 u_dom_0_U26 ( .A(n_dom_0_n11), .B(n_dom_0_n12), .Z(n_dom_0_N47) );
  XOR2_X1 u_dom_0_U25 ( .A(n_dom_0__dom_inter6_1), .B(n_dom_0_n79), .Z(
        n_dom_0_n9) );
  XOR2_X1 u_dom_0_U24 ( .A(n_dom_0_reg_pipeline), .B(n_dom_0_n78), .Z(
        n_dom_0_n10) );
  XOR2_X1 u_dom_0_U23 ( .A(n_dom_0_n9), .B(n_dom_0_n10), .Z(n_dom_0_n6) );
  XOR2_X1 u_dom_0_U22 ( .A(n_dom_0__dom_inter6_2), .B(n_dom_0_n80), .Z(
        n_dom_0_n8) );
  XOR2_X1 u_dom_0_U21 ( .A(n_dom_0_n8), .B(n_dom_0_n81), .Z(n_dom_0_n7) );
  XOR2_X1 u_dom_0_U20 ( .A(n_dom_0_n6), .B(n_dom_0_n7), .Z(n_dom_0_N48) );
  AND2_X1 u_dom_0_U19 ( .A1(io_i1_s6), .A2(io_i0_s6), .ZN(n_dom_0_N49) );
  NAND2_X1 u_dom_0_U18 ( .A1(io_i1_s1), .A2(io_i0_s0), .ZN(n_dom_0_n5) );
  XNOR2_X1 u_dom_0_U17 ( .A(p_rand_0), .B(n_dom_0_n5), .ZN(n_dom_0_N5) );
  AND2_X1 u_dom_0_U16 ( .A1(io_i1_s4), .A2(io_i0_s4), .ZN(n_dom_0_N50) );
  AND2_X1 u_dom_0_U15 ( .A1(io_i1_s3), .A2(io_i0_s3), .ZN(n_dom_0_N51) );
  AND2_X1 u_dom_0_U14 ( .A1(io_i0_s2), .A2(io_i1_s2), .ZN(n_dom_0_N52) );
  AND2_X1 u_dom_0_U13 ( .A1(io_i0_s1), .A2(io_i1_s1), .ZN(n_dom_0_N53) );
  AND2_X1 u_dom_0_U12 ( .A1(io_i0_s0), .A2(io_i1_s0), .ZN(n_dom_0_N54) );
  AND2_X1 u_dom_0_U11 ( .A1(io_i1_s5), .A2(io_i0_s5), .ZN(n_dom_0_N55) );
  NAND2_X1 u_dom_0_U10 ( .A1(io_i1_s6), .A2(io_i0_s1), .ZN(n_dom_0_n4) );
  XNOR2_X1 u_dom_0_U9 ( .A(p_rand_10), .B(n_dom_0_n4), .ZN(n_dom_0_N6) );
  NAND2_X1 u_dom_0_U8 ( .A1(io_i1_s5), .A2(io_i0_s1), .ZN(n_dom_0_n3) );
  XNOR2_X1 u_dom_0_U7 ( .A(p_rand_9), .B(n_dom_0_n3), .ZN(n_dom_0_N7) );
  NAND2_X1 u_dom_0_U6 ( .A1(io_i1_s4), .A2(io_i0_s1), .ZN(n_dom_0_n2) );
  XNOR2_X1 u_dom_0_U5 ( .A(p_rand_8), .B(n_dom_0_n2), .ZN(n_dom_0_N8) );
  NAND2_X1 u_dom_0_U4 ( .A1(io_i1_s3), .A2(io_i0_s1), .ZN(n_dom_0_n1) );
  XNOR2_X1 u_dom_0_U3 ( .A(p_rand_7), .B(n_dom_0_n1), .ZN(n_dom_0_N9) );
  DFF_X1 u_dom_0_dom_out5_reg ( .D(n_dom_0_N47), .CK(clock_0), .Q(io_o0_s5), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter5_10_reg ( .D(n_dom_0_N31), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n83) );
  DFF_X1 u_dom_0_dom_out4_reg ( .D(n_dom_0_N46), .CK(clock_0), .Q(io_o0_s4), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter4_14_reg ( .D(n_dom_0_N27), .CK(clock_0), .Q(
        n_dom_0__dom_inter4_14), .QN() );
  DFF_X1 u_dom_0_dom_out0_reg ( .D(n_dom_0_N42), .CK(clock_0), .Q(io_o0_s0), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter0_37_reg ( .D(n_dom_0_N2), .CK(clock_0), .Q(
        n_dom_0__dom_inter0_37), .QN() );
  DFF_X1 u_dom_0__dom_inter5_6_reg ( .D(n_dom_0_N32), .CK(clock_0), .Q(
        n_dom_0__dom_inter5_6), .QN() );
  DFF_X1 u_dom_0__dom_inter5_7_reg ( .D(n_dom_0_N33), .CK(clock_0), .Q(
        n_dom_0__dom_inter5_7), .QN() );
  DFF_X1 u_dom_0__dom_inter5_8_reg ( .D(n_dom_0_N34), .CK(clock_0), .Q(), .QN(
        n_dom_0_n85) );
  DFF_X1 u_dom_0__dom_inter5_9_reg ( .D(n_dom_0_N35), .CK(clock_0), .Q(), .QN(
        n_dom_0_n84) );
  DFF_X1 u_dom_0__dom_inter0_reg ( .D(n_dom_0_N0), .CK(clock_0), .Q(), .QN(
        n_dom_0_n102) );
  DFF_X1 u_dom_0_dom_out6_reg ( .D(n_dom_0_N48), .CK(clock_0), .Q(io_o0_s6), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter6_reg ( .D(n_dom_0_N36), .CK(clock_0), .Q(), .QN(
        n_dom_0_n78) );
  DFF_X1 u_dom_0__dom_inter4_12_reg ( .D(n_dom_0_N25), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n87) );
  DFF_X1 u_dom_0__dom_inter6_0_reg ( .D(n_dom_0_N37), .CK(clock_0), .Q(), .QN(
        n_dom_0_n79) );
  DFF_X1 u_dom_0__dom_inter4_15_reg ( .D(n_dom_0_N28), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n89) );
  DFF_X1 u_dom_0__dom_inter0_39_reg ( .D(n_dom_0_N4), .CK(clock_0), .Q(), .QN(
        n_dom_0_n105) );
  DFF_X1 u_dom_0__dom_inter6_1_reg ( .D(n_dom_0_N38), .CK(clock_0), .Q(
        n_dom_0__dom_inter6_1), .QN() );
  DFF_X1 u_dom_0__dom_inter6_2_reg ( .D(n_dom_0_N39), .CK(clock_0), .Q(
        n_dom_0__dom_inter6_2), .QN() );
  DFF_X1 u_dom_0__dom_inter6_3_reg ( .D(n_dom_0_N40), .CK(clock_0), .Q(), .QN(
        n_dom_0_n81) );
  DFF_X1 u_dom_0_dom_out2_reg ( .D(n_dom_0_N44), .CK(clock_0), .Q(io_o0_s2), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter2_28_reg ( .D(n_dom_0_N17), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n96) );
  DFF_X1 u_dom_0__dom_inter6_4_reg ( .D(n_dom_0_N41), .CK(clock_0), .Q(), .QN(
        n_dom_0_n80) );
  DFF_X1 u_dom_0_dom_out3_reg ( .D(n_dom_0_N45), .CK(clock_0), .Q(io_o0_s3), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter3_19_reg ( .D(n_dom_0_N20), .CK(clock_0), .Q(
        n_dom_0__dom_inter3_19), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_5_reg ( .D(n_dom_0_N55), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_5), .QN() );
  DFF_X1 u_dom_0__dom_inter4_13_reg ( .D(n_dom_0_N26), .CK(clock_0), .Q(
        n_dom_0__dom_inter4_13), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_35_reg ( .D(n_dom_0_N54), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_35), .QN() );
  DFF_X1 u_dom_0__dom_inter4_16_reg ( .D(n_dom_0_N29), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n88) );
  DFF_X1 u_dom_0_dom_out1_reg ( .D(n_dom_0_N43), .CK(clock_0), .Q(io_o0_s1), 
        .QN() );
  DFF_X1 u_dom_0__dom_inter1_reg ( .D(n_dom_0_N6), .CK(clock_0), .Q(), .QN(
        n_dom_0_n98) );
  DFF_X1 u_dom_0_reg_pipeline_29_reg ( .D(n_dom_0_N53), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_29), .QN() );
  DFF_X1 u_dom_0__dom_inter1_33_reg ( .D(n_dom_0_N10), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n101) );
  DFF_X1 u_dom_0_reg_pipeline_23_reg ( .D(n_dom_0_N52), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_23), .QN() );
  DFF_X1 u_dom_0__dom_inter2_26_reg ( .D(n_dom_0_N15), .CK(clock_0), .Q(
        n_dom_0__dom_inter2_26), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_17_reg ( .D(n_dom_0_N51), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_17), .QN() );
  DFF_X1 u_dom_0__dom_inter3_reg ( .D(n_dom_0_N18), .CK(clock_0), .Q(), .QN(
        n_dom_0_n90) );
  DFF_X1 u_dom_0_reg_pipeline_11_reg ( .D(n_dom_0_N50), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline_11), .QN() );
  DFF_X1 u_dom_0__dom_inter3_20_reg ( .D(n_dom_0_N21), .CK(clock_0), .Q(
        n_dom_0__dom_inter3_20), .QN() );
  DFF_X1 u_dom_0_reg_pipeline_reg ( .D(n_dom_0_N49), .CK(clock_0), .Q(
        n_dom_0_reg_pipeline), .QN() );
  DFF_X1 u_dom_0__dom_inter2_reg ( .D(n_dom_0_N12), .CK(clock_0), .Q(), .QN(
        n_dom_0_n94) );
  DFF_X1 u_dom_0__dom_inter5_reg ( .D(n_dom_0_N30), .CK(clock_0), .Q(), .QN(
        n_dom_0_n82) );
  DFF_X1 u_dom_0__dom_inter1_31_reg ( .D(n_dom_0_N8), .CK(clock_0), .Q(
        n_dom_0__dom_inter1_31), .QN() );
  DFF_X1 u_dom_0__dom_inter2_25_reg ( .D(n_dom_0_N14), .CK(clock_0), .Q(
        n_dom_0__dom_inter2_25), .QN() );
  DFF_X1 u_dom_0__dom_inter1_32_reg ( .D(n_dom_0_N9), .CK(clock_0), .Q(
        n_dom_0__dom_inter1_32), .QN() );
  DFF_X1 u_dom_0__dom_inter2_27_reg ( .D(n_dom_0_N16), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n97) );
  DFF_X1 u_dom_0__dom_inter1_30_reg ( .D(n_dom_0_N7), .CK(clock_0), .Q(), .QN(
        n_dom_0_n99) );
  DFF_X1 u_dom_0__dom_inter3_18_reg ( .D(n_dom_0_N19), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n91) );
  DFF_X1 u_dom_0__dom_inter0_40_reg ( .D(n_dom_0_N5), .CK(clock_0), .Q(), .QN(
        n_dom_0_n104) );
  DFF_X1 u_dom_0__dom_inter3_21_reg ( .D(n_dom_0_N22), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n93) );
  DFF_X1 u_dom_0__dom_inter0_38_reg ( .D(n_dom_0_N3), .CK(clock_0), .Q(
        n_dom_0__dom_inter0_38), .QN() );
  DFF_X1 u_dom_0__dom_inter3_22_reg ( .D(n_dom_0_N23), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n92) );
  DFF_X1 u_dom_0__dom_inter2_24_reg ( .D(n_dom_0_N13), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n95) );
  DFF_X1 u_dom_0__dom_inter4_reg ( .D(n_dom_0_N24), .CK(clock_0), .Q(), .QN(
        n_dom_0_n86) );
  DFF_X1 u_dom_0__dom_inter0_36_reg ( .D(n_dom_0_N1), .CK(clock_0), .Q(), .QN(
        n_dom_0_n103) );
  DFF_X1 u_dom_0__dom_inter1_34_reg ( .D(n_dom_0_N11), .CK(clock_0), .Q(), 
        .QN(n_dom_0_n100) );
endmodule

