
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, p_rand_0, 
        p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7, 
        p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12, p_rand_13, 
        p_rand_14, p_rand_15, p_rand_16, p_rand_17, p_rand_18, p_rand_19, 
        io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, p_rand_0, p_rand_1,
         p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7, p_rand_8,
         p_rand_9, p_rand_10, p_rand_11, p_rand_12, p_rand_13, p_rand_14,
         p_rand_15, p_rand_16, p_rand_17, p_rand_18, p_rand_19;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4;
  wire   n_hpc2_0_n75, n_hpc2_0_n74, n_hpc2_0_n73, n_hpc2_0_n72, n_hpc2_0_n71,
         n_hpc2_0_n70, n_hpc2_0_n69, n_hpc2_0_n68, n_hpc2_0_n67, n_hpc2_0_n66,
         n_hpc2_0_n65, n_hpc2_0_n64, n_hpc2_0_n63, n_hpc2_0_n62, n_hpc2_0_n61,
         n_hpc2_0_n60, n_hpc2_0_n59, n_hpc2_0_n58, n_hpc2_0_n57, n_hpc2_0_n56,
         n_hpc2_0_n55, n_hpc2_0_n54, n_hpc2_0_n53, n_hpc2_0_n52, n_hpc2_0_n51,
         n_hpc2_0_n50, n_hpc2_0_n49, n_hpc2_0_n48, n_hpc2_0_n47, n_hpc2_0_n46,
         n_hpc2_0_n45, n_hpc2_0_n44, n_hpc2_0_n43, n_hpc2_0_n42, n_hpc2_0_n41,
         n_hpc2_0_n40, n_hpc2_0_n39, n_hpc2_0_n38, n_hpc2_0_n37, n_hpc2_0_n36,
         n_hpc2_0_n35, n_hpc2_0_n34, n_hpc2_0_n33, n_hpc2_0_n32, n_hpc2_0_n31,
         n_hpc2_0_n30, n_hpc2_0_n29, n_hpc2_0_n28, n_hpc2_0_n27, n_hpc2_0_n26,
         n_hpc2_0_n25, n_hpc2_0_n24, n_hpc2_0_n23, n_hpc2_0_n22, n_hpc2_0_n21,
         n_hpc2_0_n20, n_hpc2_0_n19, n_hpc2_0_n18, n_hpc2_0_n17, n_hpc2_0_n16,
         n_hpc2_0_n15, n_hpc2_0_n14, n_hpc2_0_n13, n_hpc2_0_n12, n_hpc2_0_n11,
         n_hpc2_0_n10, n_hpc2_0_n9, n_hpc2_0_n8, n_hpc2_0_n7, n_hpc2_0_n6,
         n_hpc2_0_n5, n_hpc2_0_n4, n_hpc2_0_n3, n_hpc2_0_n2, n_hpc2_0_n1,
         n_hpc2_0_N29, n_hpc2_0_N28, n_hpc2_0_N27, n_hpc2_0_N26, n_hpc2_0_N25,
         n_hpc2_0_N24, n_hpc2_0_N23, n_hpc2_0_N22, n_hpc2_0_N21, n_hpc2_0_N20,
         n_hpc2_0_N19, n_hpc2_0_N18, n_hpc2_0_N17, n_hpc2_0_N16, n_hpc2_0_N15,
         n_hpc2_0_N14, n_hpc2_0_N13, n_hpc2_0_N12, n_hpc2_0_N11, n_hpc2_0_N10,
         n_hpc2_0_N9, n_hpc2_0_N8, n_hpc2_0_N7, n_hpc2_0_N6, n_hpc2_0_N5,
         n_hpc2_0_reg_pipeline_13, n_hpc2_0_reg_pipeline_12,
         n_hpc2_0_reg_pipeline_11, n_hpc2_0_reg_pipeline_10,
         n_hpc2_0_reg_pipeline_9, n_hpc2_0_reg_pipeline_8,
         n_hpc2_0_reg_pipeline_7, n_hpc2_0_reg_pipeline_6,
         n_hpc2_0_reg_pipeline_5, n_hpc2_0_reg_pipeline_4,
         n_hpc2_0_reg_pipeline_3, n_hpc2_0_reg_pipeline_2,
         n_hpc2_0_reg_pipeline_1, n_hpc2_0_reg_pipeline_0,
         n_hpc2_0_reg_pipeline, n_hpc2_0_N4, n_hpc2_0_N3, n_hpc2_0_N2,
         n_hpc2_0_N1, n_hpc2_0_N0, n_hpc2_0__hpc1_z41, n_hpc2_0__hpc1_z31,
         n_hpc2_0__hpc1_z21, n_hpc2_0__hpc1_z11, n_hpc2_0__hpc1_z01;

  XOR2_X1 u_hpc2_0_U87 ( .A(io_i1_s0), .B(p_rand_3), .Z(n_hpc2_0_n55) );
  XOR2_X1 u_hpc2_0_U86 ( .A(p_rand_2), .B(n_hpc2_0_n55), .Z(n_hpc2_0_n53) );
  XOR2_X1 u_hpc2_0_U85 ( .A(p_rand_1), .B(p_rand_0), .Z(n_hpc2_0_n54) );
  XOR2_X1 u_hpc2_0_U84 ( .A(n_hpc2_0_n53), .B(n_hpc2_0_n54), .Z(n_hpc2_0_N0)
         );
  XOR2_X1 u_hpc2_0_U83 ( .A(io_i1_s1), .B(p_rand_6), .Z(n_hpc2_0_n52) );
  XOR2_X1 u_hpc2_0_U82 ( .A(p_rand_5), .B(n_hpc2_0_n52), .Z(n_hpc2_0_n50) );
  XOR2_X1 u_hpc2_0_U81 ( .A(p_rand_4), .B(p_rand_0), .Z(n_hpc2_0_n51) );
  XOR2_X1 u_hpc2_0_U80 ( .A(n_hpc2_0_n50), .B(n_hpc2_0_n51), .Z(n_hpc2_0_N1)
         );
  NAND2_X1 u_hpc2_0_U79 ( .A1(n_hpc2_0_reg_pipeline_4), .A2(n_hpc2_0_n5), .ZN(
        n_hpc2_0_n49) );
  XNOR2_X1 u_hpc2_0_U78 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n49), .ZN(
        n_hpc2_0_N10) );
  AND2_X1 u_hpc2_0_U77 ( .A1(n_hpc2_0_n4), .A2(n_hpc2_0_reg_pipeline_4), .ZN(
        n_hpc2_0_N11) );
  NAND2_X1 u_hpc2_0_U76 ( .A1(n_hpc2_0_reg_pipeline_4), .A2(n_hpc2_0_n3), .ZN(
        n_hpc2_0_n48) );
  XNOR2_X1 u_hpc2_0_U75 ( .A(n_hpc2_0_reg_pipeline_5), .B(n_hpc2_0_n48), .ZN(
        n_hpc2_0_N12) );
  NAND2_X1 u_hpc2_0_U74 ( .A1(n_hpc2_0_reg_pipeline_4), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n47) );
  XNOR2_X1 u_hpc2_0_U73 ( .A(n_hpc2_0_reg_pipeline_6), .B(n_hpc2_0_n47), .ZN(
        n_hpc2_0_N13) );
  NAND2_X1 u_hpc2_0_U72 ( .A1(n_hpc2_0_reg_pipeline_4), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n46) );
  XNOR2_X1 u_hpc2_0_U71 ( .A(n_hpc2_0_reg_pipeline_7), .B(n_hpc2_0_n46), .ZN(
        n_hpc2_0_N14) );
  NAND2_X1 u_hpc2_0_U70 ( .A1(n_hpc2_0_reg_pipeline_8), .A2(n_hpc2_0_n5), .ZN(
        n_hpc2_0_n45) );
  XNOR2_X1 u_hpc2_0_U69 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n45), .ZN(
        n_hpc2_0_N15) );
  NAND2_X1 u_hpc2_0_U68 ( .A1(n_hpc2_0_reg_pipeline_8), .A2(n_hpc2_0_n4), .ZN(
        n_hpc2_0_n44) );
  XNOR2_X1 u_hpc2_0_U67 ( .A(n_hpc2_0_reg_pipeline_5), .B(n_hpc2_0_n44), .ZN(
        n_hpc2_0_N16) );
  AND2_X1 u_hpc2_0_U66 ( .A1(n_hpc2_0_n3), .A2(n_hpc2_0_reg_pipeline_8), .ZN(
        n_hpc2_0_N17) );
  NAND2_X1 u_hpc2_0_U65 ( .A1(n_hpc2_0_reg_pipeline_8), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n43) );
  XNOR2_X1 u_hpc2_0_U64 ( .A(n_hpc2_0_reg_pipeline_9), .B(n_hpc2_0_n43), .ZN(
        n_hpc2_0_N18) );
  NAND2_X1 u_hpc2_0_U63 ( .A1(n_hpc2_0_reg_pipeline_8), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n42) );
  XNOR2_X1 u_hpc2_0_U62 ( .A(n_hpc2_0_reg_pipeline_10), .B(n_hpc2_0_n42), .ZN(
        n_hpc2_0_N19) );
  XOR2_X1 u_hpc2_0_U61 ( .A(io_i1_s2), .B(p_rand_8), .Z(n_hpc2_0_n41) );
  XOR2_X1 u_hpc2_0_U60 ( .A(p_rand_7), .B(n_hpc2_0_n41), .Z(n_hpc2_0_n39) );
  XOR2_X1 u_hpc2_0_U59 ( .A(p_rand_4), .B(p_rand_1), .Z(n_hpc2_0_n40) );
  XOR2_X1 u_hpc2_0_U58 ( .A(n_hpc2_0_n39), .B(n_hpc2_0_n40), .Z(n_hpc2_0_N2)
         );
  NAND2_X1 u_hpc2_0_U57 ( .A1(n_hpc2_0_reg_pipeline_11), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n38) );
  XNOR2_X1 u_hpc2_0_U56 ( .A(n_hpc2_0_reg_pipeline_2), .B(n_hpc2_0_n38), .ZN(
        n_hpc2_0_N20) );
  NAND2_X1 u_hpc2_0_U55 ( .A1(n_hpc2_0_reg_pipeline_11), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n37) );
  XNOR2_X1 u_hpc2_0_U54 ( .A(n_hpc2_0_reg_pipeline_6), .B(n_hpc2_0_n37), .ZN(
        n_hpc2_0_N21) );
  NAND2_X1 u_hpc2_0_U53 ( .A1(n_hpc2_0_reg_pipeline_11), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n36) );
  XNOR2_X1 u_hpc2_0_U52 ( .A(n_hpc2_0_reg_pipeline_9), .B(n_hpc2_0_n36), .ZN(
        n_hpc2_0_N22) );
  AND2_X1 u_hpc2_0_U51 ( .A1(n_hpc2_0_n2), .A2(n_hpc2_0_reg_pipeline_11), .ZN(
        n_hpc2_0_N23) );
  NAND2_X1 u_hpc2_0_U50 ( .A1(n_hpc2_0_reg_pipeline_11), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n35) );
  XNOR2_X1 u_hpc2_0_U49 ( .A(n_hpc2_0_reg_pipeline_12), .B(n_hpc2_0_n35), .ZN(
        n_hpc2_0_N24) );
  NAND2_X1 u_hpc2_0_U48 ( .A1(n_hpc2_0_reg_pipeline_13), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n34) );
  XNOR2_X1 u_hpc2_0_U47 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n34), .ZN(
        n_hpc2_0_N25) );
  NAND2_X1 u_hpc2_0_U46 ( .A1(n_hpc2_0_reg_pipeline_13), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n33) );
  XNOR2_X1 u_hpc2_0_U45 ( .A(n_hpc2_0_reg_pipeline_7), .B(n_hpc2_0_n33), .ZN(
        n_hpc2_0_N26) );
  NAND2_X1 u_hpc2_0_U44 ( .A1(n_hpc2_0_reg_pipeline_13), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n32) );
  XNOR2_X1 u_hpc2_0_U43 ( .A(n_hpc2_0_reg_pipeline_10), .B(n_hpc2_0_n32), .ZN(
        n_hpc2_0_N27) );
  NAND2_X1 u_hpc2_0_U42 ( .A1(n_hpc2_0_reg_pipeline_13), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n31) );
  XNOR2_X1 u_hpc2_0_U41 ( .A(n_hpc2_0_reg_pipeline_12), .B(n_hpc2_0_n31), .ZN(
        n_hpc2_0_N28) );
  AND2_X1 u_hpc2_0_U40 ( .A1(n_hpc2_0_n1), .A2(n_hpc2_0_reg_pipeline_13), .ZN(
        n_hpc2_0_N29) );
  XOR2_X1 u_hpc2_0_U39 ( .A(io_i1_s3), .B(p_rand_9), .Z(n_hpc2_0_n30) );
  XOR2_X1 u_hpc2_0_U38 ( .A(p_rand_7), .B(n_hpc2_0_n30), .Z(n_hpc2_0_n28) );
  XOR2_X1 u_hpc2_0_U37 ( .A(p_rand_5), .B(p_rand_2), .Z(n_hpc2_0_n29) );
  XOR2_X1 u_hpc2_0_U36 ( .A(n_hpc2_0_n28), .B(n_hpc2_0_n29), .Z(n_hpc2_0_N3)
         );
  XOR2_X1 u_hpc2_0_U35 ( .A(io_i1_s4), .B(p_rand_9), .Z(n_hpc2_0_n27) );
  XOR2_X1 u_hpc2_0_U34 ( .A(p_rand_8), .B(n_hpc2_0_n27), .Z(n_hpc2_0_n25) );
  XOR2_X1 u_hpc2_0_U33 ( .A(p_rand_6), .B(p_rand_3), .Z(n_hpc2_0_n26) );
  XOR2_X1 u_hpc2_0_U32 ( .A(n_hpc2_0_n25), .B(n_hpc2_0_n26), .Z(n_hpc2_0_N4)
         );
  AND2_X1 u_hpc2_0_U31 ( .A1(n_hpc2_0_n5), .A2(n_hpc2_0_reg_pipeline), .ZN(
        n_hpc2_0_N5) );
  NAND2_X1 u_hpc2_0_U30 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n4), .ZN(
        n_hpc2_0_n24) );
  XNOR2_X1 u_hpc2_0_U29 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n24), .ZN(
        n_hpc2_0_N6) );
  NAND2_X1 u_hpc2_0_U28 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n3), .ZN(
        n_hpc2_0_n23) );
  XNOR2_X1 u_hpc2_0_U27 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n23), .ZN(
        n_hpc2_0_N7) );
  NAND2_X1 u_hpc2_0_U26 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n22) );
  XNOR2_X1 u_hpc2_0_U25 ( .A(n_hpc2_0_reg_pipeline_2), .B(n_hpc2_0_n22), .ZN(
        n_hpc2_0_N8) );
  NAND2_X1 u_hpc2_0_U24 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n21) );
  XNOR2_X1 u_hpc2_0_U23 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n21), .ZN(
        n_hpc2_0_N9) );
  XOR2_X1 u_hpc2_0_U22 ( .A(n_hpc2_0__hpc1_z01), .B(n_hpc2_0_n72), .Z(
        n_hpc2_0_n20) );
  XOR2_X1 u_hpc2_0_U21 ( .A(n_hpc2_0_n20), .B(n_hpc2_0_n73), .Z(n_hpc2_0_n18)
         );
  XOR2_X1 u_hpc2_0_U20 ( .A(n_hpc2_0_n74), .B(n_hpc2_0_n75), .Z(n_hpc2_0_n19)
         );
  XOR2_X1 u_hpc2_0_U19 ( .A(n_hpc2_0_n18), .B(n_hpc2_0_n19), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0__hpc1_z11), .B(n_hpc2_0_n68), .Z(
        n_hpc2_0_n17) );
  XOR2_X1 u_hpc2_0_U17 ( .A(n_hpc2_0_n17), .B(n_hpc2_0_n69), .Z(n_hpc2_0_n15)
         );
  XOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_n70), .B(n_hpc2_0_n71), .Z(n_hpc2_0_n16)
         );
  XOR2_X1 u_hpc2_0_U15 ( .A(n_hpc2_0_n15), .B(n_hpc2_0_n16), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0__hpc1_z21), .B(n_hpc2_0_n64), .Z(
        n_hpc2_0_n14) );
  XOR2_X1 u_hpc2_0_U13 ( .A(n_hpc2_0_n14), .B(n_hpc2_0_n65), .Z(n_hpc2_0_n12)
         );
  XOR2_X1 u_hpc2_0_U12 ( .A(n_hpc2_0_n66), .B(n_hpc2_0_n67), .Z(n_hpc2_0_n13)
         );
  XOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_n12), .B(n_hpc2_0_n13), .Z(io_o0_s2) );
  XOR2_X1 u_hpc2_0_U10 ( .A(n_hpc2_0__hpc1_z31), .B(n_hpc2_0_n60), .Z(
        n_hpc2_0_n11) );
  XOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_n11), .B(n_hpc2_0_n61), .Z(n_hpc2_0_n9) );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0_n62), .B(n_hpc2_0_n63), .Z(n_hpc2_0_n10)
         );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0_n9), .B(n_hpc2_0_n10), .Z(io_o0_s3) );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0__hpc1_z41), .B(n_hpc2_0_n56), .Z(
        n_hpc2_0_n8) );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0_n8), .B(n_hpc2_0_n57), .Z(n_hpc2_0_n6) );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0_n58), .B(n_hpc2_0_n59), .Z(n_hpc2_0_n7) );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n6), .B(n_hpc2_0_n7), .Z(io_o0_s4) );
  DFF_X1 u_hpc2_0__hpc1_z34_reg ( .D(n_hpc2_0_N24), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n63) );
  DFF_X1 u_hpc2_0__hpc1_z33_reg ( .D(n_hpc2_0_N23), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n62) );
  DFF_X1 u_hpc2_0__hpc1_z32_reg ( .D(n_hpc2_0_N22), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n61) );
  DFF_X1 u_hpc2_0__hpc1_z31_reg ( .D(n_hpc2_0_N21), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z31), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z30_reg ( .D(n_hpc2_0_N20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n60) );
  DFF_X1 u_hpc2_0__hpc1_z24_reg ( .D(n_hpc2_0_N19), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n67) );
  DFF_X1 u_hpc2_0__hpc1_z23_reg ( .D(n_hpc2_0_N18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n66) );
  DFF_X1 u_hpc2_0__hpc1_z22_reg ( .D(n_hpc2_0_N17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n65) );
  DFF_X1 u_hpc2_0__hpc1_z21_reg ( .D(n_hpc2_0_N16), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z21), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z20_reg ( .D(n_hpc2_0_N15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n64) );
  DFF_X1 u_hpc2_0__hpc1_z14_reg ( .D(n_hpc2_0_N14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n71) );
  DFF_X1 u_hpc2_0__hpc1_z13_reg ( .D(n_hpc2_0_N13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n70) );
  DFF_X1 u_hpc2_0__hpc1_z12_reg ( .D(n_hpc2_0_N12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n69) );
  DFF_X1 u_hpc2_0__hpc1_z11_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z11), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z10_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n68) );
  DFF_X1 u_hpc2_0__hpc1_z04_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n75) );
  DFF_X1 u_hpc2_0__hpc1_z03_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n74) );
  DFF_X1 u_hpc2_0__hpc1_z02_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n73) );
  DFF_X1 u_hpc2_0__hpc1_z01_reg ( .D(n_hpc2_0_N6), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z01), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z00_reg ( .D(n_hpc2_0_N5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n72) );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(io_i0_s1), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_4), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(io_i0_s0), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_8_reg ( .D(io_i0_s2), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_8), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(p_rand_11), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_1), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z43_reg ( .D(n_hpc2_0_N28), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n58) );
  DFF_X1 u_hpc2_0__hpc1_ref_v3_reg ( .D(n_hpc2_0_N3), .CK(clock_0), .Q(
        n_hpc2_0_n2), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_11_reg ( .D(io_i0_s3), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_11), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z41_reg ( .D(n_hpc2_0_N26), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z41), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v1_reg ( .D(n_hpc2_0_N1), .CK(clock_0), .Q(
        n_hpc2_0_n4), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z40_reg ( .D(n_hpc2_0_N25), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n56) );
  DFF_X1 u_hpc2_0__hpc1_z42_reg ( .D(n_hpc2_0_N27), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n57) );
  DFF_X1 u_hpc2_0__hpc1_z44_reg ( .D(n_hpc2_0_N29), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n59) );
  DFF_X1 u_hpc2_0_reg_pipeline_13_reg ( .D(io_i0_s4), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_13), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(p_rand_13), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_3), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v0_reg ( .D(n_hpc2_0_N0), .CK(clock_0), .Q(
        n_hpc2_0_n5), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(p_rand_12), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_2), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_7_reg ( .D(p_rand_16), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_7), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_12_reg ( .D(p_rand_19), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_12), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v4_reg ( .D(n_hpc2_0_N4), .CK(clock_0), .Q(
        n_hpc2_0_n1), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_6_reg ( .D(p_rand_15), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_6), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_10_reg ( .D(p_rand_18), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_10), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v2_reg ( .D(n_hpc2_0_N2), .CK(clock_0), .Q(
        n_hpc2_0_n3), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_9_reg ( .D(p_rand_17), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_9), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_5_reg ( .D(p_rand_14), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_5), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(p_rand_10), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_0), .QN() );
endmodule

