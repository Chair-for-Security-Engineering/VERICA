
module Shared_Chi3_Partial ( port_a_in, port_b_in, port_c_in, port_a_out, clk, 
        reset );
  input [1:0] port_a_in;
  input [1:0] port_b_in;
  input [1:0] port_c_in;
  input clk, reset;
  output port_a_out;
  wire   chi3_port_c_out_0_, chi3_port_c_out_1_, chi3_port_b_out_0_,
         chi3_port_b_out_1_, chi3_port_a_out_1_, chi3_st0_t2_port_a_out,
         chi3_st0_t0_port_a_out, chi3_st0_port_c_out_0_,
         chi3_st0_port_c_out_1_, chi3_st0_port_b_out_0_,
         chi3_st0_port_b_out_1_, chi3_st0_t0_n2, chi3_st0_t0_n1,
         chi3_st0_t2_n1, chi3_st0_t1_n4, chi3_st0_t1_n3, chi3_st0_t3_n2,
         chi3_st1_t2_port_a_out, chi3_st1_t0_port_a_out,
         chi3_st1_port_c_out_0_, chi3_st1_port_c_out_1_,
         chi3_st1_port_b_out_0_, chi3_st1_port_b_out_1_, chi3_st1_t0_n4,
         chi3_st1_t0_n3, chi3_st1_t2_n2, chi3_st1_t1_n4, chi3_st1_t1_n3,
         chi3_st1_t3_n2, chi3_st2_t2_port_a_out, chi3_st2_t0_port_a_out,
         chi3_st2_port_c_out_0_, chi3_st2_port_c_out_1_,
         chi3_st2_port_b_out_0_, chi3_st2_port_b_out_1_, chi3_st2_t0_n4,
         chi3_st2_t0_n3, chi3_st2_t2_n2, chi3_st2_t1_n4, chi3_st2_t1_n3,
         chi3_st2_t3_n2;
  wire   [1:0] chi3_st0_a_reg;
  wire   [1:0] chi3_st1_a_reg;
  wire   [1:0] chi3_st2_a_reg;

  DFF_X1 chi3_st0_c_reg_reg_0_ ( .D(port_c_in[0]), .CK(clk), .Q(
        chi3_st0_port_c_out_0_), .QN() );
  DFF_X1 chi3_st0_c_reg_reg_1_ ( .D(port_c_in[1]), .CK(clk), .Q(
        chi3_st0_port_c_out_1_), .QN() );
  DFF_X1 chi3_st0_b_reg_reg_0_ ( .D(port_b_in[0]), .CK(clk), .Q(
        chi3_st0_port_b_out_0_), .QN() );
  DFF_X1 chi3_st0_b_reg_reg_1_ ( .D(port_b_in[1]), .CK(clk), .Q(
        chi3_st0_port_b_out_1_), .QN() );
  DFF_X1 chi3_st0_a_reg_reg_0_ ( .D(chi3_st0_t0_port_a_out), .CK(clk), .Q(
        chi3_st0_a_reg[0]), .QN() );
  DFF_X1 chi3_st0_a_reg_reg_1_ ( .D(chi3_st0_t2_port_a_out), .CK(clk), .Q(
        chi3_st0_a_reg[1]), .QN() );
  INV_X1 chi3_st0_t0_U3 ( .A(port_c_in[1]), .ZN(chi3_st0_t0_n1) );
  NOR2_X1 chi3_st0_t0_U2 ( .A1(port_b_in[0]), .A2(chi3_st0_t0_n1), .ZN(
        chi3_st0_t0_n2) );
  XOR2_X1 chi3_st0_t0_U1 ( .A(port_a_in[0]), .B(chi3_st0_t0_n2), .Z(
        chi3_st0_t0_port_a_out) );
  NAND2_X1 chi3_st0_t2_U2 ( .A1(port_c_in[1]), .A2(port_b_in[1]), .ZN(
        chi3_st0_t2_n1) );
  XNOR2_X1 chi3_st0_t2_U1 ( .A(port_a_in[1]), .B(chi3_st0_t2_n1), .ZN(
        chi3_st0_t2_port_a_out) );
  INV_X1 chi3_st0_t1_U3 ( .A(chi3_st0_port_c_out_0_), .ZN(chi3_st0_t1_n4) );
  NOR2_X1 chi3_st0_t1_U2 ( .A1(chi3_st0_port_b_out_0_), .A2(chi3_st0_t1_n4), 
        .ZN(chi3_st0_t1_n3) );
  XOR2_X1 chi3_st0_t1_U1 ( .A(chi3_st0_a_reg[0]), .B(chi3_st0_t1_n3), .Z(
        port_a_out) );
  NAND2_X1 chi3_st0_t3_U2 ( .A1(chi3_st0_port_c_out_0_), .A2(
        chi3_st0_port_b_out_1_), .ZN(chi3_st0_t3_n2) );
  XNOR2_X1 chi3_st0_t3_U1 ( .A(chi3_st0_a_reg[1]), .B(chi3_st0_t3_n2), .ZN(
        chi3_port_a_out_1_) );
  DFF_X1 chi3_st1_c_reg_reg_0_ ( .D(port_a_in[0]), .CK(clk), .Q(
        chi3_st1_port_c_out_0_), .QN() );
  DFF_X1 chi3_st1_c_reg_reg_1_ ( .D(port_a_in[1]), .CK(clk), .Q(
        chi3_st1_port_c_out_1_), .QN() );
  DFF_X1 chi3_st1_b_reg_reg_0_ ( .D(port_c_in[0]), .CK(clk), .Q(
        chi3_st1_port_b_out_0_), .QN() );
  DFF_X1 chi3_st1_b_reg_reg_1_ ( .D(port_c_in[1]), .CK(clk), .Q(
        chi3_st1_port_b_out_1_), .QN() );
  DFF_X1 chi3_st1_a_reg_reg_0_ ( .D(chi3_st1_t0_port_a_out), .CK(clk), .Q(
        chi3_st1_a_reg[0]), .QN() );
  DFF_X1 chi3_st1_a_reg_reg_1_ ( .D(chi3_st1_t2_port_a_out), .CK(clk), .Q(
        chi3_st1_a_reg[1]), .QN() );
  INV_X1 chi3_st1_t0_U3 ( .A(port_a_in[1]), .ZN(chi3_st1_t0_n4) );
  NOR2_X1 chi3_st1_t0_U2 ( .A1(port_c_in[0]), .A2(chi3_st1_t0_n4), .ZN(
        chi3_st1_t0_n3) );
  XOR2_X1 chi3_st1_t0_U1 ( .A(port_b_in[0]), .B(chi3_st1_t0_n3), .Z(
        chi3_st1_t0_port_a_out) );
  NAND2_X1 chi3_st1_t2_U2 ( .A1(port_a_in[1]), .A2(port_c_in[1]), .ZN(
        chi3_st1_t2_n2) );
  XNOR2_X1 chi3_st1_t2_U1 ( .A(port_b_in[1]), .B(chi3_st1_t2_n2), .ZN(
        chi3_st1_t2_port_a_out) );
  INV_X1 chi3_st1_t1_U3 ( .A(chi3_st1_port_c_out_0_), .ZN(chi3_st1_t1_n4) );
  NOR2_X1 chi3_st1_t1_U2 ( .A1(chi3_st1_port_b_out_0_), .A2(chi3_st1_t1_n4), 
        .ZN(chi3_st1_t1_n3) );
  XOR2_X1 chi3_st1_t1_U1 ( .A(chi3_st1_a_reg[0]), .B(chi3_st1_t1_n3), .Z(
        chi3_port_b_out_0_) );
  NAND2_X1 chi3_st1_t3_U2 ( .A1(chi3_st1_port_c_out_0_), .A2(
        chi3_st1_port_b_out_1_), .ZN(chi3_st1_t3_n2) );
  XNOR2_X1 chi3_st1_t3_U1 ( .A(chi3_st1_a_reg[1]), .B(chi3_st1_t3_n2), .ZN(
        chi3_port_b_out_1_) );
  DFF_X1 chi3_st2_c_reg_reg_0_ ( .D(port_b_in[0]), .CK(clk), .Q(
        chi3_st2_port_c_out_0_), .QN() );
  DFF_X1 chi3_st2_c_reg_reg_1_ ( .D(port_b_in[1]), .CK(clk), .Q(
        chi3_st2_port_c_out_1_), .QN() );
  DFF_X1 chi3_st2_b_reg_reg_0_ ( .D(port_a_in[0]), .CK(clk), .Q(
        chi3_st2_port_b_out_0_), .QN() );
  DFF_X1 chi3_st2_b_reg_reg_1_ ( .D(port_a_in[1]), .CK(clk), .Q(
        chi3_st2_port_b_out_1_), .QN() );
  DFF_X1 chi3_st2_a_reg_reg_0_ ( .D(chi3_st2_t0_port_a_out), .CK(clk), .Q(
        chi3_st2_a_reg[0]), .QN() );
  DFF_X1 chi3_st2_a_reg_reg_1_ ( .D(chi3_st2_t2_port_a_out), .CK(clk), .Q(
        chi3_st2_a_reg[1]), .QN() );
  INV_X1 chi3_st2_t0_U3 ( .A(port_b_in[1]), .ZN(chi3_st2_t0_n4) );
  NOR2_X1 chi3_st2_t0_U2 ( .A1(port_a_in[0]), .A2(chi3_st2_t0_n4), .ZN(
        chi3_st2_t0_n3) );
  XOR2_X1 chi3_st2_t0_U1 ( .A(port_c_in[0]), .B(chi3_st2_t0_n3), .Z(
        chi3_st2_t0_port_a_out) );
  NAND2_X1 chi3_st2_t2_U2 ( .A1(port_b_in[1]), .A2(port_a_in[1]), .ZN(
        chi3_st2_t2_n2) );
  XNOR2_X1 chi3_st2_t2_U1 ( .A(port_c_in[1]), .B(chi3_st2_t2_n2), .ZN(
        chi3_st2_t2_port_a_out) );
  INV_X1 chi3_st2_t1_U3 ( .A(chi3_st2_port_c_out_0_), .ZN(chi3_st2_t1_n4) );
  NOR2_X1 chi3_st2_t1_U2 ( .A1(chi3_st2_port_b_out_0_), .A2(chi3_st2_t1_n4), 
        .ZN(chi3_st2_t1_n3) );
  XOR2_X1 chi3_st2_t1_U1 ( .A(chi3_st2_a_reg[0]), .B(chi3_st2_t1_n3), .Z(
        chi3_port_c_out_0_) );
  NAND2_X1 chi3_st2_t3_U2 ( .A1(chi3_st2_port_c_out_0_), .A2(
        chi3_st2_port_b_out_1_), .ZN(chi3_st2_t3_n2) );
  XNOR2_X1 chi3_st2_t3_U1 ( .A(chi3_st2_a_reg[1]), .B(chi3_st2_t3_n2), .ZN(
        chi3_port_c_out_1_) );
endmodule

