
module Sbox_opt ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i1_s0, io_i1_s1, 
        io_i2_s0, io_i2_s1, io_i3_s0, io_i3_s1, io_i4_s0, io_i4_s1, io_i5_s0, 
        io_i5_s1, io_i6_s0, io_i6_s1, io_i7_s0, io_i7_s1, io_k0_s0, io_k0_s1, 
        io_k1_s0, io_k1_s1, io_k2_s0, io_k2_s1, io_k3_s0, io_k3_s1, io_k4_s0, 
        io_k4_s1, io_k5_s0, io_k5_s1, io_k6_s0, io_k6_s1, io_k7_s0, io_k7_s1, 
        p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, 
        p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12, 
        p_rand_13, p_rand_14, p_rand_15, p_rand_16, p_rand_17, p_rand_18, 
        p_rand_19, p_rand_20, p_rand_21, p_rand_22, p_rand_23, p_rand_24, 
        p_rand_25, p_rand_26, p_rand_27, p_rand_28, p_rand_29, p_rand_30, 
        p_rand_31, p_rand_32, p_rand_33, io_o0_s0, io_o0_s1, io_o1_s0, 
        io_o1_s1, io_o2_s0, io_o2_s1, io_o3_s0, io_o3_s1, io_o4_s0, io_o4_s1, 
        io_o5_s0, io_o5_s1, io_o6_s0, io_o6_s1, io_o7_s0, io_o7_s1 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i1_s0, io_i1_s1, io_i2_s0,
         io_i2_s1, io_i3_s0, io_i3_s1, io_i4_s0, io_i4_s1, io_i5_s0, io_i5_s1,
         io_i6_s0, io_i6_s1, io_i7_s0, io_i7_s1, io_k0_s0, io_k0_s1, io_k1_s0,
         io_k1_s1, io_k2_s0, io_k2_s1, io_k3_s0, io_k3_s1, io_k4_s0, io_k4_s1,
         io_k5_s0, io_k5_s1, io_k6_s0, io_k6_s1, io_k7_s0, io_k7_s1, p_rand_0,
         p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7,
         p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12, p_rand_13,
         p_rand_14, p_rand_15, p_rand_16, p_rand_17, p_rand_18, p_rand_19,
         p_rand_20, p_rand_21, p_rand_22, p_rand_23, p_rand_24, p_rand_25,
         p_rand_26, p_rand_27, p_rand_28, p_rand_29, p_rand_30, p_rand_31,
         p_rand_32, p_rand_33;
  output io_o0_s0, io_o0_s1, io_o1_s0, io_o1_s1, io_o2_s0, io_o2_s1, io_o3_s0,
         io_o3_s1, io_o4_s0, io_o4_s1, io_o5_s0, io_o5_s1, io_o6_s0, io_o6_s1,
         io_o7_s0, io_o7_s1;
  wire   n_xor_module_1_res, n_xor_module_2_res, n_xor_module_3_res,
         n_xor_module_4_res, n_xor_module_5_res, n_xor_module_6_res,
         n_xor_module_7_res, n_xor_module_8_res, n_xor_module_9_res,
         n_xor_module_10_res, n_xor_module_11_res, n_xor_module_12_res,
         n_xor_module_13_res, n_xor_module_14_res, n_xor_module_15_res,
         n_xor_module_16_res, n_xor_module_17_res, n_xor_module_18_res,
         n_xor_module_19_res, n_xor_module_20_res, n_xor_module_21_res,
         n_xor_module_22_res, n_xor_module_23_res, n_xor_module_24_res,
         n_xor_module_25_res, n_xor_module_26_res, n_xor_module_27_res,
         n_xor_module_28_res, n_xor_module_29_res, n_xor_module_30_res,
         n_xor_module_31_res, n_xor_module_32_res, n_xor_module_33_res,
         n_xor_module_34_res, n_xor_module_35_res, n_xor_module_36_res,
         n_xor_module_37_res, n_xor_module_38_res, n_xor_module_39_res,
         n_xor_module_40_res, n_xor_module_41_res, n_xor_module_42_res,
         n_xor_module_43_res, n_xor_module_44_res, n_xor_module_45_res,
         n_xor_module_46_res, n_xor_module_47_res, n_xor_module_48_res,
         n_xor_module_49_res, n_xor_module_50_res, n_xor_module_51_res,
         n_xor_module_52_res, n_xor_module_53_res, n_xor_module_54_res,
         n_and_module_1_res, n_xor_module_55_res, n_reg_module_1_res,
         n_and_module_2_res, n_xor_module_56_res, n_reg_module_2_res,
         n_and_module_3_res, n_xor_module_57_res, n_reg_module_3_res,
         n_and_module_4_res, n_xor_module_58_res, n_reg_module_4_res,
         n_and_module_5_res, n_xor_module_59_res, n_reg_module_5_res,
         n_and_module_6_res, n_xor_module_60_res, n_reg_module_6_res,
         n_and_module_7_res, n_xor_module_61_res, n_reg_module_7_res,
         n_and_module_8_res, n_xor_module_62_res, n_reg_module_8_res,
         n_xor_module_63_res, n_xor_module_64_res, n_and_module_9_res,
         n_xor_module_65_res, n_reg_module_9_res, n_and_module_10_res,
         n_xor_module_66_res, n_reg_module_10_res, n_and_module_11_res,
         n_xor_module_67_res, n_reg_module_11_res, n_and_module_12_res,
         n_xor_module_68_res, n_reg_module_12_res, n_xor_module_69_res,
         n_xor_module_70_res, n_and_module_13_res, n_xor_module_71_res,
         n_reg_module_13_res, n_and_module_14_res, n_xor_module_72_res,
         n_reg_module_14_res, n_and_module_15_res, n_xor_module_73_res,
         n_reg_module_15_res, n_and_module_16_res, n_xor_module_74_res,
         n_reg_module_16_res, n_and_module_17_res, n_xor_module_75_res,
         n_reg_module_17_res, n_and_module_18_res, n_xor_module_76_res,
         n_reg_module_18_res, n_and_module_19_res, n_xor_module_77_res,
         n_reg_module_19_res, n_and_module_20_res, n_xor_module_78_res,
         n_reg_module_20_res, n_xor_module_79_res, n_xor_module_80_res,
         n_and_module_21_res, n_xor_module_81_res, n_reg_module_21_res,
         n_and_module_22_res, n_xor_module_82_res, n_reg_module_22_res,
         n_and_module_23_res, n_xor_module_83_res, n_reg_module_23_res,
         n_and_module_24_res, n_xor_module_84_res, n_reg_module_24_res,
         n_xor_module_85_res, n_xor_module_86_res, n_and_module_25_res,
         n_xor_module_87_res, n_reg_module_25_res, n_and_module_26_res,
         n_xor_module_88_res, n_reg_module_26_res, n_and_module_27_res,
         n_xor_module_89_res, n_reg_module_27_res, n_and_module_28_res,
         n_xor_module_90_res, n_reg_module_28_res, n_and_module_29_res,
         n_xor_module_91_res, n_reg_module_29_res, n_and_module_30_res,
         n_xor_module_92_res, n_reg_module_30_res, n_and_module_31_res,
         n_xor_module_93_res, n_reg_module_31_res, n_and_module_32_res,
         n_xor_module_94_res, n_reg_module_32_res, n_xor_module_95_res,
         n_xor_module_96_res, n_and_module_33_res, n_xor_module_97_res,
         n_reg_module_33_res, n_and_module_34_res, n_xor_module_98_res,
         n_reg_module_34_res, n_and_module_35_res, n_xor_module_99_res,
         n_reg_module_35_res, n_and_module_36_res, n_xor_module_100_res,
         n_reg_module_36_res, n_xor_module_101_res, n_xor_module_102_res,
         n_xor_module_103_res, n_xor_module_104_res, n_xor_module_105_res,
         n_xor_module_106_res, n_xor_module_107_res, n_xor_module_108_res,
         n_xor_module_109_res, n_xor_module_110_res, n_xor_module_111_res,
         n_xor_module_112_res, n_xor_module_113_res, n_xor_module_114_res,
         n_xor_module_115_res, n_xor_module_116_res, n_xor_module_117_res,
         n_xor_module_118_res, n_xor_module_119_res, n_xor_module_120_res,
         n_and_module_37_res, n_xor_module_121_res, n_reg_module_37_res,
         n_and_module_38_res, n_xor_module_122_res, n_reg_module_38_res,
         n_and_module_39_res, n_xor_module_123_res, n_reg_module_39_res,
         n_and_module_40_res, n_xor_module_124_res, n_reg_module_40_res,
         n_xor_module_125_res, n_xor_module_126_res, n_xor_module_127_res,
         n_xor_module_128_res, n_xor_module_129_res, n_xor_module_130_res,
         n_and_module_41_res, n_xor_module_131_res, n_reg_module_41_res,
         n_and_module_42_res, n_xor_module_132_res, n_reg_module_42_res,
         n_and_module_43_res, n_xor_module_133_res, n_reg_module_43_res,
         n_and_module_44_res, n_xor_module_134_res, n_reg_module_44_res,
         n_and_module_45_res, n_xor_module_135_res, n_reg_module_45_res,
         n_and_module_46_res, n_xor_module_136_res, n_reg_module_46_res,
         n_and_module_47_res, n_xor_module_137_res, n_reg_module_47_res,
         n_and_module_48_res, n_xor_module_138_res, n_reg_module_48_res,
         n_and_module_49_res, n_xor_module_139_res, n_reg_module_49_res,
         n_and_module_50_res, n_xor_module_140_res, n_reg_module_50_res,
         n_and_module_51_res, n_xor_module_141_res, n_reg_module_51_res,
         n_and_module_52_res, n_xor_module_142_res, n_reg_module_52_res,
         n_and_module_53_res, n_xor_module_143_res, n_reg_module_53_res,
         n_and_module_54_res, n_xor_module_144_res, n_reg_module_54_res,
         n_and_module_55_res, n_xor_module_145_res, n_reg_module_55_res,
         n_and_module_56_res, n_xor_module_146_res, n_reg_module_56_res,
         n_xor_module_147_res, n_xor_module_148_res, n_and_module_57_res,
         n_xor_module_149_res, n_reg_module_57_res, n_and_module_58_res,
         n_xor_module_150_res, n_reg_module_58_res, n_and_module_59_res,
         n_xor_module_151_res, n_reg_module_59_res, n_and_module_60_res,
         n_xor_module_152_res, n_reg_module_60_res, n_and_module_61_res,
         n_xor_module_153_res, n_reg_module_61_res, n_and_module_62_res,
         n_xor_module_154_res, n_reg_module_62_res, n_and_module_63_res,
         n_xor_module_155_res, n_reg_module_63_res, n_and_module_64_res,
         n_xor_module_156_res, n_reg_module_64_res, n_xor_module_157_res,
         n_xor_module_158_res, n_xor_module_159_res, n_xor_module_160_res,
         n_xor_module_161_res, n_xor_module_162_res, n_xor_module_163_res,
         n_xor_module_164_res, n_xor_module_165_res, n_xor_module_166_res,
         n_xor_module_167_res, n_xor_module_168_res, n_xor_module_169_res,
         n_xor_module_170_res, n_xor_module_171_res, n_xor_module_172_res,
         n_xor_module_173_res, n_xor_module_174_res, n_xor_module_175_res,
         n_xor_module_176_res, n_and_module_65_res, n_xor_module_177_res,
         n_reg_module_65_res, n_and_module_66_res, n_xor_module_178_res,
         n_reg_module_66_res, n_and_module_67_res, n_xor_module_179_res,
         n_reg_module_67_res, n_and_module_68_res, n_xor_module_180_res,
         n_reg_module_68_res, n_and_module_69_res, n_xor_module_181_res,
         n_reg_module_69_res, n_and_module_70_res, n_xor_module_182_res,
         n_reg_module_70_res, n_and_module_71_res, n_xor_module_183_res,
         n_reg_module_71_res, n_and_module_72_res, n_xor_module_184_res,
         n_reg_module_72_res, n_and_module_73_res, n_xor_module_185_res,
         n_reg_module_73_res, n_and_module_74_res, n_xor_module_186_res,
         n_reg_module_74_res, n_and_module_75_res, n_xor_module_187_res,
         n_reg_module_75_res, n_and_module_76_res, n_xor_module_188_res,
         n_reg_module_76_res, n_and_module_77_res, n_xor_module_189_res,
         n_reg_module_77_res, n_and_module_78_res, n_xor_module_190_res,
         n_reg_module_78_res, n_and_module_79_res, n_xor_module_191_res,
         n_reg_module_79_res, n_and_module_80_res, n_xor_module_192_res,
         n_reg_module_80_res, n_and_module_81_res, n_xor_module_193_res,
         n_reg_module_81_res, n_and_module_82_res, n_xor_module_194_res,
         n_reg_module_82_res, n_and_module_83_res, n_xor_module_195_res,
         n_reg_module_83_res, n_and_module_84_res, n_xor_module_196_res,
         n_reg_module_84_res, n_and_module_85_res, n_xor_module_197_res,
         n_reg_module_85_res, n_and_module_86_res, n_xor_module_198_res,
         n_reg_module_86_res, n_and_module_87_res, n_xor_module_199_res,
         n_reg_module_87_res, n_and_module_88_res, n_xor_module_200_res,
         n_reg_module_88_res, n_and_module_89_res, n_xor_module_201_res,
         n_reg_module_89_res, n_and_module_90_res, n_xor_module_202_res,
         n_reg_module_90_res, n_and_module_91_res, n_xor_module_203_res,
         n_reg_module_91_res, n_and_module_92_res, n_xor_module_204_res,
         n_reg_module_92_res, n_and_module_93_res, n_xor_module_205_res,
         n_reg_module_93_res, n_and_module_94_res, n_xor_module_206_res,
         n_reg_module_94_res, n_and_module_95_res, n_xor_module_207_res,
         n_reg_module_95_res, n_and_module_96_res, n_xor_module_208_res,
         n_reg_module_96_res, n_and_module_97_res, n_xor_module_209_res,
         n_reg_module_97_res, n_and_module_98_res, n_xor_module_210_res,
         n_reg_module_98_res, n_and_module_99_res, n_xor_module_211_res,
         n_reg_module_99_res, n_and_module_100_res, n_xor_module_212_res,
         n_reg_module_100_res, n_and_module_101_res, n_xor_module_213_res,
         n_reg_module_101_res, n_and_module_102_res, n_xor_module_214_res,
         n_reg_module_102_res, n_and_module_103_res, n_xor_module_215_res,
         n_reg_module_103_res, n_and_module_104_res, n_xor_module_216_res,
         n_reg_module_104_res, n_and_module_105_res, n_xor_module_217_res,
         n_reg_module_105_res, n_and_module_106_res, n_xor_module_218_res,
         n_reg_module_106_res, n_and_module_107_res, n_xor_module_219_res,
         n_reg_module_107_res, n_and_module_108_res, n_xor_module_220_res,
         n_reg_module_108_res, n_and_module_109_res, n_xor_module_221_res,
         n_reg_module_109_res, n_and_module_110_res, n_xor_module_222_res,
         n_reg_module_110_res, n_and_module_111_res, n_xor_module_223_res,
         n_reg_module_111_res, n_and_module_112_res, n_xor_module_224_res,
         n_reg_module_112_res, n_and_module_113_res, n_xor_module_225_res,
         n_reg_module_113_res, n_and_module_114_res, n_xor_module_226_res,
         n_reg_module_114_res, n_and_module_115_res, n_xor_module_227_res,
         n_reg_module_115_res, n_and_module_116_res, n_xor_module_228_res,
         n_reg_module_116_res, n_and_module_117_res, n_xor_module_229_res,
         n_reg_module_117_res, n_and_module_118_res, n_xor_module_230_res,
         n_reg_module_118_res, n_and_module_119_res, n_xor_module_231_res,
         n_reg_module_119_res, n_and_module_120_res, n_xor_module_232_res,
         n_reg_module_120_res, n_and_module_121_res, n_xor_module_233_res,
         n_reg_module_121_res, n_and_module_122_res, n_xor_module_234_res,
         n_reg_module_122_res, n_and_module_123_res, n_xor_module_235_res,
         n_reg_module_123_res, n_and_module_124_res, n_xor_module_236_res,
         n_reg_module_124_res, n_and_module_125_res, n_xor_module_237_res,
         n_reg_module_125_res, n_and_module_126_res, n_xor_module_238_res,
         n_reg_module_126_res, n_and_module_127_res, n_xor_module_239_res,
         n_reg_module_127_res, n_and_module_128_res, n_xor_module_240_res,
         n_reg_module_128_res, n_and_module_129_res, n_xor_module_241_res,
         n_reg_module_129_res, n_and_module_130_res, n_xor_module_242_res,
         n_reg_module_130_res, n_and_module_131_res, n_xor_module_243_res,
         n_reg_module_131_res, n_and_module_132_res, n_xor_module_244_res,
         n_reg_module_132_res, n_and_module_133_res, n_xor_module_245_res,
         n_reg_module_133_res, n_and_module_134_res, n_xor_module_246_res,
         n_reg_module_134_res, n_and_module_135_res, n_xor_module_247_res,
         n_reg_module_135_res, n_and_module_136_res, n_xor_module_248_res,
         n_reg_module_136_res, n_xor_module_249_res, n_xor_module_250_res,
         n_xor_module_251_res, n_xor_module_252_res, n_xor_module_253_res,
         n_xor_module_254_res, n_xor_module_255_res, n_xor_module_256_res,
         n_xor_module_257_res, n_xor_module_258_res, n_xor_module_259_res,
         n_xor_module_260_res, n_xor_module_261_res, n_xor_module_262_res,
         n_xor_module_263_res, n_xor_module_264_res, n_xor_module_265_res,
         n_xor_module_266_res, n_xor_module_267_res, n_xor_module_268_res,
         n_xor_module_269_res, n_xor_module_270_res, n_xor_module_271_res,
         n_xor_module_272_res, n_xor_module_273_res, n_xor_module_274_res,
         n_xor_module_275_res, n_xor_module_276_res, n_xor_module_277_res,
         n_xor_module_278_res, n_xor_module_279_res, n_xor_module_280_res,
         n_xor_module_281_res, n_xor_module_282_res, n_xor_module_283_res,
         n_xor_module_284_res, n_xor_module_285_res, n_xor_module_286_res,
         n_xor_module_287_res, n_xor_module_288_res, n_xor_module_289_res,
         n_xor_module_290_res, n_xor_module_291_res, n_xor_module_292_res,
         n_xor_module_293_res, n_xor_module_294_res, n_xor_module_295_res,
         n_xor_module_296_res, n_xor_module_297_res, n_xor_module_298_res,
         n_xor_module_299_res, n_xor_module_300_res, n_xor_module_301_res,
         n_xor_module_302_res, n_xor_module_303_res, n_xor_module_304_res,
         n_xor_module_305_res, n_xor_module_306_res, n_xor_module_307_res,
         n_xor_module_308_res, n_xor_module_309_res, n_xor_module_310_res,
         n_xor_module_311_res, n_xor_module_312_res, n_not_module_1_res,
         n_xor_module_313_res, n_xor_module_314_res, n_not_module_2_res,
         n_xor_module_315_res, n_xor_module_316_res, n_xor_module_317_res,
         n_xor_module_318_res, n_xor_module_319_res, n_xor_module_320_res,
         n_xor_module_321_res, n_xor_module_322_res, n_not_module_3_res,
         n_xor_module_323_res, n_xor_module_324_res, n_not_module_4_res;

  XOR2_X1 u_xor_module_1_U1 ( .A(io_i3_s0), .B(io_i0_s0), .Z(
        n_xor_module_1_res) );
  XOR2_X1 u_xor_module_2_U1 ( .A(io_i3_s1), .B(io_i0_s1), .Z(
        n_xor_module_2_res) );
  XOR2_X1 u_xor_module_3_U1 ( .A(io_i5_s0), .B(io_i0_s0), .Z(
        n_xor_module_3_res) );
  XOR2_X1 u_xor_module_4_U1 ( .A(io_i5_s1), .B(io_i0_s1), .Z(
        n_xor_module_4_res) );
  XOR2_X1 u_xor_module_5_U1 ( .A(io_i6_s0), .B(io_i0_s0), .Z(
        n_xor_module_5_res) );
  XOR2_X1 u_xor_module_6_U1 ( .A(io_i6_s1), .B(io_i0_s1), .Z(
        n_xor_module_6_res) );
  XOR2_X1 u_xor_module_7_U1 ( .A(io_i5_s0), .B(io_i3_s0), .Z(
        n_xor_module_7_res) );
  XOR2_X1 u_xor_module_8_U1 ( .A(io_i5_s1), .B(io_i3_s1), .Z(
        n_xor_module_8_res) );
  XOR2_X1 u_xor_module_9_U1 ( .A(io_i6_s0), .B(io_i4_s0), .Z(
        n_xor_module_9_res) );
  XOR2_X1 u_xor_module_10_U1 ( .A(io_i6_s1), .B(io_i4_s1), .Z(
        n_xor_module_10_res) );
  XOR2_X1 u_xor_module_11_U1 ( .A(n_xor_module_9_res), .B(n_xor_module_1_res), 
        .Z(n_xor_module_11_res) );
  XOR2_X1 u_xor_module_12_U1 ( .A(n_xor_module_10_res), .B(n_xor_module_2_res), 
        .Z(n_xor_module_12_res) );
  XOR2_X1 u_xor_module_13_U1 ( .A(io_i2_s0), .B(io_i1_s0), .Z(
        n_xor_module_13_res) );
  XOR2_X1 u_xor_module_14_U1 ( .A(io_i2_s1), .B(io_i1_s1), .Z(
        n_xor_module_14_res) );
  XOR2_X1 u_xor_module_15_U1 ( .A(n_xor_module_11_res), .B(io_i7_s0), .Z(
        n_xor_module_15_res) );
  XOR2_X1 u_xor_module_16_U1 ( .A(n_xor_module_12_res), .B(io_i7_s1), .Z(
        n_xor_module_16_res) );
  XOR2_X1 u_xor_module_17_U1 ( .A(n_xor_module_13_res), .B(io_i7_s0), .Z(
        n_xor_module_17_res) );
  XOR2_X1 u_xor_module_18_U1 ( .A(n_xor_module_14_res), .B(io_i7_s1), .Z(
        n_xor_module_18_res) );
  XOR2_X1 u_xor_module_19_U1 ( .A(n_xor_module_13_res), .B(n_xor_module_11_res), .Z(n_xor_module_19_res) );
  XOR2_X1 u_xor_module_20_U1 ( .A(n_xor_module_14_res), .B(n_xor_module_12_res), .Z(n_xor_module_20_res) );
  XOR2_X1 u_xor_module_21_U1 ( .A(io_i5_s0), .B(io_i1_s0), .Z(
        n_xor_module_21_res) );
  XOR2_X1 u_xor_module_22_U1 ( .A(io_i5_s1), .B(io_i1_s1), .Z(
        n_xor_module_22_res) );
  XOR2_X1 u_xor_module_23_U1 ( .A(io_i5_s0), .B(io_i2_s0), .Z(
        n_xor_module_23_res) );
  XOR2_X1 u_xor_module_24_U1 ( .A(io_i5_s1), .B(io_i2_s1), .Z(
        n_xor_module_24_res) );
  XOR2_X1 u_xor_module_25_U1 ( .A(n_xor_module_7_res), .B(n_xor_module_5_res), 
        .Z(n_xor_module_25_res) );
  XOR2_X1 u_xor_module_26_U1 ( .A(n_xor_module_8_res), .B(n_xor_module_6_res), 
        .Z(n_xor_module_26_res) );
  XOR2_X1 u_xor_module_27_U1 ( .A(n_xor_module_21_res), .B(n_xor_module_11_res), .Z(n_xor_module_27_res) );
  XOR2_X1 u_xor_module_28_U1 ( .A(n_xor_module_22_res), .B(n_xor_module_12_res), .Z(n_xor_module_28_res) );
  XOR2_X1 u_xor_module_29_U1 ( .A(n_xor_module_21_res), .B(n_xor_module_9_res), 
        .Z(n_xor_module_29_res) );
  XOR2_X1 u_xor_module_30_U1 ( .A(n_xor_module_22_res), .B(n_xor_module_10_res), .Z(n_xor_module_30_res) );
  XOR2_X1 u_xor_module_31_U1 ( .A(n_xor_module_23_res), .B(n_xor_module_9_res), 
        .Z(n_xor_module_31_res) );
  XOR2_X1 u_xor_module_32_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_10_res), .Z(n_xor_module_32_res) );
  XOR2_X1 u_xor_module_33_U1 ( .A(n_xor_module_31_res), .B(n_xor_module_17_res), .Z(n_xor_module_33_res) );
  XOR2_X1 u_xor_module_34_U1 ( .A(n_xor_module_32_res), .B(n_xor_module_18_res), .Z(n_xor_module_34_res) );
  XOR2_X1 u_xor_module_35_U1 ( .A(io_i7_s0), .B(io_i3_s0), .Z(
        n_xor_module_35_res) );
  XOR2_X1 u_xor_module_36_U1 ( .A(io_i7_s1), .B(io_i3_s1), .Z(
        n_xor_module_36_res) );
  XOR2_X1 u_xor_module_37_U1 ( .A(n_xor_module_35_res), .B(n_xor_module_13_res), .Z(n_xor_module_37_res) );
  XOR2_X1 u_xor_module_38_U1 ( .A(n_xor_module_36_res), .B(n_xor_module_14_res), .Z(n_xor_module_38_res) );
  XOR2_X1 u_xor_module_39_U1 ( .A(n_xor_module_37_res), .B(n_xor_module_1_res), 
        .Z(n_xor_module_39_res) );
  XOR2_X1 u_xor_module_40_U1 ( .A(n_xor_module_38_res), .B(n_xor_module_2_res), 
        .Z(n_xor_module_40_res) );
  XOR2_X1 u_xor_module_41_U1 ( .A(io_i7_s0), .B(io_i6_s0), .Z(
        n_xor_module_41_res) );
  XOR2_X1 u_xor_module_42_U1 ( .A(io_i7_s1), .B(io_i6_s1), .Z(
        n_xor_module_42_res) );
  XOR2_X1 u_xor_module_43_U1 ( .A(n_xor_module_41_res), .B(n_xor_module_13_res), .Z(n_xor_module_43_res) );
  XOR2_X1 u_xor_module_44_U1 ( .A(n_xor_module_42_res), .B(n_xor_module_14_res), .Z(n_xor_module_44_res) );
  XOR2_X1 u_xor_module_45_U1 ( .A(n_xor_module_43_res), .B(n_xor_module_3_res), 
        .Z(n_xor_module_45_res) );
  XOR2_X1 u_xor_module_46_U1 ( .A(n_xor_module_44_res), .B(n_xor_module_4_res), 
        .Z(n_xor_module_46_res) );
  XOR2_X1 u_xor_module_47_U1 ( .A(n_xor_module_19_res), .B(n_xor_module_3_res), 
        .Z(n_xor_module_47_res) );
  XOR2_X1 u_xor_module_48_U1 ( .A(n_xor_module_20_res), .B(n_xor_module_4_res), 
        .Z(n_xor_module_48_res) );
  XOR2_X1 u_xor_module_49_U1 ( .A(n_xor_module_33_res), .B(n_xor_module_39_res), .Z(n_xor_module_49_res) );
  XOR2_X1 u_xor_module_50_U1 ( .A(n_xor_module_34_res), .B(n_xor_module_40_res), .Z(n_xor_module_50_res) );
  XOR2_X1 u_xor_module_51_U1 ( .A(n_xor_module_31_res), .B(n_xor_module_5_res), 
        .Z(n_xor_module_51_res) );
  XOR2_X1 u_xor_module_52_U1 ( .A(n_xor_module_32_res), .B(n_xor_module_6_res), 
        .Z(n_xor_module_52_res) );
  XOR2_X1 u_xor_module_53_U1 ( .A(n_xor_module_23_res), .B(n_xor_module_1_res), 
        .Z(n_xor_module_53_res) );
  XOR2_X1 u_xor_module_54_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_2_res), 
        .Z(n_xor_module_54_res) );
  AND2_X1 u_and_module_1_U1 ( .A1(n_xor_module_12_res), .A2(
        n_xor_module_25_res), .ZN(n_and_module_1_res) );
  XOR2_X1 u_xor_module_55_U1 ( .A(p_rand_0), .B(n_and_module_1_res), .Z(
        n_xor_module_55_res) );
  DFF_X1 u_reg_module_1__dom_inter0_reg ( .D(n_xor_module_55_res), .CK(clock_0), .Q(n_reg_module_1_res), .QN() );
  AND2_X1 u_and_module_2_U1 ( .A1(n_xor_module_11_res), .A2(
        n_xor_module_25_res), .ZN(n_and_module_2_res) );
  XOR2_X1 u_xor_module_56_U1 ( .A(n_reg_module_1_res), .B(n_and_module_2_res), 
        .Z(n_xor_module_56_res) );
  DFF_X1 u_reg_module_2__dom_inter0_reg ( .D(n_xor_module_56_res), .CK(clock_0), .Q(n_reg_module_2_res), .QN() );
  AND2_X1 u_and_module_3_U1 ( .A1(n_xor_module_11_res), .A2(
        n_xor_module_26_res), .ZN(n_and_module_3_res) );
  XOR2_X1 u_xor_module_57_U1 ( .A(p_rand_0), .B(n_and_module_3_res), .Z(
        n_xor_module_57_res) );
  DFF_X1 u_reg_module_3__dom_inter0_reg ( .D(n_xor_module_57_res), .CK(clock_0), .Q(n_reg_module_3_res), .QN() );
  AND2_X1 u_and_module_4_U1 ( .A1(n_xor_module_12_res), .A2(
        n_xor_module_26_res), .ZN(n_and_module_4_res) );
  XOR2_X1 u_xor_module_58_U1 ( .A(n_reg_module_3_res), .B(n_and_module_4_res), 
        .Z(n_xor_module_58_res) );
  DFF_X1 u_reg_module_4__dom_inter0_reg ( .D(n_xor_module_58_res), .CK(clock_0), .Q(n_reg_module_4_res), .QN() );
  AND2_X1 u_and_module_5_U1 ( .A1(n_xor_module_16_res), .A2(
        n_xor_module_45_res), .ZN(n_and_module_5_res) );
  XOR2_X1 u_xor_module_59_U1 ( .A(p_rand_1), .B(n_and_module_5_res), .Z(
        n_xor_module_59_res) );
  DFF_X1 u_reg_module_5__dom_inter0_reg ( .D(n_xor_module_59_res), .CK(clock_0), .Q(n_reg_module_5_res), .QN() );
  AND2_X1 u_and_module_6_U1 ( .A1(n_xor_module_15_res), .A2(
        n_xor_module_45_res), .ZN(n_and_module_6_res) );
  XOR2_X1 u_xor_module_60_U1 ( .A(n_reg_module_5_res), .B(n_and_module_6_res), 
        .Z(n_xor_module_60_res) );
  DFF_X1 u_reg_module_6__dom_inter0_reg ( .D(n_xor_module_60_res), .CK(clock_0), .Q(n_reg_module_6_res), .QN() );
  AND2_X1 u_and_module_7_U1 ( .A1(n_xor_module_15_res), .A2(
        n_xor_module_46_res), .ZN(n_and_module_7_res) );
  XOR2_X1 u_xor_module_61_U1 ( .A(p_rand_1), .B(n_and_module_7_res), .Z(
        n_xor_module_61_res) );
  DFF_X1 u_reg_module_7__dom_inter0_reg ( .D(n_xor_module_61_res), .CK(clock_0), .Q(n_reg_module_7_res), .QN() );
  AND2_X1 u_and_module_8_U1 ( .A1(n_xor_module_16_res), .A2(
        n_xor_module_46_res), .ZN(n_and_module_8_res) );
  XOR2_X1 u_xor_module_62_U1 ( .A(n_reg_module_7_res), .B(n_and_module_8_res), 
        .Z(n_xor_module_62_res) );
  DFF_X1 u_reg_module_8__dom_inter0_reg ( .D(n_xor_module_62_res), .CK(clock_0), .Q(n_reg_module_8_res), .QN() );
  XOR2_X1 u_xor_module_63_U1 ( .A(n_reg_module_2_res), .B(n_xor_module_27_res), 
        .Z(n_xor_module_63_res) );
  XOR2_X1 u_xor_module_64_U1 ( .A(n_reg_module_4_res), .B(n_xor_module_28_res), 
        .Z(n_xor_module_64_res) );
  AND2_X1 u_and_module_9_U1 ( .A1(io_i7_s1), .A2(n_xor_module_37_res), .ZN(
        n_and_module_9_res) );
  XOR2_X1 u_xor_module_65_U1 ( .A(p_rand_2), .B(n_and_module_9_res), .Z(
        n_xor_module_65_res) );
  DFF_X1 u_reg_module_9__dom_inter0_reg ( .D(n_xor_module_65_res), .CK(clock_0), .Q(n_reg_module_9_res), .QN() );
  AND2_X1 u_and_module_10_U1 ( .A1(io_i7_s0), .A2(n_xor_module_37_res), .ZN(
        n_and_module_10_res) );
  XOR2_X1 u_xor_module_66_U1 ( .A(n_reg_module_9_res), .B(n_and_module_10_res), 
        .Z(n_xor_module_66_res) );
  DFF_X1 u_reg_module_10__dom_inter0_reg ( .D(n_xor_module_66_res), .CK(
        clock_0), .Q(n_reg_module_10_res), .QN() );
  AND2_X1 u_and_module_11_U1 ( .A1(io_i7_s0), .A2(n_xor_module_38_res), .ZN(
        n_and_module_11_res) );
  XOR2_X1 u_xor_module_67_U1 ( .A(p_rand_2), .B(n_and_module_11_res), .Z(
        n_xor_module_67_res) );
  DFF_X1 u_reg_module_11__dom_inter0_reg ( .D(n_xor_module_67_res), .CK(
        clock_0), .Q(n_reg_module_11_res), .QN() );
  AND2_X1 u_and_module_12_U1 ( .A1(io_i7_s1), .A2(n_xor_module_38_res), .ZN(
        n_and_module_12_res) );
  XOR2_X1 u_xor_module_68_U1 ( .A(n_reg_module_11_res), .B(n_and_module_12_res), .Z(n_xor_module_68_res) );
  DFF_X1 u_reg_module_12__dom_inter0_reg ( .D(n_xor_module_68_res), .CK(
        clock_0), .Q(n_reg_module_12_res), .QN() );
  XOR2_X1 u_xor_module_69_U1 ( .A(n_reg_module_2_res), .B(n_reg_module_10_res), 
        .Z(n_xor_module_69_res) );
  XOR2_X1 u_xor_module_70_U1 ( .A(n_reg_module_4_res), .B(n_reg_module_12_res), 
        .Z(n_xor_module_70_res) );
  AND2_X1 u_and_module_13_U1 ( .A1(n_xor_module_32_res), .A2(
        n_xor_module_5_res), .ZN(n_and_module_13_res) );
  XOR2_X1 u_xor_module_71_U1 ( .A(p_rand_3), .B(n_and_module_13_res), .Z(
        n_xor_module_71_res) );
  DFF_X1 u_reg_module_13__dom_inter0_reg ( .D(n_xor_module_71_res), .CK(
        clock_0), .Q(n_reg_module_13_res), .QN() );
  AND2_X1 u_and_module_14_U1 ( .A1(n_xor_module_31_res), .A2(
        n_xor_module_5_res), .ZN(n_and_module_14_res) );
  XOR2_X1 u_xor_module_72_U1 ( .A(n_reg_module_13_res), .B(n_and_module_14_res), .Z(n_xor_module_72_res) );
  DFF_X1 u_reg_module_14__dom_inter0_reg ( .D(n_xor_module_72_res), .CK(
        clock_0), .Q(n_reg_module_14_res), .QN() );
  AND2_X1 u_and_module_15_U1 ( .A1(n_xor_module_31_res), .A2(
        n_xor_module_6_res), .ZN(n_and_module_15_res) );
  XOR2_X1 u_xor_module_73_U1 ( .A(p_rand_3), .B(n_and_module_15_res), .Z(
        n_xor_module_73_res) );
  DFF_X1 u_reg_module_15__dom_inter0_reg ( .D(n_xor_module_73_res), .CK(
        clock_0), .Q(n_reg_module_15_res), .QN() );
  AND2_X1 u_and_module_16_U1 ( .A1(n_xor_module_32_res), .A2(
        n_xor_module_6_res), .ZN(n_and_module_16_res) );
  XOR2_X1 u_xor_module_74_U1 ( .A(n_reg_module_15_res), .B(n_and_module_16_res), .Z(n_xor_module_74_res) );
  DFF_X1 u_reg_module_16__dom_inter0_reg ( .D(n_xor_module_74_res), .CK(
        clock_0), .Q(n_reg_module_16_res), .QN() );
  AND2_X1 u_and_module_17_U1 ( .A1(n_xor_module_18_res), .A2(
        n_xor_module_43_res), .ZN(n_and_module_17_res) );
  XOR2_X1 u_xor_module_75_U1 ( .A(p_rand_4), .B(n_and_module_17_res), .Z(
        n_xor_module_75_res) );
  DFF_X1 u_reg_module_17__dom_inter0_reg ( .D(n_xor_module_75_res), .CK(
        clock_0), .Q(n_reg_module_17_res), .QN() );
  AND2_X1 u_and_module_18_U1 ( .A1(n_xor_module_17_res), .A2(
        n_xor_module_43_res), .ZN(n_and_module_18_res) );
  XOR2_X1 u_xor_module_76_U1 ( .A(n_reg_module_17_res), .B(n_and_module_18_res), .Z(n_xor_module_76_res) );
  DFF_X1 u_reg_module_18__dom_inter0_reg ( .D(n_xor_module_76_res), .CK(
        clock_0), .Q(n_reg_module_18_res), .QN() );
  AND2_X1 u_and_module_19_U1 ( .A1(n_xor_module_17_res), .A2(
        n_xor_module_44_res), .ZN(n_and_module_19_res) );
  XOR2_X1 u_xor_module_77_U1 ( .A(p_rand_4), .B(n_and_module_19_res), .Z(
        n_xor_module_77_res) );
  DFF_X1 u_reg_module_19__dom_inter0_reg ( .D(n_xor_module_77_res), .CK(
        clock_0), .Q(n_reg_module_19_res), .QN() );
  AND2_X1 u_and_module_20_U1 ( .A1(n_xor_module_18_res), .A2(
        n_xor_module_44_res), .ZN(n_and_module_20_res) );
  XOR2_X1 u_xor_module_78_U1 ( .A(n_reg_module_19_res), .B(n_and_module_20_res), .Z(n_xor_module_78_res) );
  DFF_X1 u_reg_module_20__dom_inter0_reg ( .D(n_xor_module_78_res), .CK(
        clock_0), .Q(n_reg_module_20_res), .QN() );
  XOR2_X1 u_xor_module_79_U1 ( .A(n_reg_module_14_res), .B(n_xor_module_51_res), .Z(n_xor_module_79_res) );
  XOR2_X1 u_xor_module_80_U1 ( .A(n_reg_module_16_res), .B(n_xor_module_52_res), .Z(n_xor_module_80_res) );
  AND2_X1 u_and_module_21_U1 ( .A1(n_xor_module_34_res), .A2(
        n_xor_module_39_res), .ZN(n_and_module_21_res) );
  XOR2_X1 u_xor_module_81_U1 ( .A(p_rand_5), .B(n_and_module_21_res), .Z(
        n_xor_module_81_res) );
  DFF_X1 u_reg_module_21__dom_inter0_reg ( .D(n_xor_module_81_res), .CK(
        clock_0), .Q(n_reg_module_21_res), .QN() );
  AND2_X1 u_and_module_22_U1 ( .A1(n_xor_module_33_res), .A2(
        n_xor_module_39_res), .ZN(n_and_module_22_res) );
  XOR2_X1 u_xor_module_82_U1 ( .A(n_reg_module_21_res), .B(n_and_module_22_res), .Z(n_xor_module_82_res) );
  DFF_X1 u_reg_module_22__dom_inter0_reg ( .D(n_xor_module_82_res), .CK(
        clock_0), .Q(n_reg_module_22_res), .QN() );
  AND2_X1 u_and_module_23_U1 ( .A1(n_xor_module_33_res), .A2(
        n_xor_module_40_res), .ZN(n_and_module_23_res) );
  XOR2_X1 u_xor_module_83_U1 ( .A(p_rand_5), .B(n_and_module_23_res), .Z(
        n_xor_module_83_res) );
  DFF_X1 u_reg_module_23__dom_inter0_reg ( .D(n_xor_module_83_res), .CK(
        clock_0), .Q(n_reg_module_23_res), .QN() );
  AND2_X1 u_and_module_24_U1 ( .A1(n_xor_module_34_res), .A2(
        n_xor_module_40_res), .ZN(n_and_module_24_res) );
  XOR2_X1 u_xor_module_84_U1 ( .A(n_reg_module_23_res), .B(n_and_module_24_res), .Z(n_xor_module_84_res) );
  DFF_X1 u_reg_module_24__dom_inter0_reg ( .D(n_xor_module_84_res), .CK(
        clock_0), .Q(n_reg_module_24_res), .QN() );
  XOR2_X1 u_xor_module_85_U1 ( .A(n_reg_module_14_res), .B(n_reg_module_22_res), .Z(n_xor_module_85_res) );
  XOR2_X1 u_xor_module_86_U1 ( .A(n_reg_module_16_res), .B(n_reg_module_24_res), .Z(n_xor_module_86_res) );
  AND2_X1 u_and_module_25_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_1_res), .ZN(n_and_module_25_res) );
  XOR2_X1 u_xor_module_87_U1 ( .A(p_rand_6), .B(n_and_module_25_res), .Z(
        n_xor_module_87_res) );
  DFF_X1 u_reg_module_25__dom_inter0_reg ( .D(n_xor_module_87_res), .CK(
        clock_0), .Q(n_reg_module_25_res), .QN() );
  AND2_X1 u_and_module_26_U1 ( .A1(n_xor_module_29_res), .A2(
        n_xor_module_1_res), .ZN(n_and_module_26_res) );
  XOR2_X1 u_xor_module_88_U1 ( .A(n_reg_module_25_res), .B(n_and_module_26_res), .Z(n_xor_module_88_res) );
  DFF_X1 u_reg_module_26__dom_inter0_reg ( .D(n_xor_module_88_res), .CK(
        clock_0), .Q(n_reg_module_26_res), .QN() );
  AND2_X1 u_and_module_27_U1 ( .A1(n_xor_module_29_res), .A2(
        n_xor_module_2_res), .ZN(n_and_module_27_res) );
  XOR2_X1 u_xor_module_89_U1 ( .A(p_rand_6), .B(n_and_module_27_res), .Z(
        n_xor_module_89_res) );
  DFF_X1 u_reg_module_27__dom_inter0_reg ( .D(n_xor_module_89_res), .CK(
        clock_0), .Q(n_reg_module_27_res), .QN() );
  AND2_X1 u_and_module_28_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_2_res), .ZN(n_and_module_28_res) );
  XOR2_X1 u_xor_module_90_U1 ( .A(n_reg_module_27_res), .B(n_and_module_28_res), .Z(n_xor_module_90_res) );
  DFF_X1 u_reg_module_28__dom_inter0_reg ( .D(n_xor_module_90_res), .CK(
        clock_0), .Q(n_reg_module_28_res), .QN() );
  AND2_X1 u_and_module_29_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_7_res), .ZN(n_and_module_29_res) );
  XOR2_X1 u_xor_module_91_U1 ( .A(p_rand_7), .B(n_and_module_29_res), .Z(
        n_xor_module_91_res) );
  DFF_X1 u_reg_module_29__dom_inter0_reg ( .D(n_xor_module_91_res), .CK(
        clock_0), .Q(n_reg_module_29_res), .QN() );
  AND2_X1 u_and_module_30_U1 ( .A1(n_xor_module_53_res), .A2(
        n_xor_module_7_res), .ZN(n_and_module_30_res) );
  XOR2_X1 u_xor_module_92_U1 ( .A(n_reg_module_29_res), .B(n_and_module_30_res), .Z(n_xor_module_92_res) );
  DFF_X1 u_reg_module_30__dom_inter0_reg ( .D(n_xor_module_92_res), .CK(
        clock_0), .Q(n_reg_module_30_res), .QN() );
  AND2_X1 u_and_module_31_U1 ( .A1(n_xor_module_53_res), .A2(
        n_xor_module_8_res), .ZN(n_and_module_31_res) );
  XOR2_X1 u_xor_module_93_U1 ( .A(p_rand_7), .B(n_and_module_31_res), .Z(
        n_xor_module_93_res) );
  DFF_X1 u_reg_module_31__dom_inter0_reg ( .D(n_xor_module_93_res), .CK(
        clock_0), .Q(n_reg_module_31_res), .QN() );
  AND2_X1 u_and_module_32_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_8_res), .ZN(n_and_module_32_res) );
  XOR2_X1 u_xor_module_94_U1 ( .A(n_reg_module_31_res), .B(n_and_module_32_res), .Z(n_xor_module_94_res) );
  DFF_X1 u_reg_module_32__dom_inter0_reg ( .D(n_xor_module_94_res), .CK(
        clock_0), .Q(n_reg_module_32_res), .QN() );
  XOR2_X1 u_xor_module_95_U1 ( .A(n_reg_module_26_res), .B(n_reg_module_30_res), .Z(n_xor_module_95_res) );
  XOR2_X1 u_xor_module_96_U1 ( .A(n_reg_module_28_res), .B(n_reg_module_32_res), .Z(n_xor_module_96_res) );
  AND2_X1 u_and_module_33_U1 ( .A1(n_xor_module_20_res), .A2(
        n_xor_module_3_res), .ZN(n_and_module_33_res) );
  XOR2_X1 u_xor_module_97_U1 ( .A(p_rand_8), .B(n_and_module_33_res), .Z(
        n_xor_module_97_res) );
  DFF_X1 u_reg_module_33__dom_inter0_reg ( .D(n_xor_module_97_res), .CK(
        clock_0), .Q(n_reg_module_33_res), .QN() );
  AND2_X1 u_and_module_34_U1 ( .A1(n_xor_module_19_res), .A2(
        n_xor_module_3_res), .ZN(n_and_module_34_res) );
  XOR2_X1 u_xor_module_98_U1 ( .A(n_reg_module_33_res), .B(n_and_module_34_res), .Z(n_xor_module_98_res) );
  DFF_X1 u_reg_module_34__dom_inter0_reg ( .D(n_xor_module_98_res), .CK(
        clock_0), .Q(n_reg_module_34_res), .QN() );
  AND2_X1 u_and_module_35_U1 ( .A1(n_xor_module_19_res), .A2(
        n_xor_module_4_res), .ZN(n_and_module_35_res) );
  XOR2_X1 u_xor_module_99_U1 ( .A(p_rand_8), .B(n_and_module_35_res), .Z(
        n_xor_module_99_res) );
  DFF_X1 u_reg_module_35__dom_inter0_reg ( .D(n_xor_module_99_res), .CK(
        clock_0), .Q(n_reg_module_35_res), .QN() );
  AND2_X1 u_and_module_36_U1 ( .A1(n_xor_module_20_res), .A2(
        n_xor_module_4_res), .ZN(n_and_module_36_res) );
  XOR2_X1 u_xor_module_100_U1 ( .A(n_reg_module_35_res), .B(
        n_and_module_36_res), .Z(n_xor_module_100_res) );
  DFF_X1 u_reg_module_36__dom_inter0_reg ( .D(n_xor_module_100_res), .CK(
        clock_0), .Q(n_reg_module_36_res), .QN() );
  XOR2_X1 u_xor_module_101_U1 ( .A(n_reg_module_26_res), .B(
        n_reg_module_34_res), .Z(n_xor_module_101_res) );
  XOR2_X1 u_xor_module_102_U1 ( .A(n_reg_module_28_res), .B(
        n_reg_module_36_res), .Z(n_xor_module_102_res) );
  XOR2_X1 u_xor_module_103_U1 ( .A(n_reg_module_6_res), .B(n_xor_module_63_res), .Z(n_xor_module_103_res) );
  XOR2_X1 u_xor_module_104_U1 ( .A(n_reg_module_8_res), .B(n_xor_module_64_res), .Z(n_xor_module_104_res) );
  XOR2_X1 u_xor_module_105_U1 ( .A(n_xor_module_47_res), .B(
        n_xor_module_69_res), .Z(n_xor_module_105_res) );
  XOR2_X1 u_xor_module_106_U1 ( .A(n_xor_module_48_res), .B(
        n_xor_module_70_res), .Z(n_xor_module_106_res) );
  XOR2_X1 u_xor_module_107_U1 ( .A(n_reg_module_18_res), .B(
        n_xor_module_79_res), .Z(n_xor_module_107_res) );
  XOR2_X1 u_xor_module_108_U1 ( .A(n_reg_module_20_res), .B(
        n_xor_module_80_res), .Z(n_xor_module_108_res) );
  XOR2_X1 u_xor_module_109_U1 ( .A(n_xor_module_101_res), .B(
        n_xor_module_85_res), .Z(n_xor_module_109_res) );
  XOR2_X1 u_xor_module_110_U1 ( .A(n_xor_module_102_res), .B(
        n_xor_module_86_res), .Z(n_xor_module_110_res) );
  XOR2_X1 u_xor_module_111_U1 ( .A(n_xor_module_95_res), .B(
        n_xor_module_103_res), .Z(n_xor_module_111_res) );
  XOR2_X1 u_xor_module_112_U1 ( .A(n_xor_module_96_res), .B(
        n_xor_module_104_res), .Z(n_xor_module_112_res) );
  XOR2_X1 u_xor_module_113_U1 ( .A(n_xor_module_101_res), .B(
        n_xor_module_105_res), .Z(n_xor_module_113_res) );
  XOR2_X1 u_xor_module_114_U1 ( .A(n_xor_module_102_res), .B(
        n_xor_module_106_res), .Z(n_xor_module_114_res) );
  XOR2_X1 u_xor_module_115_U1 ( .A(n_xor_module_95_res), .B(
        n_xor_module_107_res), .Z(n_xor_module_115_res) );
  XOR2_X1 u_xor_module_116_U1 ( .A(n_xor_module_96_res), .B(
        n_xor_module_108_res), .Z(n_xor_module_116_res) );
  XOR2_X1 u_xor_module_117_U1 ( .A(n_xor_module_49_res), .B(
        n_xor_module_109_res), .Z(n_xor_module_117_res) );
  XOR2_X1 u_xor_module_118_U1 ( .A(n_xor_module_50_res), .B(
        n_xor_module_110_res), .Z(n_xor_module_118_res) );
  XOR2_X1 u_xor_module_119_U1 ( .A(n_xor_module_117_res), .B(
        n_xor_module_115_res), .Z(n_xor_module_119_res) );
  XOR2_X1 u_xor_module_120_U1 ( .A(n_xor_module_118_res), .B(
        n_xor_module_116_res), .Z(n_xor_module_120_res) );
  AND2_X1 u_and_module_37_U1 ( .A1(n_xor_module_112_res), .A2(
        n_xor_module_115_res), .ZN(n_and_module_37_res) );
  XOR2_X1 u_xor_module_121_U1 ( .A(p_rand_9), .B(n_and_module_37_res), .Z(
        n_xor_module_121_res) );
  DFF_X1 u_reg_module_37__dom_inter0_reg ( .D(n_xor_module_121_res), .CK(
        clock_0), .Q(n_reg_module_37_res), .QN() );
  AND2_X1 u_and_module_38_U1 ( .A1(n_xor_module_111_res), .A2(
        n_xor_module_115_res), .ZN(n_and_module_38_res) );
  XOR2_X1 u_xor_module_122_U1 ( .A(n_reg_module_37_res), .B(
        n_and_module_38_res), .Z(n_xor_module_122_res) );
  DFF_X1 u_reg_module_38__dom_inter0_reg ( .D(n_xor_module_122_res), .CK(
        clock_0), .Q(n_reg_module_38_res), .QN() );
  AND2_X1 u_and_module_39_U1 ( .A1(n_xor_module_111_res), .A2(
        n_xor_module_116_res), .ZN(n_and_module_39_res) );
  XOR2_X1 u_xor_module_123_U1 ( .A(p_rand_9), .B(n_and_module_39_res), .Z(
        n_xor_module_123_res) );
  DFF_X1 u_reg_module_39__dom_inter0_reg ( .D(n_xor_module_123_res), .CK(
        clock_0), .Q(n_reg_module_39_res), .QN() );
  AND2_X1 u_and_module_40_U1 ( .A1(n_xor_module_112_res), .A2(
        n_xor_module_116_res), .ZN(n_and_module_40_res) );
  XOR2_X1 u_xor_module_124_U1 ( .A(n_reg_module_39_res), .B(
        n_and_module_40_res), .Z(n_xor_module_124_res) );
  DFF_X1 u_reg_module_40__dom_inter0_reg ( .D(n_xor_module_124_res), .CK(
        clock_0), .Q(n_reg_module_40_res), .QN() );
  XOR2_X1 u_xor_module_125_U1 ( .A(n_reg_module_38_res), .B(
        n_xor_module_113_res), .Z(n_xor_module_125_res) );
  XOR2_X1 u_xor_module_126_U1 ( .A(n_reg_module_40_res), .B(
        n_xor_module_114_res), .Z(n_xor_module_126_res) );
  XOR2_X1 u_xor_module_127_U1 ( .A(n_xor_module_113_res), .B(
        n_xor_module_111_res), .Z(n_xor_module_127_res) );
  XOR2_X1 u_xor_module_128_U1 ( .A(n_xor_module_114_res), .B(
        n_xor_module_112_res), .Z(n_xor_module_128_res) );
  XOR2_X1 u_xor_module_129_U1 ( .A(n_reg_module_38_res), .B(
        n_xor_module_117_res), .Z(n_xor_module_129_res) );
  XOR2_X1 u_xor_module_130_U1 ( .A(n_reg_module_40_res), .B(
        n_xor_module_118_res), .Z(n_xor_module_130_res) );
  AND2_X1 u_and_module_41_U1 ( .A1(n_xor_module_128_res), .A2(
        n_xor_module_129_res), .ZN(n_and_module_41_res) );
  XOR2_X1 u_xor_module_131_U1 ( .A(p_rand_10), .B(n_and_module_41_res), .Z(
        n_xor_module_131_res) );
  DFF_X1 u_reg_module_41__dom_inter0_reg ( .D(n_xor_module_131_res), .CK(
        clock_0), .Q(n_reg_module_41_res), .QN() );
  AND2_X1 u_and_module_42_U1 ( .A1(n_xor_module_127_res), .A2(
        n_xor_module_129_res), .ZN(n_and_module_42_res) );
  XOR2_X1 u_xor_module_132_U1 ( .A(n_reg_module_41_res), .B(
        n_and_module_42_res), .Z(n_xor_module_132_res) );
  DFF_X1 u_reg_module_42__dom_inter0_reg ( .D(n_xor_module_132_res), .CK(
        clock_0), .Q(n_reg_module_42_res), .QN() );
  AND2_X1 u_and_module_43_U1 ( .A1(n_xor_module_127_res), .A2(
        n_xor_module_130_res), .ZN(n_and_module_43_res) );
  XOR2_X1 u_xor_module_133_U1 ( .A(p_rand_10), .B(n_and_module_43_res), .Z(
        n_xor_module_133_res) );
  DFF_X1 u_reg_module_43__dom_inter0_reg ( .D(n_xor_module_133_res), .CK(
        clock_0), .Q(n_reg_module_43_res), .QN() );
  AND2_X1 u_and_module_44_U1 ( .A1(n_xor_module_128_res), .A2(
        n_xor_module_130_res), .ZN(n_and_module_44_res) );
  XOR2_X1 u_xor_module_134_U1 ( .A(n_reg_module_43_res), .B(
        n_and_module_44_res), .Z(n_xor_module_134_res) );
  DFF_X1 u_reg_module_44__dom_inter0_reg ( .D(n_xor_module_134_res), .CK(
        clock_0), .Q(n_reg_module_44_res), .QN() );
  AND2_X1 u_and_module_45_U1 ( .A1(n_xor_module_120_res), .A2(
        n_xor_module_125_res), .ZN(n_and_module_45_res) );
  XOR2_X1 u_xor_module_135_U1 ( .A(p_rand_11), .B(n_and_module_45_res), .Z(
        n_xor_module_135_res) );
  DFF_X1 u_reg_module_45__dom_inter0_reg ( .D(n_xor_module_135_res), .CK(
        clock_0), .Q(n_reg_module_45_res), .QN() );
  AND2_X1 u_and_module_46_U1 ( .A1(n_xor_module_119_res), .A2(
        n_xor_module_125_res), .ZN(n_and_module_46_res) );
  XOR2_X1 u_xor_module_136_U1 ( .A(n_reg_module_45_res), .B(
        n_and_module_46_res), .Z(n_xor_module_136_res) );
  DFF_X1 u_reg_module_46__dom_inter0_reg ( .D(n_xor_module_136_res), .CK(
        clock_0), .Q(n_reg_module_46_res), .QN() );
  AND2_X1 u_and_module_47_U1 ( .A1(n_xor_module_119_res), .A2(
        n_xor_module_126_res), .ZN(n_and_module_47_res) );
  XOR2_X1 u_xor_module_137_U1 ( .A(p_rand_11), .B(n_and_module_47_res), .Z(
        n_xor_module_137_res) );
  DFF_X1 u_reg_module_47__dom_inter0_reg ( .D(n_xor_module_137_res), .CK(
        clock_0), .Q(n_reg_module_47_res), .QN() );
  AND2_X1 u_and_module_48_U1 ( .A1(n_xor_module_120_res), .A2(
        n_xor_module_126_res), .ZN(n_and_module_48_res) );
  XOR2_X1 u_xor_module_138_U1 ( .A(n_reg_module_47_res), .B(
        n_and_module_48_res), .Z(n_xor_module_138_res) );
  DFF_X1 u_reg_module_48__dom_inter0_reg ( .D(n_xor_module_138_res), .CK(
        clock_0), .Q(n_reg_module_48_res), .QN() );
  AND2_X1 u_and_module_49_U1 ( .A1(n_xor_module_118_res), .A2(
        n_xor_module_111_res), .ZN(n_and_module_49_res) );
  XOR2_X1 u_xor_module_139_U1 ( .A(p_rand_12), .B(n_and_module_49_res), .Z(
        n_xor_module_139_res) );
  DFF_X1 u_reg_module_49__dom_inter0_reg ( .D(n_xor_module_139_res), .CK(
        clock_0), .Q(n_reg_module_49_res), .QN() );
  AND2_X1 u_and_module_50_U1 ( .A1(n_xor_module_117_res), .A2(
        n_xor_module_111_res), .ZN(n_and_module_50_res) );
  XOR2_X1 u_xor_module_140_U1 ( .A(n_reg_module_49_res), .B(
        n_and_module_50_res), .Z(n_xor_module_140_res) );
  DFF_X1 u_reg_module_50__dom_inter0_reg ( .D(n_xor_module_140_res), .CK(
        clock_0), .Q(n_reg_module_50_res), .QN() );
  AND2_X1 u_and_module_51_U1 ( .A1(n_xor_module_117_res), .A2(
        n_xor_module_112_res), .ZN(n_and_module_51_res) );
  XOR2_X1 u_xor_module_141_U1 ( .A(p_rand_12), .B(n_and_module_51_res), .Z(
        n_xor_module_141_res) );
  DFF_X1 u_reg_module_51__dom_inter0_reg ( .D(n_xor_module_141_res), .CK(
        clock_0), .Q(n_reg_module_51_res), .QN() );
  AND2_X1 u_and_module_52_U1 ( .A1(n_xor_module_118_res), .A2(
        n_xor_module_112_res), .ZN(n_and_module_52_res) );
  XOR2_X1 u_xor_module_142_U1 ( .A(n_reg_module_51_res), .B(
        n_and_module_52_res), .Z(n_xor_module_142_res) );
  DFF_X1 u_reg_module_52__dom_inter0_reg ( .D(n_xor_module_142_res), .CK(
        clock_0), .Q(n_reg_module_52_res), .QN() );
  AND2_X1 u_and_module_53_U1 ( .A1(n_reg_module_52_res), .A2(
        n_xor_module_127_res), .ZN(n_and_module_53_res) );
  XOR2_X1 u_xor_module_143_U1 ( .A(p_rand_13), .B(n_and_module_53_res), .Z(
        n_xor_module_143_res) );
  DFF_X1 u_reg_module_53__dom_inter0_reg ( .D(n_xor_module_143_res), .CK(
        clock_0), .Q(n_reg_module_53_res), .QN() );
  AND2_X1 u_and_module_54_U1 ( .A1(n_reg_module_50_res), .A2(
        n_xor_module_127_res), .ZN(n_and_module_54_res) );
  XOR2_X1 u_xor_module_144_U1 ( .A(n_reg_module_53_res), .B(
        n_and_module_54_res), .Z(n_xor_module_144_res) );
  DFF_X1 u_reg_module_54__dom_inter0_reg ( .D(n_xor_module_144_res), .CK(
        clock_0), .Q(n_reg_module_54_res), .QN() );
  AND2_X1 u_and_module_55_U1 ( .A1(n_reg_module_50_res), .A2(
        n_xor_module_128_res), .ZN(n_and_module_55_res) );
  XOR2_X1 u_xor_module_145_U1 ( .A(p_rand_13), .B(n_and_module_55_res), .Z(
        n_xor_module_145_res) );
  DFF_X1 u_reg_module_55__dom_inter0_reg ( .D(n_xor_module_145_res), .CK(
        clock_0), .Q(n_reg_module_55_res), .QN() );
  AND2_X1 u_and_module_56_U1 ( .A1(n_reg_module_52_res), .A2(
        n_xor_module_128_res), .ZN(n_and_module_56_res) );
  XOR2_X1 u_xor_module_146_U1 ( .A(n_reg_module_55_res), .B(
        n_and_module_56_res), .Z(n_xor_module_146_res) );
  DFF_X1 u_reg_module_56__dom_inter0_reg ( .D(n_xor_module_146_res), .CK(
        clock_0), .Q(n_reg_module_56_res), .QN() );
  XOR2_X1 u_xor_module_147_U1 ( .A(n_reg_module_38_res), .B(
        n_xor_module_127_res), .Z(n_xor_module_147_res) );
  XOR2_X1 u_xor_module_148_U1 ( .A(n_reg_module_40_res), .B(
        n_xor_module_128_res), .Z(n_xor_module_148_res) );
  AND2_X1 u_and_module_57_U1 ( .A1(n_xor_module_116_res), .A2(
        n_xor_module_113_res), .ZN(n_and_module_57_res) );
  XOR2_X1 u_xor_module_149_U1 ( .A(p_rand_14), .B(n_and_module_57_res), .Z(
        n_xor_module_149_res) );
  DFF_X1 u_reg_module_57__dom_inter0_reg ( .D(n_xor_module_149_res), .CK(
        clock_0), .Q(n_reg_module_57_res), .QN() );
  AND2_X1 u_and_module_58_U1 ( .A1(n_xor_module_115_res), .A2(
        n_xor_module_113_res), .ZN(n_and_module_58_res) );
  XOR2_X1 u_xor_module_150_U1 ( .A(n_reg_module_57_res), .B(
        n_and_module_58_res), .Z(n_xor_module_150_res) );
  DFF_X1 u_reg_module_58__dom_inter0_reg ( .D(n_xor_module_150_res), .CK(
        clock_0), .Q(n_reg_module_58_res), .QN() );
  AND2_X1 u_and_module_59_U1 ( .A1(n_xor_module_115_res), .A2(
        n_xor_module_114_res), .ZN(n_and_module_59_res) );
  XOR2_X1 u_xor_module_151_U1 ( .A(p_rand_14), .B(n_and_module_59_res), .Z(
        n_xor_module_151_res) );
  DFF_X1 u_reg_module_59__dom_inter0_reg ( .D(n_xor_module_151_res), .CK(
        clock_0), .Q(n_reg_module_59_res), .QN() );
  AND2_X1 u_and_module_60_U1 ( .A1(n_xor_module_116_res), .A2(
        n_xor_module_114_res), .ZN(n_and_module_60_res) );
  XOR2_X1 u_xor_module_152_U1 ( .A(n_reg_module_59_res), .B(
        n_and_module_60_res), .Z(n_xor_module_152_res) );
  DFF_X1 u_reg_module_60__dom_inter0_reg ( .D(n_xor_module_152_res), .CK(
        clock_0), .Q(n_reg_module_60_res), .QN() );
  AND2_X1 u_and_module_61_U1 ( .A1(n_reg_module_60_res), .A2(
        n_xor_module_119_res), .ZN(n_and_module_61_res) );
  XOR2_X1 u_xor_module_153_U1 ( .A(p_rand_15), .B(n_and_module_61_res), .Z(
        n_xor_module_153_res) );
  DFF_X1 u_reg_module_61__dom_inter0_reg ( .D(n_xor_module_153_res), .CK(
        clock_0), .Q(n_reg_module_61_res), .QN() );
  AND2_X1 u_and_module_62_U1 ( .A1(n_reg_module_58_res), .A2(
        n_xor_module_119_res), .ZN(n_and_module_62_res) );
  XOR2_X1 u_xor_module_154_U1 ( .A(n_reg_module_61_res), .B(
        n_and_module_62_res), .Z(n_xor_module_154_res) );
  DFF_X1 u_reg_module_62__dom_inter0_reg ( .D(n_xor_module_154_res), .CK(
        clock_0), .Q(n_reg_module_62_res), .QN() );
  AND2_X1 u_and_module_63_U1 ( .A1(n_reg_module_58_res), .A2(
        n_xor_module_120_res), .ZN(n_and_module_63_res) );
  XOR2_X1 u_xor_module_155_U1 ( .A(p_rand_15), .B(n_and_module_63_res), .Z(
        n_xor_module_155_res) );
  DFF_X1 u_reg_module_63__dom_inter0_reg ( .D(n_xor_module_155_res), .CK(
        clock_0), .Q(n_reg_module_63_res), .QN() );
  AND2_X1 u_and_module_64_U1 ( .A1(n_reg_module_60_res), .A2(
        n_xor_module_120_res), .ZN(n_and_module_64_res) );
  XOR2_X1 u_xor_module_156_U1 ( .A(n_reg_module_63_res), .B(
        n_and_module_64_res), .Z(n_xor_module_156_res) );
  DFF_X1 u_reg_module_64__dom_inter0_reg ( .D(n_xor_module_156_res), .CK(
        clock_0), .Q(n_reg_module_64_res), .QN() );
  XOR2_X1 u_xor_module_157_U1 ( .A(n_reg_module_38_res), .B(
        n_xor_module_119_res), .Z(n_xor_module_157_res) );
  XOR2_X1 u_xor_module_158_U1 ( .A(n_reg_module_40_res), .B(
        n_xor_module_120_res), .Z(n_xor_module_158_res) );
  XOR2_X1 u_xor_module_159_U1 ( .A(n_reg_module_42_res), .B(
        n_xor_module_113_res), .Z(n_xor_module_159_res) );
  XOR2_X1 u_xor_module_160_U1 ( .A(n_reg_module_44_res), .B(
        n_xor_module_114_res), .Z(n_xor_module_160_res) );
  XOR2_X1 u_xor_module_161_U1 ( .A(n_xor_module_147_res), .B(
        n_reg_module_54_res), .Z(n_xor_module_161_res) );
  XOR2_X1 u_xor_module_162_U1 ( .A(n_xor_module_148_res), .B(
        n_reg_module_56_res), .Z(n_xor_module_162_res) );
  XOR2_X1 u_xor_module_163_U1 ( .A(n_reg_module_46_res), .B(
        n_xor_module_117_res), .Z(n_xor_module_163_res) );
  XOR2_X1 u_xor_module_164_U1 ( .A(n_reg_module_48_res), .B(
        n_xor_module_118_res), .Z(n_xor_module_164_res) );
  XOR2_X1 u_xor_module_165_U1 ( .A(n_xor_module_157_res), .B(
        n_reg_module_62_res), .Z(n_xor_module_165_res) );
  XOR2_X1 u_xor_module_166_U1 ( .A(n_xor_module_158_res), .B(
        n_reg_module_64_res), .Z(n_xor_module_166_res) );
  XOR2_X1 u_xor_module_167_U1 ( .A(n_xor_module_165_res), .B(
        n_xor_module_161_res), .Z(n_xor_module_167_res) );
  XOR2_X1 u_xor_module_168_U1 ( .A(n_xor_module_166_res), .B(
        n_xor_module_162_res), .Z(n_xor_module_168_res) );
  XOR2_X1 u_xor_module_169_U1 ( .A(n_xor_module_163_res), .B(
        n_xor_module_159_res), .Z(n_xor_module_169_res) );
  XOR2_X1 u_xor_module_170_U1 ( .A(n_xor_module_164_res), .B(
        n_xor_module_160_res), .Z(n_xor_module_170_res) );
  XOR2_X1 u_xor_module_171_U1 ( .A(n_xor_module_161_res), .B(
        n_xor_module_159_res), .Z(n_xor_module_171_res) );
  XOR2_X1 u_xor_module_172_U1 ( .A(n_xor_module_162_res), .B(
        n_xor_module_160_res), .Z(n_xor_module_172_res) );
  XOR2_X1 u_xor_module_173_U1 ( .A(n_xor_module_165_res), .B(
        n_xor_module_163_res), .Z(n_xor_module_173_res) );
  XOR2_X1 u_xor_module_174_U1 ( .A(n_xor_module_166_res), .B(
        n_xor_module_164_res), .Z(n_xor_module_174_res) );
  XOR2_X1 u_xor_module_175_U1 ( .A(n_xor_module_167_res), .B(
        n_xor_module_169_res), .Z(n_xor_module_175_res) );
  XOR2_X1 u_xor_module_176_U1 ( .A(n_xor_module_168_res), .B(
        n_xor_module_170_res), .Z(n_xor_module_176_res) );
  AND2_X1 u_and_module_65_U1 ( .A1(n_xor_module_12_res), .A2(
        n_xor_module_173_res), .ZN(n_and_module_65_res) );
  XOR2_X1 u_xor_module_177_U1 ( .A(p_rand_16), .B(n_and_module_65_res), .Z(
        n_xor_module_177_res) );
  DFF_X1 u_reg_module_65__dom_inter0_reg ( .D(n_xor_module_177_res), .CK(
        clock_0), .Q(n_reg_module_65_res), .QN() );
  AND2_X1 u_and_module_66_U1 ( .A1(n_xor_module_11_res), .A2(
        n_xor_module_173_res), .ZN(n_and_module_66_res) );
  XOR2_X1 u_xor_module_178_U1 ( .A(n_reg_module_65_res), .B(
        n_and_module_66_res), .Z(n_xor_module_178_res) );
  DFF_X1 u_reg_module_66__dom_inter0_reg ( .D(n_xor_module_178_res), .CK(
        clock_0), .Q(n_reg_module_66_res), .QN() );
  AND2_X1 u_and_module_67_U1 ( .A1(n_xor_module_11_res), .A2(
        n_xor_module_174_res), .ZN(n_and_module_67_res) );
  XOR2_X1 u_xor_module_179_U1 ( .A(p_rand_16), .B(n_and_module_67_res), .Z(
        n_xor_module_179_res) );
  DFF_X1 u_reg_module_67__dom_inter0_reg ( .D(n_xor_module_179_res), .CK(
        clock_0), .Q(n_reg_module_67_res), .QN() );
  AND2_X1 u_and_module_68_U1 ( .A1(n_xor_module_12_res), .A2(
        n_xor_module_174_res), .ZN(n_and_module_68_res) );
  XOR2_X1 u_xor_module_180_U1 ( .A(n_reg_module_67_res), .B(
        n_and_module_68_res), .Z(n_xor_module_180_res) );
  DFF_X1 u_reg_module_68__dom_inter0_reg ( .D(n_xor_module_180_res), .CK(
        clock_0), .Q(n_reg_module_68_res), .QN() );
  AND2_X1 u_and_module_69_U1 ( .A1(n_xor_module_16_res), .A2(
        n_xor_module_165_res), .ZN(n_and_module_69_res) );
  XOR2_X1 u_xor_module_181_U1 ( .A(p_rand_17), .B(n_and_module_69_res), .Z(
        n_xor_module_181_res) );
  DFF_X1 u_reg_module_69__dom_inter0_reg ( .D(n_xor_module_181_res), .CK(
        clock_0), .Q(n_reg_module_69_res), .QN() );
  AND2_X1 u_and_module_70_U1 ( .A1(n_xor_module_15_res), .A2(
        n_xor_module_165_res), .ZN(n_and_module_70_res) );
  XOR2_X1 u_xor_module_182_U1 ( .A(n_reg_module_69_res), .B(
        n_and_module_70_res), .Z(n_xor_module_182_res) );
  DFF_X1 u_reg_module_70__dom_inter0_reg ( .D(n_xor_module_182_res), .CK(
        clock_0), .Q(n_reg_module_70_res), .QN() );
  AND2_X1 u_and_module_71_U1 ( .A1(n_xor_module_15_res), .A2(
        n_xor_module_166_res), .ZN(n_and_module_71_res) );
  XOR2_X1 u_xor_module_183_U1 ( .A(p_rand_17), .B(n_and_module_71_res), .Z(
        n_xor_module_183_res) );
  DFF_X1 u_reg_module_71__dom_inter0_reg ( .D(n_xor_module_183_res), .CK(
        clock_0), .Q(n_reg_module_71_res), .QN() );
  AND2_X1 u_and_module_72_U1 ( .A1(n_xor_module_16_res), .A2(
        n_xor_module_166_res), .ZN(n_and_module_72_res) );
  XOR2_X1 u_xor_module_184_U1 ( .A(n_reg_module_71_res), .B(
        n_and_module_72_res), .Z(n_xor_module_184_res) );
  DFF_X1 u_reg_module_72__dom_inter0_reg ( .D(n_xor_module_184_res), .CK(
        clock_0), .Q(n_reg_module_72_res), .QN() );
  AND2_X1 u_and_module_73_U1 ( .A1(io_i7_s1), .A2(n_xor_module_163_res), .ZN(
        n_and_module_73_res) );
  XOR2_X1 u_xor_module_185_U1 ( .A(p_rand_18), .B(n_and_module_73_res), .Z(
        n_xor_module_185_res) );
  DFF_X1 u_reg_module_73__dom_inter0_reg ( .D(n_xor_module_185_res), .CK(
        clock_0), .Q(n_reg_module_73_res), .QN() );
  AND2_X1 u_and_module_74_U1 ( .A1(io_i7_s0), .A2(n_xor_module_163_res), .ZN(
        n_and_module_74_res) );
  XOR2_X1 u_xor_module_186_U1 ( .A(n_reg_module_73_res), .B(
        n_and_module_74_res), .Z(n_xor_module_186_res) );
  DFF_X1 u_reg_module_74__dom_inter0_reg ( .D(n_xor_module_186_res), .CK(
        clock_0), .Q(n_reg_module_74_res), .QN() );
  AND2_X1 u_and_module_75_U1 ( .A1(io_i7_s0), .A2(n_xor_module_164_res), .ZN(
        n_and_module_75_res) );
  XOR2_X1 u_xor_module_187_U1 ( .A(p_rand_18), .B(n_and_module_75_res), .Z(
        n_xor_module_187_res) );
  DFF_X1 u_reg_module_75__dom_inter0_reg ( .D(n_xor_module_187_res), .CK(
        clock_0), .Q(n_reg_module_75_res), .QN() );
  AND2_X1 u_and_module_76_U1 ( .A1(io_i7_s1), .A2(n_xor_module_164_res), .ZN(
        n_and_module_76_res) );
  XOR2_X1 u_xor_module_188_U1 ( .A(n_reg_module_75_res), .B(
        n_and_module_76_res), .Z(n_xor_module_188_res) );
  DFF_X1 u_reg_module_76__dom_inter0_reg ( .D(n_xor_module_188_res), .CK(
        clock_0), .Q(n_reg_module_76_res), .QN() );
  AND2_X1 u_and_module_77_U1 ( .A1(n_xor_module_32_res), .A2(
        n_xor_module_171_res), .ZN(n_and_module_77_res) );
  XOR2_X1 u_xor_module_189_U1 ( .A(p_rand_19), .B(n_and_module_77_res), .Z(
        n_xor_module_189_res) );
  DFF_X1 u_reg_module_77__dom_inter0_reg ( .D(n_xor_module_189_res), .CK(
        clock_0), .Q(n_reg_module_77_res), .QN() );
  AND2_X1 u_and_module_78_U1 ( .A1(n_xor_module_31_res), .A2(
        n_xor_module_171_res), .ZN(n_and_module_78_res) );
  XOR2_X1 u_xor_module_190_U1 ( .A(n_reg_module_77_res), .B(
        n_and_module_78_res), .Z(n_xor_module_190_res) );
  DFF_X1 u_reg_module_78__dom_inter0_reg ( .D(n_xor_module_190_res), .CK(
        clock_0), .Q(n_reg_module_78_res), .QN() );
  AND2_X1 u_and_module_79_U1 ( .A1(n_xor_module_31_res), .A2(
        n_xor_module_172_res), .ZN(n_and_module_79_res) );
  XOR2_X1 u_xor_module_191_U1 ( .A(p_rand_19), .B(n_and_module_79_res), .Z(
        n_xor_module_191_res) );
  DFF_X1 u_reg_module_79__dom_inter0_reg ( .D(n_xor_module_191_res), .CK(
        clock_0), .Q(n_reg_module_79_res), .QN() );
  AND2_X1 u_and_module_80_U1 ( .A1(n_xor_module_32_res), .A2(
        n_xor_module_172_res), .ZN(n_and_module_80_res) );
  XOR2_X1 u_xor_module_192_U1 ( .A(n_reg_module_79_res), .B(
        n_and_module_80_res), .Z(n_xor_module_192_res) );
  DFF_X1 u_reg_module_80__dom_inter0_reg ( .D(n_xor_module_192_res), .CK(
        clock_0), .Q(n_reg_module_80_res), .QN() );
  AND2_X1 u_and_module_81_U1 ( .A1(n_xor_module_18_res), .A2(
        n_xor_module_161_res), .ZN(n_and_module_81_res) );
  XOR2_X1 u_xor_module_193_U1 ( .A(p_rand_20), .B(n_and_module_81_res), .Z(
        n_xor_module_193_res) );
  DFF_X1 u_reg_module_81__dom_inter0_reg ( .D(n_xor_module_193_res), .CK(
        clock_0), .Q(n_reg_module_81_res), .QN() );
  AND2_X1 u_and_module_82_U1 ( .A1(n_xor_module_17_res), .A2(
        n_xor_module_161_res), .ZN(n_and_module_82_res) );
  XOR2_X1 u_xor_module_194_U1 ( .A(n_reg_module_81_res), .B(
        n_and_module_82_res), .Z(n_xor_module_194_res) );
  DFF_X1 u_reg_module_82__dom_inter0_reg ( .D(n_xor_module_194_res), .CK(
        clock_0), .Q(n_reg_module_82_res), .QN() );
  AND2_X1 u_and_module_83_U1 ( .A1(n_xor_module_17_res), .A2(
        n_xor_module_162_res), .ZN(n_and_module_83_res) );
  XOR2_X1 u_xor_module_195_U1 ( .A(p_rand_20), .B(n_and_module_83_res), .Z(
        n_xor_module_195_res) );
  DFF_X1 u_reg_module_83__dom_inter0_reg ( .D(n_xor_module_195_res), .CK(
        clock_0), .Q(n_reg_module_83_res), .QN() );
  AND2_X1 u_and_module_84_U1 ( .A1(n_xor_module_18_res), .A2(
        n_xor_module_162_res), .ZN(n_and_module_84_res) );
  XOR2_X1 u_xor_module_196_U1 ( .A(n_reg_module_83_res), .B(
        n_and_module_84_res), .Z(n_xor_module_196_res) );
  DFF_X1 u_reg_module_84__dom_inter0_reg ( .D(n_xor_module_196_res), .CK(
        clock_0), .Q(n_reg_module_84_res), .QN() );
  AND2_X1 u_and_module_85_U1 ( .A1(n_xor_module_34_res), .A2(
        n_xor_module_159_res), .ZN(n_and_module_85_res) );
  XOR2_X1 u_xor_module_197_U1 ( .A(p_rand_21), .B(n_and_module_85_res), .Z(
        n_xor_module_197_res) );
  DFF_X1 u_reg_module_85__dom_inter0_reg ( .D(n_xor_module_197_res), .CK(
        clock_0), .Q(n_reg_module_85_res), .QN() );
  AND2_X1 u_and_module_86_U1 ( .A1(n_xor_module_33_res), .A2(
        n_xor_module_159_res), .ZN(n_and_module_86_res) );
  XOR2_X1 u_xor_module_198_U1 ( .A(n_reg_module_85_res), .B(
        n_and_module_86_res), .Z(n_xor_module_198_res) );
  DFF_X1 u_reg_module_86__dom_inter0_reg ( .D(n_xor_module_198_res), .CK(
        clock_0), .Q(n_reg_module_86_res), .QN() );
  AND2_X1 u_and_module_87_U1 ( .A1(n_xor_module_33_res), .A2(
        n_xor_module_160_res), .ZN(n_and_module_87_res) );
  XOR2_X1 u_xor_module_199_U1 ( .A(p_rand_21), .B(n_and_module_87_res), .Z(
        n_xor_module_199_res) );
  DFF_X1 u_reg_module_87__dom_inter0_reg ( .D(n_xor_module_199_res), .CK(
        clock_0), .Q(n_reg_module_87_res), .QN() );
  AND2_X1 u_and_module_88_U1 ( .A1(n_xor_module_34_res), .A2(
        n_xor_module_160_res), .ZN(n_and_module_88_res) );
  XOR2_X1 u_xor_module_200_U1 ( .A(n_reg_module_87_res), .B(
        n_and_module_88_res), .Z(n_xor_module_200_res) );
  DFF_X1 u_reg_module_88__dom_inter0_reg ( .D(n_xor_module_200_res), .CK(
        clock_0), .Q(n_reg_module_88_res), .QN() );
  AND2_X1 u_and_module_89_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_169_res), .ZN(n_and_module_89_res) );
  XOR2_X1 u_xor_module_201_U1 ( .A(p_rand_22), .B(n_and_module_89_res), .Z(
        n_xor_module_201_res) );
  DFF_X1 u_reg_module_89__dom_inter0_reg ( .D(n_xor_module_201_res), .CK(
        clock_0), .Q(n_reg_module_89_res), .QN() );
  AND2_X1 u_and_module_90_U1 ( .A1(n_xor_module_29_res), .A2(
        n_xor_module_169_res), .ZN(n_and_module_90_res) );
  XOR2_X1 u_xor_module_202_U1 ( .A(n_reg_module_89_res), .B(
        n_and_module_90_res), .Z(n_xor_module_202_res) );
  DFF_X1 u_reg_module_90__dom_inter0_reg ( .D(n_xor_module_202_res), .CK(
        clock_0), .Q(n_reg_module_90_res), .QN() );
  AND2_X1 u_and_module_91_U1 ( .A1(n_xor_module_29_res), .A2(
        n_xor_module_170_res), .ZN(n_and_module_91_res) );
  XOR2_X1 u_xor_module_203_U1 ( .A(p_rand_22), .B(n_and_module_91_res), .Z(
        n_xor_module_203_res) );
  DFF_X1 u_reg_module_91__dom_inter0_reg ( .D(n_xor_module_203_res), .CK(
        clock_0), .Q(n_reg_module_91_res), .QN() );
  AND2_X1 u_and_module_92_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_170_res), .ZN(n_and_module_92_res) );
  XOR2_X1 u_xor_module_204_U1 ( .A(n_reg_module_91_res), .B(
        n_and_module_92_res), .Z(n_xor_module_204_res) );
  DFF_X1 u_reg_module_92__dom_inter0_reg ( .D(n_xor_module_204_res), .CK(
        clock_0), .Q(n_reg_module_92_res), .QN() );
  AND2_X1 u_and_module_93_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_175_res), .ZN(n_and_module_93_res) );
  XOR2_X1 u_xor_module_205_U1 ( .A(p_rand_23), .B(n_and_module_93_res), .Z(
        n_xor_module_205_res) );
  DFF_X1 u_reg_module_93__dom_inter0_reg ( .D(n_xor_module_205_res), .CK(
        clock_0), .Q(n_reg_module_93_res), .QN() );
  AND2_X1 u_and_module_94_U1 ( .A1(n_xor_module_53_res), .A2(
        n_xor_module_175_res), .ZN(n_and_module_94_res) );
  XOR2_X1 u_xor_module_206_U1 ( .A(n_reg_module_93_res), .B(
        n_and_module_94_res), .Z(n_xor_module_206_res) );
  DFF_X1 u_reg_module_94__dom_inter0_reg ( .D(n_xor_module_206_res), .CK(
        clock_0), .Q(n_reg_module_94_res), .QN() );
  AND2_X1 u_and_module_95_U1 ( .A1(n_xor_module_53_res), .A2(
        n_xor_module_176_res), .ZN(n_and_module_95_res) );
  XOR2_X1 u_xor_module_207_U1 ( .A(p_rand_23), .B(n_and_module_95_res), .Z(
        n_xor_module_207_res) );
  DFF_X1 u_reg_module_95__dom_inter0_reg ( .D(n_xor_module_207_res), .CK(
        clock_0), .Q(n_reg_module_95_res), .QN() );
  AND2_X1 u_and_module_96_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_176_res), .ZN(n_and_module_96_res) );
  XOR2_X1 u_xor_module_208_U1 ( .A(n_reg_module_95_res), .B(
        n_and_module_96_res), .Z(n_xor_module_208_res) );
  DFF_X1 u_reg_module_96__dom_inter0_reg ( .D(n_xor_module_208_res), .CK(
        clock_0), .Q(n_reg_module_96_res), .QN() );
  AND2_X1 u_and_module_97_U1 ( .A1(n_xor_module_20_res), .A2(
        n_xor_module_167_res), .ZN(n_and_module_97_res) );
  XOR2_X1 u_xor_module_209_U1 ( .A(p_rand_24), .B(n_and_module_97_res), .Z(
        n_xor_module_209_res) );
  DFF_X1 u_reg_module_97__dom_inter0_reg ( .D(n_xor_module_209_res), .CK(
        clock_0), .Q(n_reg_module_97_res), .QN() );
  AND2_X1 u_and_module_98_U1 ( .A1(n_xor_module_19_res), .A2(
        n_xor_module_167_res), .ZN(n_and_module_98_res) );
  XOR2_X1 u_xor_module_210_U1 ( .A(n_reg_module_97_res), .B(
        n_and_module_98_res), .Z(n_xor_module_210_res) );
  DFF_X1 u_reg_module_98__dom_inter0_reg ( .D(n_xor_module_210_res), .CK(
        clock_0), .Q(n_reg_module_98_res), .QN() );
  AND2_X1 u_and_module_99_U1 ( .A1(n_xor_module_19_res), .A2(
        n_xor_module_168_res), .ZN(n_and_module_99_res) );
  XOR2_X1 u_xor_module_211_U1 ( .A(p_rand_24), .B(n_and_module_99_res), .Z(
        n_xor_module_211_res) );
  DFF_X1 u_reg_module_99__dom_inter0_reg ( .D(n_xor_module_211_res), .CK(
        clock_0), .Q(n_reg_module_99_res), .QN() );
  AND2_X1 u_and_module_100_U1 ( .A1(n_xor_module_20_res), .A2(
        n_xor_module_168_res), .ZN(n_and_module_100_res) );
  XOR2_X1 u_xor_module_212_U1 ( .A(n_reg_module_99_res), .B(
        n_and_module_100_res), .Z(n_xor_module_212_res) );
  DFF_X1 u_reg_module_100__dom_inter0_reg ( .D(n_xor_module_212_res), .CK(
        clock_0), .Q(n_reg_module_100_res), .QN() );
  AND2_X1 u_and_module_101_U1 ( .A1(n_xor_module_26_res), .A2(
        n_xor_module_173_res), .ZN(n_and_module_101_res) );
  XOR2_X1 u_xor_module_213_U1 ( .A(p_rand_25), .B(n_and_module_101_res), .Z(
        n_xor_module_213_res) );
  DFF_X1 u_reg_module_101__dom_inter0_reg ( .D(n_xor_module_213_res), .CK(
        clock_0), .Q(n_reg_module_101_res), .QN() );
  AND2_X1 u_and_module_102_U1 ( .A1(n_xor_module_25_res), .A2(
        n_xor_module_173_res), .ZN(n_and_module_102_res) );
  XOR2_X1 u_xor_module_214_U1 ( .A(n_reg_module_101_res), .B(
        n_and_module_102_res), .Z(n_xor_module_214_res) );
  DFF_X1 u_reg_module_102__dom_inter0_reg ( .D(n_xor_module_214_res), .CK(
        clock_0), .Q(n_reg_module_102_res), .QN() );
  AND2_X1 u_and_module_103_U1 ( .A1(n_xor_module_25_res), .A2(
        n_xor_module_174_res), .ZN(n_and_module_103_res) );
  XOR2_X1 u_xor_module_215_U1 ( .A(p_rand_25), .B(n_and_module_103_res), .Z(
        n_xor_module_215_res) );
  DFF_X1 u_reg_module_103__dom_inter0_reg ( .D(n_xor_module_215_res), .CK(
        clock_0), .Q(n_reg_module_103_res), .QN() );
  AND2_X1 u_and_module_104_U1 ( .A1(n_xor_module_26_res), .A2(
        n_xor_module_174_res), .ZN(n_and_module_104_res) );
  XOR2_X1 u_xor_module_216_U1 ( .A(n_reg_module_103_res), .B(
        n_and_module_104_res), .Z(n_xor_module_216_res) );
  DFF_X1 u_reg_module_104__dom_inter0_reg ( .D(n_xor_module_216_res), .CK(
        clock_0), .Q(n_reg_module_104_res), .QN() );
  AND2_X1 u_and_module_105_U1 ( .A1(n_xor_module_46_res), .A2(
        n_xor_module_165_res), .ZN(n_and_module_105_res) );
  XOR2_X1 u_xor_module_217_U1 ( .A(p_rand_26), .B(n_and_module_105_res), .Z(
        n_xor_module_217_res) );
  DFF_X1 u_reg_module_105__dom_inter0_reg ( .D(n_xor_module_217_res), .CK(
        clock_0), .Q(n_reg_module_105_res), .QN() );
  AND2_X1 u_and_module_106_U1 ( .A1(n_xor_module_45_res), .A2(
        n_xor_module_165_res), .ZN(n_and_module_106_res) );
  XOR2_X1 u_xor_module_218_U1 ( .A(n_reg_module_105_res), .B(
        n_and_module_106_res), .Z(n_xor_module_218_res) );
  DFF_X1 u_reg_module_106__dom_inter0_reg ( .D(n_xor_module_218_res), .CK(
        clock_0), .Q(n_reg_module_106_res), .QN() );
  AND2_X1 u_and_module_107_U1 ( .A1(n_xor_module_45_res), .A2(
        n_xor_module_166_res), .ZN(n_and_module_107_res) );
  XOR2_X1 u_xor_module_219_U1 ( .A(p_rand_26), .B(n_and_module_107_res), .Z(
        n_xor_module_219_res) );
  DFF_X1 u_reg_module_107__dom_inter0_reg ( .D(n_xor_module_219_res), .CK(
        clock_0), .Q(n_reg_module_107_res), .QN() );
  AND2_X1 u_and_module_108_U1 ( .A1(n_xor_module_46_res), .A2(
        n_xor_module_166_res), .ZN(n_and_module_108_res) );
  XOR2_X1 u_xor_module_220_U1 ( .A(n_reg_module_107_res), .B(
        n_and_module_108_res), .Z(n_xor_module_220_res) );
  DFF_X1 u_reg_module_108__dom_inter0_reg ( .D(n_xor_module_220_res), .CK(
        clock_0), .Q(n_reg_module_108_res), .QN() );
  AND2_X1 u_and_module_109_U1 ( .A1(n_xor_module_38_res), .A2(
        n_xor_module_163_res), .ZN(n_and_module_109_res) );
  XOR2_X1 u_xor_module_221_U1 ( .A(p_rand_27), .B(n_and_module_109_res), .Z(
        n_xor_module_221_res) );
  DFF_X1 u_reg_module_109__dom_inter0_reg ( .D(n_xor_module_221_res), .CK(
        clock_0), .Q(n_reg_module_109_res), .QN() );
  AND2_X1 u_and_module_110_U1 ( .A1(n_xor_module_37_res), .A2(
        n_xor_module_163_res), .ZN(n_and_module_110_res) );
  XOR2_X1 u_xor_module_222_U1 ( .A(n_reg_module_109_res), .B(
        n_and_module_110_res), .Z(n_xor_module_222_res) );
  DFF_X1 u_reg_module_110__dom_inter0_reg ( .D(n_xor_module_222_res), .CK(
        clock_0), .Q(n_reg_module_110_res), .QN() );
  AND2_X1 u_and_module_111_U1 ( .A1(n_xor_module_37_res), .A2(
        n_xor_module_164_res), .ZN(n_and_module_111_res) );
  XOR2_X1 u_xor_module_223_U1 ( .A(p_rand_27), .B(n_and_module_111_res), .Z(
        n_xor_module_223_res) );
  DFF_X1 u_reg_module_111__dom_inter0_reg ( .D(n_xor_module_223_res), .CK(
        clock_0), .Q(n_reg_module_111_res), .QN() );
  AND2_X1 u_and_module_112_U1 ( .A1(n_xor_module_38_res), .A2(
        n_xor_module_164_res), .ZN(n_and_module_112_res) );
  XOR2_X1 u_xor_module_224_U1 ( .A(n_reg_module_111_res), .B(
        n_and_module_112_res), .Z(n_xor_module_224_res) );
  DFF_X1 u_reg_module_112__dom_inter0_reg ( .D(n_xor_module_224_res), .CK(
        clock_0), .Q(n_reg_module_112_res), .QN() );
  AND2_X1 u_and_module_113_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_171_res), .ZN(n_and_module_113_res) );
  XOR2_X1 u_xor_module_225_U1 ( .A(p_rand_28), .B(n_and_module_113_res), .Z(
        n_xor_module_225_res) );
  DFF_X1 u_reg_module_113__dom_inter0_reg ( .D(n_xor_module_225_res), .CK(
        clock_0), .Q(n_reg_module_113_res), .QN() );
  AND2_X1 u_and_module_114_U1 ( .A1(n_xor_module_5_res), .A2(
        n_xor_module_171_res), .ZN(n_and_module_114_res) );
  XOR2_X1 u_xor_module_226_U1 ( .A(n_reg_module_113_res), .B(
        n_and_module_114_res), .Z(n_xor_module_226_res) );
  DFF_X1 u_reg_module_114__dom_inter0_reg ( .D(n_xor_module_226_res), .CK(
        clock_0), .Q(n_reg_module_114_res), .QN() );
  AND2_X1 u_and_module_115_U1 ( .A1(n_xor_module_5_res), .A2(
        n_xor_module_172_res), .ZN(n_and_module_115_res) );
  XOR2_X1 u_xor_module_227_U1 ( .A(p_rand_28), .B(n_and_module_115_res), .Z(
        n_xor_module_227_res) );
  DFF_X1 u_reg_module_115__dom_inter0_reg ( .D(n_xor_module_227_res), .CK(
        clock_0), .Q(n_reg_module_115_res), .QN() );
  AND2_X1 u_and_module_116_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_172_res), .ZN(n_and_module_116_res) );
  XOR2_X1 u_xor_module_228_U1 ( .A(n_reg_module_115_res), .B(
        n_and_module_116_res), .Z(n_xor_module_228_res) );
  DFF_X1 u_reg_module_116__dom_inter0_reg ( .D(n_xor_module_228_res), .CK(
        clock_0), .Q(n_reg_module_116_res), .QN() );
  AND2_X1 u_and_module_117_U1 ( .A1(n_xor_module_44_res), .A2(
        n_xor_module_161_res), .ZN(n_and_module_117_res) );
  XOR2_X1 u_xor_module_229_U1 ( .A(p_rand_29), .B(n_and_module_117_res), .Z(
        n_xor_module_229_res) );
  DFF_X1 u_reg_module_117__dom_inter0_reg ( .D(n_xor_module_229_res), .CK(
        clock_0), .Q(n_reg_module_117_res), .QN() );
  AND2_X1 u_and_module_118_U1 ( .A1(n_xor_module_43_res), .A2(
        n_xor_module_161_res), .ZN(n_and_module_118_res) );
  XOR2_X1 u_xor_module_230_U1 ( .A(n_reg_module_117_res), .B(
        n_and_module_118_res), .Z(n_xor_module_230_res) );
  DFF_X1 u_reg_module_118__dom_inter0_reg ( .D(n_xor_module_230_res), .CK(
        clock_0), .Q(n_reg_module_118_res), .QN() );
  AND2_X1 u_and_module_119_U1 ( .A1(n_xor_module_43_res), .A2(
        n_xor_module_162_res), .ZN(n_and_module_119_res) );
  XOR2_X1 u_xor_module_231_U1 ( .A(p_rand_29), .B(n_and_module_119_res), .Z(
        n_xor_module_231_res) );
  DFF_X1 u_reg_module_119__dom_inter0_reg ( .D(n_xor_module_231_res), .CK(
        clock_0), .Q(n_reg_module_119_res), .QN() );
  AND2_X1 u_and_module_120_U1 ( .A1(n_xor_module_44_res), .A2(
        n_xor_module_162_res), .ZN(n_and_module_120_res) );
  XOR2_X1 u_xor_module_232_U1 ( .A(n_reg_module_119_res), .B(
        n_and_module_120_res), .Z(n_xor_module_232_res) );
  DFF_X1 u_reg_module_120__dom_inter0_reg ( .D(n_xor_module_232_res), .CK(
        clock_0), .Q(n_reg_module_120_res), .QN() );
  AND2_X1 u_and_module_121_U1 ( .A1(n_xor_module_40_res), .A2(
        n_xor_module_159_res), .ZN(n_and_module_121_res) );
  XOR2_X1 u_xor_module_233_U1 ( .A(p_rand_30), .B(n_and_module_121_res), .Z(
        n_xor_module_233_res) );
  DFF_X1 u_reg_module_121__dom_inter0_reg ( .D(n_xor_module_233_res), .CK(
        clock_0), .Q(n_reg_module_121_res), .QN() );
  AND2_X1 u_and_module_122_U1 ( .A1(n_xor_module_39_res), .A2(
        n_xor_module_159_res), .ZN(n_and_module_122_res) );
  XOR2_X1 u_xor_module_234_U1 ( .A(n_reg_module_121_res), .B(
        n_and_module_122_res), .Z(n_xor_module_234_res) );
  DFF_X1 u_reg_module_122__dom_inter0_reg ( .D(n_xor_module_234_res), .CK(
        clock_0), .Q(n_reg_module_122_res), .QN() );
  AND2_X1 u_and_module_123_U1 ( .A1(n_xor_module_39_res), .A2(
        n_xor_module_160_res), .ZN(n_and_module_123_res) );
  XOR2_X1 u_xor_module_235_U1 ( .A(p_rand_30), .B(n_and_module_123_res), .Z(
        n_xor_module_235_res) );
  DFF_X1 u_reg_module_123__dom_inter0_reg ( .D(n_xor_module_235_res), .CK(
        clock_0), .Q(n_reg_module_123_res), .QN() );
  AND2_X1 u_and_module_124_U1 ( .A1(n_xor_module_40_res), .A2(
        n_xor_module_160_res), .ZN(n_and_module_124_res) );
  XOR2_X1 u_xor_module_236_U1 ( .A(n_reg_module_123_res), .B(
        n_and_module_124_res), .Z(n_xor_module_236_res) );
  DFF_X1 u_reg_module_124__dom_inter0_reg ( .D(n_xor_module_236_res), .CK(
        clock_0), .Q(n_reg_module_124_res), .QN() );
  AND2_X1 u_and_module_125_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_169_res), .ZN(n_and_module_125_res) );
  XOR2_X1 u_xor_module_237_U1 ( .A(p_rand_31), .B(n_and_module_125_res), .Z(
        n_xor_module_237_res) );
  DFF_X1 u_reg_module_125__dom_inter0_reg ( .D(n_xor_module_237_res), .CK(
        clock_0), .Q(n_reg_module_125_res), .QN() );
  AND2_X1 u_and_module_126_U1 ( .A1(n_xor_module_1_res), .A2(
        n_xor_module_169_res), .ZN(n_and_module_126_res) );
  XOR2_X1 u_xor_module_238_U1 ( .A(n_reg_module_125_res), .B(
        n_and_module_126_res), .Z(n_xor_module_238_res) );
  DFF_X1 u_reg_module_126__dom_inter0_reg ( .D(n_xor_module_238_res), .CK(
        clock_0), .Q(n_reg_module_126_res), .QN() );
  AND2_X1 u_and_module_127_U1 ( .A1(n_xor_module_1_res), .A2(
        n_xor_module_170_res), .ZN(n_and_module_127_res) );
  XOR2_X1 u_xor_module_239_U1 ( .A(p_rand_31), .B(n_and_module_127_res), .Z(
        n_xor_module_239_res) );
  DFF_X1 u_reg_module_127__dom_inter0_reg ( .D(n_xor_module_239_res), .CK(
        clock_0), .Q(n_reg_module_127_res), .QN() );
  AND2_X1 u_and_module_128_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_170_res), .ZN(n_and_module_128_res) );
  XOR2_X1 u_xor_module_240_U1 ( .A(n_reg_module_127_res), .B(
        n_and_module_128_res), .Z(n_xor_module_240_res) );
  DFF_X1 u_reg_module_128__dom_inter0_reg ( .D(n_xor_module_240_res), .CK(
        clock_0), .Q(n_reg_module_128_res), .QN() );
  AND2_X1 u_and_module_129_U1 ( .A1(n_xor_module_8_res), .A2(
        n_xor_module_175_res), .ZN(n_and_module_129_res) );
  XOR2_X1 u_xor_module_241_U1 ( .A(p_rand_32), .B(n_and_module_129_res), .Z(
        n_xor_module_241_res) );
  DFF_X1 u_reg_module_129__dom_inter0_reg ( .D(n_xor_module_241_res), .CK(
        clock_0), .Q(n_reg_module_129_res), .QN() );
  AND2_X1 u_and_module_130_U1 ( .A1(n_xor_module_7_res), .A2(
        n_xor_module_175_res), .ZN(n_and_module_130_res) );
  XOR2_X1 u_xor_module_242_U1 ( .A(n_reg_module_129_res), .B(
        n_and_module_130_res), .Z(n_xor_module_242_res) );
  DFF_X1 u_reg_module_130__dom_inter0_reg ( .D(n_xor_module_242_res), .CK(
        clock_0), .Q(n_reg_module_130_res), .QN() );
  AND2_X1 u_and_module_131_U1 ( .A1(n_xor_module_7_res), .A2(
        n_xor_module_176_res), .ZN(n_and_module_131_res) );
  XOR2_X1 u_xor_module_243_U1 ( .A(p_rand_32), .B(n_and_module_131_res), .Z(
        n_xor_module_243_res) );
  DFF_X1 u_reg_module_131__dom_inter0_reg ( .D(n_xor_module_243_res), .CK(
        clock_0), .Q(n_reg_module_131_res), .QN() );
  AND2_X1 u_and_module_132_U1 ( .A1(n_xor_module_8_res), .A2(
        n_xor_module_176_res), .ZN(n_and_module_132_res) );
  XOR2_X1 u_xor_module_244_U1 ( .A(n_reg_module_131_res), .B(
        n_and_module_132_res), .Z(n_xor_module_244_res) );
  DFF_X1 u_reg_module_132__dom_inter0_reg ( .D(n_xor_module_244_res), .CK(
        clock_0), .Q(n_reg_module_132_res), .QN() );
  AND2_X1 u_and_module_133_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_167_res), .ZN(n_and_module_133_res) );
  XOR2_X1 u_xor_module_245_U1 ( .A(p_rand_33), .B(n_and_module_133_res), .Z(
        n_xor_module_245_res) );
  DFF_X1 u_reg_module_133__dom_inter0_reg ( .D(n_xor_module_245_res), .CK(
        clock_0), .Q(n_reg_module_133_res), .QN() );
  AND2_X1 u_and_module_134_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_167_res), .ZN(n_and_module_134_res) );
  XOR2_X1 u_xor_module_246_U1 ( .A(n_reg_module_133_res), .B(
        n_and_module_134_res), .Z(n_xor_module_246_res) );
  DFF_X1 u_reg_module_134__dom_inter0_reg ( .D(n_xor_module_246_res), .CK(
        clock_0), .Q(n_reg_module_134_res), .QN() );
  AND2_X1 u_and_module_135_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_168_res), .ZN(n_and_module_135_res) );
  XOR2_X1 u_xor_module_247_U1 ( .A(p_rand_33), .B(n_and_module_135_res), .Z(
        n_xor_module_247_res) );
  DFF_X1 u_reg_module_135__dom_inter0_reg ( .D(n_xor_module_247_res), .CK(
        clock_0), .Q(n_reg_module_135_res), .QN() );
  AND2_X1 u_and_module_136_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_168_res), .ZN(n_and_module_136_res) );
  XOR2_X1 u_xor_module_248_U1 ( .A(n_reg_module_135_res), .B(
        n_and_module_136_res), .Z(n_xor_module_248_res) );
  DFF_X1 u_reg_module_136__dom_inter0_reg ( .D(n_xor_module_248_res), .CK(
        clock_0), .Q(n_reg_module_136_res), .QN() );
  XOR2_X1 u_xor_module_249_U1 ( .A(n_reg_module_130_res), .B(
        n_reg_module_126_res), .Z(n_xor_module_249_res) );
  XOR2_X1 u_xor_module_250_U1 ( .A(n_reg_module_132_res), .B(
        n_reg_module_128_res), .Z(n_xor_module_250_res) );
  XOR2_X1 u_xor_module_251_U1 ( .A(n_reg_module_106_res), .B(
        n_reg_module_82_res), .Z(n_xor_module_251_res) );
  XOR2_X1 u_xor_module_252_U1 ( .A(n_reg_module_108_res), .B(
        n_reg_module_84_res), .Z(n_xor_module_252_res) );
  XOR2_X1 u_xor_module_253_U1 ( .A(n_reg_module_74_res), .B(
        n_reg_module_66_res), .Z(n_xor_module_253_res) );
  XOR2_X1 u_xor_module_254_U1 ( .A(n_reg_module_76_res), .B(
        n_reg_module_68_res), .Z(n_xor_module_254_res) );
  XOR2_X1 u_xor_module_255_U1 ( .A(n_reg_module_102_res), .B(
        n_reg_module_70_res), .Z(n_xor_module_255_res) );
  XOR2_X1 u_xor_module_256_U1 ( .A(n_reg_module_104_res), .B(
        n_reg_module_72_res), .Z(n_xor_module_256_res) );
  XOR2_X1 u_xor_module_257_U1 ( .A(n_reg_module_114_res), .B(
        n_reg_module_98_res), .Z(n_xor_module_257_res) );
  XOR2_X1 u_xor_module_258_U1 ( .A(n_reg_module_116_res), .B(
        n_reg_module_100_res), .Z(n_xor_module_258_res) );
  XOR2_X1 u_xor_module_259_U1 ( .A(n_reg_module_126_res), .B(
        n_reg_module_78_res), .Z(n_xor_module_259_res) );
  XOR2_X1 u_xor_module_260_U1 ( .A(n_reg_module_128_res), .B(
        n_reg_module_80_res), .Z(n_xor_module_260_res) );
  XOR2_X1 u_xor_module_261_U1 ( .A(n_xor_module_259_res), .B(
        n_reg_module_130_res), .Z(n_xor_module_261_res) );
  XOR2_X1 u_xor_module_262_U1 ( .A(n_xor_module_260_res), .B(
        n_reg_module_132_res), .Z(n_xor_module_262_res) );
  XOR2_X1 u_xor_module_263_U1 ( .A(n_xor_module_255_res), .B(
        n_reg_module_66_res), .Z(n_xor_module_263_res) );
  XOR2_X1 u_xor_module_264_U1 ( .A(n_xor_module_256_res), .B(
        n_reg_module_68_res), .Z(n_xor_module_264_res) );
  XOR2_X1 u_xor_module_265_U1 ( .A(n_reg_module_118_res), .B(
        n_reg_module_86_res), .Z(n_xor_module_265_res) );
  XOR2_X1 u_xor_module_266_U1 ( .A(n_reg_module_120_res), .B(
        n_reg_module_88_res), .Z(n_xor_module_266_res) );
  XOR2_X1 u_xor_module_267_U1 ( .A(n_reg_module_94_res), .B(
        n_reg_module_90_res), .Z(n_xor_module_267_res) );
  XOR2_X1 u_xor_module_268_U1 ( .A(n_reg_module_96_res), .B(
        n_reg_module_92_res), .Z(n_xor_module_268_res) );
  XOR2_X1 u_xor_module_269_U1 ( .A(n_xor_module_257_res), .B(
        n_reg_module_94_res), .Z(n_xor_module_269_res) );
  XOR2_X1 u_xor_module_270_U1 ( .A(n_xor_module_258_res), .B(
        n_reg_module_96_res), .Z(n_xor_module_270_res) );
  XOR2_X1 u_xor_module_271_U1 ( .A(n_xor_module_253_res), .B(
        n_reg_module_122_res), .Z(n_xor_module_271_res) );
  XOR2_X1 u_xor_module_272_U1 ( .A(n_xor_module_254_res), .B(
        n_reg_module_124_res), .Z(n_xor_module_272_res) );
  XOR2_X1 u_xor_module_273_U1 ( .A(n_reg_module_86_res), .B(
        n_reg_module_74_res), .Z(n_xor_module_273_res) );
  XOR2_X1 u_xor_module_274_U1 ( .A(n_reg_module_88_res), .B(
        n_reg_module_76_res), .Z(n_xor_module_274_res) );
  XOR2_X1 u_xor_module_275_U1 ( .A(n_xor_module_249_res), .B(
        n_reg_module_82_res), .Z(n_xor_module_275_res) );
  XOR2_X1 u_xor_module_276_U1 ( .A(n_xor_module_250_res), .B(
        n_reg_module_84_res), .Z(n_xor_module_276_res) );
  XOR2_X1 u_xor_module_277_U1 ( .A(n_reg_module_126_res), .B(
        n_reg_module_90_res), .Z(n_xor_module_277_res) );
  XOR2_X1 u_xor_module_278_U1 ( .A(n_reg_module_128_res), .B(
        n_reg_module_92_res), .Z(n_xor_module_278_res) );
  XOR2_X1 u_xor_module_279_U1 ( .A(n_xor_module_251_res), .B(
        n_reg_module_102_res), .Z(n_xor_module_279_res) );
  XOR2_X1 u_xor_module_280_U1 ( .A(n_xor_module_252_res), .B(
        n_reg_module_104_res), .Z(n_xor_module_280_res) );
  XOR2_X1 u_xor_module_281_U1 ( .A(n_xor_module_249_res), .B(
        n_reg_module_106_res), .Z(n_xor_module_281_res) );
  XOR2_X1 u_xor_module_282_U1 ( .A(n_xor_module_250_res), .B(
        n_reg_module_108_res), .Z(n_xor_module_282_res) );
  XOR2_X1 u_xor_module_283_U1 ( .A(n_xor_module_251_res), .B(
        n_reg_module_110_res), .Z(n_xor_module_283_res) );
  XOR2_X1 u_xor_module_284_U1 ( .A(n_xor_module_252_res), .B(
        n_reg_module_112_res), .Z(n_xor_module_284_res) );
  XOR2_X1 u_xor_module_285_U1 ( .A(n_xor_module_265_res), .B(
        n_reg_module_114_res), .Z(n_xor_module_285_res) );
  XOR2_X1 u_xor_module_286_U1 ( .A(n_xor_module_266_res), .B(
        n_reg_module_116_res), .Z(n_xor_module_286_res) );
  XOR2_X1 u_xor_module_287_U1 ( .A(n_xor_module_257_res), .B(
        n_reg_module_134_res), .Z(n_xor_module_287_res) );
  XOR2_X1 u_xor_module_288_U1 ( .A(n_xor_module_258_res), .B(
        n_reg_module_136_res), .Z(n_xor_module_288_res) );
  XOR2_X1 u_xor_module_289_U1 ( .A(n_xor_module_251_res), .B(
        n_xor_module_249_res), .Z(n_xor_module_289_res) );
  XOR2_X1 u_xor_module_290_U1 ( .A(n_xor_module_252_res), .B(
        n_xor_module_250_res), .Z(n_xor_module_290_res) );
  XOR2_X1 u_xor_module_291_U1 ( .A(n_xor_module_263_res), .B(
        n_xor_module_251_res), .Z(n_xor_module_291_res) );
  XOR2_X1 u_xor_module_292_U1 ( .A(n_xor_module_264_res), .B(
        n_xor_module_252_res), .Z(n_xor_module_292_res) );
  XOR2_X1 u_xor_module_293_U1 ( .A(n_xor_module_273_res), .B(
        n_xor_module_255_res), .Z(n_xor_module_293_res) );
  XOR2_X1 u_xor_module_294_U1 ( .A(n_xor_module_274_res), .B(
        n_xor_module_256_res), .Z(n_xor_module_294_res) );
  XOR2_X1 u_xor_module_295_U1 ( .A(n_xor_module_253_res), .B(
        n_xor_module_285_res), .Z(n_xor_module_295_res) );
  XOR2_X1 u_xor_module_296_U1 ( .A(n_xor_module_254_res), .B(
        n_xor_module_286_res), .Z(n_xor_module_296_res) );
  XOR2_X1 u_xor_module_297_U1 ( .A(n_xor_module_267_res), .B(
        n_xor_module_279_res), .Z(n_xor_module_297_res) );
  XOR2_X1 u_xor_module_298_U1 ( .A(n_xor_module_268_res), .B(
        n_xor_module_280_res), .Z(n_xor_module_298_res) );
  XOR2_X1 u_xor_module_299_U1 ( .A(n_xor_module_269_res), .B(
        n_xor_module_261_res), .Z(n_xor_module_299_res) );
  XOR2_X1 u_xor_module_300_U1 ( .A(n_xor_module_270_res), .B(
        n_xor_module_262_res), .Z(n_xor_module_300_res) );
  XOR2_X1 u_xor_module_301_U1 ( .A(n_xor_module_267_res), .B(
        n_xor_module_263_res), .Z(n_xor_module_301_res) );
  XOR2_X1 u_xor_module_302_U1 ( .A(n_xor_module_268_res), .B(
        n_xor_module_264_res), .Z(n_xor_module_302_res) );
  XOR2_X1 u_xor_module_303_U1 ( .A(n_xor_module_269_res), .B(
        n_xor_module_265_res), .Z(n_xor_module_303_res) );
  XOR2_X1 u_xor_module_304_U1 ( .A(n_xor_module_270_res), .B(
        n_xor_module_266_res), .Z(n_xor_module_304_res) );
  XOR2_X1 u_xor_module_305_U1 ( .A(n_xor_module_277_res), .B(
        n_xor_module_271_res), .Z(n_xor_module_305_res) );
  XOR2_X1 u_xor_module_306_U1 ( .A(n_xor_module_278_res), .B(
        n_xor_module_272_res), .Z(n_xor_module_306_res) );
  XOR2_X1 u_xor_module_307_U1 ( .A(n_xor_module_283_res), .B(
        n_xor_module_271_res), .Z(n_xor_module_307_res) );
  XOR2_X1 u_xor_module_308_U1 ( .A(n_xor_module_284_res), .B(
        n_xor_module_272_res), .Z(n_xor_module_308_res) );
  XOR2_X1 u_xor_module_309_U1 ( .A(n_xor_module_297_res), .B(
        n_xor_module_261_res), .Z(n_xor_module_309_res) );
  XOR2_X1 u_xor_module_310_U1 ( .A(n_xor_module_298_res), .B(
        n_xor_module_262_res), .Z(n_xor_module_310_res) );
  XOR2_X1 u_xor_module_311_U1 ( .A(n_xor_module_301_res), .B(
        n_xor_module_281_res), .Z(n_xor_module_311_res) );
  XOR2_X1 u_xor_module_312_U1 ( .A(n_xor_module_302_res), .B(
        n_xor_module_282_res), .Z(n_xor_module_312_res) );
  INV_X1 u_not_module_1_U1 ( .A(n_xor_module_311_res), .ZN(n_not_module_1_res)
         );
  XOR2_X1 u_xor_module_313_U1 ( .A(n_xor_module_305_res), .B(
        n_xor_module_287_res), .Z(n_xor_module_313_res) );
  XOR2_X1 u_xor_module_314_U1 ( .A(n_xor_module_306_res), .B(
        n_xor_module_288_res), .Z(n_xor_module_314_res) );
  INV_X1 u_not_module_2_U1 ( .A(n_xor_module_313_res), .ZN(n_not_module_2_res)
         );
  XOR2_X1 u_xor_module_315_U1 ( .A(n_xor_module_291_res), .B(
        n_xor_module_261_res), .Z(n_xor_module_315_res) );
  XOR2_X1 u_xor_module_316_U1 ( .A(n_xor_module_292_res), .B(
        n_xor_module_262_res), .Z(n_xor_module_316_res) );
  XOR2_X1 u_xor_module_317_U1 ( .A(n_xor_module_293_res), .B(
        n_xor_module_289_res), .Z(n_xor_module_317_res) );
  XOR2_X1 u_xor_module_318_U1 ( .A(n_xor_module_294_res), .B(
        n_xor_module_290_res), .Z(n_xor_module_318_res) );
  XOR2_X1 u_xor_module_319_U1 ( .A(n_xor_module_307_res), .B(
        n_xor_module_299_res), .Z(n_xor_module_319_res) );
  XOR2_X1 u_xor_module_320_U1 ( .A(n_xor_module_308_res), .B(
        n_xor_module_300_res), .Z(n_xor_module_320_res) );
  XOR2_X1 u_xor_module_321_U1 ( .A(n_xor_module_303_res), .B(
        n_xor_module_275_res), .Z(n_xor_module_321_res) );
  XOR2_X1 u_xor_module_322_U1 ( .A(n_xor_module_304_res), .B(
        n_xor_module_276_res), .Z(n_xor_module_322_res) );
  INV_X1 u_not_module_3_U1 ( .A(n_xor_module_321_res), .ZN(n_not_module_3_res)
         );
  XOR2_X1 u_xor_module_323_U1 ( .A(n_xor_module_295_res), .B(
        n_xor_module_261_res), .Z(n_xor_module_323_res) );
  XOR2_X1 u_xor_module_324_U1 ( .A(n_xor_module_296_res), .B(
        n_xor_module_262_res), .Z(n_xor_module_324_res) );
  INV_X1 u_not_module_4_U1 ( .A(n_xor_module_323_res), .ZN(n_not_module_4_res)
         );
  XOR2_X1 u_xor_module_325_U1 ( .A(io_k0_s0), .B(n_xor_module_309_res), .Z(
        io_o0_s0) );
  XOR2_X1 u_xor_module_326_U1 ( .A(io_k0_s1), .B(n_xor_module_310_res), .Z(
        io_o0_s1) );
  XOR2_X1 u_xor_module_327_U1 ( .A(io_k1_s0), .B(n_not_module_1_res), .Z(
        io_o1_s0) );
  XOR2_X1 u_xor_module_328_U1 ( .A(io_k1_s1), .B(n_xor_module_312_res), .Z(
        io_o1_s1) );
  XOR2_X1 u_xor_module_329_U1 ( .A(io_k2_s0), .B(n_not_module_2_res), .Z(
        io_o2_s0) );
  XOR2_X1 u_xor_module_330_U1 ( .A(io_k2_s1), .B(n_xor_module_314_res), .Z(
        io_o2_s1) );
  XOR2_X1 u_xor_module_331_U1 ( .A(io_k3_s0), .B(n_xor_module_315_res), .Z(
        io_o3_s0) );
  XOR2_X1 u_xor_module_332_U1 ( .A(io_k3_s1), .B(n_xor_module_316_res), .Z(
        io_o3_s1) );
  XOR2_X1 u_xor_module_333_U1 ( .A(io_k4_s0), .B(n_xor_module_317_res), .Z(
        io_o4_s0) );
  XOR2_X1 u_xor_module_334_U1 ( .A(io_k4_s1), .B(n_xor_module_318_res), .Z(
        io_o4_s1) );
  XOR2_X1 u_xor_module_335_U1 ( .A(io_k5_s0), .B(n_xor_module_319_res), .Z(
        io_o5_s0) );
  XOR2_X1 u_xor_module_336_U1 ( .A(io_k5_s1), .B(n_xor_module_320_res), .Z(
        io_o5_s1) );
  XOR2_X1 u_xor_module_337_U1 ( .A(io_k6_s0), .B(n_not_module_3_res), .Z(
        io_o6_s0) );
  XOR2_X1 u_xor_module_338_U1 ( .A(io_k6_s1), .B(n_xor_module_322_res), .Z(
        io_o6_s1) );
  XOR2_X1 u_xor_module_339_U1 ( .A(io_k7_s0), .B(n_not_module_4_res), .Z(
        io_o7_s0) );
  XOR2_X1 u_xor_module_340_U1 ( .A(io_k7_s1), .B(n_xor_module_324_res), .Z(
        io_o7_s1) );
endmodule

