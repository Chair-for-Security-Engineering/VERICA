
module KeyAddition ( clock, reset, io_state, io_key, io_out );
  input [3:0] io_state;
  input [3:0] io_key;
  output [3:0] io_out;
  input clock, reset;


  XOR2_X1 U5 ( .A(io_state[3]), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 U6 ( .A(io_state[2]), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 U7 ( .A(io_state[1]), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 U8 ( .A(io_state[0]), .B(io_key[0]), .Z(io_out[0]) );
endmodule

