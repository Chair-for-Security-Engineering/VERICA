
module CINI3 ( port_a_0, port_a_1, port_a_2, port_a_3, port_b_0, port_b_1, 
        port_b_2, port_b_3, port_c_0, port_c_1, port_c_2, port_c_3, 
        port_rand_ref, port_rand_mul, clk, reset );
  input [6:0] port_a_0;
  input [6:0] port_a_1;
  input [6:0] port_a_2;
  input [6:0] port_a_3;
  input [6:0] port_b_0;
  input [6:0] port_b_1;
  input [6:0] port_b_2;
  input [6:0] port_b_3;
  output [6:0] port_c_0;
  output [6:0] port_c_1;
  output [6:0] port_c_2;
  output [6:0] port_c_3;
  input [5:0] port_rand_ref;
  input [5:0] port_rand_mul;
  input clk, reset;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, ref_1_n76, ref_1_n75,
         ref_1_n74, ref_1_n73, ref_1_n72, ref_1_n71, ref_1_n70, ref_1_n69,
         ref_1_n68, ref_1_n67, ref_1_n66, ref_1_n65, ref_1_n64, ref_1_n63,
         ref_1_n62, ref_1_n61, ref_1_n60, ref_1_n59, ref_1_n58, ref_1_n57,
         ref_1_n56, ref_1_n55, ref_1_n54, ref_1_n53, ref_1_n52, ref_1_n51,
         ref_1_n50, ref_1_n49, ref_1_n48, ref_1_n47, ref_1_n46, ref_1_n45,
         ref_1_n44, ref_1_n43, ref_1_n42, ref_1_n41, ref_1_n40, ref_1_n39,
         ref_1_n38, ref_1_n37, ref_1_n36, ref_1_n35, ref_1_n34, ref_1_n33,
         ref_1_n32, ref_1_n31, ref_1_n30, ref_1_n29, ref_1_n28, ref_1_n27,
         ref_1_n26, ref_1_n25, ref_1_n24, ref_1_n23, ref_1_n22, ref_1_n21,
         ref_1_n20, ref_1_n19, ref_1_n18, ref_1_n17, ref_1_n16, ref_1_n15,
         ref_1_n14, ref_1_n13, ref_1_n12, ref_1_n11, ref_1_n10, ref_1_n9,
         ref_1_n8, ref_1_n7, ref_1_n6, ref_1_n5, ref_1_n4, ref_1_n3, ref_1_n2,
         ref_1_n1, ref_1_maj_223_port_o, ref_1_maj_222_port_o,
         ref_1_maj_221_port_o, ref_1_maj_220_port_o, ref_1_maj_219_port_o,
         ref_1_maj_218_port_o, ref_1_maj_217_port_o, ref_1_maj_216_port_o,
         ref_1_maj_215_port_o, ref_1_maj_214_port_o, ref_1_maj_213_port_o,
         ref_1_maj_212_port_o, ref_1_maj_211_port_o, ref_1_maj_210_port_o,
         ref_1_maj_209_port_o, ref_1_maj_208_port_o, ref_1_maj_207_port_o,
         ref_1_maj_206_port_o, ref_1_maj_205_port_o, ref_1_maj_204_port_o,
         ref_1_maj_203_port_o, ref_1_maj_202_port_o, ref_1_maj_201_port_o,
         ref_1_maj_200_port_o, ref_1_maj_199_port_o, ref_1_maj_198_port_o,
         ref_1_maj_197_port_o, ref_1_maj_196_port_o, ref_1_maj_195_port_o,
         ref_1_maj_194_port_o, ref_1_maj_193_port_o, ref_1_maj_192_port_o,
         ref_1_maj_191_port_o, ref_1_maj_190_port_o, ref_1_maj_189_port_o,
         ref_1_maj_188_port_o, ref_1_maj_187_port_o, ref_1_maj_186_port_o,
         ref_1_maj_185_port_o, ref_1_maj_184_port_o, ref_1_maj_183_port_o,
         ref_1_maj_182_port_o, ref_1_maj_181_port_o, ref_1_maj_180_port_o,
         ref_1_maj_179_port_o, ref_1_maj_178_port_o, ref_1_maj_177_port_o,
         ref_1_maj_176_port_o, ref_1_maj_175_port_o, ref_1_maj_174_port_o,
         ref_1_maj_173_port_o, ref_1_maj_172_port_o, ref_1_maj_171_port_o,
         ref_1_maj_170_port_o, ref_1_maj_169_port_o, ref_1_maj_168_port_o,
         ref_1_maj_167_port_o, ref_1_maj_166_port_o, ref_1_maj_165_port_o,
         ref_1_maj_164_port_o, ref_1_maj_163_port_o, ref_1_maj_162_port_o,
         ref_1_maj_161_port_o, ref_1_maj_160_port_o, ref_1_maj_159_port_o,
         ref_1_maj_158_port_o, ref_1_maj_157_port_o, ref_1_maj_156_port_o,
         ref_1_maj_155_port_o, ref_1_maj_154_port_o, ref_1_maj_153_port_o,
         ref_1_maj_152_port_o, ref_1_maj_151_port_o, ref_1_maj_150_port_o,
         ref_1_maj_149_port_o, ref_1_maj_148_port_o, ref_1_maj_147_port_o,
         ref_1_maj_146_port_o, ref_1_maj_145_port_o, ref_1_maj_144_port_o,
         ref_1_maj_143_port_o, ref_1_maj_142_port_o, ref_1_maj_141_port_o,
         ref_1_maj_140_port_o, ref_1_maj_139_port_o, ref_1_maj_138_port_o,
         ref_1_maj_137_port_o, ref_1_maj_136_port_o, ref_1_maj_135_port_o,
         ref_1_maj_134_port_o, ref_1_maj_133_port_o, ref_1_maj_132_port_o,
         ref_1_maj_131_port_o, ref_1_maj_130_port_o, ref_1_maj_129_port_o,
         ref_1_maj_128_port_o, ref_1_maj_127_port_o, ref_1_maj_126_port_o,
         ref_1_maj_125_port_o, ref_1_maj_124_port_o, ref_1_refreshed_3_0_,
         ref_1_refreshed_3_1_, ref_1_refreshed_3_2_, ref_1_refreshed_3_3_,
         ref_1_refreshed_3_4_, ref_1_refreshed_3_5_, ref_1_refreshed_3_6_,
         ref_1_maj_123_port_o, ref_1_maj_122_port_o, ref_1_maj_121_port_o,
         ref_1_maj_120_port_o, ref_1_refreshed_2_0_, ref_1_refreshed_2_1_,
         ref_1_refreshed_2_2_, ref_1_refreshed_2_3_, ref_1_refreshed_2_4_,
         ref_1_refreshed_2_5_, ref_1_refreshed_2_6_, ref_1_maj_119_port_o,
         ref_1_maj_118_port_o, ref_1_maj_117_port_o, ref_1_maj_116_port_o,
         ref_1_refreshed_1_0_, ref_1_refreshed_1_1_, ref_1_refreshed_1_2_,
         ref_1_refreshed_1_3_, ref_1_refreshed_1_4_, ref_1_refreshed_1_5_,
         ref_1_refreshed_1_6_, ref_1_maj_115_port_o, ref_1_maj_114_port_o,
         ref_1_maj_113_port_o, ref_1_maj_112_port_o, ref_1_refreshed_0_0_,
         ref_1_refreshed_0_1_, ref_1_refreshed_0_2_, ref_1_refreshed_0_3_,
         ref_1_refreshed_0_4_, ref_1_refreshed_0_5_, ref_1_refreshed_0_6_,
         ref_1_simpleXor_166_port_z, ref_1_simpleXor_165_port_z,
         ref_1_simpleXor_163_port_z, ref_1_simpleXor_162_port_z,
         ref_1_simpleXor_160_port_z, ref_1_simpleXor_159_port_z,
         ref_1_simpleXor_157_port_z, ref_1_simpleXor_156_port_z,
         ref_1_simpleXor_154_port_z, ref_1_simpleXor_153_port_z,
         ref_1_simpleXor_151_port_z, ref_1_simpleXor_150_port_z,
         ref_1_simpleXor_148_port_z, ref_1_simpleXor_147_port_z,
         ref_1_simpleXor_145_port_z, ref_1_simpleXor_144_port_z,
         ref_1_simpleXor_142_port_z, ref_1_simpleXor_141_port_z,
         ref_1_simpleXor_139_port_z, ref_1_simpleXor_138_port_z,
         ref_1_simpleXor_136_port_z, ref_1_simpleXor_135_port_z,
         ref_1_simpleXor_133_port_z, ref_1_simpleXor_132_port_z,
         ref_1_simpleXor_130_port_z, ref_1_simpleXor_129_port_z,
         ref_1_simpleXor_127_port_z, ref_1_simpleXor_126_port_z,
         ref_1_simpleXor_124_port_z, ref_1_simpleXor_123_port_z,
         ref_1_simpleXor_121_port_z, ref_1_simpleXor_120_port_z,
         ref_1_simpleXor_118_port_z, ref_1_simpleXor_117_port_z,
         ref_1_simpleXor_115_port_z, ref_1_simpleXor_114_port_z,
         ref_1_simpleXor_112_port_z, ref_1_simpleXor_111_port_z,
         ref_1_simpleXor_109_port_z, ref_1_simpleXor_108_port_z,
         ref_1_simpleXor_106_port_z, ref_1_simpleXor_105_port_z,
         ref_1_simpleXor_103_port_z, ref_1_simpleXor_102_port_z,
         ref_1_simpleXor_100_port_z, ref_1_simpleXor_99_port_z,
         ref_1_simpleXor_97_port_z, ref_1_simpleXor_96_port_z,
         ref_1_simpleXor_94_port_z, ref_1_simpleXor_93_port_z,
         ref_1_simpleXor_91_port_z, ref_1_simpleXor_90_port_z,
         ref_1_simpleXor_88_port_z, ref_1_simpleXor_87_port_z,
         ref_1_simpleXor_85_port_z, ref_1_simpleXor_84_port_z,
         ref_1_maj_112_n17, ref_1_maj_112_n16, ref_1_maj_112_n15,
         ref_1_maj_112_n14, ref_1_maj_112_n13, ref_1_maj_112_n12,
         ref_1_maj_112_n11, ref_1_maj_112_n10, ref_1_maj_112_n9,
         ref_1_maj_112_n8, ref_1_maj_112_n7, ref_1_maj_112_n6,
         ref_1_maj_112_n5, ref_1_maj_112_n4, ref_1_maj_112_n3,
         ref_1_maj_112_n2, ref_1_maj_112_n1, ref_1_maj_113_n34,
         ref_1_maj_113_n33, ref_1_maj_113_n32, ref_1_maj_113_n31,
         ref_1_maj_113_n30, ref_1_maj_113_n29, ref_1_maj_113_n28,
         ref_1_maj_113_n27, ref_1_maj_113_n26, ref_1_maj_113_n25,
         ref_1_maj_113_n24, ref_1_maj_113_n23, ref_1_maj_113_n22,
         ref_1_maj_113_n21, ref_1_maj_113_n20, ref_1_maj_113_n19,
         ref_1_maj_113_n18, ref_1_maj_114_n34, ref_1_maj_114_n33,
         ref_1_maj_114_n32, ref_1_maj_114_n31, ref_1_maj_114_n30,
         ref_1_maj_114_n29, ref_1_maj_114_n28, ref_1_maj_114_n27,
         ref_1_maj_114_n26, ref_1_maj_114_n25, ref_1_maj_114_n24,
         ref_1_maj_114_n23, ref_1_maj_114_n22, ref_1_maj_114_n21,
         ref_1_maj_114_n20, ref_1_maj_114_n19, ref_1_maj_114_n18,
         ref_1_maj_115_n34, ref_1_maj_115_n33, ref_1_maj_115_n32,
         ref_1_maj_115_n31, ref_1_maj_115_n30, ref_1_maj_115_n29,
         ref_1_maj_115_n28, ref_1_maj_115_n27, ref_1_maj_115_n26,
         ref_1_maj_115_n25, ref_1_maj_115_n24, ref_1_maj_115_n23,
         ref_1_maj_115_n22, ref_1_maj_115_n21, ref_1_maj_115_n20,
         ref_1_maj_115_n19, ref_1_maj_115_n18, ref_1_maj_116_n34,
         ref_1_maj_116_n33, ref_1_maj_116_n32, ref_1_maj_116_n31,
         ref_1_maj_116_n30, ref_1_maj_116_n29, ref_1_maj_116_n28,
         ref_1_maj_116_n27, ref_1_maj_116_n26, ref_1_maj_116_n25,
         ref_1_maj_116_n24, ref_1_maj_116_n23, ref_1_maj_116_n22,
         ref_1_maj_116_n21, ref_1_maj_116_n20, ref_1_maj_116_n19,
         ref_1_maj_116_n18, ref_1_maj_117_n34, ref_1_maj_117_n33,
         ref_1_maj_117_n32, ref_1_maj_117_n31, ref_1_maj_117_n30,
         ref_1_maj_117_n29, ref_1_maj_117_n28, ref_1_maj_117_n27,
         ref_1_maj_117_n26, ref_1_maj_117_n25, ref_1_maj_117_n24,
         ref_1_maj_117_n23, ref_1_maj_117_n22, ref_1_maj_117_n21,
         ref_1_maj_117_n20, ref_1_maj_117_n19, ref_1_maj_117_n18,
         ref_1_maj_118_n34, ref_1_maj_118_n33, ref_1_maj_118_n32,
         ref_1_maj_118_n31, ref_1_maj_118_n30, ref_1_maj_118_n29,
         ref_1_maj_118_n28, ref_1_maj_118_n27, ref_1_maj_118_n26,
         ref_1_maj_118_n25, ref_1_maj_118_n24, ref_1_maj_118_n23,
         ref_1_maj_118_n22, ref_1_maj_118_n21, ref_1_maj_118_n20,
         ref_1_maj_118_n19, ref_1_maj_118_n18, ref_1_maj_119_n34,
         ref_1_maj_119_n33, ref_1_maj_119_n32, ref_1_maj_119_n31,
         ref_1_maj_119_n30, ref_1_maj_119_n29, ref_1_maj_119_n28,
         ref_1_maj_119_n27, ref_1_maj_119_n26, ref_1_maj_119_n25,
         ref_1_maj_119_n24, ref_1_maj_119_n23, ref_1_maj_119_n22,
         ref_1_maj_119_n21, ref_1_maj_119_n20, ref_1_maj_119_n19,
         ref_1_maj_119_n18, ref_1_maj_120_n34, ref_1_maj_120_n33,
         ref_1_maj_120_n32, ref_1_maj_120_n31, ref_1_maj_120_n30,
         ref_1_maj_120_n29, ref_1_maj_120_n28, ref_1_maj_120_n27,
         ref_1_maj_120_n26, ref_1_maj_120_n25, ref_1_maj_120_n24,
         ref_1_maj_120_n23, ref_1_maj_120_n22, ref_1_maj_120_n21,
         ref_1_maj_120_n20, ref_1_maj_120_n19, ref_1_maj_120_n18,
         ref_1_maj_121_n34, ref_1_maj_121_n33, ref_1_maj_121_n32,
         ref_1_maj_121_n31, ref_1_maj_121_n30, ref_1_maj_121_n29,
         ref_1_maj_121_n28, ref_1_maj_121_n27, ref_1_maj_121_n26,
         ref_1_maj_121_n25, ref_1_maj_121_n24, ref_1_maj_121_n23,
         ref_1_maj_121_n22, ref_1_maj_121_n21, ref_1_maj_121_n20,
         ref_1_maj_121_n19, ref_1_maj_121_n18, ref_1_maj_122_n34,
         ref_1_maj_122_n33, ref_1_maj_122_n32, ref_1_maj_122_n31,
         ref_1_maj_122_n30, ref_1_maj_122_n29, ref_1_maj_122_n28,
         ref_1_maj_122_n27, ref_1_maj_122_n26, ref_1_maj_122_n25,
         ref_1_maj_122_n24, ref_1_maj_122_n23, ref_1_maj_122_n22,
         ref_1_maj_122_n21, ref_1_maj_122_n20, ref_1_maj_122_n19,
         ref_1_maj_122_n18, ref_1_maj_123_n34, ref_1_maj_123_n33,
         ref_1_maj_123_n32, ref_1_maj_123_n31, ref_1_maj_123_n30,
         ref_1_maj_123_n29, ref_1_maj_123_n28, ref_1_maj_123_n27,
         ref_1_maj_123_n26, ref_1_maj_123_n25, ref_1_maj_123_n24,
         ref_1_maj_123_n23, ref_1_maj_123_n22, ref_1_maj_123_n21,
         ref_1_maj_123_n20, ref_1_maj_123_n19, ref_1_maj_123_n18,
         ref_1_maj_124_n34, ref_1_maj_124_n33, ref_1_maj_124_n32,
         ref_1_maj_124_n31, ref_1_maj_124_n30, ref_1_maj_124_n29,
         ref_1_maj_124_n28, ref_1_maj_124_n27, ref_1_maj_124_n26,
         ref_1_maj_124_n25, ref_1_maj_124_n24, ref_1_maj_124_n23,
         ref_1_maj_124_n22, ref_1_maj_124_n21, ref_1_maj_124_n20,
         ref_1_maj_124_n19, ref_1_maj_124_n18, ref_1_maj_125_n34,
         ref_1_maj_125_n33, ref_1_maj_125_n32, ref_1_maj_125_n31,
         ref_1_maj_125_n30, ref_1_maj_125_n29, ref_1_maj_125_n28,
         ref_1_maj_125_n27, ref_1_maj_125_n26, ref_1_maj_125_n25,
         ref_1_maj_125_n24, ref_1_maj_125_n23, ref_1_maj_125_n22,
         ref_1_maj_125_n21, ref_1_maj_125_n20, ref_1_maj_125_n19,
         ref_1_maj_125_n18, ref_1_maj_126_n34, ref_1_maj_126_n33,
         ref_1_maj_126_n32, ref_1_maj_126_n31, ref_1_maj_126_n30,
         ref_1_maj_126_n29, ref_1_maj_126_n28, ref_1_maj_126_n27,
         ref_1_maj_126_n26, ref_1_maj_126_n25, ref_1_maj_126_n24,
         ref_1_maj_126_n23, ref_1_maj_126_n22, ref_1_maj_126_n21,
         ref_1_maj_126_n20, ref_1_maj_126_n19, ref_1_maj_126_n18,
         ref_1_maj_127_n34, ref_1_maj_127_n33, ref_1_maj_127_n32,
         ref_1_maj_127_n31, ref_1_maj_127_n30, ref_1_maj_127_n29,
         ref_1_maj_127_n28, ref_1_maj_127_n27, ref_1_maj_127_n26,
         ref_1_maj_127_n25, ref_1_maj_127_n24, ref_1_maj_127_n23,
         ref_1_maj_127_n22, ref_1_maj_127_n21, ref_1_maj_127_n20,
         ref_1_maj_127_n19, ref_1_maj_127_n18, ref_1_maj_128_n34,
         ref_1_maj_128_n33, ref_1_maj_128_n32, ref_1_maj_128_n31,
         ref_1_maj_128_n30, ref_1_maj_128_n29, ref_1_maj_128_n28,
         ref_1_maj_128_n27, ref_1_maj_128_n26, ref_1_maj_128_n25,
         ref_1_maj_128_n24, ref_1_maj_128_n23, ref_1_maj_128_n22,
         ref_1_maj_128_n21, ref_1_maj_128_n20, ref_1_maj_128_n19,
         ref_1_maj_128_n18, ref_1_maj_129_n34, ref_1_maj_129_n33,
         ref_1_maj_129_n32, ref_1_maj_129_n31, ref_1_maj_129_n30,
         ref_1_maj_129_n29, ref_1_maj_129_n28, ref_1_maj_129_n27,
         ref_1_maj_129_n26, ref_1_maj_129_n25, ref_1_maj_129_n24,
         ref_1_maj_129_n23, ref_1_maj_129_n22, ref_1_maj_129_n21,
         ref_1_maj_129_n20, ref_1_maj_129_n19, ref_1_maj_129_n18,
         ref_1_maj_130_n34, ref_1_maj_130_n33, ref_1_maj_130_n32,
         ref_1_maj_130_n31, ref_1_maj_130_n30, ref_1_maj_130_n29,
         ref_1_maj_130_n28, ref_1_maj_130_n27, ref_1_maj_130_n26,
         ref_1_maj_130_n25, ref_1_maj_130_n24, ref_1_maj_130_n23,
         ref_1_maj_130_n22, ref_1_maj_130_n21, ref_1_maj_130_n20,
         ref_1_maj_130_n19, ref_1_maj_130_n18, ref_1_maj_131_n34,
         ref_1_maj_131_n33, ref_1_maj_131_n32, ref_1_maj_131_n31,
         ref_1_maj_131_n30, ref_1_maj_131_n29, ref_1_maj_131_n28,
         ref_1_maj_131_n27, ref_1_maj_131_n26, ref_1_maj_131_n25,
         ref_1_maj_131_n24, ref_1_maj_131_n23, ref_1_maj_131_n22,
         ref_1_maj_131_n21, ref_1_maj_131_n20, ref_1_maj_131_n19,
         ref_1_maj_131_n18, ref_1_maj_132_n34, ref_1_maj_132_n33,
         ref_1_maj_132_n32, ref_1_maj_132_n31, ref_1_maj_132_n30,
         ref_1_maj_132_n29, ref_1_maj_132_n28, ref_1_maj_132_n27,
         ref_1_maj_132_n26, ref_1_maj_132_n25, ref_1_maj_132_n24,
         ref_1_maj_132_n23, ref_1_maj_132_n22, ref_1_maj_132_n21,
         ref_1_maj_132_n20, ref_1_maj_132_n19, ref_1_maj_132_n18,
         ref_1_maj_133_n34, ref_1_maj_133_n33, ref_1_maj_133_n32,
         ref_1_maj_133_n31, ref_1_maj_133_n30, ref_1_maj_133_n29,
         ref_1_maj_133_n28, ref_1_maj_133_n27, ref_1_maj_133_n26,
         ref_1_maj_133_n25, ref_1_maj_133_n24, ref_1_maj_133_n23,
         ref_1_maj_133_n22, ref_1_maj_133_n21, ref_1_maj_133_n20,
         ref_1_maj_133_n19, ref_1_maj_133_n18, ref_1_maj_134_n34,
         ref_1_maj_134_n33, ref_1_maj_134_n32, ref_1_maj_134_n31,
         ref_1_maj_134_n30, ref_1_maj_134_n29, ref_1_maj_134_n28,
         ref_1_maj_134_n27, ref_1_maj_134_n26, ref_1_maj_134_n25,
         ref_1_maj_134_n24, ref_1_maj_134_n23, ref_1_maj_134_n22,
         ref_1_maj_134_n21, ref_1_maj_134_n20, ref_1_maj_134_n19,
         ref_1_maj_134_n18, ref_1_maj_135_n34, ref_1_maj_135_n33,
         ref_1_maj_135_n32, ref_1_maj_135_n31, ref_1_maj_135_n30,
         ref_1_maj_135_n29, ref_1_maj_135_n28, ref_1_maj_135_n27,
         ref_1_maj_135_n26, ref_1_maj_135_n25, ref_1_maj_135_n24,
         ref_1_maj_135_n23, ref_1_maj_135_n22, ref_1_maj_135_n21,
         ref_1_maj_135_n20, ref_1_maj_135_n19, ref_1_maj_135_n18,
         ref_1_maj_136_n34, ref_1_maj_136_n33, ref_1_maj_136_n32,
         ref_1_maj_136_n31, ref_1_maj_136_n30, ref_1_maj_136_n29,
         ref_1_maj_136_n28, ref_1_maj_136_n27, ref_1_maj_136_n26,
         ref_1_maj_136_n25, ref_1_maj_136_n24, ref_1_maj_136_n23,
         ref_1_maj_136_n22, ref_1_maj_136_n21, ref_1_maj_136_n20,
         ref_1_maj_136_n19, ref_1_maj_136_n18, ref_1_maj_137_n34,
         ref_1_maj_137_n33, ref_1_maj_137_n32, ref_1_maj_137_n31,
         ref_1_maj_137_n30, ref_1_maj_137_n29, ref_1_maj_137_n28,
         ref_1_maj_137_n27, ref_1_maj_137_n26, ref_1_maj_137_n25,
         ref_1_maj_137_n24, ref_1_maj_137_n23, ref_1_maj_137_n22,
         ref_1_maj_137_n21, ref_1_maj_137_n20, ref_1_maj_137_n19,
         ref_1_maj_137_n18, ref_1_maj_138_n34, ref_1_maj_138_n33,
         ref_1_maj_138_n32, ref_1_maj_138_n31, ref_1_maj_138_n30,
         ref_1_maj_138_n29, ref_1_maj_138_n28, ref_1_maj_138_n27,
         ref_1_maj_138_n26, ref_1_maj_138_n25, ref_1_maj_138_n24,
         ref_1_maj_138_n23, ref_1_maj_138_n22, ref_1_maj_138_n21,
         ref_1_maj_138_n20, ref_1_maj_138_n19, ref_1_maj_138_n18,
         ref_1_maj_139_n34, ref_1_maj_139_n33, ref_1_maj_139_n32,
         ref_1_maj_139_n31, ref_1_maj_139_n30, ref_1_maj_139_n29,
         ref_1_maj_139_n28, ref_1_maj_139_n27, ref_1_maj_139_n26,
         ref_1_maj_139_n25, ref_1_maj_139_n24, ref_1_maj_139_n23,
         ref_1_maj_139_n22, ref_1_maj_139_n21, ref_1_maj_139_n20,
         ref_1_maj_139_n19, ref_1_maj_139_n18, ref_1_maj_140_n34,
         ref_1_maj_140_n33, ref_1_maj_140_n32, ref_1_maj_140_n31,
         ref_1_maj_140_n30, ref_1_maj_140_n29, ref_1_maj_140_n28,
         ref_1_maj_140_n27, ref_1_maj_140_n26, ref_1_maj_140_n25,
         ref_1_maj_140_n24, ref_1_maj_140_n23, ref_1_maj_140_n22,
         ref_1_maj_140_n21, ref_1_maj_140_n20, ref_1_maj_140_n19,
         ref_1_maj_140_n18, ref_1_maj_141_n34, ref_1_maj_141_n33,
         ref_1_maj_141_n32, ref_1_maj_141_n31, ref_1_maj_141_n30,
         ref_1_maj_141_n29, ref_1_maj_141_n28, ref_1_maj_141_n27,
         ref_1_maj_141_n26, ref_1_maj_141_n25, ref_1_maj_141_n24,
         ref_1_maj_141_n23, ref_1_maj_141_n22, ref_1_maj_141_n21,
         ref_1_maj_141_n20, ref_1_maj_141_n19, ref_1_maj_141_n18,
         ref_1_maj_142_n34, ref_1_maj_142_n33, ref_1_maj_142_n32,
         ref_1_maj_142_n31, ref_1_maj_142_n30, ref_1_maj_142_n29,
         ref_1_maj_142_n28, ref_1_maj_142_n27, ref_1_maj_142_n26,
         ref_1_maj_142_n25, ref_1_maj_142_n24, ref_1_maj_142_n23,
         ref_1_maj_142_n22, ref_1_maj_142_n21, ref_1_maj_142_n20,
         ref_1_maj_142_n19, ref_1_maj_142_n18, ref_1_maj_143_n34,
         ref_1_maj_143_n33, ref_1_maj_143_n32, ref_1_maj_143_n31,
         ref_1_maj_143_n30, ref_1_maj_143_n29, ref_1_maj_143_n28,
         ref_1_maj_143_n27, ref_1_maj_143_n26, ref_1_maj_143_n25,
         ref_1_maj_143_n24, ref_1_maj_143_n23, ref_1_maj_143_n22,
         ref_1_maj_143_n21, ref_1_maj_143_n20, ref_1_maj_143_n19,
         ref_1_maj_143_n18, ref_1_maj_144_n34, ref_1_maj_144_n33,
         ref_1_maj_144_n32, ref_1_maj_144_n31, ref_1_maj_144_n30,
         ref_1_maj_144_n29, ref_1_maj_144_n28, ref_1_maj_144_n27,
         ref_1_maj_144_n26, ref_1_maj_144_n25, ref_1_maj_144_n24,
         ref_1_maj_144_n23, ref_1_maj_144_n22, ref_1_maj_144_n21,
         ref_1_maj_144_n20, ref_1_maj_144_n19, ref_1_maj_144_n18,
         ref_1_maj_145_n34, ref_1_maj_145_n33, ref_1_maj_145_n32,
         ref_1_maj_145_n31, ref_1_maj_145_n30, ref_1_maj_145_n29,
         ref_1_maj_145_n28, ref_1_maj_145_n27, ref_1_maj_145_n26,
         ref_1_maj_145_n25, ref_1_maj_145_n24, ref_1_maj_145_n23,
         ref_1_maj_145_n22, ref_1_maj_145_n21, ref_1_maj_145_n20,
         ref_1_maj_145_n19, ref_1_maj_145_n18, ref_1_maj_146_n34,
         ref_1_maj_146_n33, ref_1_maj_146_n32, ref_1_maj_146_n31,
         ref_1_maj_146_n30, ref_1_maj_146_n29, ref_1_maj_146_n28,
         ref_1_maj_146_n27, ref_1_maj_146_n26, ref_1_maj_146_n25,
         ref_1_maj_146_n24, ref_1_maj_146_n23, ref_1_maj_146_n22,
         ref_1_maj_146_n21, ref_1_maj_146_n20, ref_1_maj_146_n19,
         ref_1_maj_146_n18, ref_1_maj_147_n34, ref_1_maj_147_n33,
         ref_1_maj_147_n32, ref_1_maj_147_n31, ref_1_maj_147_n30,
         ref_1_maj_147_n29, ref_1_maj_147_n28, ref_1_maj_147_n27,
         ref_1_maj_147_n26, ref_1_maj_147_n25, ref_1_maj_147_n24,
         ref_1_maj_147_n23, ref_1_maj_147_n22, ref_1_maj_147_n21,
         ref_1_maj_147_n20, ref_1_maj_147_n19, ref_1_maj_147_n18,
         ref_1_maj_148_n34, ref_1_maj_148_n33, ref_1_maj_148_n32,
         ref_1_maj_148_n31, ref_1_maj_148_n30, ref_1_maj_148_n29,
         ref_1_maj_148_n28, ref_1_maj_148_n27, ref_1_maj_148_n26,
         ref_1_maj_148_n25, ref_1_maj_148_n24, ref_1_maj_148_n23,
         ref_1_maj_148_n22, ref_1_maj_148_n21, ref_1_maj_148_n20,
         ref_1_maj_148_n19, ref_1_maj_148_n18, ref_1_maj_149_n34,
         ref_1_maj_149_n33, ref_1_maj_149_n32, ref_1_maj_149_n31,
         ref_1_maj_149_n30, ref_1_maj_149_n29, ref_1_maj_149_n28,
         ref_1_maj_149_n27, ref_1_maj_149_n26, ref_1_maj_149_n25,
         ref_1_maj_149_n24, ref_1_maj_149_n23, ref_1_maj_149_n22,
         ref_1_maj_149_n21, ref_1_maj_149_n20, ref_1_maj_149_n19,
         ref_1_maj_149_n18, ref_1_maj_150_n34, ref_1_maj_150_n33,
         ref_1_maj_150_n32, ref_1_maj_150_n31, ref_1_maj_150_n30,
         ref_1_maj_150_n29, ref_1_maj_150_n28, ref_1_maj_150_n27,
         ref_1_maj_150_n26, ref_1_maj_150_n25, ref_1_maj_150_n24,
         ref_1_maj_150_n23, ref_1_maj_150_n22, ref_1_maj_150_n21,
         ref_1_maj_150_n20, ref_1_maj_150_n19, ref_1_maj_150_n18,
         ref_1_maj_151_n34, ref_1_maj_151_n33, ref_1_maj_151_n32,
         ref_1_maj_151_n31, ref_1_maj_151_n30, ref_1_maj_151_n29,
         ref_1_maj_151_n28, ref_1_maj_151_n27, ref_1_maj_151_n26,
         ref_1_maj_151_n25, ref_1_maj_151_n24, ref_1_maj_151_n23,
         ref_1_maj_151_n22, ref_1_maj_151_n21, ref_1_maj_151_n20,
         ref_1_maj_151_n19, ref_1_maj_151_n18, ref_1_maj_152_n34,
         ref_1_maj_152_n33, ref_1_maj_152_n32, ref_1_maj_152_n31,
         ref_1_maj_152_n30, ref_1_maj_152_n29, ref_1_maj_152_n28,
         ref_1_maj_152_n27, ref_1_maj_152_n26, ref_1_maj_152_n25,
         ref_1_maj_152_n24, ref_1_maj_152_n23, ref_1_maj_152_n22,
         ref_1_maj_152_n21, ref_1_maj_152_n20, ref_1_maj_152_n19,
         ref_1_maj_152_n18, ref_1_maj_153_n34, ref_1_maj_153_n33,
         ref_1_maj_153_n32, ref_1_maj_153_n31, ref_1_maj_153_n30,
         ref_1_maj_153_n29, ref_1_maj_153_n28, ref_1_maj_153_n27,
         ref_1_maj_153_n26, ref_1_maj_153_n25, ref_1_maj_153_n24,
         ref_1_maj_153_n23, ref_1_maj_153_n22, ref_1_maj_153_n21,
         ref_1_maj_153_n20, ref_1_maj_153_n19, ref_1_maj_153_n18,
         ref_1_maj_154_n34, ref_1_maj_154_n33, ref_1_maj_154_n32,
         ref_1_maj_154_n31, ref_1_maj_154_n30, ref_1_maj_154_n29,
         ref_1_maj_154_n28, ref_1_maj_154_n27, ref_1_maj_154_n26,
         ref_1_maj_154_n25, ref_1_maj_154_n24, ref_1_maj_154_n23,
         ref_1_maj_154_n22, ref_1_maj_154_n21, ref_1_maj_154_n20,
         ref_1_maj_154_n19, ref_1_maj_154_n18, ref_1_maj_155_n34,
         ref_1_maj_155_n33, ref_1_maj_155_n32, ref_1_maj_155_n31,
         ref_1_maj_155_n30, ref_1_maj_155_n29, ref_1_maj_155_n28,
         ref_1_maj_155_n27, ref_1_maj_155_n26, ref_1_maj_155_n25,
         ref_1_maj_155_n24, ref_1_maj_155_n23, ref_1_maj_155_n22,
         ref_1_maj_155_n21, ref_1_maj_155_n20, ref_1_maj_155_n19,
         ref_1_maj_155_n18, ref_1_maj_156_n34, ref_1_maj_156_n33,
         ref_1_maj_156_n32, ref_1_maj_156_n31, ref_1_maj_156_n30,
         ref_1_maj_156_n29, ref_1_maj_156_n28, ref_1_maj_156_n27,
         ref_1_maj_156_n26, ref_1_maj_156_n25, ref_1_maj_156_n24,
         ref_1_maj_156_n23, ref_1_maj_156_n22, ref_1_maj_156_n21,
         ref_1_maj_156_n20, ref_1_maj_156_n19, ref_1_maj_156_n18,
         ref_1_maj_157_n34, ref_1_maj_157_n33, ref_1_maj_157_n32,
         ref_1_maj_157_n31, ref_1_maj_157_n30, ref_1_maj_157_n29,
         ref_1_maj_157_n28, ref_1_maj_157_n27, ref_1_maj_157_n26,
         ref_1_maj_157_n25, ref_1_maj_157_n24, ref_1_maj_157_n23,
         ref_1_maj_157_n22, ref_1_maj_157_n21, ref_1_maj_157_n20,
         ref_1_maj_157_n19, ref_1_maj_157_n18, ref_1_maj_158_n34,
         ref_1_maj_158_n33, ref_1_maj_158_n32, ref_1_maj_158_n31,
         ref_1_maj_158_n30, ref_1_maj_158_n29, ref_1_maj_158_n28,
         ref_1_maj_158_n27, ref_1_maj_158_n26, ref_1_maj_158_n25,
         ref_1_maj_158_n24, ref_1_maj_158_n23, ref_1_maj_158_n22,
         ref_1_maj_158_n21, ref_1_maj_158_n20, ref_1_maj_158_n19,
         ref_1_maj_158_n18, ref_1_maj_159_n34, ref_1_maj_159_n33,
         ref_1_maj_159_n32, ref_1_maj_159_n31, ref_1_maj_159_n30,
         ref_1_maj_159_n29, ref_1_maj_159_n28, ref_1_maj_159_n27,
         ref_1_maj_159_n26, ref_1_maj_159_n25, ref_1_maj_159_n24,
         ref_1_maj_159_n23, ref_1_maj_159_n22, ref_1_maj_159_n21,
         ref_1_maj_159_n20, ref_1_maj_159_n19, ref_1_maj_159_n18,
         ref_1_maj_160_n34, ref_1_maj_160_n33, ref_1_maj_160_n32,
         ref_1_maj_160_n31, ref_1_maj_160_n30, ref_1_maj_160_n29,
         ref_1_maj_160_n28, ref_1_maj_160_n27, ref_1_maj_160_n26,
         ref_1_maj_160_n25, ref_1_maj_160_n24, ref_1_maj_160_n23,
         ref_1_maj_160_n22, ref_1_maj_160_n21, ref_1_maj_160_n20,
         ref_1_maj_160_n19, ref_1_maj_160_n18, ref_1_maj_161_n34,
         ref_1_maj_161_n33, ref_1_maj_161_n32, ref_1_maj_161_n31,
         ref_1_maj_161_n30, ref_1_maj_161_n29, ref_1_maj_161_n28,
         ref_1_maj_161_n27, ref_1_maj_161_n26, ref_1_maj_161_n25,
         ref_1_maj_161_n24, ref_1_maj_161_n23, ref_1_maj_161_n22,
         ref_1_maj_161_n21, ref_1_maj_161_n20, ref_1_maj_161_n19,
         ref_1_maj_161_n18, ref_1_maj_162_n34, ref_1_maj_162_n33,
         ref_1_maj_162_n32, ref_1_maj_162_n31, ref_1_maj_162_n30,
         ref_1_maj_162_n29, ref_1_maj_162_n28, ref_1_maj_162_n27,
         ref_1_maj_162_n26, ref_1_maj_162_n25, ref_1_maj_162_n24,
         ref_1_maj_162_n23, ref_1_maj_162_n22, ref_1_maj_162_n21,
         ref_1_maj_162_n20, ref_1_maj_162_n19, ref_1_maj_162_n18,
         ref_1_maj_163_n34, ref_1_maj_163_n33, ref_1_maj_163_n32,
         ref_1_maj_163_n31, ref_1_maj_163_n30, ref_1_maj_163_n29,
         ref_1_maj_163_n28, ref_1_maj_163_n27, ref_1_maj_163_n26,
         ref_1_maj_163_n25, ref_1_maj_163_n24, ref_1_maj_163_n23,
         ref_1_maj_163_n22, ref_1_maj_163_n21, ref_1_maj_163_n20,
         ref_1_maj_163_n19, ref_1_maj_163_n18, ref_1_maj_164_n34,
         ref_1_maj_164_n33, ref_1_maj_164_n32, ref_1_maj_164_n31,
         ref_1_maj_164_n30, ref_1_maj_164_n29, ref_1_maj_164_n28,
         ref_1_maj_164_n27, ref_1_maj_164_n26, ref_1_maj_164_n25,
         ref_1_maj_164_n24, ref_1_maj_164_n23, ref_1_maj_164_n22,
         ref_1_maj_164_n21, ref_1_maj_164_n20, ref_1_maj_164_n19,
         ref_1_maj_164_n18, ref_1_maj_165_n34, ref_1_maj_165_n33,
         ref_1_maj_165_n32, ref_1_maj_165_n31, ref_1_maj_165_n30,
         ref_1_maj_165_n29, ref_1_maj_165_n28, ref_1_maj_165_n27,
         ref_1_maj_165_n26, ref_1_maj_165_n25, ref_1_maj_165_n24,
         ref_1_maj_165_n23, ref_1_maj_165_n22, ref_1_maj_165_n21,
         ref_1_maj_165_n20, ref_1_maj_165_n19, ref_1_maj_165_n18,
         ref_1_maj_166_n34, ref_1_maj_166_n33, ref_1_maj_166_n32,
         ref_1_maj_166_n31, ref_1_maj_166_n30, ref_1_maj_166_n29,
         ref_1_maj_166_n28, ref_1_maj_166_n27, ref_1_maj_166_n26,
         ref_1_maj_166_n25, ref_1_maj_166_n24, ref_1_maj_166_n23,
         ref_1_maj_166_n22, ref_1_maj_166_n21, ref_1_maj_166_n20,
         ref_1_maj_166_n19, ref_1_maj_166_n18, ref_1_maj_167_n34,
         ref_1_maj_167_n33, ref_1_maj_167_n32, ref_1_maj_167_n31,
         ref_1_maj_167_n30, ref_1_maj_167_n29, ref_1_maj_167_n28,
         ref_1_maj_167_n27, ref_1_maj_167_n26, ref_1_maj_167_n25,
         ref_1_maj_167_n24, ref_1_maj_167_n23, ref_1_maj_167_n22,
         ref_1_maj_167_n21, ref_1_maj_167_n20, ref_1_maj_167_n19,
         ref_1_maj_167_n18, ref_1_maj_168_n34, ref_1_maj_168_n33,
         ref_1_maj_168_n32, ref_1_maj_168_n31, ref_1_maj_168_n30,
         ref_1_maj_168_n29, ref_1_maj_168_n28, ref_1_maj_168_n27,
         ref_1_maj_168_n26, ref_1_maj_168_n25, ref_1_maj_168_n24,
         ref_1_maj_168_n23, ref_1_maj_168_n22, ref_1_maj_168_n21,
         ref_1_maj_168_n20, ref_1_maj_168_n19, ref_1_maj_168_n18,
         ref_1_maj_169_n34, ref_1_maj_169_n33, ref_1_maj_169_n32,
         ref_1_maj_169_n31, ref_1_maj_169_n30, ref_1_maj_169_n29,
         ref_1_maj_169_n28, ref_1_maj_169_n27, ref_1_maj_169_n26,
         ref_1_maj_169_n25, ref_1_maj_169_n24, ref_1_maj_169_n23,
         ref_1_maj_169_n22, ref_1_maj_169_n21, ref_1_maj_169_n20,
         ref_1_maj_169_n19, ref_1_maj_169_n18, ref_1_maj_170_n34,
         ref_1_maj_170_n33, ref_1_maj_170_n32, ref_1_maj_170_n31,
         ref_1_maj_170_n30, ref_1_maj_170_n29, ref_1_maj_170_n28,
         ref_1_maj_170_n27, ref_1_maj_170_n26, ref_1_maj_170_n25,
         ref_1_maj_170_n24, ref_1_maj_170_n23, ref_1_maj_170_n22,
         ref_1_maj_170_n21, ref_1_maj_170_n20, ref_1_maj_170_n19,
         ref_1_maj_170_n18, ref_1_maj_171_n34, ref_1_maj_171_n33,
         ref_1_maj_171_n32, ref_1_maj_171_n31, ref_1_maj_171_n30,
         ref_1_maj_171_n29, ref_1_maj_171_n28, ref_1_maj_171_n27,
         ref_1_maj_171_n26, ref_1_maj_171_n25, ref_1_maj_171_n24,
         ref_1_maj_171_n23, ref_1_maj_171_n22, ref_1_maj_171_n21,
         ref_1_maj_171_n20, ref_1_maj_171_n19, ref_1_maj_171_n18,
         ref_1_maj_172_n34, ref_1_maj_172_n33, ref_1_maj_172_n32,
         ref_1_maj_172_n31, ref_1_maj_172_n30, ref_1_maj_172_n29,
         ref_1_maj_172_n28, ref_1_maj_172_n27, ref_1_maj_172_n26,
         ref_1_maj_172_n25, ref_1_maj_172_n24, ref_1_maj_172_n23,
         ref_1_maj_172_n22, ref_1_maj_172_n21, ref_1_maj_172_n20,
         ref_1_maj_172_n19, ref_1_maj_172_n18, ref_1_maj_173_n34,
         ref_1_maj_173_n33, ref_1_maj_173_n32, ref_1_maj_173_n31,
         ref_1_maj_173_n30, ref_1_maj_173_n29, ref_1_maj_173_n28,
         ref_1_maj_173_n27, ref_1_maj_173_n26, ref_1_maj_173_n25,
         ref_1_maj_173_n24, ref_1_maj_173_n23, ref_1_maj_173_n22,
         ref_1_maj_173_n21, ref_1_maj_173_n20, ref_1_maj_173_n19,
         ref_1_maj_173_n18, ref_1_maj_174_n34, ref_1_maj_174_n33,
         ref_1_maj_174_n32, ref_1_maj_174_n31, ref_1_maj_174_n30,
         ref_1_maj_174_n29, ref_1_maj_174_n28, ref_1_maj_174_n27,
         ref_1_maj_174_n26, ref_1_maj_174_n25, ref_1_maj_174_n24,
         ref_1_maj_174_n23, ref_1_maj_174_n22, ref_1_maj_174_n21,
         ref_1_maj_174_n20, ref_1_maj_174_n19, ref_1_maj_174_n18,
         ref_1_maj_175_n34, ref_1_maj_175_n33, ref_1_maj_175_n32,
         ref_1_maj_175_n31, ref_1_maj_175_n30, ref_1_maj_175_n29,
         ref_1_maj_175_n28, ref_1_maj_175_n27, ref_1_maj_175_n26,
         ref_1_maj_175_n25, ref_1_maj_175_n24, ref_1_maj_175_n23,
         ref_1_maj_175_n22, ref_1_maj_175_n21, ref_1_maj_175_n20,
         ref_1_maj_175_n19, ref_1_maj_175_n18, ref_1_maj_176_n34,
         ref_1_maj_176_n33, ref_1_maj_176_n32, ref_1_maj_176_n31,
         ref_1_maj_176_n30, ref_1_maj_176_n29, ref_1_maj_176_n28,
         ref_1_maj_176_n27, ref_1_maj_176_n26, ref_1_maj_176_n25,
         ref_1_maj_176_n24, ref_1_maj_176_n23, ref_1_maj_176_n22,
         ref_1_maj_176_n21, ref_1_maj_176_n20, ref_1_maj_176_n19,
         ref_1_maj_176_n18, ref_1_maj_177_n34, ref_1_maj_177_n33,
         ref_1_maj_177_n32, ref_1_maj_177_n31, ref_1_maj_177_n30,
         ref_1_maj_177_n29, ref_1_maj_177_n28, ref_1_maj_177_n27,
         ref_1_maj_177_n26, ref_1_maj_177_n25, ref_1_maj_177_n24,
         ref_1_maj_177_n23, ref_1_maj_177_n22, ref_1_maj_177_n21,
         ref_1_maj_177_n20, ref_1_maj_177_n19, ref_1_maj_177_n18,
         ref_1_maj_178_n34, ref_1_maj_178_n33, ref_1_maj_178_n32,
         ref_1_maj_178_n31, ref_1_maj_178_n30, ref_1_maj_178_n29,
         ref_1_maj_178_n28, ref_1_maj_178_n27, ref_1_maj_178_n26,
         ref_1_maj_178_n25, ref_1_maj_178_n24, ref_1_maj_178_n23,
         ref_1_maj_178_n22, ref_1_maj_178_n21, ref_1_maj_178_n20,
         ref_1_maj_178_n19, ref_1_maj_178_n18, ref_1_maj_179_n34,
         ref_1_maj_179_n33, ref_1_maj_179_n32, ref_1_maj_179_n31,
         ref_1_maj_179_n30, ref_1_maj_179_n29, ref_1_maj_179_n28,
         ref_1_maj_179_n27, ref_1_maj_179_n26, ref_1_maj_179_n25,
         ref_1_maj_179_n24, ref_1_maj_179_n23, ref_1_maj_179_n22,
         ref_1_maj_179_n21, ref_1_maj_179_n20, ref_1_maj_179_n19,
         ref_1_maj_179_n18, ref_1_maj_180_n34, ref_1_maj_180_n33,
         ref_1_maj_180_n32, ref_1_maj_180_n31, ref_1_maj_180_n30,
         ref_1_maj_180_n29, ref_1_maj_180_n28, ref_1_maj_180_n27,
         ref_1_maj_180_n26, ref_1_maj_180_n25, ref_1_maj_180_n24,
         ref_1_maj_180_n23, ref_1_maj_180_n22, ref_1_maj_180_n21,
         ref_1_maj_180_n20, ref_1_maj_180_n19, ref_1_maj_180_n18,
         ref_1_maj_181_n34, ref_1_maj_181_n33, ref_1_maj_181_n32,
         ref_1_maj_181_n31, ref_1_maj_181_n30, ref_1_maj_181_n29,
         ref_1_maj_181_n28, ref_1_maj_181_n27, ref_1_maj_181_n26,
         ref_1_maj_181_n25, ref_1_maj_181_n24, ref_1_maj_181_n23,
         ref_1_maj_181_n22, ref_1_maj_181_n21, ref_1_maj_181_n20,
         ref_1_maj_181_n19, ref_1_maj_181_n18, ref_1_maj_182_n34,
         ref_1_maj_182_n33, ref_1_maj_182_n32, ref_1_maj_182_n31,
         ref_1_maj_182_n30, ref_1_maj_182_n29, ref_1_maj_182_n28,
         ref_1_maj_182_n27, ref_1_maj_182_n26, ref_1_maj_182_n25,
         ref_1_maj_182_n24, ref_1_maj_182_n23, ref_1_maj_182_n22,
         ref_1_maj_182_n21, ref_1_maj_182_n20, ref_1_maj_182_n19,
         ref_1_maj_182_n18, ref_1_maj_183_n34, ref_1_maj_183_n33,
         ref_1_maj_183_n32, ref_1_maj_183_n31, ref_1_maj_183_n30,
         ref_1_maj_183_n29, ref_1_maj_183_n28, ref_1_maj_183_n27,
         ref_1_maj_183_n26, ref_1_maj_183_n25, ref_1_maj_183_n24,
         ref_1_maj_183_n23, ref_1_maj_183_n22, ref_1_maj_183_n21,
         ref_1_maj_183_n20, ref_1_maj_183_n19, ref_1_maj_183_n18,
         ref_1_maj_184_n34, ref_1_maj_184_n33, ref_1_maj_184_n32,
         ref_1_maj_184_n31, ref_1_maj_184_n30, ref_1_maj_184_n29,
         ref_1_maj_184_n28, ref_1_maj_184_n27, ref_1_maj_184_n26,
         ref_1_maj_184_n25, ref_1_maj_184_n24, ref_1_maj_184_n23,
         ref_1_maj_184_n22, ref_1_maj_184_n21, ref_1_maj_184_n20,
         ref_1_maj_184_n19, ref_1_maj_184_n18, ref_1_maj_185_n34,
         ref_1_maj_185_n33, ref_1_maj_185_n32, ref_1_maj_185_n31,
         ref_1_maj_185_n30, ref_1_maj_185_n29, ref_1_maj_185_n28,
         ref_1_maj_185_n27, ref_1_maj_185_n26, ref_1_maj_185_n25,
         ref_1_maj_185_n24, ref_1_maj_185_n23, ref_1_maj_185_n22,
         ref_1_maj_185_n21, ref_1_maj_185_n20, ref_1_maj_185_n19,
         ref_1_maj_185_n18, ref_1_maj_186_n34, ref_1_maj_186_n33,
         ref_1_maj_186_n32, ref_1_maj_186_n31, ref_1_maj_186_n30,
         ref_1_maj_186_n29, ref_1_maj_186_n28, ref_1_maj_186_n27,
         ref_1_maj_186_n26, ref_1_maj_186_n25, ref_1_maj_186_n24,
         ref_1_maj_186_n23, ref_1_maj_186_n22, ref_1_maj_186_n21,
         ref_1_maj_186_n20, ref_1_maj_186_n19, ref_1_maj_186_n18,
         ref_1_maj_187_n34, ref_1_maj_187_n33, ref_1_maj_187_n32,
         ref_1_maj_187_n31, ref_1_maj_187_n30, ref_1_maj_187_n29,
         ref_1_maj_187_n28, ref_1_maj_187_n27, ref_1_maj_187_n26,
         ref_1_maj_187_n25, ref_1_maj_187_n24, ref_1_maj_187_n23,
         ref_1_maj_187_n22, ref_1_maj_187_n21, ref_1_maj_187_n20,
         ref_1_maj_187_n19, ref_1_maj_187_n18, ref_1_maj_188_n34,
         ref_1_maj_188_n33, ref_1_maj_188_n32, ref_1_maj_188_n31,
         ref_1_maj_188_n30, ref_1_maj_188_n29, ref_1_maj_188_n28,
         ref_1_maj_188_n27, ref_1_maj_188_n26, ref_1_maj_188_n25,
         ref_1_maj_188_n24, ref_1_maj_188_n23, ref_1_maj_188_n22,
         ref_1_maj_188_n21, ref_1_maj_188_n20, ref_1_maj_188_n19,
         ref_1_maj_188_n18, ref_1_maj_189_n34, ref_1_maj_189_n33,
         ref_1_maj_189_n32, ref_1_maj_189_n31, ref_1_maj_189_n30,
         ref_1_maj_189_n29, ref_1_maj_189_n28, ref_1_maj_189_n27,
         ref_1_maj_189_n26, ref_1_maj_189_n25, ref_1_maj_189_n24,
         ref_1_maj_189_n23, ref_1_maj_189_n22, ref_1_maj_189_n21,
         ref_1_maj_189_n20, ref_1_maj_189_n19, ref_1_maj_189_n18,
         ref_1_maj_190_n34, ref_1_maj_190_n33, ref_1_maj_190_n32,
         ref_1_maj_190_n31, ref_1_maj_190_n30, ref_1_maj_190_n29,
         ref_1_maj_190_n28, ref_1_maj_190_n27, ref_1_maj_190_n26,
         ref_1_maj_190_n25, ref_1_maj_190_n24, ref_1_maj_190_n23,
         ref_1_maj_190_n22, ref_1_maj_190_n21, ref_1_maj_190_n20,
         ref_1_maj_190_n19, ref_1_maj_190_n18, ref_1_maj_191_n34,
         ref_1_maj_191_n33, ref_1_maj_191_n32, ref_1_maj_191_n31,
         ref_1_maj_191_n30, ref_1_maj_191_n29, ref_1_maj_191_n28,
         ref_1_maj_191_n27, ref_1_maj_191_n26, ref_1_maj_191_n25,
         ref_1_maj_191_n24, ref_1_maj_191_n23, ref_1_maj_191_n22,
         ref_1_maj_191_n21, ref_1_maj_191_n20, ref_1_maj_191_n19,
         ref_1_maj_191_n18, ref_1_maj_192_n34, ref_1_maj_192_n33,
         ref_1_maj_192_n32, ref_1_maj_192_n31, ref_1_maj_192_n30,
         ref_1_maj_192_n29, ref_1_maj_192_n28, ref_1_maj_192_n27,
         ref_1_maj_192_n26, ref_1_maj_192_n25, ref_1_maj_192_n24,
         ref_1_maj_192_n23, ref_1_maj_192_n22, ref_1_maj_192_n21,
         ref_1_maj_192_n20, ref_1_maj_192_n19, ref_1_maj_192_n18,
         ref_1_maj_193_n34, ref_1_maj_193_n33, ref_1_maj_193_n32,
         ref_1_maj_193_n31, ref_1_maj_193_n30, ref_1_maj_193_n29,
         ref_1_maj_193_n28, ref_1_maj_193_n27, ref_1_maj_193_n26,
         ref_1_maj_193_n25, ref_1_maj_193_n24, ref_1_maj_193_n23,
         ref_1_maj_193_n22, ref_1_maj_193_n21, ref_1_maj_193_n20,
         ref_1_maj_193_n19, ref_1_maj_193_n18, ref_1_maj_194_n34,
         ref_1_maj_194_n33, ref_1_maj_194_n32, ref_1_maj_194_n31,
         ref_1_maj_194_n30, ref_1_maj_194_n29, ref_1_maj_194_n28,
         ref_1_maj_194_n27, ref_1_maj_194_n26, ref_1_maj_194_n25,
         ref_1_maj_194_n24, ref_1_maj_194_n23, ref_1_maj_194_n22,
         ref_1_maj_194_n21, ref_1_maj_194_n20, ref_1_maj_194_n19,
         ref_1_maj_194_n18, ref_1_maj_195_n34, ref_1_maj_195_n33,
         ref_1_maj_195_n32, ref_1_maj_195_n31, ref_1_maj_195_n30,
         ref_1_maj_195_n29, ref_1_maj_195_n28, ref_1_maj_195_n27,
         ref_1_maj_195_n26, ref_1_maj_195_n25, ref_1_maj_195_n24,
         ref_1_maj_195_n23, ref_1_maj_195_n22, ref_1_maj_195_n21,
         ref_1_maj_195_n20, ref_1_maj_195_n19, ref_1_maj_195_n18,
         ref_1_maj_196_n34, ref_1_maj_196_n33, ref_1_maj_196_n32,
         ref_1_maj_196_n31, ref_1_maj_196_n30, ref_1_maj_196_n29,
         ref_1_maj_196_n28, ref_1_maj_196_n27, ref_1_maj_196_n26,
         ref_1_maj_196_n25, ref_1_maj_196_n24, ref_1_maj_196_n23,
         ref_1_maj_196_n22, ref_1_maj_196_n21, ref_1_maj_196_n20,
         ref_1_maj_196_n19, ref_1_maj_196_n18, ref_1_maj_197_n34,
         ref_1_maj_197_n33, ref_1_maj_197_n32, ref_1_maj_197_n31,
         ref_1_maj_197_n30, ref_1_maj_197_n29, ref_1_maj_197_n28,
         ref_1_maj_197_n27, ref_1_maj_197_n26, ref_1_maj_197_n25,
         ref_1_maj_197_n24, ref_1_maj_197_n23, ref_1_maj_197_n22,
         ref_1_maj_197_n21, ref_1_maj_197_n20, ref_1_maj_197_n19,
         ref_1_maj_197_n18, ref_1_maj_198_n34, ref_1_maj_198_n33,
         ref_1_maj_198_n32, ref_1_maj_198_n31, ref_1_maj_198_n30,
         ref_1_maj_198_n29, ref_1_maj_198_n28, ref_1_maj_198_n27,
         ref_1_maj_198_n26, ref_1_maj_198_n25, ref_1_maj_198_n24,
         ref_1_maj_198_n23, ref_1_maj_198_n22, ref_1_maj_198_n21,
         ref_1_maj_198_n20, ref_1_maj_198_n19, ref_1_maj_198_n18,
         ref_1_maj_199_n34, ref_1_maj_199_n33, ref_1_maj_199_n32,
         ref_1_maj_199_n31, ref_1_maj_199_n30, ref_1_maj_199_n29,
         ref_1_maj_199_n28, ref_1_maj_199_n27, ref_1_maj_199_n26,
         ref_1_maj_199_n25, ref_1_maj_199_n24, ref_1_maj_199_n23,
         ref_1_maj_199_n22, ref_1_maj_199_n21, ref_1_maj_199_n20,
         ref_1_maj_199_n19, ref_1_maj_199_n18, ref_1_maj_200_n34,
         ref_1_maj_200_n33, ref_1_maj_200_n32, ref_1_maj_200_n31,
         ref_1_maj_200_n30, ref_1_maj_200_n29, ref_1_maj_200_n28,
         ref_1_maj_200_n27, ref_1_maj_200_n26, ref_1_maj_200_n25,
         ref_1_maj_200_n24, ref_1_maj_200_n23, ref_1_maj_200_n22,
         ref_1_maj_200_n21, ref_1_maj_200_n20, ref_1_maj_200_n19,
         ref_1_maj_200_n18, ref_1_maj_201_n34, ref_1_maj_201_n33,
         ref_1_maj_201_n32, ref_1_maj_201_n31, ref_1_maj_201_n30,
         ref_1_maj_201_n29, ref_1_maj_201_n28, ref_1_maj_201_n27,
         ref_1_maj_201_n26, ref_1_maj_201_n25, ref_1_maj_201_n24,
         ref_1_maj_201_n23, ref_1_maj_201_n22, ref_1_maj_201_n21,
         ref_1_maj_201_n20, ref_1_maj_201_n19, ref_1_maj_201_n18,
         ref_1_maj_202_n34, ref_1_maj_202_n33, ref_1_maj_202_n32,
         ref_1_maj_202_n31, ref_1_maj_202_n30, ref_1_maj_202_n29,
         ref_1_maj_202_n28, ref_1_maj_202_n27, ref_1_maj_202_n26,
         ref_1_maj_202_n25, ref_1_maj_202_n24, ref_1_maj_202_n23,
         ref_1_maj_202_n22, ref_1_maj_202_n21, ref_1_maj_202_n20,
         ref_1_maj_202_n19, ref_1_maj_202_n18, ref_1_maj_203_n34,
         ref_1_maj_203_n33, ref_1_maj_203_n32, ref_1_maj_203_n31,
         ref_1_maj_203_n30, ref_1_maj_203_n29, ref_1_maj_203_n28,
         ref_1_maj_203_n27, ref_1_maj_203_n26, ref_1_maj_203_n25,
         ref_1_maj_203_n24, ref_1_maj_203_n23, ref_1_maj_203_n22,
         ref_1_maj_203_n21, ref_1_maj_203_n20, ref_1_maj_203_n19,
         ref_1_maj_203_n18, ref_1_maj_204_n34, ref_1_maj_204_n33,
         ref_1_maj_204_n32, ref_1_maj_204_n31, ref_1_maj_204_n30,
         ref_1_maj_204_n29, ref_1_maj_204_n28, ref_1_maj_204_n27,
         ref_1_maj_204_n26, ref_1_maj_204_n25, ref_1_maj_204_n24,
         ref_1_maj_204_n23, ref_1_maj_204_n22, ref_1_maj_204_n21,
         ref_1_maj_204_n20, ref_1_maj_204_n19, ref_1_maj_204_n18,
         ref_1_maj_205_n34, ref_1_maj_205_n33, ref_1_maj_205_n32,
         ref_1_maj_205_n31, ref_1_maj_205_n30, ref_1_maj_205_n29,
         ref_1_maj_205_n28, ref_1_maj_205_n27, ref_1_maj_205_n26,
         ref_1_maj_205_n25, ref_1_maj_205_n24, ref_1_maj_205_n23,
         ref_1_maj_205_n22, ref_1_maj_205_n21, ref_1_maj_205_n20,
         ref_1_maj_205_n19, ref_1_maj_205_n18, ref_1_maj_206_n34,
         ref_1_maj_206_n33, ref_1_maj_206_n32, ref_1_maj_206_n31,
         ref_1_maj_206_n30, ref_1_maj_206_n29, ref_1_maj_206_n28,
         ref_1_maj_206_n27, ref_1_maj_206_n26, ref_1_maj_206_n25,
         ref_1_maj_206_n24, ref_1_maj_206_n23, ref_1_maj_206_n22,
         ref_1_maj_206_n21, ref_1_maj_206_n20, ref_1_maj_206_n19,
         ref_1_maj_206_n18, ref_1_maj_207_n34, ref_1_maj_207_n33,
         ref_1_maj_207_n32, ref_1_maj_207_n31, ref_1_maj_207_n30,
         ref_1_maj_207_n29, ref_1_maj_207_n28, ref_1_maj_207_n27,
         ref_1_maj_207_n26, ref_1_maj_207_n25, ref_1_maj_207_n24,
         ref_1_maj_207_n23, ref_1_maj_207_n22, ref_1_maj_207_n21,
         ref_1_maj_207_n20, ref_1_maj_207_n19, ref_1_maj_207_n18,
         ref_1_maj_208_n34, ref_1_maj_208_n33, ref_1_maj_208_n32,
         ref_1_maj_208_n31, ref_1_maj_208_n30, ref_1_maj_208_n29,
         ref_1_maj_208_n28, ref_1_maj_208_n27, ref_1_maj_208_n26,
         ref_1_maj_208_n25, ref_1_maj_208_n24, ref_1_maj_208_n23,
         ref_1_maj_208_n22, ref_1_maj_208_n21, ref_1_maj_208_n20,
         ref_1_maj_208_n19, ref_1_maj_208_n18, ref_1_maj_209_n34,
         ref_1_maj_209_n33, ref_1_maj_209_n32, ref_1_maj_209_n31,
         ref_1_maj_209_n30, ref_1_maj_209_n29, ref_1_maj_209_n28,
         ref_1_maj_209_n27, ref_1_maj_209_n26, ref_1_maj_209_n25,
         ref_1_maj_209_n24, ref_1_maj_209_n23, ref_1_maj_209_n22,
         ref_1_maj_209_n21, ref_1_maj_209_n20, ref_1_maj_209_n19,
         ref_1_maj_209_n18, ref_1_maj_210_n34, ref_1_maj_210_n33,
         ref_1_maj_210_n32, ref_1_maj_210_n31, ref_1_maj_210_n30,
         ref_1_maj_210_n29, ref_1_maj_210_n28, ref_1_maj_210_n27,
         ref_1_maj_210_n26, ref_1_maj_210_n25, ref_1_maj_210_n24,
         ref_1_maj_210_n23, ref_1_maj_210_n22, ref_1_maj_210_n21,
         ref_1_maj_210_n20, ref_1_maj_210_n19, ref_1_maj_210_n18,
         ref_1_maj_211_n34, ref_1_maj_211_n33, ref_1_maj_211_n32,
         ref_1_maj_211_n31, ref_1_maj_211_n30, ref_1_maj_211_n29,
         ref_1_maj_211_n28, ref_1_maj_211_n27, ref_1_maj_211_n26,
         ref_1_maj_211_n25, ref_1_maj_211_n24, ref_1_maj_211_n23,
         ref_1_maj_211_n22, ref_1_maj_211_n21, ref_1_maj_211_n20,
         ref_1_maj_211_n19, ref_1_maj_211_n18, ref_1_maj_212_n34,
         ref_1_maj_212_n33, ref_1_maj_212_n32, ref_1_maj_212_n31,
         ref_1_maj_212_n30, ref_1_maj_212_n29, ref_1_maj_212_n28,
         ref_1_maj_212_n27, ref_1_maj_212_n26, ref_1_maj_212_n25,
         ref_1_maj_212_n24, ref_1_maj_212_n23, ref_1_maj_212_n22,
         ref_1_maj_212_n21, ref_1_maj_212_n20, ref_1_maj_212_n19,
         ref_1_maj_212_n18, ref_1_maj_213_n34, ref_1_maj_213_n33,
         ref_1_maj_213_n32, ref_1_maj_213_n31, ref_1_maj_213_n30,
         ref_1_maj_213_n29, ref_1_maj_213_n28, ref_1_maj_213_n27,
         ref_1_maj_213_n26, ref_1_maj_213_n25, ref_1_maj_213_n24,
         ref_1_maj_213_n23, ref_1_maj_213_n22, ref_1_maj_213_n21,
         ref_1_maj_213_n20, ref_1_maj_213_n19, ref_1_maj_213_n18,
         ref_1_maj_214_n34, ref_1_maj_214_n33, ref_1_maj_214_n32,
         ref_1_maj_214_n31, ref_1_maj_214_n30, ref_1_maj_214_n29,
         ref_1_maj_214_n28, ref_1_maj_214_n27, ref_1_maj_214_n26,
         ref_1_maj_214_n25, ref_1_maj_214_n24, ref_1_maj_214_n23,
         ref_1_maj_214_n22, ref_1_maj_214_n21, ref_1_maj_214_n20,
         ref_1_maj_214_n19, ref_1_maj_214_n18, ref_1_maj_215_n34,
         ref_1_maj_215_n33, ref_1_maj_215_n32, ref_1_maj_215_n31,
         ref_1_maj_215_n30, ref_1_maj_215_n29, ref_1_maj_215_n28,
         ref_1_maj_215_n27, ref_1_maj_215_n26, ref_1_maj_215_n25,
         ref_1_maj_215_n24, ref_1_maj_215_n23, ref_1_maj_215_n22,
         ref_1_maj_215_n21, ref_1_maj_215_n20, ref_1_maj_215_n19,
         ref_1_maj_215_n18, ref_1_maj_216_n34, ref_1_maj_216_n33,
         ref_1_maj_216_n32, ref_1_maj_216_n31, ref_1_maj_216_n30,
         ref_1_maj_216_n29, ref_1_maj_216_n28, ref_1_maj_216_n27,
         ref_1_maj_216_n26, ref_1_maj_216_n25, ref_1_maj_216_n24,
         ref_1_maj_216_n23, ref_1_maj_216_n22, ref_1_maj_216_n21,
         ref_1_maj_216_n20, ref_1_maj_216_n19, ref_1_maj_216_n18,
         ref_1_maj_217_n34, ref_1_maj_217_n33, ref_1_maj_217_n32,
         ref_1_maj_217_n31, ref_1_maj_217_n30, ref_1_maj_217_n29,
         ref_1_maj_217_n28, ref_1_maj_217_n27, ref_1_maj_217_n26,
         ref_1_maj_217_n25, ref_1_maj_217_n24, ref_1_maj_217_n23,
         ref_1_maj_217_n22, ref_1_maj_217_n21, ref_1_maj_217_n20,
         ref_1_maj_217_n19, ref_1_maj_217_n18, ref_1_maj_218_n34,
         ref_1_maj_218_n33, ref_1_maj_218_n32, ref_1_maj_218_n31,
         ref_1_maj_218_n30, ref_1_maj_218_n29, ref_1_maj_218_n28,
         ref_1_maj_218_n27, ref_1_maj_218_n26, ref_1_maj_218_n25,
         ref_1_maj_218_n24, ref_1_maj_218_n23, ref_1_maj_218_n22,
         ref_1_maj_218_n21, ref_1_maj_218_n20, ref_1_maj_218_n19,
         ref_1_maj_218_n18, ref_1_maj_219_n34, ref_1_maj_219_n33,
         ref_1_maj_219_n32, ref_1_maj_219_n31, ref_1_maj_219_n30,
         ref_1_maj_219_n29, ref_1_maj_219_n28, ref_1_maj_219_n27,
         ref_1_maj_219_n26, ref_1_maj_219_n25, ref_1_maj_219_n24,
         ref_1_maj_219_n23, ref_1_maj_219_n22, ref_1_maj_219_n21,
         ref_1_maj_219_n20, ref_1_maj_219_n19, ref_1_maj_219_n18,
         ref_1_maj_220_n34, ref_1_maj_220_n33, ref_1_maj_220_n32,
         ref_1_maj_220_n31, ref_1_maj_220_n30, ref_1_maj_220_n29,
         ref_1_maj_220_n28, ref_1_maj_220_n27, ref_1_maj_220_n26,
         ref_1_maj_220_n25, ref_1_maj_220_n24, ref_1_maj_220_n23,
         ref_1_maj_220_n22, ref_1_maj_220_n21, ref_1_maj_220_n20,
         ref_1_maj_220_n19, ref_1_maj_220_n18, ref_1_maj_221_n34,
         ref_1_maj_221_n33, ref_1_maj_221_n32, ref_1_maj_221_n31,
         ref_1_maj_221_n30, ref_1_maj_221_n29, ref_1_maj_221_n28,
         ref_1_maj_221_n27, ref_1_maj_221_n26, ref_1_maj_221_n25,
         ref_1_maj_221_n24, ref_1_maj_221_n23, ref_1_maj_221_n22,
         ref_1_maj_221_n21, ref_1_maj_221_n20, ref_1_maj_221_n19,
         ref_1_maj_221_n18, ref_1_maj_222_n34, ref_1_maj_222_n33,
         ref_1_maj_222_n32, ref_1_maj_222_n31, ref_1_maj_222_n30,
         ref_1_maj_222_n29, ref_1_maj_222_n28, ref_1_maj_222_n27,
         ref_1_maj_222_n26, ref_1_maj_222_n25, ref_1_maj_222_n24,
         ref_1_maj_222_n23, ref_1_maj_222_n22, ref_1_maj_222_n21,
         ref_1_maj_222_n20, ref_1_maj_222_n19, ref_1_maj_222_n18,
         ref_1_maj_223_n34, ref_1_maj_223_n33, ref_1_maj_223_n32,
         ref_1_maj_223_n31, ref_1_maj_223_n30, ref_1_maj_223_n29,
         ref_1_maj_223_n28, ref_1_maj_223_n27, ref_1_maj_223_n26,
         ref_1_maj_223_n25, ref_1_maj_223_n24, ref_1_maj_223_n23,
         ref_1_maj_223_n22, ref_1_maj_223_n21, ref_1_maj_223_n20,
         ref_1_maj_223_n19, ref_1_maj_223_n18;
  wire   [6:0] ref_1_port_o_0_0;
  wire   [6:0] ref_1_port_o_0_1;
  wire   [6:0] ref_1_port_o_0_2;
  wire   [6:0] ref_1_port_o_0_3;
  wire   [6:0] ref_1_port_o_1_0;
  wire   [6:0] ref_1_port_o_1_1;
  wire   [6:0] ref_1_port_o_1_2;
  wire   [6:0] ref_1_port_o_1_3;
  wire   [6:0] ref_1_port_o_2_0;
  wire   [6:0] ref_1_port_o_2_1;
  wire   [6:0] ref_1_port_o_2_2;
  wire   [6:0] ref_1_port_o_2_3;
  wire   [6:0] ref_1_port_o_3_0;
  wire   [6:0] ref_1_port_o_3_1;
  wire   [6:0] ref_1_port_o_3_2;
  wire   [6:0] ref_1_port_o_3_3;
  wire   [6:0] temp_0_0;
  wire   [6:0] mult_ab_0_1;
  wire   [6:0] mult_ab_0_2;
  wire   [6:0] mult_ab_0_3;
  wire   [6:0] temp_0_1;
  wire   [6:0] mult_ab_1_0;
  wire   [6:0] mult_ab_1_2;
  wire   [6:0] mult_ab_1_3;
  wire   [6:0] temp_0_2;
  wire   [6:0] mult_ab_2_0;
  wire   [6:0] mult_ab_2_1;
  wire   [6:0] mult_ab_2_3;
  wire   [6:0] temp_0_3;
  wire   [6:0] mult_ab_3_0;
  wire   [6:0] mult_ab_3_1;
  wire   [6:0] mult_ab_3_2;

  DFF_X1 mult_ab_0_0_reg_6_ ( .D(N96), .CK(clk), .Q(temp_0_0[6]), .QN() );
  DFF_X1 mult_ab_0_0_reg_5_ ( .D(N80), .CK(clk), .Q(temp_0_0[5]), .QN() );
  DFF_X1 mult_ab_0_0_reg_4_ ( .D(N64), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 mult_ab_0_0_reg_3_ ( .D(N48), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 mult_ab_0_0_reg_2_ ( .D(N32), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 mult_ab_0_0_reg_1_ ( .D(N16), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 mult_ab_0_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 mult_ab_3_3_reg_6_ ( .D(N111), .CK(clk), .Q(temp_0_3[6]), .QN() );
  DFF_X1 mult_ab_3_3_reg_5_ ( .D(N95), .CK(clk), .Q(temp_0_3[5]), .QN() );
  DFF_X1 mult_ab_3_3_reg_4_ ( .D(N79), .CK(clk), .Q(temp_0_3[4]), .QN() );
  DFF_X1 mult_ab_3_3_reg_3_ ( .D(N63), .CK(clk), .Q(temp_0_3[3]), .QN() );
  DFF_X1 mult_ab_3_3_reg_2_ ( .D(N47), .CK(clk), .Q(temp_0_3[2]), .QN() );
  DFF_X1 mult_ab_3_3_reg_1_ ( .D(N31), .CK(clk), .Q(temp_0_3[1]), .QN() );
  DFF_X1 mult_ab_3_3_reg_0_ ( .D(N15), .CK(clk), .Q(temp_0_3[0]), .QN() );
  DFF_X1 mult_ab_0_1_reg_6_ ( .D(N97), .CK(clk), .Q(mult_ab_0_1[6]), .QN() );
  DFF_X1 mult_ab_0_1_reg_5_ ( .D(N81), .CK(clk), .Q(mult_ab_0_1[5]), .QN() );
  DFF_X1 mult_ab_0_1_reg_4_ ( .D(N65), .CK(clk), .Q(mult_ab_0_1[4]), .QN() );
  DFF_X1 mult_ab_0_1_reg_3_ ( .D(N49), .CK(clk), .Q(mult_ab_0_1[3]), .QN() );
  DFF_X1 mult_ab_0_1_reg_2_ ( .D(N33), .CK(clk), .Q(mult_ab_0_1[2]), .QN() );
  DFF_X1 mult_ab_0_1_reg_1_ ( .D(N17), .CK(clk), .Q(mult_ab_0_1[1]), .QN() );
  DFF_X1 mult_ab_0_1_reg_0_ ( .D(N1), .CK(clk), .Q(mult_ab_0_1[0]), .QN() );
  DFF_X1 mult_ab_0_2_reg_6_ ( .D(N98), .CK(clk), .Q(mult_ab_0_2[6]), .QN() );
  DFF_X1 mult_ab_0_2_reg_5_ ( .D(N82), .CK(clk), .Q(mult_ab_0_2[5]), .QN() );
  DFF_X1 mult_ab_0_2_reg_4_ ( .D(N66), .CK(clk), .Q(mult_ab_0_2[4]), .QN() );
  DFF_X1 mult_ab_0_2_reg_3_ ( .D(N50), .CK(clk), .Q(mult_ab_0_2[3]), .QN() );
  DFF_X1 mult_ab_0_2_reg_2_ ( .D(N34), .CK(clk), .Q(mult_ab_0_2[2]), .QN() );
  DFF_X1 mult_ab_0_2_reg_1_ ( .D(N18), .CK(clk), .Q(mult_ab_0_2[1]), .QN() );
  DFF_X1 mult_ab_0_2_reg_0_ ( .D(N2), .CK(clk), .Q(mult_ab_0_2[0]), .QN() );
  DFF_X1 mult_ab_2_3_reg_6_ ( .D(N107), .CK(clk), .Q(mult_ab_2_3[6]), .QN() );
  DFF_X1 mult_ab_2_3_reg_5_ ( .D(N91), .CK(clk), .Q(mult_ab_2_3[5]), .QN() );
  DFF_X1 mult_ab_2_3_reg_4_ ( .D(N75), .CK(clk), .Q(mult_ab_2_3[4]), .QN() );
  DFF_X1 mult_ab_2_3_reg_3_ ( .D(N59), .CK(clk), .Q(mult_ab_2_3[3]), .QN() );
  DFF_X1 mult_ab_2_3_reg_2_ ( .D(N43), .CK(clk), .Q(mult_ab_2_3[2]), .QN() );
  DFF_X1 mult_ab_2_3_reg_1_ ( .D(N27), .CK(clk), .Q(mult_ab_2_3[1]), .QN() );
  DFF_X1 mult_ab_2_3_reg_0_ ( .D(N11), .CK(clk), .Q(mult_ab_2_3[0]), .QN() );
  DFF_X1 mult_ab_1_3_reg_6_ ( .D(N103), .CK(clk), .Q(mult_ab_1_3[6]), .QN() );
  DFF_X1 mult_ab_1_3_reg_5_ ( .D(N87), .CK(clk), .Q(mult_ab_1_3[5]), .QN() );
  DFF_X1 mult_ab_1_3_reg_4_ ( .D(N71), .CK(clk), .Q(mult_ab_1_3[4]), .QN() );
  DFF_X1 mult_ab_1_3_reg_3_ ( .D(N55), .CK(clk), .Q(mult_ab_1_3[3]), .QN() );
  DFF_X1 mult_ab_1_3_reg_2_ ( .D(N39), .CK(clk), .Q(mult_ab_1_3[2]), .QN() );
  DFF_X1 mult_ab_1_3_reg_1_ ( .D(N23), .CK(clk), .Q(mult_ab_1_3[1]), .QN() );
  DFF_X1 mult_ab_1_3_reg_0_ ( .D(N7), .CK(clk), .Q(mult_ab_1_3[0]), .QN() );
  DFF_X1 mult_ab_0_3_reg_6_ ( .D(N99), .CK(clk), .Q(mult_ab_0_3[6]), .QN() );
  DFF_X1 mult_ab_0_3_reg_5_ ( .D(N83), .CK(clk), .Q(mult_ab_0_3[5]), .QN() );
  DFF_X1 mult_ab_0_3_reg_4_ ( .D(N67), .CK(clk), .Q(mult_ab_0_3[4]), .QN() );
  DFF_X1 mult_ab_0_3_reg_3_ ( .D(N51), .CK(clk), .Q(mult_ab_0_3[3]), .QN() );
  DFF_X1 mult_ab_0_3_reg_2_ ( .D(N35), .CK(clk), .Q(mult_ab_0_3[2]), .QN() );
  DFF_X1 mult_ab_0_3_reg_1_ ( .D(N19), .CK(clk), .Q(mult_ab_0_3[1]), .QN() );
  DFF_X1 mult_ab_0_3_reg_0_ ( .D(N3), .CK(clk), .Q(mult_ab_0_3[0]), .QN() );
  DFF_X1 mult_ab_3_1_reg_6_ ( .D(N109), .CK(clk), .Q(mult_ab_3_1[6]), .QN() );
  DFF_X1 mult_ab_3_1_reg_5_ ( .D(N93), .CK(clk), .Q(mult_ab_3_1[5]), .QN() );
  DFF_X1 mult_ab_3_1_reg_4_ ( .D(N77), .CK(clk), .Q(mult_ab_3_1[4]), .QN() );
  DFF_X1 mult_ab_3_1_reg_3_ ( .D(N61), .CK(clk), .Q(mult_ab_3_1[3]), .QN() );
  DFF_X1 mult_ab_3_1_reg_2_ ( .D(N45), .CK(clk), .Q(mult_ab_3_1[2]), .QN() );
  DFF_X1 mult_ab_3_1_reg_1_ ( .D(N29), .CK(clk), .Q(mult_ab_3_1[1]), .QN() );
  DFF_X1 mult_ab_3_1_reg_0_ ( .D(N13), .CK(clk), .Q(mult_ab_3_1[0]), .QN() );
  DFF_X1 mult_ab_1_1_reg_6_ ( .D(N101), .CK(clk), .Q(temp_0_1[6]), .QN() );
  DFF_X1 mult_ab_1_1_reg_5_ ( .D(N85), .CK(clk), .Q(temp_0_1[5]), .QN() );
  DFF_X1 mult_ab_1_1_reg_4_ ( .D(N69), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 mult_ab_1_1_reg_3_ ( .D(N53), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 mult_ab_1_1_reg_2_ ( .D(N37), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 mult_ab_1_1_reg_1_ ( .D(N21), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 mult_ab_1_1_reg_0_ ( .D(N5), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 mult_ab_3_0_reg_6_ ( .D(N108), .CK(clk), .Q(mult_ab_3_0[6]), .QN() );
  DFF_X1 mult_ab_3_0_reg_5_ ( .D(N92), .CK(clk), .Q(mult_ab_3_0[5]), .QN() );
  DFF_X1 mult_ab_3_0_reg_4_ ( .D(N76), .CK(clk), .Q(mult_ab_3_0[4]), .QN() );
  DFF_X1 mult_ab_3_0_reg_3_ ( .D(N60), .CK(clk), .Q(mult_ab_3_0[3]), .QN() );
  DFF_X1 mult_ab_3_0_reg_2_ ( .D(N44), .CK(clk), .Q(mult_ab_3_0[2]), .QN() );
  DFF_X1 mult_ab_3_0_reg_1_ ( .D(N28), .CK(clk), .Q(mult_ab_3_0[1]), .QN() );
  DFF_X1 mult_ab_3_0_reg_0_ ( .D(N12), .CK(clk), .Q(mult_ab_3_0[0]), .QN() );
  DFF_X1 mult_ab_2_2_reg_6_ ( .D(N106), .CK(clk), .Q(temp_0_2[6]), .QN() );
  DFF_X1 mult_ab_2_2_reg_5_ ( .D(N90), .CK(clk), .Q(temp_0_2[5]), .QN() );
  DFF_X1 mult_ab_2_2_reg_4_ ( .D(N74), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 mult_ab_2_2_reg_3_ ( .D(N58), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 mult_ab_2_2_reg_2_ ( .D(N42), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 mult_ab_2_2_reg_1_ ( .D(N26), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 mult_ab_2_2_reg_0_ ( .D(N10), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 mult_ab_3_2_reg_6_ ( .D(N110), .CK(clk), .Q(mult_ab_3_2[6]), .QN() );
  DFF_X1 mult_ab_3_2_reg_5_ ( .D(N94), .CK(clk), .Q(mult_ab_3_2[5]), .QN() );
  DFF_X1 mult_ab_3_2_reg_4_ ( .D(N78), .CK(clk), .Q(mult_ab_3_2[4]), .QN() );
  DFF_X1 mult_ab_3_2_reg_3_ ( .D(N62), .CK(clk), .Q(mult_ab_3_2[3]), .QN() );
  DFF_X1 mult_ab_3_2_reg_2_ ( .D(N46), .CK(clk), .Q(mult_ab_3_2[2]), .QN() );
  DFF_X1 mult_ab_3_2_reg_1_ ( .D(N30), .CK(clk), .Q(mult_ab_3_2[1]), .QN() );
  DFF_X1 mult_ab_3_2_reg_0_ ( .D(N14), .CK(clk), .Q(mult_ab_3_2[0]), .QN() );
  DFF_X1 mult_ab_1_2_reg_6_ ( .D(N102), .CK(clk), .Q(mult_ab_1_2[6]), .QN() );
  DFF_X1 mult_ab_1_2_reg_5_ ( .D(N86), .CK(clk), .Q(mult_ab_1_2[5]), .QN() );
  DFF_X1 mult_ab_1_2_reg_4_ ( .D(N70), .CK(clk), .Q(mult_ab_1_2[4]), .QN() );
  DFF_X1 mult_ab_1_2_reg_3_ ( .D(N54), .CK(clk), .Q(mult_ab_1_2[3]), .QN() );
  DFF_X1 mult_ab_1_2_reg_2_ ( .D(N38), .CK(clk), .Q(mult_ab_1_2[2]), .QN() );
  DFF_X1 mult_ab_1_2_reg_1_ ( .D(N22), .CK(clk), .Q(mult_ab_1_2[1]), .QN() );
  DFF_X1 mult_ab_1_2_reg_0_ ( .D(N6), .CK(clk), .Q(mult_ab_1_2[0]), .QN() );
  DFF_X1 mult_ab_2_0_reg_6_ ( .D(N104), .CK(clk), .Q(mult_ab_2_0[6]), .QN() );
  DFF_X1 mult_ab_2_0_reg_5_ ( .D(N88), .CK(clk), .Q(mult_ab_2_0[5]), .QN() );
  DFF_X1 mult_ab_2_0_reg_4_ ( .D(N72), .CK(clk), .Q(mult_ab_2_0[4]), .QN() );
  DFF_X1 mult_ab_2_0_reg_3_ ( .D(N56), .CK(clk), .Q(mult_ab_2_0[3]), .QN() );
  DFF_X1 mult_ab_2_0_reg_2_ ( .D(N40), .CK(clk), .Q(mult_ab_2_0[2]), .QN() );
  DFF_X1 mult_ab_2_0_reg_1_ ( .D(N24), .CK(clk), .Q(mult_ab_2_0[1]), .QN() );
  DFF_X1 mult_ab_2_0_reg_0_ ( .D(N8), .CK(clk), .Q(mult_ab_2_0[0]), .QN() );
  DFF_X1 mult_ab_2_1_reg_6_ ( .D(N105), .CK(clk), .Q(mult_ab_2_1[6]), .QN() );
  DFF_X1 mult_ab_2_1_reg_5_ ( .D(N89), .CK(clk), .Q(mult_ab_2_1[5]), .QN() );
  DFF_X1 mult_ab_2_1_reg_4_ ( .D(N73), .CK(clk), .Q(mult_ab_2_1[4]), .QN() );
  DFF_X1 mult_ab_2_1_reg_3_ ( .D(N57), .CK(clk), .Q(mult_ab_2_1[3]), .QN() );
  DFF_X1 mult_ab_2_1_reg_2_ ( .D(N41), .CK(clk), .Q(mult_ab_2_1[2]), .QN() );
  DFF_X1 mult_ab_2_1_reg_1_ ( .D(N25), .CK(clk), .Q(mult_ab_2_1[1]), .QN() );
  DFF_X1 mult_ab_2_1_reg_0_ ( .D(N9), .CK(clk), .Q(mult_ab_2_1[0]), .QN() );
  DFF_X1 mult_ab_1_0_reg_6_ ( .D(N100), .CK(clk), .Q(mult_ab_1_0[6]), .QN() );
  DFF_X1 mult_ab_1_0_reg_5_ ( .D(N84), .CK(clk), .Q(mult_ab_1_0[5]), .QN() );
  DFF_X1 mult_ab_1_0_reg_4_ ( .D(N68), .CK(clk), .Q(mult_ab_1_0[4]), .QN() );
  DFF_X1 mult_ab_1_0_reg_3_ ( .D(N52), .CK(clk), .Q(mult_ab_1_0[3]), .QN() );
  DFF_X1 mult_ab_1_0_reg_2_ ( .D(N36), .CK(clk), .Q(mult_ab_1_0[2]), .QN() );
  DFF_X1 mult_ab_1_0_reg_1_ ( .D(N20), .CK(clk), .Q(mult_ab_1_0[1]), .QN() );
  DFF_X1 mult_ab_1_0_reg_0_ ( .D(N4), .CK(clk), .Q(mult_ab_1_0[0]), .QN() );
  XNOR2_X1 U283 ( .A(port_rand_mul[0]), .B(n106), .ZN(N4) );
  NAND2_X1 U284 ( .A1(ref_1_port_o_1_0[0]), .A2(port_a_1[0]), .ZN(n106) );
  XNOR2_X1 U285 ( .A(port_rand_mul[0]), .B(n122), .ZN(N20) );
  NAND2_X1 U286 ( .A1(ref_1_port_o_1_0[1]), .A2(port_a_1[1]), .ZN(n122) );
  XNOR2_X1 U287 ( .A(port_rand_mul[0]), .B(n109), .ZN(N36) );
  NAND2_X1 U288 ( .A1(ref_1_port_o_1_0[2]), .A2(port_a_1[2]), .ZN(n109) );
  XNOR2_X1 U289 ( .A(port_rand_mul[0]), .B(n96), .ZN(N52) );
  NAND2_X1 U290 ( .A1(ref_1_port_o_1_0[3]), .A2(port_a_1[3]), .ZN(n96) );
  XNOR2_X1 U291 ( .A(port_rand_mul[0]), .B(n83), .ZN(N68) );
  NAND2_X1 U292 ( .A1(ref_1_port_o_1_0[4]), .A2(port_a_1[4]), .ZN(n83) );
  XNOR2_X1 U293 ( .A(port_rand_mul[0]), .B(n69), .ZN(N84) );
  NAND2_X1 U294 ( .A1(ref_1_port_o_1_0[5]), .A2(port_a_1[5]), .ZN(n69) );
  XNOR2_X1 U295 ( .A(port_rand_mul[0]), .B(n139), .ZN(N100) );
  NAND2_X1 U296 ( .A1(ref_1_port_o_1_0[6]), .A2(port_a_1[6]), .ZN(n139) );
  XNOR2_X1 U297 ( .A(port_rand_mul[3]), .B(n64), .ZN(N9) );
  NAND2_X1 U298 ( .A1(ref_1_port_o_2_1[0]), .A2(port_a_2[0]), .ZN(n64) );
  XNOR2_X1 U299 ( .A(port_rand_mul[3]), .B(n118), .ZN(N25) );
  NAND2_X1 U300 ( .A1(ref_1_port_o_2_1[1]), .A2(port_a_2[1]), .ZN(n118) );
  XNOR2_X1 U301 ( .A(port_rand_mul[3]), .B(n104), .ZN(N41) );
  NAND2_X1 U302 ( .A1(ref_1_port_o_2_1[2]), .A2(port_a_2[2]), .ZN(n104) );
  XNOR2_X1 U303 ( .A(port_rand_mul[3]), .B(n92), .ZN(N57) );
  NAND2_X1 U304 ( .A1(ref_1_port_o_2_1[3]), .A2(port_a_2[3]), .ZN(n92) );
  XNOR2_X1 U305 ( .A(port_rand_mul[3]), .B(n78), .ZN(N73) );
  NAND2_X1 U306 ( .A1(ref_1_port_o_2_1[4]), .A2(port_a_2[4]), .ZN(n78) );
  XNOR2_X1 U307 ( .A(port_rand_mul[3]), .B(n65), .ZN(N89) );
  NAND2_X1 U308 ( .A1(ref_1_port_o_2_1[5]), .A2(port_a_2[5]), .ZN(n65) );
  XNOR2_X1 U309 ( .A(port_rand_mul[3]), .B(n135), .ZN(N105) );
  NAND2_X1 U310 ( .A1(ref_1_port_o_2_1[6]), .A2(port_a_2[6]), .ZN(n135) );
  XNOR2_X1 U311 ( .A(port_rand_mul[1]), .B(n73), .ZN(N8) );
  NAND2_X1 U312 ( .A1(ref_1_port_o_2_0[0]), .A2(port_a_2[0]), .ZN(n73) );
  XNOR2_X1 U313 ( .A(port_rand_mul[1]), .B(n119), .ZN(N24) );
  NAND2_X1 U314 ( .A1(ref_1_port_o_2_0[1]), .A2(port_a_2[1]), .ZN(n119) );
  XNOR2_X1 U315 ( .A(port_rand_mul[1]), .B(n105), .ZN(N40) );
  NAND2_X1 U316 ( .A1(ref_1_port_o_2_0[2]), .A2(port_a_2[2]), .ZN(n105) );
  XNOR2_X1 U317 ( .A(port_rand_mul[1]), .B(n93), .ZN(N56) );
  NAND2_X1 U318 ( .A1(ref_1_port_o_2_0[3]), .A2(port_a_2[3]), .ZN(n93) );
  XNOR2_X1 U319 ( .A(port_rand_mul[1]), .B(n79), .ZN(N72) );
  NAND2_X1 U320 ( .A1(ref_1_port_o_2_0[4]), .A2(port_a_2[4]), .ZN(n79) );
  XNOR2_X1 U321 ( .A(port_rand_mul[1]), .B(n66), .ZN(N88) );
  NAND2_X1 U322 ( .A1(ref_1_port_o_2_0[5]), .A2(port_a_2[5]), .ZN(n66) );
  XNOR2_X1 U323 ( .A(port_rand_mul[1]), .B(n136), .ZN(N104) );
  NAND2_X1 U324 ( .A1(ref_1_port_o_2_0[6]), .A2(port_a_2[6]), .ZN(n136) );
  XNOR2_X1 U325 ( .A(port_rand_mul[3]), .B(n90), .ZN(N6) );
  NAND2_X1 U326 ( .A1(ref_1_port_o_1_2[0]), .A2(port_a_1[0]), .ZN(n90) );
  XNOR2_X1 U327 ( .A(port_rand_mul[3]), .B(n121), .ZN(N22) );
  NAND2_X1 U328 ( .A1(ref_1_port_o_1_2[1]), .A2(port_a_1[1]), .ZN(n121) );
  XNOR2_X1 U329 ( .A(port_rand_mul[3]), .B(n108), .ZN(N38) );
  NAND2_X1 U330 ( .A1(ref_1_port_o_1_2[2]), .A2(port_a_1[2]), .ZN(n108) );
  XNOR2_X1 U331 ( .A(port_rand_mul[3]), .B(n95), .ZN(N54) );
  NAND2_X1 U332 ( .A1(ref_1_port_o_1_2[3]), .A2(port_a_1[3]), .ZN(n95) );
  XNOR2_X1 U333 ( .A(port_rand_mul[3]), .B(n81), .ZN(N70) );
  NAND2_X1 U334 ( .A1(ref_1_port_o_1_2[4]), .A2(port_a_1[4]), .ZN(n81) );
  XNOR2_X1 U335 ( .A(port_rand_mul[3]), .B(n68), .ZN(N86) );
  NAND2_X1 U336 ( .A1(ref_1_port_o_1_2[5]), .A2(port_a_1[5]), .ZN(n68) );
  XNOR2_X1 U337 ( .A(port_rand_mul[3]), .B(n138), .ZN(N102) );
  NAND2_X1 U338 ( .A1(ref_1_port_o_1_2[6]), .A2(port_a_1[6]), .ZN(n138) );
  XNOR2_X1 U339 ( .A(port_rand_mul[5]), .B(n127), .ZN(N14) );
  NAND2_X1 U340 ( .A1(ref_1_port_o_3_2[0]), .A2(port_a_3[0]), .ZN(n127) );
  XNOR2_X1 U341 ( .A(port_rand_mul[5]), .B(n113), .ZN(N30) );
  NAND2_X1 U342 ( .A1(ref_1_port_o_3_2[1]), .A2(port_a_3[1]), .ZN(n113) );
  XNOR2_X1 U343 ( .A(port_rand_mul[5]), .B(n100), .ZN(N46) );
  NAND2_X1 U344 ( .A1(ref_1_port_o_3_2[2]), .A2(port_a_3[2]), .ZN(n100) );
  XNOR2_X1 U345 ( .A(port_rand_mul[5]), .B(n87), .ZN(N62) );
  NAND2_X1 U346 ( .A1(ref_1_port_o_3_2[3]), .A2(port_a_3[3]), .ZN(n87) );
  XNOR2_X1 U347 ( .A(port_rand_mul[5]), .B(n74), .ZN(N78) );
  NAND2_X1 U348 ( .A1(ref_1_port_o_3_2[4]), .A2(port_a_3[4]), .ZN(n74) );
  XNOR2_X1 U349 ( .A(port_rand_mul[5]), .B(n60), .ZN(N94) );
  NAND2_X1 U350 ( .A1(ref_1_port_o_3_2[5]), .A2(port_a_3[5]), .ZN(n60) );
  XNOR2_X1 U351 ( .A(port_rand_mul[5]), .B(n130), .ZN(N110) );
  NAND2_X1 U352 ( .A1(ref_1_port_o_3_2[6]), .A2(port_a_3[6]), .ZN(n130) );
  XNOR2_X1 U353 ( .A(port_rand_mul[2]), .B(n129), .ZN(N12) );
  NAND2_X1 U354 ( .A1(ref_1_port_o_3_0[0]), .A2(port_a_3[0]), .ZN(n129) );
  XNOR2_X1 U355 ( .A(port_rand_mul[2]), .B(n116), .ZN(N28) );
  NAND2_X1 U356 ( .A1(ref_1_port_o_3_0[1]), .A2(port_a_3[1]), .ZN(n116) );
  XNOR2_X1 U357 ( .A(port_rand_mul[2]), .B(n102), .ZN(N44) );
  NAND2_X1 U358 ( .A1(ref_1_port_o_3_0[2]), .A2(port_a_3[2]), .ZN(n102) );
  XNOR2_X1 U359 ( .A(port_rand_mul[2]), .B(n89), .ZN(N60) );
  NAND2_X1 U360 ( .A1(ref_1_port_o_3_0[3]), .A2(port_a_3[3]), .ZN(n89) );
  XNOR2_X1 U361 ( .A(port_rand_mul[2]), .B(n76), .ZN(N76) );
  NAND2_X1 U362 ( .A1(ref_1_port_o_3_0[4]), .A2(port_a_3[4]), .ZN(n76) );
  XNOR2_X1 U363 ( .A(port_rand_mul[2]), .B(n62), .ZN(N92) );
  NAND2_X1 U364 ( .A1(ref_1_port_o_3_0[5]), .A2(port_a_3[5]), .ZN(n62) );
  XNOR2_X1 U365 ( .A(port_rand_mul[2]), .B(n133), .ZN(N108) );
  NAND2_X1 U366 ( .A1(ref_1_port_o_3_0[6]), .A2(port_a_3[6]), .ZN(n133) );
  XNOR2_X1 U367 ( .A(port_rand_mul[4]), .B(n128), .ZN(N13) );
  NAND2_X1 U368 ( .A1(ref_1_port_o_3_1[0]), .A2(port_a_3[0]), .ZN(n128) );
  XNOR2_X1 U369 ( .A(port_rand_mul[4]), .B(n115), .ZN(N29) );
  NAND2_X1 U370 ( .A1(ref_1_port_o_3_1[1]), .A2(port_a_3[1]), .ZN(n115) );
  XNOR2_X1 U371 ( .A(port_rand_mul[4]), .B(n101), .ZN(N45) );
  NAND2_X1 U372 ( .A1(ref_1_port_o_3_1[2]), .A2(port_a_3[2]), .ZN(n101) );
  XNOR2_X1 U373 ( .A(port_rand_mul[4]), .B(n88), .ZN(N61) );
  NAND2_X1 U374 ( .A1(ref_1_port_o_3_1[3]), .A2(port_a_3[3]), .ZN(n88) );
  XNOR2_X1 U375 ( .A(port_rand_mul[4]), .B(n75), .ZN(N77) );
  NAND2_X1 U376 ( .A1(ref_1_port_o_3_1[4]), .A2(port_a_3[4]), .ZN(n75) );
  XNOR2_X1 U377 ( .A(port_rand_mul[4]), .B(n61), .ZN(N93) );
  NAND2_X1 U378 ( .A1(ref_1_port_o_3_1[5]), .A2(port_a_3[5]), .ZN(n61) );
  XNOR2_X1 U379 ( .A(port_rand_mul[4]), .B(n132), .ZN(N109) );
  NAND2_X1 U380 ( .A1(ref_1_port_o_3_1[6]), .A2(port_a_3[6]), .ZN(n132) );
  XNOR2_X1 U381 ( .A(port_rand_mul[2]), .B(n114), .ZN(N3) );
  NAND2_X1 U382 ( .A1(ref_1_port_o_0_3[0]), .A2(port_a_0[0]), .ZN(n114) );
  XNOR2_X1 U383 ( .A(port_rand_mul[2]), .B(n124), .ZN(N19) );
  NAND2_X1 U384 ( .A1(ref_1_port_o_0_3[1]), .A2(port_a_0[1]), .ZN(n124) );
  XNOR2_X1 U385 ( .A(port_rand_mul[2]), .B(n110), .ZN(N35) );
  NAND2_X1 U386 ( .A1(ref_1_port_o_0_3[2]), .A2(port_a_0[2]), .ZN(n110) );
  XNOR2_X1 U387 ( .A(port_rand_mul[2]), .B(n97), .ZN(N51) );
  NAND2_X1 U388 ( .A1(ref_1_port_o_0_3[3]), .A2(port_a_0[3]), .ZN(n97) );
  XNOR2_X1 U389 ( .A(port_rand_mul[2]), .B(n84), .ZN(N67) );
  NAND2_X1 U390 ( .A1(ref_1_port_o_0_3[4]), .A2(port_a_0[4]), .ZN(n84) );
  XNOR2_X1 U391 ( .A(port_rand_mul[2]), .B(n70), .ZN(N83) );
  NAND2_X1 U392 ( .A1(ref_1_port_o_0_3[5]), .A2(port_a_0[5]), .ZN(n70) );
  XNOR2_X1 U393 ( .A(port_rand_mul[2]), .B(n57), .ZN(N99) );
  NAND2_X1 U394 ( .A1(ref_1_port_o_0_3[6]), .A2(port_a_0[6]), .ZN(n57) );
  XNOR2_X1 U395 ( .A(port_rand_mul[4]), .B(n82), .ZN(N7) );
  NAND2_X1 U396 ( .A1(ref_1_port_o_1_3[0]), .A2(port_a_1[0]), .ZN(n82) );
  XNOR2_X1 U397 ( .A(port_rand_mul[4]), .B(n120), .ZN(N23) );
  NAND2_X1 U398 ( .A1(ref_1_port_o_1_3[1]), .A2(port_a_1[1]), .ZN(n120) );
  XNOR2_X1 U399 ( .A(port_rand_mul[4]), .B(n107), .ZN(N39) );
  NAND2_X1 U400 ( .A1(ref_1_port_o_1_3[2]), .A2(port_a_1[2]), .ZN(n107) );
  XNOR2_X1 U401 ( .A(port_rand_mul[4]), .B(n94), .ZN(N55) );
  NAND2_X1 U402 ( .A1(ref_1_port_o_1_3[3]), .A2(port_a_1[3]), .ZN(n94) );
  XNOR2_X1 U403 ( .A(port_rand_mul[4]), .B(n80), .ZN(N71) );
  NAND2_X1 U404 ( .A1(ref_1_port_o_1_3[4]), .A2(port_a_1[4]), .ZN(n80) );
  XNOR2_X1 U405 ( .A(port_rand_mul[4]), .B(n67), .ZN(N87) );
  NAND2_X1 U406 ( .A1(ref_1_port_o_1_3[5]), .A2(port_a_1[5]), .ZN(n67) );
  XNOR2_X1 U407 ( .A(port_rand_mul[4]), .B(n137), .ZN(N103) );
  NAND2_X1 U408 ( .A1(ref_1_port_o_1_3[6]), .A2(port_a_1[6]), .ZN(n137) );
  XNOR2_X1 U409 ( .A(port_rand_mul[5]), .B(n131), .ZN(N11) );
  NAND2_X1 U410 ( .A1(ref_1_port_o_2_3[0]), .A2(port_a_2[0]), .ZN(n131) );
  XNOR2_X1 U411 ( .A(port_rand_mul[5]), .B(n117), .ZN(N27) );
  NAND2_X1 U412 ( .A1(ref_1_port_o_2_3[1]), .A2(port_a_2[1]), .ZN(n117) );
  XNOR2_X1 U413 ( .A(port_rand_mul[5]), .B(n103), .ZN(N43) );
  NAND2_X1 U414 ( .A1(ref_1_port_o_2_3[2]), .A2(port_a_2[2]), .ZN(n103) );
  XNOR2_X1 U415 ( .A(port_rand_mul[5]), .B(n91), .ZN(N59) );
  NAND2_X1 U416 ( .A1(ref_1_port_o_2_3[3]), .A2(port_a_2[3]), .ZN(n91) );
  XNOR2_X1 U417 ( .A(port_rand_mul[5]), .B(n77), .ZN(N75) );
  NAND2_X1 U418 ( .A1(ref_1_port_o_2_3[4]), .A2(port_a_2[4]), .ZN(n77) );
  XNOR2_X1 U419 ( .A(port_rand_mul[5]), .B(n63), .ZN(N91) );
  NAND2_X1 U420 ( .A1(ref_1_port_o_2_3[5]), .A2(port_a_2[5]), .ZN(n63) );
  XNOR2_X1 U421 ( .A(port_rand_mul[5]), .B(n134), .ZN(N107) );
  NAND2_X1 U422 ( .A1(ref_1_port_o_2_3[6]), .A2(port_a_2[6]), .ZN(n134) );
  XNOR2_X1 U423 ( .A(port_rand_mul[1]), .B(n123), .ZN(N2) );
  NAND2_X1 U424 ( .A1(ref_1_port_o_0_2[0]), .A2(port_a_0[0]), .ZN(n123) );
  XNOR2_X1 U425 ( .A(port_rand_mul[1]), .B(n125), .ZN(N18) );
  NAND2_X1 U426 ( .A1(ref_1_port_o_0_2[1]), .A2(port_a_0[1]), .ZN(n125) );
  XNOR2_X1 U427 ( .A(port_rand_mul[1]), .B(n111), .ZN(N34) );
  NAND2_X1 U428 ( .A1(ref_1_port_o_0_2[2]), .A2(port_a_0[2]), .ZN(n111) );
  XNOR2_X1 U429 ( .A(port_rand_mul[1]), .B(n98), .ZN(N50) );
  NAND2_X1 U430 ( .A1(ref_1_port_o_0_2[3]), .A2(port_a_0[3]), .ZN(n98) );
  XNOR2_X1 U431 ( .A(port_rand_mul[1]), .B(n85), .ZN(N66) );
  NAND2_X1 U432 ( .A1(ref_1_port_o_0_2[4]), .A2(port_a_0[4]), .ZN(n85) );
  XNOR2_X1 U433 ( .A(port_rand_mul[1]), .B(n71), .ZN(N82) );
  NAND2_X1 U434 ( .A1(ref_1_port_o_0_2[5]), .A2(port_a_0[5]), .ZN(n71) );
  XNOR2_X1 U435 ( .A(port_rand_mul[1]), .B(n58), .ZN(N98) );
  NAND2_X1 U436 ( .A1(ref_1_port_o_0_2[6]), .A2(port_a_0[6]), .ZN(n58) );
  XNOR2_X1 U437 ( .A(port_rand_mul[0]), .B(n140), .ZN(N1) );
  NAND2_X1 U438 ( .A1(ref_1_port_o_0_1[0]), .A2(port_a_0[0]), .ZN(n140) );
  XNOR2_X1 U439 ( .A(port_rand_mul[0]), .B(n126), .ZN(N17) );
  NAND2_X1 U440 ( .A1(ref_1_port_o_0_1[1]), .A2(port_a_0[1]), .ZN(n126) );
  XNOR2_X1 U441 ( .A(port_rand_mul[0]), .B(n112), .ZN(N33) );
  NAND2_X1 U442 ( .A1(ref_1_port_o_0_1[2]), .A2(port_a_0[2]), .ZN(n112) );
  XNOR2_X1 U443 ( .A(port_rand_mul[0]), .B(n99), .ZN(N49) );
  NAND2_X1 U444 ( .A1(ref_1_port_o_0_1[3]), .A2(port_a_0[3]), .ZN(n99) );
  XNOR2_X1 U445 ( .A(port_rand_mul[0]), .B(n86), .ZN(N65) );
  NAND2_X1 U446 ( .A1(ref_1_port_o_0_1[4]), .A2(port_a_0[4]), .ZN(n86) );
  XNOR2_X1 U447 ( .A(port_rand_mul[0]), .B(n72), .ZN(N81) );
  NAND2_X1 U448 ( .A1(ref_1_port_o_0_1[5]), .A2(port_a_0[5]), .ZN(n72) );
  XNOR2_X1 U449 ( .A(port_rand_mul[0]), .B(n59), .ZN(N97) );
  NAND2_X1 U450 ( .A1(ref_1_port_o_0_1[6]), .A2(port_a_0[6]), .ZN(n59) );
  AND2_X1 U451 ( .A1(ref_1_port_o_2_2[0]), .A2(port_a_2[0]), .ZN(N10) );
  AND2_X1 U452 ( .A1(ref_1_port_o_2_2[1]), .A2(port_a_2[1]), .ZN(N26) );
  AND2_X1 U453 ( .A1(ref_1_port_o_2_2[2]), .A2(port_a_2[2]), .ZN(N42) );
  AND2_X1 U454 ( .A1(ref_1_port_o_2_2[3]), .A2(port_a_2[3]), .ZN(N58) );
  AND2_X1 U455 ( .A1(ref_1_port_o_2_2[4]), .A2(port_a_2[4]), .ZN(N74) );
  AND2_X1 U456 ( .A1(ref_1_port_o_2_2[5]), .A2(port_a_2[5]), .ZN(N90) );
  AND2_X1 U457 ( .A1(ref_1_port_o_2_2[6]), .A2(port_a_2[6]), .ZN(N106) );
  AND2_X1 U458 ( .A1(ref_1_port_o_1_1[0]), .A2(port_a_1[0]), .ZN(N5) );
  AND2_X1 U459 ( .A1(ref_1_port_o_1_1[1]), .A2(port_a_1[1]), .ZN(N21) );
  AND2_X1 U460 ( .A1(ref_1_port_o_1_1[2]), .A2(port_a_1[2]), .ZN(N37) );
  AND2_X1 U461 ( .A1(ref_1_port_o_1_1[3]), .A2(port_a_1[3]), .ZN(N53) );
  AND2_X1 U462 ( .A1(ref_1_port_o_1_1[4]), .A2(port_a_1[4]), .ZN(N69) );
  AND2_X1 U463 ( .A1(ref_1_port_o_1_1[5]), .A2(port_a_1[5]), .ZN(N85) );
  AND2_X1 U464 ( .A1(ref_1_port_o_1_1[6]), .A2(port_a_1[6]), .ZN(N101) );
  AND2_X1 U465 ( .A1(ref_1_port_o_3_3[0]), .A2(port_a_3[0]), .ZN(N15) );
  AND2_X1 U466 ( .A1(ref_1_port_o_3_3[1]), .A2(port_a_3[1]), .ZN(N31) );
  AND2_X1 U467 ( .A1(ref_1_port_o_3_3[2]), .A2(port_a_3[2]), .ZN(N47) );
  AND2_X1 U468 ( .A1(ref_1_port_o_3_3[3]), .A2(port_a_3[3]), .ZN(N63) );
  AND2_X1 U469 ( .A1(ref_1_port_o_3_3[4]), .A2(port_a_3[4]), .ZN(N79) );
  AND2_X1 U470 ( .A1(ref_1_port_o_3_3[5]), .A2(port_a_3[5]), .ZN(N95) );
  AND2_X1 U471 ( .A1(ref_1_port_o_3_3[6]), .A2(port_a_3[6]), .ZN(N111) );
  AND2_X1 U472 ( .A1(ref_1_port_o_0_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U473 ( .A1(ref_1_port_o_0_0[1]), .A2(port_a_0[1]), .ZN(N16) );
  AND2_X1 U474 ( .A1(ref_1_port_o_0_0[2]), .A2(port_a_0[2]), .ZN(N32) );
  AND2_X1 U475 ( .A1(ref_1_port_o_0_0[3]), .A2(port_a_0[3]), .ZN(N48) );
  AND2_X1 U476 ( .A1(ref_1_port_o_0_0[4]), .A2(port_a_0[4]), .ZN(N64) );
  AND2_X1 U477 ( .A1(ref_1_port_o_0_0[5]), .A2(port_a_0[5]), .ZN(N80) );
  AND2_X1 U478 ( .A1(ref_1_port_o_0_0[6]), .A2(port_a_0[6]), .ZN(N96) );
  XOR2_X1 U479 ( .A(n13), .B(n14), .Z(port_c_3[0]) );
  XNOR2_X1 U480 ( .A(temp_0_3[0]), .B(mult_ab_3_2[0]), .ZN(n13) );
  XNOR2_X1 U481 ( .A(mult_ab_3_1[0]), .B(mult_ab_3_0[0]), .ZN(n14) );
  XOR2_X1 U482 ( .A(n11), .B(n12), .Z(port_c_3[1]) );
  XNOR2_X1 U483 ( .A(temp_0_3[1]), .B(mult_ab_3_2[1]), .ZN(n11) );
  XNOR2_X1 U484 ( .A(mult_ab_3_1[1]), .B(mult_ab_3_0[1]), .ZN(n12) );
  XOR2_X1 U485 ( .A(n9), .B(n10), .Z(port_c_3[2]) );
  XNOR2_X1 U486 ( .A(temp_0_3[2]), .B(mult_ab_3_2[2]), .ZN(n9) );
  XNOR2_X1 U487 ( .A(mult_ab_3_1[2]), .B(mult_ab_3_0[2]), .ZN(n10) );
  XOR2_X1 U488 ( .A(n7), .B(n8), .Z(port_c_3[3]) );
  XNOR2_X1 U489 ( .A(temp_0_3[3]), .B(mult_ab_3_2[3]), .ZN(n7) );
  XNOR2_X1 U490 ( .A(mult_ab_3_1[3]), .B(mult_ab_3_0[3]), .ZN(n8) );
  XOR2_X1 U491 ( .A(n5), .B(n6), .Z(port_c_3[4]) );
  XNOR2_X1 U492 ( .A(temp_0_3[4]), .B(mult_ab_3_2[4]), .ZN(n5) );
  XNOR2_X1 U493 ( .A(mult_ab_3_1[4]), .B(mult_ab_3_0[4]), .ZN(n6) );
  XOR2_X1 U494 ( .A(n3), .B(n4), .Z(port_c_3[5]) );
  XNOR2_X1 U495 ( .A(temp_0_3[5]), .B(mult_ab_3_2[5]), .ZN(n3) );
  XNOR2_X1 U496 ( .A(mult_ab_3_1[5]), .B(mult_ab_3_0[5]), .ZN(n4) );
  XOR2_X1 U497 ( .A(n1), .B(n2), .Z(port_c_3[6]) );
  XNOR2_X1 U498 ( .A(temp_0_3[6]), .B(mult_ab_3_2[6]), .ZN(n1) );
  XNOR2_X1 U499 ( .A(mult_ab_3_1[6]), .B(mult_ab_3_0[6]), .ZN(n2) );
  XOR2_X1 U500 ( .A(n27), .B(n28), .Z(port_c_2[0]) );
  XNOR2_X1 U501 ( .A(temp_0_2[0]), .B(mult_ab_2_3[0]), .ZN(n27) );
  XNOR2_X1 U502 ( .A(mult_ab_2_1[0]), .B(mult_ab_2_0[0]), .ZN(n28) );
  XOR2_X1 U503 ( .A(n25), .B(n26), .Z(port_c_2[1]) );
  XNOR2_X1 U504 ( .A(temp_0_2[1]), .B(mult_ab_2_3[1]), .ZN(n25) );
  XNOR2_X1 U505 ( .A(mult_ab_2_1[1]), .B(mult_ab_2_0[1]), .ZN(n26) );
  XOR2_X1 U506 ( .A(n23), .B(n24), .Z(port_c_2[2]) );
  XNOR2_X1 U507 ( .A(temp_0_2[2]), .B(mult_ab_2_3[2]), .ZN(n23) );
  XNOR2_X1 U508 ( .A(mult_ab_2_1[2]), .B(mult_ab_2_0[2]), .ZN(n24) );
  XOR2_X1 U509 ( .A(n21), .B(n22), .Z(port_c_2[3]) );
  XNOR2_X1 U510 ( .A(temp_0_2[3]), .B(mult_ab_2_3[3]), .ZN(n21) );
  XNOR2_X1 U511 ( .A(mult_ab_2_1[3]), .B(mult_ab_2_0[3]), .ZN(n22) );
  XOR2_X1 U512 ( .A(n19), .B(n20), .Z(port_c_2[4]) );
  XNOR2_X1 U513 ( .A(temp_0_2[4]), .B(mult_ab_2_3[4]), .ZN(n19) );
  XNOR2_X1 U514 ( .A(mult_ab_2_1[4]), .B(mult_ab_2_0[4]), .ZN(n20) );
  XOR2_X1 U515 ( .A(n17), .B(n18), .Z(port_c_2[5]) );
  XNOR2_X1 U516 ( .A(temp_0_2[5]), .B(mult_ab_2_3[5]), .ZN(n17) );
  XNOR2_X1 U517 ( .A(mult_ab_2_1[5]), .B(mult_ab_2_0[5]), .ZN(n18) );
  XOR2_X1 U518 ( .A(n15), .B(n16), .Z(port_c_2[6]) );
  XNOR2_X1 U519 ( .A(temp_0_2[6]), .B(mult_ab_2_3[6]), .ZN(n15) );
  XNOR2_X1 U520 ( .A(mult_ab_2_1[6]), .B(mult_ab_2_0[6]), .ZN(n16) );
  XOR2_X1 U521 ( .A(n41), .B(n42), .Z(port_c_1[0]) );
  XNOR2_X1 U522 ( .A(temp_0_1[0]), .B(mult_ab_1_3[0]), .ZN(n41) );
  XNOR2_X1 U523 ( .A(mult_ab_1_2[0]), .B(mult_ab_1_0[0]), .ZN(n42) );
  XOR2_X1 U524 ( .A(n39), .B(n40), .Z(port_c_1[1]) );
  XNOR2_X1 U525 ( .A(temp_0_1[1]), .B(mult_ab_1_3[1]), .ZN(n39) );
  XNOR2_X1 U526 ( .A(mult_ab_1_2[1]), .B(mult_ab_1_0[1]), .ZN(n40) );
  XOR2_X1 U527 ( .A(n37), .B(n38), .Z(port_c_1[2]) );
  XNOR2_X1 U528 ( .A(temp_0_1[2]), .B(mult_ab_1_3[2]), .ZN(n37) );
  XNOR2_X1 U529 ( .A(mult_ab_1_2[2]), .B(mult_ab_1_0[2]), .ZN(n38) );
  XOR2_X1 U530 ( .A(n35), .B(n36), .Z(port_c_1[3]) );
  XNOR2_X1 U531 ( .A(temp_0_1[3]), .B(mult_ab_1_3[3]), .ZN(n35) );
  XNOR2_X1 U532 ( .A(mult_ab_1_2[3]), .B(mult_ab_1_0[3]), .ZN(n36) );
  XOR2_X1 U533 ( .A(n33), .B(n34), .Z(port_c_1[4]) );
  XNOR2_X1 U534 ( .A(temp_0_1[4]), .B(mult_ab_1_3[4]), .ZN(n33) );
  XNOR2_X1 U535 ( .A(mult_ab_1_2[4]), .B(mult_ab_1_0[4]), .ZN(n34) );
  XOR2_X1 U536 ( .A(n31), .B(n32), .Z(port_c_1[5]) );
  XNOR2_X1 U537 ( .A(temp_0_1[5]), .B(mult_ab_1_3[5]), .ZN(n31) );
  XNOR2_X1 U538 ( .A(mult_ab_1_2[5]), .B(mult_ab_1_0[5]), .ZN(n32) );
  XOR2_X1 U539 ( .A(n29), .B(n30), .Z(port_c_1[6]) );
  XNOR2_X1 U540 ( .A(temp_0_1[6]), .B(mult_ab_1_3[6]), .ZN(n29) );
  XNOR2_X1 U541 ( .A(mult_ab_1_2[6]), .B(mult_ab_1_0[6]), .ZN(n30) );
  XOR2_X1 U542 ( .A(n55), .B(n56), .Z(port_c_0[0]) );
  XNOR2_X1 U543 ( .A(temp_0_0[0]), .B(mult_ab_0_3[0]), .ZN(n55) );
  XNOR2_X1 U544 ( .A(mult_ab_0_2[0]), .B(mult_ab_0_1[0]), .ZN(n56) );
  XOR2_X1 U545 ( .A(n53), .B(n54), .Z(port_c_0[1]) );
  XNOR2_X1 U546 ( .A(temp_0_0[1]), .B(mult_ab_0_3[1]), .ZN(n53) );
  XNOR2_X1 U547 ( .A(mult_ab_0_2[1]), .B(mult_ab_0_1[1]), .ZN(n54) );
  XOR2_X1 U548 ( .A(n51), .B(n52), .Z(port_c_0[2]) );
  XNOR2_X1 U549 ( .A(temp_0_0[2]), .B(mult_ab_0_3[2]), .ZN(n51) );
  XNOR2_X1 U550 ( .A(mult_ab_0_2[2]), .B(mult_ab_0_1[2]), .ZN(n52) );
  XOR2_X1 U551 ( .A(n49), .B(n50), .Z(port_c_0[3]) );
  XNOR2_X1 U552 ( .A(temp_0_0[3]), .B(mult_ab_0_3[3]), .ZN(n49) );
  XNOR2_X1 U553 ( .A(mult_ab_0_2[3]), .B(mult_ab_0_1[3]), .ZN(n50) );
  XOR2_X1 U554 ( .A(n47), .B(n48), .Z(port_c_0[4]) );
  XNOR2_X1 U555 ( .A(temp_0_0[4]), .B(mult_ab_0_3[4]), .ZN(n47) );
  XNOR2_X1 U556 ( .A(mult_ab_0_2[4]), .B(mult_ab_0_1[4]), .ZN(n48) );
  XOR2_X1 U557 ( .A(n45), .B(n46), .Z(port_c_0[5]) );
  XNOR2_X1 U558 ( .A(temp_0_0[5]), .B(mult_ab_0_3[5]), .ZN(n45) );
  XNOR2_X1 U559 ( .A(mult_ab_0_2[5]), .B(mult_ab_0_1[5]), .ZN(n46) );
  XOR2_X1 U560 ( .A(n43), .B(n44), .Z(port_c_0[6]) );
  XNOR2_X1 U561 ( .A(temp_0_0[6]), .B(mult_ab_0_3[6]), .ZN(n43) );
  XNOR2_X1 U562 ( .A(mult_ab_0_2[6]), .B(mult_ab_0_1[6]), .ZN(n44) );
  BUF_X1 ref_1_U78 ( .A(ref_1_refreshed_0_6_), .Z(ref_1_n76) );
  BUF_X1 ref_1_U77 ( .A(ref_1_refreshed_1_6_), .Z(ref_1_n57) );
  BUF_X1 ref_1_U76 ( .A(ref_1_refreshed_2_6_), .Z(ref_1_n38) );
  BUF_X1 ref_1_U75 ( .A(ref_1_refreshed_3_6_), .Z(ref_1_n19) );
  BUF_X1 ref_1_U74 ( .A(ref_1_refreshed_0_5_), .Z(ref_1_n75) );
  BUF_X1 ref_1_U73 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n66) );
  BUF_X1 ref_1_U72 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n60) );
  BUF_X1 ref_1_U71 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n63) );
  BUF_X1 ref_1_U70 ( .A(ref_1_refreshed_0_5_), .Z(ref_1_n74) );
  BUF_X1 ref_1_U69 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n69) );
  BUF_X1 ref_1_U68 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n72) );
  BUF_X1 ref_1_U67 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n65) );
  BUF_X1 ref_1_U66 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n59) );
  BUF_X1 ref_1_U65 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n62) );
  BUF_X1 ref_1_U64 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n68) );
  BUF_X1 ref_1_U63 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n71) );
  BUF_X1 ref_1_U62 ( .A(ref_1_refreshed_0_2_), .Z(ref_1_n64) );
  BUF_X1 ref_1_U61 ( .A(ref_1_refreshed_0_0_), .Z(ref_1_n58) );
  BUF_X1 ref_1_U60 ( .A(ref_1_refreshed_0_1_), .Z(ref_1_n61) );
  BUF_X1 ref_1_U59 ( .A(ref_1_refreshed_0_5_), .Z(ref_1_n73) );
  BUF_X1 ref_1_U58 ( .A(ref_1_refreshed_0_3_), .Z(ref_1_n67) );
  BUF_X1 ref_1_U57 ( .A(ref_1_refreshed_0_4_), .Z(ref_1_n70) );
  BUF_X1 ref_1_U56 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n41) );
  BUF_X1 ref_1_U55 ( .A(ref_1_refreshed_1_5_), .Z(ref_1_n56) );
  BUF_X1 ref_1_U54 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n50) );
  BUF_X1 ref_1_U53 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n47) );
  BUF_X1 ref_1_U52 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n40) );
  BUF_X1 ref_1_U51 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n44) );
  BUF_X1 ref_1_U50 ( .A(ref_1_refreshed_1_5_), .Z(ref_1_n55) );
  BUF_X1 ref_1_U49 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n49) );
  BUF_X1 ref_1_U48 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n53) );
  BUF_X1 ref_1_U47 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n46) );
  BUF_X1 ref_1_U46 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n43) );
  BUF_X1 ref_1_U45 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n52) );
  BUF_X1 ref_1_U44 ( .A(ref_1_refreshed_1_2_), .Z(ref_1_n45) );
  BUF_X1 ref_1_U43 ( .A(ref_1_refreshed_1_0_), .Z(ref_1_n39) );
  BUF_X1 ref_1_U42 ( .A(ref_1_refreshed_1_1_), .Z(ref_1_n42) );
  BUF_X1 ref_1_U41 ( .A(ref_1_refreshed_1_5_), .Z(ref_1_n54) );
  BUF_X1 ref_1_U40 ( .A(ref_1_refreshed_1_3_), .Z(ref_1_n48) );
  BUF_X1 ref_1_U39 ( .A(ref_1_refreshed_1_4_), .Z(ref_1_n51) );
  BUF_X1 ref_1_U38 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n34) );
  BUF_X1 ref_1_U37 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n28) );
  BUF_X1 ref_1_U36 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n22) );
  BUF_X1 ref_1_U35 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n25) );
  BUF_X1 ref_1_U34 ( .A(ref_1_refreshed_2_5_), .Z(ref_1_n37) );
  BUF_X1 ref_1_U33 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n31) );
  BUF_X1 ref_1_U32 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n33) );
  BUF_X1 ref_1_U31 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n27) );
  BUF_X1 ref_1_U30 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n21) );
  BUF_X1 ref_1_U29 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n24) );
  BUF_X1 ref_1_U28 ( .A(ref_1_refreshed_2_5_), .Z(ref_1_n36) );
  BUF_X1 ref_1_U27 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n30) );
  BUF_X1 ref_1_U26 ( .A(ref_1_refreshed_2_2_), .Z(ref_1_n26) );
  BUF_X1 ref_1_U25 ( .A(ref_1_refreshed_2_0_), .Z(ref_1_n20) );
  BUF_X1 ref_1_U24 ( .A(ref_1_refreshed_2_1_), .Z(ref_1_n23) );
  BUF_X1 ref_1_U23 ( .A(ref_1_refreshed_2_5_), .Z(ref_1_n35) );
  BUF_X1 ref_1_U22 ( .A(ref_1_refreshed_2_3_), .Z(ref_1_n29) );
  BUF_X1 ref_1_U21 ( .A(ref_1_refreshed_2_4_), .Z(ref_1_n32) );
  BUF_X1 ref_1_U20 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n9) );
  BUF_X1 ref_1_U19 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n3) );
  BUF_X1 ref_1_U18 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n6) );
  BUF_X1 ref_1_U17 ( .A(ref_1_refreshed_3_5_), .Z(ref_1_n18) );
  BUF_X1 ref_1_U16 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n12) );
  BUF_X1 ref_1_U15 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n15) );
  BUF_X1 ref_1_U14 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n8) );
  BUF_X1 ref_1_U13 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n2) );
  BUF_X1 ref_1_U12 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n5) );
  BUF_X1 ref_1_U11 ( .A(ref_1_refreshed_3_5_), .Z(ref_1_n17) );
  BUF_X1 ref_1_U10 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n11) );
  BUF_X1 ref_1_U9 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n14) );
  BUF_X1 ref_1_U8 ( .A(ref_1_refreshed_3_2_), .Z(ref_1_n7) );
  BUF_X1 ref_1_U7 ( .A(ref_1_refreshed_3_0_), .Z(ref_1_n1) );
  BUF_X1 ref_1_U6 ( .A(ref_1_refreshed_3_1_), .Z(ref_1_n4) );
  BUF_X1 ref_1_U5 ( .A(ref_1_refreshed_3_5_), .Z(ref_1_n16) );
  BUF_X1 ref_1_U4 ( .A(ref_1_refreshed_3_3_), .Z(ref_1_n10) );
  BUF_X1 ref_1_U3 ( .A(ref_1_refreshed_3_4_), .Z(ref_1_n13) );
  DFF_X1 ref_1_reg_out_3_3_reg_0_ ( .D(ref_1_maj_127_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_1_ ( .D(ref_1_maj_143_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_2_ ( .D(ref_1_maj_159_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_3_ ( .D(ref_1_maj_175_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_4_ ( .D(ref_1_maj_191_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_5_ ( .D(ref_1_maj_207_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[5]), .QN() );
  DFF_X1 ref_1_reg_out_3_3_reg_6_ ( .D(ref_1_maj_223_port_o), .CK(clk), .Q(
        ref_1_port_o_3_3[6]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_0_ ( .D(ref_1_maj_126_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_1_ ( .D(ref_1_maj_142_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_2_ ( .D(ref_1_maj_158_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_3_ ( .D(ref_1_maj_174_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_4_ ( .D(ref_1_maj_190_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_5_ ( .D(ref_1_maj_206_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[5]), .QN() );
  DFF_X1 ref_1_reg_out_3_2_reg_6_ ( .D(ref_1_maj_222_port_o), .CK(clk), .Q(
        ref_1_port_o_3_2[6]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_0_ ( .D(ref_1_maj_125_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_1_ ( .D(ref_1_maj_141_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_2_ ( .D(ref_1_maj_157_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_3_ ( .D(ref_1_maj_173_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_4_ ( .D(ref_1_maj_189_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_5_ ( .D(ref_1_maj_205_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[5]), .QN() );
  DFF_X1 ref_1_reg_out_3_1_reg_6_ ( .D(ref_1_maj_221_port_o), .CK(clk), .Q(
        ref_1_port_o_3_1[6]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_0_ ( .D(ref_1_maj_124_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_1_ ( .D(ref_1_maj_140_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_2_ ( .D(ref_1_maj_156_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_3_ ( .D(ref_1_maj_172_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_4_ ( .D(ref_1_maj_188_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_5_ ( .D(ref_1_maj_204_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[5]), .QN() );
  DFF_X1 ref_1_reg_out_3_0_reg_6_ ( .D(ref_1_maj_220_port_o), .CK(clk), .Q(
        ref_1_port_o_3_0[6]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_0_ ( .D(ref_1_maj_123_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_1_ ( .D(ref_1_maj_139_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_2_ ( .D(ref_1_maj_155_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_3_ ( .D(ref_1_maj_171_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_4_ ( .D(ref_1_maj_187_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_5_ ( .D(ref_1_maj_203_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[5]), .QN() );
  DFF_X1 ref_1_reg_out_2_3_reg_6_ ( .D(ref_1_maj_219_port_o), .CK(clk), .Q(
        ref_1_port_o_2_3[6]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_0_ ( .D(ref_1_maj_122_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_1_ ( .D(ref_1_maj_138_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_2_ ( .D(ref_1_maj_154_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_3_ ( .D(ref_1_maj_170_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_4_ ( .D(ref_1_maj_186_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_5_ ( .D(ref_1_maj_202_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[5]), .QN() );
  DFF_X1 ref_1_reg_out_2_2_reg_6_ ( .D(ref_1_maj_218_port_o), .CK(clk), .Q(
        ref_1_port_o_2_2[6]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_0_ ( .D(ref_1_maj_121_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_1_ ( .D(ref_1_maj_137_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_2_ ( .D(ref_1_maj_153_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_3_ ( .D(ref_1_maj_169_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_4_ ( .D(ref_1_maj_185_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_5_ ( .D(ref_1_maj_201_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[5]), .QN() );
  DFF_X1 ref_1_reg_out_2_1_reg_6_ ( .D(ref_1_maj_217_port_o), .CK(clk), .Q(
        ref_1_port_o_2_1[6]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_0_ ( .D(ref_1_maj_120_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_1_ ( .D(ref_1_maj_136_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_2_ ( .D(ref_1_maj_152_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_3_ ( .D(ref_1_maj_168_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_4_ ( .D(ref_1_maj_184_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_5_ ( .D(ref_1_maj_200_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[5]), .QN() );
  DFF_X1 ref_1_reg_out_2_0_reg_6_ ( .D(ref_1_maj_216_port_o), .CK(clk), .Q(
        ref_1_port_o_2_0[6]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_0_ ( .D(ref_1_maj_119_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_1_ ( .D(ref_1_maj_135_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_2_ ( .D(ref_1_maj_151_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_3_ ( .D(ref_1_maj_167_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_4_ ( .D(ref_1_maj_183_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_5_ ( .D(ref_1_maj_199_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[5]), .QN() );
  DFF_X1 ref_1_reg_out_1_3_reg_6_ ( .D(ref_1_maj_215_port_o), .CK(clk), .Q(
        ref_1_port_o_1_3[6]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_0_ ( .D(ref_1_maj_118_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_1_ ( .D(ref_1_maj_134_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_2_ ( .D(ref_1_maj_150_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_3_ ( .D(ref_1_maj_166_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_4_ ( .D(ref_1_maj_182_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_5_ ( .D(ref_1_maj_198_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[5]), .QN() );
  DFF_X1 ref_1_reg_out_1_2_reg_6_ ( .D(ref_1_maj_214_port_o), .CK(clk), .Q(
        ref_1_port_o_1_2[6]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_0_ ( .D(ref_1_maj_117_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_1_ ( .D(ref_1_maj_133_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_2_ ( .D(ref_1_maj_149_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_3_ ( .D(ref_1_maj_165_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_4_ ( .D(ref_1_maj_181_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_5_ ( .D(ref_1_maj_197_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[5]), .QN() );
  DFF_X1 ref_1_reg_out_1_1_reg_6_ ( .D(ref_1_maj_213_port_o), .CK(clk), .Q(
        ref_1_port_o_1_1[6]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_0_ ( .D(ref_1_maj_116_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_1_ ( .D(ref_1_maj_132_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_2_ ( .D(ref_1_maj_148_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_3_ ( .D(ref_1_maj_164_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_4_ ( .D(ref_1_maj_180_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_5_ ( .D(ref_1_maj_196_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[5]), .QN() );
  DFF_X1 ref_1_reg_out_1_0_reg_6_ ( .D(ref_1_maj_212_port_o), .CK(clk), .Q(
        ref_1_port_o_1_0[6]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_0_ ( .D(ref_1_maj_115_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_1_ ( .D(ref_1_maj_131_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_2_ ( .D(ref_1_maj_147_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_3_ ( .D(ref_1_maj_163_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_4_ ( .D(ref_1_maj_179_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_5_ ( .D(ref_1_maj_195_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[5]), .QN() );
  DFF_X1 ref_1_reg_out_0_3_reg_6_ ( .D(ref_1_maj_211_port_o), .CK(clk), .Q(
        ref_1_port_o_0_3[6]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_0_ ( .D(ref_1_maj_114_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_1_ ( .D(ref_1_maj_130_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_2_ ( .D(ref_1_maj_146_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_3_ ( .D(ref_1_maj_162_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_4_ ( .D(ref_1_maj_178_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_5_ ( .D(ref_1_maj_194_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[5]), .QN() );
  DFF_X1 ref_1_reg_out_0_2_reg_6_ ( .D(ref_1_maj_210_port_o), .CK(clk), .Q(
        ref_1_port_o_0_2[6]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_0_ ( .D(ref_1_maj_113_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_1_ ( .D(ref_1_maj_129_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_2_ ( .D(ref_1_maj_145_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_3_ ( .D(ref_1_maj_161_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_4_ ( .D(ref_1_maj_177_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_5_ ( .D(ref_1_maj_193_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[5]), .QN() );
  DFF_X1 ref_1_reg_out_0_1_reg_6_ ( .D(ref_1_maj_209_port_o), .CK(clk), .Q(
        ref_1_port_o_0_1[6]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_0_ ( .D(ref_1_maj_112_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[0]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_1_ ( .D(ref_1_maj_128_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[1]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_2_ ( .D(ref_1_maj_144_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[2]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_3_ ( .D(ref_1_maj_160_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[3]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_4_ ( .D(ref_1_maj_176_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[4]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_5_ ( .D(ref_1_maj_192_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[5]), .QN() );
  DFF_X1 ref_1_reg_out_0_0_reg_6_ ( .D(ref_1_maj_208_port_o), .CK(clk), .Q(
        ref_1_port_o_0_0[6]), .QN() );
  XOR2_X1 ref_1_simpleXor_84_U1 ( .A(port_rand_ref[0]), .B(port_b_0[0]), .Z(
        ref_1_simpleXor_84_port_z) );
  XOR2_X1 ref_1_simpleXor_85_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_84_port_z), .Z(ref_1_simpleXor_85_port_z) );
  XOR2_X1 ref_1_simpleXor_86_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_85_port_z), .Z(ref_1_refreshed_0_0_) );
  XOR2_X1 ref_1_simpleXor_87_U1 ( .A(port_rand_ref[0]), .B(port_b_1[0]), .Z(
        ref_1_simpleXor_87_port_z) );
  XOR2_X1 ref_1_simpleXor_88_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_87_port_z), .Z(ref_1_simpleXor_88_port_z) );
  XOR2_X1 ref_1_simpleXor_89_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_88_port_z), .Z(ref_1_refreshed_1_0_) );
  XOR2_X1 ref_1_simpleXor_90_U1 ( .A(port_rand_ref[1]), .B(port_b_2[0]), .Z(
        ref_1_simpleXor_90_port_z) );
  XOR2_X1 ref_1_simpleXor_91_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_90_port_z), .Z(ref_1_simpleXor_91_port_z) );
  XOR2_X1 ref_1_simpleXor_92_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_91_port_z), .Z(ref_1_refreshed_2_0_) );
  XOR2_X1 ref_1_simpleXor_93_U1 ( .A(port_rand_ref[2]), .B(port_b_3[0]), .Z(
        ref_1_simpleXor_93_port_z) );
  XOR2_X1 ref_1_simpleXor_94_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_93_port_z), .Z(ref_1_simpleXor_94_port_z) );
  XOR2_X1 ref_1_simpleXor_95_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_94_port_z), .Z(ref_1_refreshed_3_0_) );
  XOR2_X1 ref_1_simpleXor_96_U1 ( .A(port_rand_ref[0]), .B(port_b_0[1]), .Z(
        ref_1_simpleXor_96_port_z) );
  XOR2_X1 ref_1_simpleXor_97_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_96_port_z), .Z(ref_1_simpleXor_97_port_z) );
  XOR2_X1 ref_1_simpleXor_98_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_97_port_z), .Z(ref_1_refreshed_0_1_) );
  XOR2_X1 ref_1_simpleXor_99_U1 ( .A(port_rand_ref[0]), .B(port_b_1[1]), .Z(
        ref_1_simpleXor_99_port_z) );
  XOR2_X1 ref_1_simpleXor_100_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_99_port_z), .Z(ref_1_simpleXor_100_port_z) );
  XOR2_X1 ref_1_simpleXor_101_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_100_port_z), .Z(ref_1_refreshed_1_1_) );
  XOR2_X1 ref_1_simpleXor_102_U1 ( .A(port_rand_ref[1]), .B(port_b_2[1]), .Z(
        ref_1_simpleXor_102_port_z) );
  XOR2_X1 ref_1_simpleXor_103_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_102_port_z), .Z(ref_1_simpleXor_103_port_z) );
  XOR2_X1 ref_1_simpleXor_104_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_103_port_z), .Z(ref_1_refreshed_2_1_) );
  XOR2_X1 ref_1_simpleXor_105_U1 ( .A(port_rand_ref[2]), .B(port_b_3[1]), .Z(
        ref_1_simpleXor_105_port_z) );
  XOR2_X1 ref_1_simpleXor_106_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_105_port_z), .Z(ref_1_simpleXor_106_port_z) );
  XOR2_X1 ref_1_simpleXor_107_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_106_port_z), .Z(ref_1_refreshed_3_1_) );
  XOR2_X1 ref_1_simpleXor_108_U1 ( .A(port_rand_ref[0]), .B(port_b_0[2]), .Z(
        ref_1_simpleXor_108_port_z) );
  XOR2_X1 ref_1_simpleXor_109_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_108_port_z), .Z(ref_1_simpleXor_109_port_z) );
  XOR2_X1 ref_1_simpleXor_110_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_109_port_z), .Z(ref_1_refreshed_0_2_) );
  XOR2_X1 ref_1_simpleXor_111_U1 ( .A(port_rand_ref[0]), .B(port_b_1[2]), .Z(
        ref_1_simpleXor_111_port_z) );
  XOR2_X1 ref_1_simpleXor_112_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_111_port_z), .Z(ref_1_simpleXor_112_port_z) );
  XOR2_X1 ref_1_simpleXor_113_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_112_port_z), .Z(ref_1_refreshed_1_2_) );
  XOR2_X1 ref_1_simpleXor_114_U1 ( .A(port_rand_ref[1]), .B(port_b_2[2]), .Z(
        ref_1_simpleXor_114_port_z) );
  XOR2_X1 ref_1_simpleXor_115_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_114_port_z), .Z(ref_1_simpleXor_115_port_z) );
  XOR2_X1 ref_1_simpleXor_116_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_115_port_z), .Z(ref_1_refreshed_2_2_) );
  XOR2_X1 ref_1_simpleXor_117_U1 ( .A(port_rand_ref[2]), .B(port_b_3[2]), .Z(
        ref_1_simpleXor_117_port_z) );
  XOR2_X1 ref_1_simpleXor_118_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_117_port_z), .Z(ref_1_simpleXor_118_port_z) );
  XOR2_X1 ref_1_simpleXor_119_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_118_port_z), .Z(ref_1_refreshed_3_2_) );
  XOR2_X1 ref_1_simpleXor_120_U1 ( .A(port_rand_ref[0]), .B(port_b_0[3]), .Z(
        ref_1_simpleXor_120_port_z) );
  XOR2_X1 ref_1_simpleXor_121_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_120_port_z), .Z(ref_1_simpleXor_121_port_z) );
  XOR2_X1 ref_1_simpleXor_122_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_121_port_z), .Z(ref_1_refreshed_0_3_) );
  XOR2_X1 ref_1_simpleXor_123_U1 ( .A(port_rand_ref[0]), .B(port_b_1[3]), .Z(
        ref_1_simpleXor_123_port_z) );
  XOR2_X1 ref_1_simpleXor_124_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_123_port_z), .Z(ref_1_simpleXor_124_port_z) );
  XOR2_X1 ref_1_simpleXor_125_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_124_port_z), .Z(ref_1_refreshed_1_3_) );
  XOR2_X1 ref_1_simpleXor_126_U1 ( .A(port_rand_ref[1]), .B(port_b_2[3]), .Z(
        ref_1_simpleXor_126_port_z) );
  XOR2_X1 ref_1_simpleXor_127_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_126_port_z), .Z(ref_1_simpleXor_127_port_z) );
  XOR2_X1 ref_1_simpleXor_128_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_127_port_z), .Z(ref_1_refreshed_2_3_) );
  XOR2_X1 ref_1_simpleXor_129_U1 ( .A(port_rand_ref[2]), .B(port_b_3[3]), .Z(
        ref_1_simpleXor_129_port_z) );
  XOR2_X1 ref_1_simpleXor_130_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_129_port_z), .Z(ref_1_simpleXor_130_port_z) );
  XOR2_X1 ref_1_simpleXor_131_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_130_port_z), .Z(ref_1_refreshed_3_3_) );
  XOR2_X1 ref_1_simpleXor_132_U1 ( .A(port_rand_ref[0]), .B(port_b_0[4]), .Z(
        ref_1_simpleXor_132_port_z) );
  XOR2_X1 ref_1_simpleXor_133_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_132_port_z), .Z(ref_1_simpleXor_133_port_z) );
  XOR2_X1 ref_1_simpleXor_134_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_133_port_z), .Z(ref_1_refreshed_0_4_) );
  XOR2_X1 ref_1_simpleXor_135_U1 ( .A(port_rand_ref[0]), .B(port_b_1[4]), .Z(
        ref_1_simpleXor_135_port_z) );
  XOR2_X1 ref_1_simpleXor_136_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_135_port_z), .Z(ref_1_simpleXor_136_port_z) );
  XOR2_X1 ref_1_simpleXor_137_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_136_port_z), .Z(ref_1_refreshed_1_4_) );
  XOR2_X1 ref_1_simpleXor_138_U1 ( .A(port_rand_ref[1]), .B(port_b_2[4]), .Z(
        ref_1_simpleXor_138_port_z) );
  XOR2_X1 ref_1_simpleXor_139_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_138_port_z), .Z(ref_1_simpleXor_139_port_z) );
  XOR2_X1 ref_1_simpleXor_140_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_139_port_z), .Z(ref_1_refreshed_2_4_) );
  XOR2_X1 ref_1_simpleXor_141_U1 ( .A(port_rand_ref[2]), .B(port_b_3[4]), .Z(
        ref_1_simpleXor_141_port_z) );
  XOR2_X1 ref_1_simpleXor_142_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_141_port_z), .Z(ref_1_simpleXor_142_port_z) );
  XOR2_X1 ref_1_simpleXor_143_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_142_port_z), .Z(ref_1_refreshed_3_4_) );
  XOR2_X1 ref_1_simpleXor_144_U1 ( .A(port_rand_ref[0]), .B(port_b_0[5]), .Z(
        ref_1_simpleXor_144_port_z) );
  XOR2_X1 ref_1_simpleXor_145_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_144_port_z), .Z(ref_1_simpleXor_145_port_z) );
  XOR2_X1 ref_1_simpleXor_146_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_145_port_z), .Z(ref_1_refreshed_0_5_) );
  XOR2_X1 ref_1_simpleXor_147_U1 ( .A(port_rand_ref[0]), .B(port_b_1[5]), .Z(
        ref_1_simpleXor_147_port_z) );
  XOR2_X1 ref_1_simpleXor_148_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_147_port_z), .Z(ref_1_simpleXor_148_port_z) );
  XOR2_X1 ref_1_simpleXor_149_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_148_port_z), .Z(ref_1_refreshed_1_5_) );
  XOR2_X1 ref_1_simpleXor_150_U1 ( .A(port_rand_ref[1]), .B(port_b_2[5]), .Z(
        ref_1_simpleXor_150_port_z) );
  XOR2_X1 ref_1_simpleXor_151_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_150_port_z), .Z(ref_1_simpleXor_151_port_z) );
  XOR2_X1 ref_1_simpleXor_152_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_151_port_z), .Z(ref_1_refreshed_2_5_) );
  XOR2_X1 ref_1_simpleXor_153_U1 ( .A(port_rand_ref[2]), .B(port_b_3[5]), .Z(
        ref_1_simpleXor_153_port_z) );
  XOR2_X1 ref_1_simpleXor_154_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_153_port_z), .Z(ref_1_simpleXor_154_port_z) );
  XOR2_X1 ref_1_simpleXor_155_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_154_port_z), .Z(ref_1_refreshed_3_5_) );
  XOR2_X1 ref_1_simpleXor_156_U1 ( .A(port_rand_ref[0]), .B(port_b_0[6]), .Z(
        ref_1_simpleXor_156_port_z) );
  XOR2_X1 ref_1_simpleXor_157_U1 ( .A(port_rand_ref[1]), .B(
        ref_1_simpleXor_156_port_z), .Z(ref_1_simpleXor_157_port_z) );
  XOR2_X1 ref_1_simpleXor_158_U1 ( .A(port_rand_ref[2]), .B(
        ref_1_simpleXor_157_port_z), .Z(ref_1_refreshed_0_6_) );
  XOR2_X1 ref_1_simpleXor_159_U1 ( .A(port_rand_ref[0]), .B(port_b_1[6]), .Z(
        ref_1_simpleXor_159_port_z) );
  XOR2_X1 ref_1_simpleXor_160_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_159_port_z), .Z(ref_1_simpleXor_160_port_z) );
  XOR2_X1 ref_1_simpleXor_161_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_160_port_z), .Z(ref_1_refreshed_1_6_) );
  XOR2_X1 ref_1_simpleXor_162_U1 ( .A(port_rand_ref[1]), .B(port_b_2[6]), .Z(
        ref_1_simpleXor_162_port_z) );
  XOR2_X1 ref_1_simpleXor_163_U1 ( .A(port_rand_ref[3]), .B(
        ref_1_simpleXor_162_port_z), .Z(ref_1_simpleXor_163_port_z) );
  XOR2_X1 ref_1_simpleXor_164_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_163_port_z), .Z(ref_1_refreshed_2_6_) );
  XOR2_X1 ref_1_simpleXor_165_U1 ( .A(port_rand_ref[2]), .B(port_b_3[6]), .Z(
        ref_1_simpleXor_165_port_z) );
  XOR2_X1 ref_1_simpleXor_166_U1 ( .A(port_rand_ref[4]), .B(
        ref_1_simpleXor_165_port_z), .Z(ref_1_simpleXor_166_port_z) );
  XOR2_X1 ref_1_simpleXor_167_U1 ( .A(port_rand_ref[5]), .B(
        ref_1_simpleXor_166_port_z), .Z(ref_1_refreshed_3_6_) );
  OR2_X1 ref_1_maj_112_U19 ( .A1(ref_1_maj_112_n8), .A2(ref_1_maj_112_n9), 
        .ZN(ref_1_maj_112_n7) );
  NAND2_X1 ref_1_maj_112_U18 ( .A1(ref_1_maj_112_n9), .A2(ref_1_maj_112_n8), 
        .ZN(ref_1_maj_112_n5) );
  NAND2_X1 ref_1_maj_112_U17 ( .A1(ref_1_refreshed_0_6_), .A2(ref_1_maj_112_n7), .ZN(ref_1_maj_112_n6) );
  NAND2_X1 ref_1_maj_112_U16 ( .A1(ref_1_maj_112_n5), .A2(ref_1_maj_112_n6), 
        .ZN(ref_1_maj_112_n4) );
  NAND2_X1 ref_1_maj_112_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_112_n10), .ZN(
        ref_1_maj_112_n17) );
  NAND2_X1 ref_1_maj_112_U14 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_112_n16) );
  NAND2_X1 ref_1_maj_112_U13 ( .A1(ref_1_maj_112_n16), .A2(ref_1_maj_112_n17), 
        .ZN(ref_1_maj_112_n13) );
  NAND2_X1 ref_1_maj_112_U12 ( .A1(ref_1_refreshed_0_2_), .A2(
        ref_1_maj_112_n11), .ZN(ref_1_maj_112_n15) );
  NAND2_X1 ref_1_maj_112_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_112_n14) );
  NAND2_X1 ref_1_maj_112_U10 ( .A1(ref_1_maj_112_n14), .A2(ref_1_maj_112_n15), 
        .ZN(ref_1_maj_112_n12) );
  XOR2_X1 ref_1_maj_112_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_112_n11), 
        .Z(ref_1_maj_112_n9) );
  XOR2_X1 ref_1_maj_112_U8 ( .A(ref_1_n75), .B(ref_1_maj_112_n10), .Z(
        ref_1_maj_112_n8) );
  XOR2_X1 ref_1_maj_112_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), .Z(ref_1_maj_112_n11) );
  XOR2_X1 ref_1_maj_112_U6 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), .Z(ref_1_maj_112_n10) );
  OR2_X1 ref_1_maj_112_U5 ( .A1(ref_1_maj_112_n12), .A2(ref_1_maj_112_n13), 
        .ZN(ref_1_maj_112_n3) );
  NAND2_X1 ref_1_maj_112_U4 ( .A1(ref_1_maj_112_n13), .A2(ref_1_maj_112_n12), 
        .ZN(ref_1_maj_112_n1) );
  NAND2_X1 ref_1_maj_112_U3 ( .A1(ref_1_maj_112_n3), .A2(ref_1_maj_112_n4), 
        .ZN(ref_1_maj_112_n2) );
  NAND2_X1 ref_1_maj_112_U2 ( .A1(ref_1_maj_112_n1), .A2(ref_1_maj_112_n2), 
        .ZN(ref_1_maj_112_port_o) );
  OR2_X1 ref_1_maj_113_U19 ( .A1(ref_1_maj_113_n27), .A2(ref_1_maj_113_n26), 
        .ZN(ref_1_maj_113_n28) );
  NAND2_X1 ref_1_maj_113_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_113_n28), .ZN(
        ref_1_maj_113_n29) );
  NAND2_X1 ref_1_maj_113_U17 ( .A1(ref_1_maj_113_n26), .A2(ref_1_maj_113_n27), 
        .ZN(ref_1_maj_113_n30) );
  NAND2_X1 ref_1_maj_113_U16 ( .A1(ref_1_maj_113_n30), .A2(ref_1_maj_113_n29), 
        .ZN(ref_1_maj_113_n31) );
  NAND2_X1 ref_1_maj_113_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_113_n25), .ZN(
        ref_1_maj_113_n18) );
  NAND2_X1 ref_1_maj_113_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_113_n19) );
  NAND2_X1 ref_1_maj_113_U13 ( .A1(ref_1_maj_113_n19), .A2(ref_1_maj_113_n18), 
        .ZN(ref_1_maj_113_n22) );
  NAND2_X1 ref_1_maj_113_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_113_n24), .ZN(
        ref_1_maj_113_n20) );
  NAND2_X1 ref_1_maj_113_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_113_n21) );
  NAND2_X1 ref_1_maj_113_U10 ( .A1(ref_1_maj_113_n21), .A2(ref_1_maj_113_n20), 
        .ZN(ref_1_maj_113_n23) );
  XOR2_X1 ref_1_maj_113_U9 ( .A(ref_1_n64), .B(ref_1_maj_113_n24), .Z(
        ref_1_maj_113_n26) );
  XOR2_X1 ref_1_maj_113_U8 ( .A(ref_1_n73), .B(ref_1_maj_113_n25), .Z(
        ref_1_maj_113_n27) );
  XOR2_X1 ref_1_maj_113_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_113_n24) );
  XOR2_X1 ref_1_maj_113_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_113_n25) );
  OR2_X1 ref_1_maj_113_U5 ( .A1(ref_1_maj_113_n23), .A2(ref_1_maj_113_n22), 
        .ZN(ref_1_maj_113_n32) );
  NAND2_X1 ref_1_maj_113_U4 ( .A1(ref_1_maj_113_n22), .A2(ref_1_maj_113_n23), 
        .ZN(ref_1_maj_113_n34) );
  NAND2_X1 ref_1_maj_113_U3 ( .A1(ref_1_maj_113_n32), .A2(ref_1_maj_113_n31), 
        .ZN(ref_1_maj_113_n33) );
  NAND2_X1 ref_1_maj_113_U2 ( .A1(ref_1_maj_113_n34), .A2(ref_1_maj_113_n33), 
        .ZN(ref_1_maj_113_port_o) );
  OR2_X1 ref_1_maj_114_U19 ( .A1(ref_1_maj_114_n27), .A2(ref_1_maj_114_n26), 
        .ZN(ref_1_maj_114_n28) );
  NAND2_X1 ref_1_maj_114_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_114_n28), .ZN(
        ref_1_maj_114_n29) );
  NAND2_X1 ref_1_maj_114_U17 ( .A1(ref_1_maj_114_n26), .A2(ref_1_maj_114_n27), 
        .ZN(ref_1_maj_114_n30) );
  NAND2_X1 ref_1_maj_114_U16 ( .A1(ref_1_maj_114_n30), .A2(ref_1_maj_114_n29), 
        .ZN(ref_1_maj_114_n31) );
  NAND2_X1 ref_1_maj_114_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_114_n25), .ZN(
        ref_1_maj_114_n18) );
  NAND2_X1 ref_1_maj_114_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_114_n19) );
  NAND2_X1 ref_1_maj_114_U13 ( .A1(ref_1_maj_114_n19), .A2(ref_1_maj_114_n18), 
        .ZN(ref_1_maj_114_n22) );
  NAND2_X1 ref_1_maj_114_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_114_n24), .ZN(
        ref_1_maj_114_n20) );
  NAND2_X1 ref_1_maj_114_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_114_n21) );
  NAND2_X1 ref_1_maj_114_U10 ( .A1(ref_1_maj_114_n21), .A2(ref_1_maj_114_n20), 
        .ZN(ref_1_maj_114_n23) );
  XOR2_X1 ref_1_maj_114_U9 ( .A(ref_1_n64), .B(ref_1_maj_114_n24), .Z(
        ref_1_maj_114_n26) );
  XOR2_X1 ref_1_maj_114_U8 ( .A(ref_1_n73), .B(ref_1_maj_114_n25), .Z(
        ref_1_maj_114_n27) );
  XOR2_X1 ref_1_maj_114_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_114_n24) );
  XOR2_X1 ref_1_maj_114_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_114_n25) );
  OR2_X1 ref_1_maj_114_U5 ( .A1(ref_1_maj_114_n23), .A2(ref_1_maj_114_n22), 
        .ZN(ref_1_maj_114_n32) );
  NAND2_X1 ref_1_maj_114_U4 ( .A1(ref_1_maj_114_n22), .A2(ref_1_maj_114_n23), 
        .ZN(ref_1_maj_114_n34) );
  NAND2_X1 ref_1_maj_114_U3 ( .A1(ref_1_maj_114_n32), .A2(ref_1_maj_114_n31), 
        .ZN(ref_1_maj_114_n33) );
  NAND2_X1 ref_1_maj_114_U2 ( .A1(ref_1_maj_114_n34), .A2(ref_1_maj_114_n33), 
        .ZN(ref_1_maj_114_port_o) );
  OR2_X1 ref_1_maj_115_U19 ( .A1(ref_1_maj_115_n27), .A2(ref_1_maj_115_n26), 
        .ZN(ref_1_maj_115_n28) );
  NAND2_X1 ref_1_maj_115_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_115_n28), .ZN(
        ref_1_maj_115_n29) );
  NAND2_X1 ref_1_maj_115_U17 ( .A1(ref_1_maj_115_n26), .A2(ref_1_maj_115_n27), 
        .ZN(ref_1_maj_115_n30) );
  NAND2_X1 ref_1_maj_115_U16 ( .A1(ref_1_maj_115_n30), .A2(ref_1_maj_115_n29), 
        .ZN(ref_1_maj_115_n31) );
  NAND2_X1 ref_1_maj_115_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_115_n25), .ZN(
        ref_1_maj_115_n18) );
  NAND2_X1 ref_1_maj_115_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_115_n19) );
  NAND2_X1 ref_1_maj_115_U13 ( .A1(ref_1_maj_115_n19), .A2(ref_1_maj_115_n18), 
        .ZN(ref_1_maj_115_n22) );
  NAND2_X1 ref_1_maj_115_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_115_n24), .ZN(
        ref_1_maj_115_n20) );
  NAND2_X1 ref_1_maj_115_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_115_n21) );
  NAND2_X1 ref_1_maj_115_U10 ( .A1(ref_1_maj_115_n21), .A2(ref_1_maj_115_n20), 
        .ZN(ref_1_maj_115_n23) );
  XOR2_X1 ref_1_maj_115_U9 ( .A(ref_1_n64), .B(ref_1_maj_115_n24), .Z(
        ref_1_maj_115_n26) );
  XOR2_X1 ref_1_maj_115_U8 ( .A(ref_1_n73), .B(ref_1_maj_115_n25), .Z(
        ref_1_maj_115_n27) );
  XOR2_X1 ref_1_maj_115_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_115_n24) );
  XOR2_X1 ref_1_maj_115_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_115_n25) );
  OR2_X1 ref_1_maj_115_U5 ( .A1(ref_1_maj_115_n23), .A2(ref_1_maj_115_n22), 
        .ZN(ref_1_maj_115_n32) );
  NAND2_X1 ref_1_maj_115_U4 ( .A1(ref_1_maj_115_n22), .A2(ref_1_maj_115_n23), 
        .ZN(ref_1_maj_115_n34) );
  NAND2_X1 ref_1_maj_115_U3 ( .A1(ref_1_maj_115_n32), .A2(ref_1_maj_115_n31), 
        .ZN(ref_1_maj_115_n33) );
  NAND2_X1 ref_1_maj_115_U2 ( .A1(ref_1_maj_115_n34), .A2(ref_1_maj_115_n33), 
        .ZN(ref_1_maj_115_port_o) );
  OR2_X1 ref_1_maj_116_U19 ( .A1(ref_1_maj_116_n27), .A2(ref_1_maj_116_n26), 
        .ZN(ref_1_maj_116_n28) );
  NAND2_X1 ref_1_maj_116_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_116_n28), .ZN(
        ref_1_maj_116_n29) );
  NAND2_X1 ref_1_maj_116_U17 ( .A1(ref_1_maj_116_n26), .A2(ref_1_maj_116_n27), 
        .ZN(ref_1_maj_116_n30) );
  NAND2_X1 ref_1_maj_116_U16 ( .A1(ref_1_maj_116_n30), .A2(ref_1_maj_116_n29), 
        .ZN(ref_1_maj_116_n31) );
  NAND2_X1 ref_1_maj_116_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_116_n25), .ZN(
        ref_1_maj_116_n18) );
  NAND2_X1 ref_1_maj_116_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_116_n19) );
  NAND2_X1 ref_1_maj_116_U13 ( .A1(ref_1_maj_116_n19), .A2(ref_1_maj_116_n18), 
        .ZN(ref_1_maj_116_n22) );
  NAND2_X1 ref_1_maj_116_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_116_n24), .ZN(
        ref_1_maj_116_n20) );
  NAND2_X1 ref_1_maj_116_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_116_n21) );
  NAND2_X1 ref_1_maj_116_U10 ( .A1(ref_1_maj_116_n21), .A2(ref_1_maj_116_n20), 
        .ZN(ref_1_maj_116_n23) );
  XOR2_X1 ref_1_maj_116_U9 ( .A(ref_1_n45), .B(ref_1_maj_116_n24), .Z(
        ref_1_maj_116_n26) );
  XOR2_X1 ref_1_maj_116_U8 ( .A(ref_1_n54), .B(ref_1_maj_116_n25), .Z(
        ref_1_maj_116_n27) );
  XOR2_X1 ref_1_maj_116_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_116_n24) );
  XOR2_X1 ref_1_maj_116_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_116_n25) );
  OR2_X1 ref_1_maj_116_U5 ( .A1(ref_1_maj_116_n23), .A2(ref_1_maj_116_n22), 
        .ZN(ref_1_maj_116_n32) );
  NAND2_X1 ref_1_maj_116_U4 ( .A1(ref_1_maj_116_n22), .A2(ref_1_maj_116_n23), 
        .ZN(ref_1_maj_116_n34) );
  NAND2_X1 ref_1_maj_116_U3 ( .A1(ref_1_maj_116_n32), .A2(ref_1_maj_116_n31), 
        .ZN(ref_1_maj_116_n33) );
  NAND2_X1 ref_1_maj_116_U2 ( .A1(ref_1_maj_116_n34), .A2(ref_1_maj_116_n33), 
        .ZN(ref_1_maj_116_port_o) );
  OR2_X1 ref_1_maj_117_U19 ( .A1(ref_1_maj_117_n27), .A2(ref_1_maj_117_n26), 
        .ZN(ref_1_maj_117_n28) );
  NAND2_X1 ref_1_maj_117_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_117_n28), .ZN(
        ref_1_maj_117_n29) );
  NAND2_X1 ref_1_maj_117_U17 ( .A1(ref_1_maj_117_n26), .A2(ref_1_maj_117_n27), 
        .ZN(ref_1_maj_117_n30) );
  NAND2_X1 ref_1_maj_117_U16 ( .A1(ref_1_maj_117_n30), .A2(ref_1_maj_117_n29), 
        .ZN(ref_1_maj_117_n31) );
  NAND2_X1 ref_1_maj_117_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_117_n25), .ZN(
        ref_1_maj_117_n18) );
  NAND2_X1 ref_1_maj_117_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_117_n19) );
  NAND2_X1 ref_1_maj_117_U13 ( .A1(ref_1_maj_117_n19), .A2(ref_1_maj_117_n18), 
        .ZN(ref_1_maj_117_n22) );
  NAND2_X1 ref_1_maj_117_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_117_n24), .ZN(
        ref_1_maj_117_n20) );
  NAND2_X1 ref_1_maj_117_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_117_n21) );
  NAND2_X1 ref_1_maj_117_U10 ( .A1(ref_1_maj_117_n21), .A2(ref_1_maj_117_n20), 
        .ZN(ref_1_maj_117_n23) );
  XOR2_X1 ref_1_maj_117_U9 ( .A(ref_1_n45), .B(ref_1_maj_117_n24), .Z(
        ref_1_maj_117_n26) );
  XOR2_X1 ref_1_maj_117_U8 ( .A(ref_1_n54), .B(ref_1_maj_117_n25), .Z(
        ref_1_maj_117_n27) );
  XOR2_X1 ref_1_maj_117_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_117_n24) );
  XOR2_X1 ref_1_maj_117_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_117_n25) );
  OR2_X1 ref_1_maj_117_U5 ( .A1(ref_1_maj_117_n23), .A2(ref_1_maj_117_n22), 
        .ZN(ref_1_maj_117_n32) );
  NAND2_X1 ref_1_maj_117_U4 ( .A1(ref_1_maj_117_n22), .A2(ref_1_maj_117_n23), 
        .ZN(ref_1_maj_117_n34) );
  NAND2_X1 ref_1_maj_117_U3 ( .A1(ref_1_maj_117_n32), .A2(ref_1_maj_117_n31), 
        .ZN(ref_1_maj_117_n33) );
  NAND2_X1 ref_1_maj_117_U2 ( .A1(ref_1_maj_117_n34), .A2(ref_1_maj_117_n33), 
        .ZN(ref_1_maj_117_port_o) );
  OR2_X1 ref_1_maj_118_U19 ( .A1(ref_1_maj_118_n27), .A2(ref_1_maj_118_n26), 
        .ZN(ref_1_maj_118_n28) );
  NAND2_X1 ref_1_maj_118_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_118_n28), .ZN(
        ref_1_maj_118_n29) );
  NAND2_X1 ref_1_maj_118_U17 ( .A1(ref_1_maj_118_n26), .A2(ref_1_maj_118_n27), 
        .ZN(ref_1_maj_118_n30) );
  NAND2_X1 ref_1_maj_118_U16 ( .A1(ref_1_maj_118_n30), .A2(ref_1_maj_118_n29), 
        .ZN(ref_1_maj_118_n31) );
  NAND2_X1 ref_1_maj_118_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_118_n25), .ZN(
        ref_1_maj_118_n18) );
  NAND2_X1 ref_1_maj_118_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_118_n19) );
  NAND2_X1 ref_1_maj_118_U13 ( .A1(ref_1_maj_118_n19), .A2(ref_1_maj_118_n18), 
        .ZN(ref_1_maj_118_n22) );
  NAND2_X1 ref_1_maj_118_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_118_n24), .ZN(
        ref_1_maj_118_n20) );
  NAND2_X1 ref_1_maj_118_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_118_n21) );
  NAND2_X1 ref_1_maj_118_U10 ( .A1(ref_1_maj_118_n21), .A2(ref_1_maj_118_n20), 
        .ZN(ref_1_maj_118_n23) );
  XOR2_X1 ref_1_maj_118_U9 ( .A(ref_1_n45), .B(ref_1_maj_118_n24), .Z(
        ref_1_maj_118_n26) );
  XOR2_X1 ref_1_maj_118_U8 ( .A(ref_1_n54), .B(ref_1_maj_118_n25), .Z(
        ref_1_maj_118_n27) );
  XOR2_X1 ref_1_maj_118_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_118_n24) );
  XOR2_X1 ref_1_maj_118_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_118_n25) );
  OR2_X1 ref_1_maj_118_U5 ( .A1(ref_1_maj_118_n23), .A2(ref_1_maj_118_n22), 
        .ZN(ref_1_maj_118_n32) );
  NAND2_X1 ref_1_maj_118_U4 ( .A1(ref_1_maj_118_n22), .A2(ref_1_maj_118_n23), 
        .ZN(ref_1_maj_118_n34) );
  NAND2_X1 ref_1_maj_118_U3 ( .A1(ref_1_maj_118_n32), .A2(ref_1_maj_118_n31), 
        .ZN(ref_1_maj_118_n33) );
  NAND2_X1 ref_1_maj_118_U2 ( .A1(ref_1_maj_118_n34), .A2(ref_1_maj_118_n33), 
        .ZN(ref_1_maj_118_port_o) );
  OR2_X1 ref_1_maj_119_U19 ( .A1(ref_1_maj_119_n27), .A2(ref_1_maj_119_n26), 
        .ZN(ref_1_maj_119_n28) );
  NAND2_X1 ref_1_maj_119_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_119_n28), .ZN(
        ref_1_maj_119_n29) );
  NAND2_X1 ref_1_maj_119_U17 ( .A1(ref_1_maj_119_n26), .A2(ref_1_maj_119_n27), 
        .ZN(ref_1_maj_119_n30) );
  NAND2_X1 ref_1_maj_119_U16 ( .A1(ref_1_maj_119_n30), .A2(ref_1_maj_119_n29), 
        .ZN(ref_1_maj_119_n31) );
  NAND2_X1 ref_1_maj_119_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_119_n25), .ZN(
        ref_1_maj_119_n18) );
  NAND2_X1 ref_1_maj_119_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_119_n19) );
  NAND2_X1 ref_1_maj_119_U13 ( .A1(ref_1_maj_119_n19), .A2(ref_1_maj_119_n18), 
        .ZN(ref_1_maj_119_n22) );
  NAND2_X1 ref_1_maj_119_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_119_n24), .ZN(
        ref_1_maj_119_n20) );
  NAND2_X1 ref_1_maj_119_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_119_n21) );
  NAND2_X1 ref_1_maj_119_U10 ( .A1(ref_1_maj_119_n21), .A2(ref_1_maj_119_n20), 
        .ZN(ref_1_maj_119_n23) );
  XOR2_X1 ref_1_maj_119_U9 ( .A(ref_1_n45), .B(ref_1_maj_119_n24), .Z(
        ref_1_maj_119_n26) );
  XOR2_X1 ref_1_maj_119_U8 ( .A(ref_1_n54), .B(ref_1_maj_119_n25), .Z(
        ref_1_maj_119_n27) );
  XOR2_X1 ref_1_maj_119_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_119_n24) );
  XOR2_X1 ref_1_maj_119_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_119_n25) );
  OR2_X1 ref_1_maj_119_U5 ( .A1(ref_1_maj_119_n23), .A2(ref_1_maj_119_n22), 
        .ZN(ref_1_maj_119_n32) );
  NAND2_X1 ref_1_maj_119_U4 ( .A1(ref_1_maj_119_n22), .A2(ref_1_maj_119_n23), 
        .ZN(ref_1_maj_119_n34) );
  NAND2_X1 ref_1_maj_119_U3 ( .A1(ref_1_maj_119_n32), .A2(ref_1_maj_119_n31), 
        .ZN(ref_1_maj_119_n33) );
  NAND2_X1 ref_1_maj_119_U2 ( .A1(ref_1_maj_119_n34), .A2(ref_1_maj_119_n33), 
        .ZN(ref_1_maj_119_port_o) );
  OR2_X1 ref_1_maj_120_U19 ( .A1(ref_1_maj_120_n27), .A2(ref_1_maj_120_n26), 
        .ZN(ref_1_maj_120_n28) );
  NAND2_X1 ref_1_maj_120_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_120_n28), .ZN(
        ref_1_maj_120_n29) );
  NAND2_X1 ref_1_maj_120_U17 ( .A1(ref_1_maj_120_n26), .A2(ref_1_maj_120_n27), 
        .ZN(ref_1_maj_120_n30) );
  NAND2_X1 ref_1_maj_120_U16 ( .A1(ref_1_maj_120_n30), .A2(ref_1_maj_120_n29), 
        .ZN(ref_1_maj_120_n31) );
  NAND2_X1 ref_1_maj_120_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_120_n25), .ZN(
        ref_1_maj_120_n18) );
  NAND2_X1 ref_1_maj_120_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_120_n19) );
  NAND2_X1 ref_1_maj_120_U13 ( .A1(ref_1_maj_120_n19), .A2(ref_1_maj_120_n18), 
        .ZN(ref_1_maj_120_n22) );
  NAND2_X1 ref_1_maj_120_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_120_n24), .ZN(
        ref_1_maj_120_n20) );
  NAND2_X1 ref_1_maj_120_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_120_n21) );
  NAND2_X1 ref_1_maj_120_U10 ( .A1(ref_1_maj_120_n21), .A2(ref_1_maj_120_n20), 
        .ZN(ref_1_maj_120_n23) );
  XOR2_X1 ref_1_maj_120_U9 ( .A(ref_1_n26), .B(ref_1_maj_120_n24), .Z(
        ref_1_maj_120_n26) );
  XOR2_X1 ref_1_maj_120_U8 ( .A(ref_1_n35), .B(ref_1_maj_120_n25), .Z(
        ref_1_maj_120_n27) );
  XOR2_X1 ref_1_maj_120_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_120_n24) );
  XOR2_X1 ref_1_maj_120_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_120_n25) );
  OR2_X1 ref_1_maj_120_U5 ( .A1(ref_1_maj_120_n23), .A2(ref_1_maj_120_n22), 
        .ZN(ref_1_maj_120_n32) );
  NAND2_X1 ref_1_maj_120_U4 ( .A1(ref_1_maj_120_n22), .A2(ref_1_maj_120_n23), 
        .ZN(ref_1_maj_120_n34) );
  NAND2_X1 ref_1_maj_120_U3 ( .A1(ref_1_maj_120_n32), .A2(ref_1_maj_120_n31), 
        .ZN(ref_1_maj_120_n33) );
  NAND2_X1 ref_1_maj_120_U2 ( .A1(ref_1_maj_120_n34), .A2(ref_1_maj_120_n33), 
        .ZN(ref_1_maj_120_port_o) );
  OR2_X1 ref_1_maj_121_U19 ( .A1(ref_1_maj_121_n27), .A2(ref_1_maj_121_n26), 
        .ZN(ref_1_maj_121_n28) );
  NAND2_X1 ref_1_maj_121_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_121_n28), .ZN(
        ref_1_maj_121_n29) );
  NAND2_X1 ref_1_maj_121_U17 ( .A1(ref_1_maj_121_n26), .A2(ref_1_maj_121_n27), 
        .ZN(ref_1_maj_121_n30) );
  NAND2_X1 ref_1_maj_121_U16 ( .A1(ref_1_maj_121_n30), .A2(ref_1_maj_121_n29), 
        .ZN(ref_1_maj_121_n31) );
  NAND2_X1 ref_1_maj_121_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_121_n25), .ZN(
        ref_1_maj_121_n18) );
  NAND2_X1 ref_1_maj_121_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_121_n19) );
  NAND2_X1 ref_1_maj_121_U13 ( .A1(ref_1_maj_121_n19), .A2(ref_1_maj_121_n18), 
        .ZN(ref_1_maj_121_n22) );
  NAND2_X1 ref_1_maj_121_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_121_n24), .ZN(
        ref_1_maj_121_n20) );
  NAND2_X1 ref_1_maj_121_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_121_n21) );
  NAND2_X1 ref_1_maj_121_U10 ( .A1(ref_1_maj_121_n21), .A2(ref_1_maj_121_n20), 
        .ZN(ref_1_maj_121_n23) );
  XOR2_X1 ref_1_maj_121_U9 ( .A(ref_1_n26), .B(ref_1_maj_121_n24), .Z(
        ref_1_maj_121_n26) );
  XOR2_X1 ref_1_maj_121_U8 ( .A(ref_1_n35), .B(ref_1_maj_121_n25), .Z(
        ref_1_maj_121_n27) );
  XOR2_X1 ref_1_maj_121_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_121_n24) );
  XOR2_X1 ref_1_maj_121_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_121_n25) );
  OR2_X1 ref_1_maj_121_U5 ( .A1(ref_1_maj_121_n23), .A2(ref_1_maj_121_n22), 
        .ZN(ref_1_maj_121_n32) );
  NAND2_X1 ref_1_maj_121_U4 ( .A1(ref_1_maj_121_n22), .A2(ref_1_maj_121_n23), 
        .ZN(ref_1_maj_121_n34) );
  NAND2_X1 ref_1_maj_121_U3 ( .A1(ref_1_maj_121_n32), .A2(ref_1_maj_121_n31), 
        .ZN(ref_1_maj_121_n33) );
  NAND2_X1 ref_1_maj_121_U2 ( .A1(ref_1_maj_121_n34), .A2(ref_1_maj_121_n33), 
        .ZN(ref_1_maj_121_port_o) );
  OR2_X1 ref_1_maj_122_U19 ( .A1(ref_1_maj_122_n27), .A2(ref_1_maj_122_n26), 
        .ZN(ref_1_maj_122_n28) );
  NAND2_X1 ref_1_maj_122_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_122_n28), .ZN(
        ref_1_maj_122_n29) );
  NAND2_X1 ref_1_maj_122_U17 ( .A1(ref_1_maj_122_n26), .A2(ref_1_maj_122_n27), 
        .ZN(ref_1_maj_122_n30) );
  NAND2_X1 ref_1_maj_122_U16 ( .A1(ref_1_maj_122_n30), .A2(ref_1_maj_122_n29), 
        .ZN(ref_1_maj_122_n31) );
  NAND2_X1 ref_1_maj_122_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_122_n25), .ZN(
        ref_1_maj_122_n18) );
  NAND2_X1 ref_1_maj_122_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_122_n19) );
  NAND2_X1 ref_1_maj_122_U13 ( .A1(ref_1_maj_122_n19), .A2(ref_1_maj_122_n18), 
        .ZN(ref_1_maj_122_n22) );
  NAND2_X1 ref_1_maj_122_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_122_n24), .ZN(
        ref_1_maj_122_n20) );
  NAND2_X1 ref_1_maj_122_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_122_n21) );
  NAND2_X1 ref_1_maj_122_U10 ( .A1(ref_1_maj_122_n21), .A2(ref_1_maj_122_n20), 
        .ZN(ref_1_maj_122_n23) );
  XOR2_X1 ref_1_maj_122_U9 ( .A(ref_1_n26), .B(ref_1_maj_122_n24), .Z(
        ref_1_maj_122_n26) );
  XOR2_X1 ref_1_maj_122_U8 ( .A(ref_1_n35), .B(ref_1_maj_122_n25), .Z(
        ref_1_maj_122_n27) );
  XOR2_X1 ref_1_maj_122_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_122_n24) );
  XOR2_X1 ref_1_maj_122_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_122_n25) );
  OR2_X1 ref_1_maj_122_U5 ( .A1(ref_1_maj_122_n23), .A2(ref_1_maj_122_n22), 
        .ZN(ref_1_maj_122_n32) );
  NAND2_X1 ref_1_maj_122_U4 ( .A1(ref_1_maj_122_n22), .A2(ref_1_maj_122_n23), 
        .ZN(ref_1_maj_122_n34) );
  NAND2_X1 ref_1_maj_122_U3 ( .A1(ref_1_maj_122_n32), .A2(ref_1_maj_122_n31), 
        .ZN(ref_1_maj_122_n33) );
  NAND2_X1 ref_1_maj_122_U2 ( .A1(ref_1_maj_122_n34), .A2(ref_1_maj_122_n33), 
        .ZN(ref_1_maj_122_port_o) );
  OR2_X1 ref_1_maj_123_U19 ( .A1(ref_1_maj_123_n27), .A2(ref_1_maj_123_n26), 
        .ZN(ref_1_maj_123_n28) );
  NAND2_X1 ref_1_maj_123_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_123_n28), .ZN(
        ref_1_maj_123_n29) );
  NAND2_X1 ref_1_maj_123_U17 ( .A1(ref_1_maj_123_n26), .A2(ref_1_maj_123_n27), 
        .ZN(ref_1_maj_123_n30) );
  NAND2_X1 ref_1_maj_123_U16 ( .A1(ref_1_maj_123_n30), .A2(ref_1_maj_123_n29), 
        .ZN(ref_1_maj_123_n31) );
  NAND2_X1 ref_1_maj_123_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_123_n25), .ZN(
        ref_1_maj_123_n18) );
  NAND2_X1 ref_1_maj_123_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_123_n19) );
  NAND2_X1 ref_1_maj_123_U13 ( .A1(ref_1_maj_123_n19), .A2(ref_1_maj_123_n18), 
        .ZN(ref_1_maj_123_n22) );
  NAND2_X1 ref_1_maj_123_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_123_n24), .ZN(
        ref_1_maj_123_n20) );
  NAND2_X1 ref_1_maj_123_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_123_n21) );
  NAND2_X1 ref_1_maj_123_U10 ( .A1(ref_1_maj_123_n21), .A2(ref_1_maj_123_n20), 
        .ZN(ref_1_maj_123_n23) );
  XOR2_X1 ref_1_maj_123_U9 ( .A(ref_1_n26), .B(ref_1_maj_123_n24), .Z(
        ref_1_maj_123_n26) );
  XOR2_X1 ref_1_maj_123_U8 ( .A(ref_1_n35), .B(ref_1_maj_123_n25), .Z(
        ref_1_maj_123_n27) );
  XOR2_X1 ref_1_maj_123_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_123_n24) );
  XOR2_X1 ref_1_maj_123_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_123_n25) );
  OR2_X1 ref_1_maj_123_U5 ( .A1(ref_1_maj_123_n23), .A2(ref_1_maj_123_n22), 
        .ZN(ref_1_maj_123_n32) );
  NAND2_X1 ref_1_maj_123_U4 ( .A1(ref_1_maj_123_n22), .A2(ref_1_maj_123_n23), 
        .ZN(ref_1_maj_123_n34) );
  NAND2_X1 ref_1_maj_123_U3 ( .A1(ref_1_maj_123_n32), .A2(ref_1_maj_123_n31), 
        .ZN(ref_1_maj_123_n33) );
  NAND2_X1 ref_1_maj_123_U2 ( .A1(ref_1_maj_123_n34), .A2(ref_1_maj_123_n33), 
        .ZN(ref_1_maj_123_port_o) );
  OR2_X1 ref_1_maj_124_U19 ( .A1(ref_1_maj_124_n27), .A2(ref_1_maj_124_n26), 
        .ZN(ref_1_maj_124_n28) );
  NAND2_X1 ref_1_maj_124_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_124_n28), .ZN(
        ref_1_maj_124_n29) );
  NAND2_X1 ref_1_maj_124_U17 ( .A1(ref_1_maj_124_n26), .A2(ref_1_maj_124_n27), 
        .ZN(ref_1_maj_124_n30) );
  NAND2_X1 ref_1_maj_124_U16 ( .A1(ref_1_maj_124_n30), .A2(ref_1_maj_124_n29), 
        .ZN(ref_1_maj_124_n31) );
  NAND2_X1 ref_1_maj_124_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_124_n25), .ZN(
        ref_1_maj_124_n18) );
  NAND2_X1 ref_1_maj_124_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_124_n19) );
  NAND2_X1 ref_1_maj_124_U13 ( .A1(ref_1_maj_124_n19), .A2(ref_1_maj_124_n18), 
        .ZN(ref_1_maj_124_n22) );
  NAND2_X1 ref_1_maj_124_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_124_n24), .ZN(
        ref_1_maj_124_n20) );
  NAND2_X1 ref_1_maj_124_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_124_n21) );
  NAND2_X1 ref_1_maj_124_U10 ( .A1(ref_1_maj_124_n21), .A2(ref_1_maj_124_n20), 
        .ZN(ref_1_maj_124_n23) );
  XOR2_X1 ref_1_maj_124_U9 ( .A(ref_1_n7), .B(ref_1_maj_124_n24), .Z(
        ref_1_maj_124_n26) );
  XOR2_X1 ref_1_maj_124_U8 ( .A(ref_1_n16), .B(ref_1_maj_124_n25), .Z(
        ref_1_maj_124_n27) );
  XOR2_X1 ref_1_maj_124_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_124_n24)
         );
  XOR2_X1 ref_1_maj_124_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_124_n25) );
  OR2_X1 ref_1_maj_124_U5 ( .A1(ref_1_maj_124_n23), .A2(ref_1_maj_124_n22), 
        .ZN(ref_1_maj_124_n32) );
  NAND2_X1 ref_1_maj_124_U4 ( .A1(ref_1_maj_124_n22), .A2(ref_1_maj_124_n23), 
        .ZN(ref_1_maj_124_n34) );
  NAND2_X1 ref_1_maj_124_U3 ( .A1(ref_1_maj_124_n32), .A2(ref_1_maj_124_n31), 
        .ZN(ref_1_maj_124_n33) );
  NAND2_X1 ref_1_maj_124_U2 ( .A1(ref_1_maj_124_n34), .A2(ref_1_maj_124_n33), 
        .ZN(ref_1_maj_124_port_o) );
  OR2_X1 ref_1_maj_125_U19 ( .A1(ref_1_maj_125_n27), .A2(ref_1_maj_125_n26), 
        .ZN(ref_1_maj_125_n28) );
  NAND2_X1 ref_1_maj_125_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_125_n28), .ZN(
        ref_1_maj_125_n29) );
  NAND2_X1 ref_1_maj_125_U17 ( .A1(ref_1_maj_125_n26), .A2(ref_1_maj_125_n27), 
        .ZN(ref_1_maj_125_n30) );
  NAND2_X1 ref_1_maj_125_U16 ( .A1(ref_1_maj_125_n30), .A2(ref_1_maj_125_n29), 
        .ZN(ref_1_maj_125_n31) );
  NAND2_X1 ref_1_maj_125_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_125_n25), .ZN(
        ref_1_maj_125_n18) );
  NAND2_X1 ref_1_maj_125_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_125_n19) );
  NAND2_X1 ref_1_maj_125_U13 ( .A1(ref_1_maj_125_n19), .A2(ref_1_maj_125_n18), 
        .ZN(ref_1_maj_125_n22) );
  NAND2_X1 ref_1_maj_125_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_125_n24), .ZN(
        ref_1_maj_125_n20) );
  NAND2_X1 ref_1_maj_125_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_125_n21) );
  NAND2_X1 ref_1_maj_125_U10 ( .A1(ref_1_maj_125_n21), .A2(ref_1_maj_125_n20), 
        .ZN(ref_1_maj_125_n23) );
  XOR2_X1 ref_1_maj_125_U9 ( .A(ref_1_n7), .B(ref_1_maj_125_n24), .Z(
        ref_1_maj_125_n26) );
  XOR2_X1 ref_1_maj_125_U8 ( .A(ref_1_n16), .B(ref_1_maj_125_n25), .Z(
        ref_1_maj_125_n27) );
  XOR2_X1 ref_1_maj_125_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_125_n24)
         );
  XOR2_X1 ref_1_maj_125_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_125_n25) );
  OR2_X1 ref_1_maj_125_U5 ( .A1(ref_1_maj_125_n23), .A2(ref_1_maj_125_n22), 
        .ZN(ref_1_maj_125_n32) );
  NAND2_X1 ref_1_maj_125_U4 ( .A1(ref_1_maj_125_n22), .A2(ref_1_maj_125_n23), 
        .ZN(ref_1_maj_125_n34) );
  NAND2_X1 ref_1_maj_125_U3 ( .A1(ref_1_maj_125_n32), .A2(ref_1_maj_125_n31), 
        .ZN(ref_1_maj_125_n33) );
  NAND2_X1 ref_1_maj_125_U2 ( .A1(ref_1_maj_125_n34), .A2(ref_1_maj_125_n33), 
        .ZN(ref_1_maj_125_port_o) );
  OR2_X1 ref_1_maj_126_U19 ( .A1(ref_1_maj_126_n27), .A2(ref_1_maj_126_n26), 
        .ZN(ref_1_maj_126_n28) );
  NAND2_X1 ref_1_maj_126_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_126_n28), .ZN(
        ref_1_maj_126_n29) );
  NAND2_X1 ref_1_maj_126_U17 ( .A1(ref_1_maj_126_n26), .A2(ref_1_maj_126_n27), 
        .ZN(ref_1_maj_126_n30) );
  NAND2_X1 ref_1_maj_126_U16 ( .A1(ref_1_maj_126_n30), .A2(ref_1_maj_126_n29), 
        .ZN(ref_1_maj_126_n31) );
  NAND2_X1 ref_1_maj_126_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_126_n25), .ZN(
        ref_1_maj_126_n18) );
  NAND2_X1 ref_1_maj_126_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_126_n19) );
  NAND2_X1 ref_1_maj_126_U13 ( .A1(ref_1_maj_126_n19), .A2(ref_1_maj_126_n18), 
        .ZN(ref_1_maj_126_n22) );
  NAND2_X1 ref_1_maj_126_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_126_n24), .ZN(
        ref_1_maj_126_n20) );
  NAND2_X1 ref_1_maj_126_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_126_n21) );
  NAND2_X1 ref_1_maj_126_U10 ( .A1(ref_1_maj_126_n21), .A2(ref_1_maj_126_n20), 
        .ZN(ref_1_maj_126_n23) );
  XOR2_X1 ref_1_maj_126_U9 ( .A(ref_1_n7), .B(ref_1_maj_126_n24), .Z(
        ref_1_maj_126_n26) );
  XOR2_X1 ref_1_maj_126_U8 ( .A(ref_1_n16), .B(ref_1_maj_126_n25), .Z(
        ref_1_maj_126_n27) );
  XOR2_X1 ref_1_maj_126_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_126_n24)
         );
  XOR2_X1 ref_1_maj_126_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_126_n25) );
  OR2_X1 ref_1_maj_126_U5 ( .A1(ref_1_maj_126_n23), .A2(ref_1_maj_126_n22), 
        .ZN(ref_1_maj_126_n32) );
  NAND2_X1 ref_1_maj_126_U4 ( .A1(ref_1_maj_126_n22), .A2(ref_1_maj_126_n23), 
        .ZN(ref_1_maj_126_n34) );
  NAND2_X1 ref_1_maj_126_U3 ( .A1(ref_1_maj_126_n32), .A2(ref_1_maj_126_n31), 
        .ZN(ref_1_maj_126_n33) );
  NAND2_X1 ref_1_maj_126_U2 ( .A1(ref_1_maj_126_n34), .A2(ref_1_maj_126_n33), 
        .ZN(ref_1_maj_126_port_o) );
  OR2_X1 ref_1_maj_127_U19 ( .A1(ref_1_maj_127_n27), .A2(ref_1_maj_127_n26), 
        .ZN(ref_1_maj_127_n28) );
  NAND2_X1 ref_1_maj_127_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_127_n28), .ZN(
        ref_1_maj_127_n29) );
  NAND2_X1 ref_1_maj_127_U17 ( .A1(ref_1_maj_127_n26), .A2(ref_1_maj_127_n27), 
        .ZN(ref_1_maj_127_n30) );
  NAND2_X1 ref_1_maj_127_U16 ( .A1(ref_1_maj_127_n30), .A2(ref_1_maj_127_n29), 
        .ZN(ref_1_maj_127_n31) );
  NAND2_X1 ref_1_maj_127_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_127_n25), .ZN(
        ref_1_maj_127_n18) );
  NAND2_X1 ref_1_maj_127_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_127_n19) );
  NAND2_X1 ref_1_maj_127_U13 ( .A1(ref_1_maj_127_n19), .A2(ref_1_maj_127_n18), 
        .ZN(ref_1_maj_127_n22) );
  NAND2_X1 ref_1_maj_127_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_127_n24), .ZN(
        ref_1_maj_127_n20) );
  NAND2_X1 ref_1_maj_127_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_127_n21) );
  NAND2_X1 ref_1_maj_127_U10 ( .A1(ref_1_maj_127_n21), .A2(ref_1_maj_127_n20), 
        .ZN(ref_1_maj_127_n23) );
  XOR2_X1 ref_1_maj_127_U9 ( .A(ref_1_n7), .B(ref_1_maj_127_n24), .Z(
        ref_1_maj_127_n26) );
  XOR2_X1 ref_1_maj_127_U8 ( .A(ref_1_n16), .B(ref_1_maj_127_n25), .Z(
        ref_1_maj_127_n27) );
  XOR2_X1 ref_1_maj_127_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_127_n24)
         );
  XOR2_X1 ref_1_maj_127_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_127_n25) );
  OR2_X1 ref_1_maj_127_U5 ( .A1(ref_1_maj_127_n23), .A2(ref_1_maj_127_n22), 
        .ZN(ref_1_maj_127_n32) );
  NAND2_X1 ref_1_maj_127_U4 ( .A1(ref_1_maj_127_n22), .A2(ref_1_maj_127_n23), 
        .ZN(ref_1_maj_127_n34) );
  NAND2_X1 ref_1_maj_127_U3 ( .A1(ref_1_maj_127_n32), .A2(ref_1_maj_127_n31), 
        .ZN(ref_1_maj_127_n33) );
  NAND2_X1 ref_1_maj_127_U2 ( .A1(ref_1_maj_127_n34), .A2(ref_1_maj_127_n33), 
        .ZN(ref_1_maj_127_port_o) );
  OR2_X1 ref_1_maj_128_U19 ( .A1(ref_1_maj_128_n27), .A2(ref_1_maj_128_n26), 
        .ZN(ref_1_maj_128_n28) );
  NAND2_X1 ref_1_maj_128_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_128_n28), .ZN(
        ref_1_maj_128_n29) );
  NAND2_X1 ref_1_maj_128_U17 ( .A1(ref_1_maj_128_n26), .A2(ref_1_maj_128_n27), 
        .ZN(ref_1_maj_128_n30) );
  NAND2_X1 ref_1_maj_128_U16 ( .A1(ref_1_maj_128_n30), .A2(ref_1_maj_128_n29), 
        .ZN(ref_1_maj_128_n31) );
  NAND2_X1 ref_1_maj_128_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_128_n25), .ZN(
        ref_1_maj_128_n18) );
  NAND2_X1 ref_1_maj_128_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_128_n19) );
  NAND2_X1 ref_1_maj_128_U13 ( .A1(ref_1_maj_128_n19), .A2(ref_1_maj_128_n18), 
        .ZN(ref_1_maj_128_n22) );
  NAND2_X1 ref_1_maj_128_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_128_n24), .ZN(
        ref_1_maj_128_n20) );
  NAND2_X1 ref_1_maj_128_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_128_n21) );
  NAND2_X1 ref_1_maj_128_U10 ( .A1(ref_1_maj_128_n21), .A2(ref_1_maj_128_n20), 
        .ZN(ref_1_maj_128_n23) );
  XOR2_X1 ref_1_maj_128_U9 ( .A(ref_1_n64), .B(ref_1_maj_128_n24), .Z(
        ref_1_maj_128_n26) );
  XOR2_X1 ref_1_maj_128_U8 ( .A(ref_1_n73), .B(ref_1_maj_128_n25), .Z(
        ref_1_maj_128_n27) );
  XOR2_X1 ref_1_maj_128_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_128_n24) );
  XOR2_X1 ref_1_maj_128_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_128_n25) );
  OR2_X1 ref_1_maj_128_U5 ( .A1(ref_1_maj_128_n23), .A2(ref_1_maj_128_n22), 
        .ZN(ref_1_maj_128_n32) );
  NAND2_X1 ref_1_maj_128_U4 ( .A1(ref_1_maj_128_n22), .A2(ref_1_maj_128_n23), 
        .ZN(ref_1_maj_128_n34) );
  NAND2_X1 ref_1_maj_128_U3 ( .A1(ref_1_maj_128_n32), .A2(ref_1_maj_128_n31), 
        .ZN(ref_1_maj_128_n33) );
  NAND2_X1 ref_1_maj_128_U2 ( .A1(ref_1_maj_128_n34), .A2(ref_1_maj_128_n33), 
        .ZN(ref_1_maj_128_port_o) );
  OR2_X1 ref_1_maj_129_U19 ( .A1(ref_1_maj_129_n27), .A2(ref_1_maj_129_n26), 
        .ZN(ref_1_maj_129_n28) );
  NAND2_X1 ref_1_maj_129_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_129_n28), .ZN(
        ref_1_maj_129_n29) );
  NAND2_X1 ref_1_maj_129_U17 ( .A1(ref_1_maj_129_n26), .A2(ref_1_maj_129_n27), 
        .ZN(ref_1_maj_129_n30) );
  NAND2_X1 ref_1_maj_129_U16 ( .A1(ref_1_maj_129_n30), .A2(ref_1_maj_129_n29), 
        .ZN(ref_1_maj_129_n31) );
  NAND2_X1 ref_1_maj_129_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_129_n25), .ZN(
        ref_1_maj_129_n18) );
  NAND2_X1 ref_1_maj_129_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_129_n19) );
  NAND2_X1 ref_1_maj_129_U13 ( .A1(ref_1_maj_129_n19), .A2(ref_1_maj_129_n18), 
        .ZN(ref_1_maj_129_n22) );
  NAND2_X1 ref_1_maj_129_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_129_n24), .ZN(
        ref_1_maj_129_n20) );
  NAND2_X1 ref_1_maj_129_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_129_n21) );
  NAND2_X1 ref_1_maj_129_U10 ( .A1(ref_1_maj_129_n21), .A2(ref_1_maj_129_n20), 
        .ZN(ref_1_maj_129_n23) );
  XOR2_X1 ref_1_maj_129_U9 ( .A(ref_1_n64), .B(ref_1_maj_129_n24), .Z(
        ref_1_maj_129_n26) );
  XOR2_X1 ref_1_maj_129_U8 ( .A(ref_1_n73), .B(ref_1_maj_129_n25), .Z(
        ref_1_maj_129_n27) );
  XOR2_X1 ref_1_maj_129_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_129_n24) );
  XOR2_X1 ref_1_maj_129_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_129_n25) );
  OR2_X1 ref_1_maj_129_U5 ( .A1(ref_1_maj_129_n23), .A2(ref_1_maj_129_n22), 
        .ZN(ref_1_maj_129_n32) );
  NAND2_X1 ref_1_maj_129_U4 ( .A1(ref_1_maj_129_n22), .A2(ref_1_maj_129_n23), 
        .ZN(ref_1_maj_129_n34) );
  NAND2_X1 ref_1_maj_129_U3 ( .A1(ref_1_maj_129_n32), .A2(ref_1_maj_129_n31), 
        .ZN(ref_1_maj_129_n33) );
  NAND2_X1 ref_1_maj_129_U2 ( .A1(ref_1_maj_129_n34), .A2(ref_1_maj_129_n33), 
        .ZN(ref_1_maj_129_port_o) );
  OR2_X1 ref_1_maj_130_U19 ( .A1(ref_1_maj_130_n27), .A2(ref_1_maj_130_n26), 
        .ZN(ref_1_maj_130_n28) );
  NAND2_X1 ref_1_maj_130_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_130_n28), .ZN(
        ref_1_maj_130_n29) );
  NAND2_X1 ref_1_maj_130_U17 ( .A1(ref_1_maj_130_n26), .A2(ref_1_maj_130_n27), 
        .ZN(ref_1_maj_130_n30) );
  NAND2_X1 ref_1_maj_130_U16 ( .A1(ref_1_maj_130_n30), .A2(ref_1_maj_130_n29), 
        .ZN(ref_1_maj_130_n31) );
  NAND2_X1 ref_1_maj_130_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_130_n25), .ZN(
        ref_1_maj_130_n18) );
  NAND2_X1 ref_1_maj_130_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_130_n19) );
  NAND2_X1 ref_1_maj_130_U13 ( .A1(ref_1_maj_130_n19), .A2(ref_1_maj_130_n18), 
        .ZN(ref_1_maj_130_n22) );
  NAND2_X1 ref_1_maj_130_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_130_n24), .ZN(
        ref_1_maj_130_n20) );
  NAND2_X1 ref_1_maj_130_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_130_n21) );
  NAND2_X1 ref_1_maj_130_U10 ( .A1(ref_1_maj_130_n21), .A2(ref_1_maj_130_n20), 
        .ZN(ref_1_maj_130_n23) );
  XOR2_X1 ref_1_maj_130_U9 ( .A(ref_1_n64), .B(ref_1_maj_130_n24), .Z(
        ref_1_maj_130_n26) );
  XOR2_X1 ref_1_maj_130_U8 ( .A(ref_1_n73), .B(ref_1_maj_130_n25), .Z(
        ref_1_maj_130_n27) );
  XOR2_X1 ref_1_maj_130_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_130_n24) );
  XOR2_X1 ref_1_maj_130_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_130_n25) );
  OR2_X1 ref_1_maj_130_U5 ( .A1(ref_1_maj_130_n23), .A2(ref_1_maj_130_n22), 
        .ZN(ref_1_maj_130_n32) );
  NAND2_X1 ref_1_maj_130_U4 ( .A1(ref_1_maj_130_n22), .A2(ref_1_maj_130_n23), 
        .ZN(ref_1_maj_130_n34) );
  NAND2_X1 ref_1_maj_130_U3 ( .A1(ref_1_maj_130_n32), .A2(ref_1_maj_130_n31), 
        .ZN(ref_1_maj_130_n33) );
  NAND2_X1 ref_1_maj_130_U2 ( .A1(ref_1_maj_130_n34), .A2(ref_1_maj_130_n33), 
        .ZN(ref_1_maj_130_port_o) );
  OR2_X1 ref_1_maj_131_U19 ( .A1(ref_1_maj_131_n27), .A2(ref_1_maj_131_n26), 
        .ZN(ref_1_maj_131_n28) );
  NAND2_X1 ref_1_maj_131_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_131_n28), .ZN(
        ref_1_maj_131_n29) );
  NAND2_X1 ref_1_maj_131_U17 ( .A1(ref_1_maj_131_n26), .A2(ref_1_maj_131_n27), 
        .ZN(ref_1_maj_131_n30) );
  NAND2_X1 ref_1_maj_131_U16 ( .A1(ref_1_maj_131_n30), .A2(ref_1_maj_131_n29), 
        .ZN(ref_1_maj_131_n31) );
  NAND2_X1 ref_1_maj_131_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_131_n25), .ZN(
        ref_1_maj_131_n18) );
  NAND2_X1 ref_1_maj_131_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_131_n19) );
  NAND2_X1 ref_1_maj_131_U13 ( .A1(ref_1_maj_131_n19), .A2(ref_1_maj_131_n18), 
        .ZN(ref_1_maj_131_n22) );
  NAND2_X1 ref_1_maj_131_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_131_n24), .ZN(
        ref_1_maj_131_n20) );
  NAND2_X1 ref_1_maj_131_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_131_n21) );
  NAND2_X1 ref_1_maj_131_U10 ( .A1(ref_1_maj_131_n21), .A2(ref_1_maj_131_n20), 
        .ZN(ref_1_maj_131_n23) );
  XOR2_X1 ref_1_maj_131_U9 ( .A(ref_1_n64), .B(ref_1_maj_131_n24), .Z(
        ref_1_maj_131_n26) );
  XOR2_X1 ref_1_maj_131_U8 ( .A(ref_1_n73), .B(ref_1_maj_131_n25), .Z(
        ref_1_maj_131_n27) );
  XOR2_X1 ref_1_maj_131_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_131_n24) );
  XOR2_X1 ref_1_maj_131_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_131_n25) );
  OR2_X1 ref_1_maj_131_U5 ( .A1(ref_1_maj_131_n23), .A2(ref_1_maj_131_n22), 
        .ZN(ref_1_maj_131_n32) );
  NAND2_X1 ref_1_maj_131_U4 ( .A1(ref_1_maj_131_n22), .A2(ref_1_maj_131_n23), 
        .ZN(ref_1_maj_131_n34) );
  NAND2_X1 ref_1_maj_131_U3 ( .A1(ref_1_maj_131_n32), .A2(ref_1_maj_131_n31), 
        .ZN(ref_1_maj_131_n33) );
  NAND2_X1 ref_1_maj_131_U2 ( .A1(ref_1_maj_131_n34), .A2(ref_1_maj_131_n33), 
        .ZN(ref_1_maj_131_port_o) );
  OR2_X1 ref_1_maj_132_U19 ( .A1(ref_1_maj_132_n27), .A2(ref_1_maj_132_n26), 
        .ZN(ref_1_maj_132_n28) );
  NAND2_X1 ref_1_maj_132_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_132_n28), .ZN(
        ref_1_maj_132_n29) );
  NAND2_X1 ref_1_maj_132_U17 ( .A1(ref_1_maj_132_n26), .A2(ref_1_maj_132_n27), 
        .ZN(ref_1_maj_132_n30) );
  NAND2_X1 ref_1_maj_132_U16 ( .A1(ref_1_maj_132_n30), .A2(ref_1_maj_132_n29), 
        .ZN(ref_1_maj_132_n31) );
  NAND2_X1 ref_1_maj_132_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_132_n25), .ZN(
        ref_1_maj_132_n18) );
  NAND2_X1 ref_1_maj_132_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_132_n19) );
  NAND2_X1 ref_1_maj_132_U13 ( .A1(ref_1_maj_132_n19), .A2(ref_1_maj_132_n18), 
        .ZN(ref_1_maj_132_n22) );
  NAND2_X1 ref_1_maj_132_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_132_n24), .ZN(
        ref_1_maj_132_n20) );
  NAND2_X1 ref_1_maj_132_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_132_n21) );
  NAND2_X1 ref_1_maj_132_U10 ( .A1(ref_1_maj_132_n21), .A2(ref_1_maj_132_n20), 
        .ZN(ref_1_maj_132_n23) );
  XOR2_X1 ref_1_maj_132_U9 ( .A(ref_1_n45), .B(ref_1_maj_132_n24), .Z(
        ref_1_maj_132_n26) );
  XOR2_X1 ref_1_maj_132_U8 ( .A(ref_1_n54), .B(ref_1_maj_132_n25), .Z(
        ref_1_maj_132_n27) );
  XOR2_X1 ref_1_maj_132_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_132_n24) );
  XOR2_X1 ref_1_maj_132_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_132_n25) );
  OR2_X1 ref_1_maj_132_U5 ( .A1(ref_1_maj_132_n23), .A2(ref_1_maj_132_n22), 
        .ZN(ref_1_maj_132_n32) );
  NAND2_X1 ref_1_maj_132_U4 ( .A1(ref_1_maj_132_n22), .A2(ref_1_maj_132_n23), 
        .ZN(ref_1_maj_132_n34) );
  NAND2_X1 ref_1_maj_132_U3 ( .A1(ref_1_maj_132_n32), .A2(ref_1_maj_132_n31), 
        .ZN(ref_1_maj_132_n33) );
  NAND2_X1 ref_1_maj_132_U2 ( .A1(ref_1_maj_132_n34), .A2(ref_1_maj_132_n33), 
        .ZN(ref_1_maj_132_port_o) );
  OR2_X1 ref_1_maj_133_U19 ( .A1(ref_1_maj_133_n27), .A2(ref_1_maj_133_n26), 
        .ZN(ref_1_maj_133_n28) );
  NAND2_X1 ref_1_maj_133_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_133_n28), .ZN(
        ref_1_maj_133_n29) );
  NAND2_X1 ref_1_maj_133_U17 ( .A1(ref_1_maj_133_n26), .A2(ref_1_maj_133_n27), 
        .ZN(ref_1_maj_133_n30) );
  NAND2_X1 ref_1_maj_133_U16 ( .A1(ref_1_maj_133_n30), .A2(ref_1_maj_133_n29), 
        .ZN(ref_1_maj_133_n31) );
  NAND2_X1 ref_1_maj_133_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_133_n25), .ZN(
        ref_1_maj_133_n18) );
  NAND2_X1 ref_1_maj_133_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_133_n19) );
  NAND2_X1 ref_1_maj_133_U13 ( .A1(ref_1_maj_133_n19), .A2(ref_1_maj_133_n18), 
        .ZN(ref_1_maj_133_n22) );
  NAND2_X1 ref_1_maj_133_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_133_n24), .ZN(
        ref_1_maj_133_n20) );
  NAND2_X1 ref_1_maj_133_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_133_n21) );
  NAND2_X1 ref_1_maj_133_U10 ( .A1(ref_1_maj_133_n21), .A2(ref_1_maj_133_n20), 
        .ZN(ref_1_maj_133_n23) );
  XOR2_X1 ref_1_maj_133_U9 ( .A(ref_1_n45), .B(ref_1_maj_133_n24), .Z(
        ref_1_maj_133_n26) );
  XOR2_X1 ref_1_maj_133_U8 ( .A(ref_1_n54), .B(ref_1_maj_133_n25), .Z(
        ref_1_maj_133_n27) );
  XOR2_X1 ref_1_maj_133_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_133_n24) );
  XOR2_X1 ref_1_maj_133_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_133_n25) );
  OR2_X1 ref_1_maj_133_U5 ( .A1(ref_1_maj_133_n23), .A2(ref_1_maj_133_n22), 
        .ZN(ref_1_maj_133_n32) );
  NAND2_X1 ref_1_maj_133_U4 ( .A1(ref_1_maj_133_n22), .A2(ref_1_maj_133_n23), 
        .ZN(ref_1_maj_133_n34) );
  NAND2_X1 ref_1_maj_133_U3 ( .A1(ref_1_maj_133_n32), .A2(ref_1_maj_133_n31), 
        .ZN(ref_1_maj_133_n33) );
  NAND2_X1 ref_1_maj_133_U2 ( .A1(ref_1_maj_133_n34), .A2(ref_1_maj_133_n33), 
        .ZN(ref_1_maj_133_port_o) );
  OR2_X1 ref_1_maj_134_U19 ( .A1(ref_1_maj_134_n27), .A2(ref_1_maj_134_n26), 
        .ZN(ref_1_maj_134_n28) );
  NAND2_X1 ref_1_maj_134_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_134_n28), .ZN(
        ref_1_maj_134_n29) );
  NAND2_X1 ref_1_maj_134_U17 ( .A1(ref_1_maj_134_n26), .A2(ref_1_maj_134_n27), 
        .ZN(ref_1_maj_134_n30) );
  NAND2_X1 ref_1_maj_134_U16 ( .A1(ref_1_maj_134_n30), .A2(ref_1_maj_134_n29), 
        .ZN(ref_1_maj_134_n31) );
  NAND2_X1 ref_1_maj_134_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_134_n25), .ZN(
        ref_1_maj_134_n18) );
  NAND2_X1 ref_1_maj_134_U14 ( .A1(ref_1_n48), .A2(ref_1_n51), .ZN(
        ref_1_maj_134_n19) );
  NAND2_X1 ref_1_maj_134_U13 ( .A1(ref_1_maj_134_n19), .A2(ref_1_maj_134_n18), 
        .ZN(ref_1_maj_134_n22) );
  NAND2_X1 ref_1_maj_134_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_134_n24), .ZN(
        ref_1_maj_134_n20) );
  NAND2_X1 ref_1_maj_134_U11 ( .A1(ref_1_n39), .A2(ref_1_n42), .ZN(
        ref_1_maj_134_n21) );
  NAND2_X1 ref_1_maj_134_U10 ( .A1(ref_1_maj_134_n21), .A2(ref_1_maj_134_n20), 
        .ZN(ref_1_maj_134_n23) );
  XOR2_X1 ref_1_maj_134_U9 ( .A(ref_1_n45), .B(ref_1_maj_134_n24), .Z(
        ref_1_maj_134_n26) );
  XOR2_X1 ref_1_maj_134_U8 ( .A(ref_1_n54), .B(ref_1_maj_134_n25), .Z(
        ref_1_maj_134_n27) );
  XOR2_X1 ref_1_maj_134_U7 ( .A(ref_1_n39), .B(ref_1_n42), .Z(
        ref_1_maj_134_n24) );
  XOR2_X1 ref_1_maj_134_U6 ( .A(ref_1_n48), .B(ref_1_n51), .Z(
        ref_1_maj_134_n25) );
  OR2_X1 ref_1_maj_134_U5 ( .A1(ref_1_maj_134_n23), .A2(ref_1_maj_134_n22), 
        .ZN(ref_1_maj_134_n32) );
  NAND2_X1 ref_1_maj_134_U4 ( .A1(ref_1_maj_134_n22), .A2(ref_1_maj_134_n23), 
        .ZN(ref_1_maj_134_n34) );
  NAND2_X1 ref_1_maj_134_U3 ( .A1(ref_1_maj_134_n32), .A2(ref_1_maj_134_n31), 
        .ZN(ref_1_maj_134_n33) );
  NAND2_X1 ref_1_maj_134_U2 ( .A1(ref_1_maj_134_n34), .A2(ref_1_maj_134_n33), 
        .ZN(ref_1_maj_134_port_o) );
  OR2_X1 ref_1_maj_135_U19 ( .A1(ref_1_maj_135_n27), .A2(ref_1_maj_135_n26), 
        .ZN(ref_1_maj_135_n28) );
  NAND2_X1 ref_1_maj_135_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_135_n28), .ZN(
        ref_1_maj_135_n29) );
  NAND2_X1 ref_1_maj_135_U17 ( .A1(ref_1_maj_135_n26), .A2(ref_1_maj_135_n27), 
        .ZN(ref_1_maj_135_n30) );
  NAND2_X1 ref_1_maj_135_U16 ( .A1(ref_1_maj_135_n30), .A2(ref_1_maj_135_n29), 
        .ZN(ref_1_maj_135_n31) );
  NAND2_X1 ref_1_maj_135_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_135_n25), .ZN(
        ref_1_maj_135_n18) );
  NAND2_X1 ref_1_maj_135_U14 ( .A1(ref_1_n48), .A2(ref_1_n52), .ZN(
        ref_1_maj_135_n19) );
  NAND2_X1 ref_1_maj_135_U13 ( .A1(ref_1_maj_135_n19), .A2(ref_1_maj_135_n18), 
        .ZN(ref_1_maj_135_n22) );
  NAND2_X1 ref_1_maj_135_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_135_n24), .ZN(
        ref_1_maj_135_n20) );
  NAND2_X1 ref_1_maj_135_U11 ( .A1(ref_1_n39), .A2(ref_1_n43), .ZN(
        ref_1_maj_135_n21) );
  NAND2_X1 ref_1_maj_135_U10 ( .A1(ref_1_maj_135_n21), .A2(ref_1_maj_135_n20), 
        .ZN(ref_1_maj_135_n23) );
  XOR2_X1 ref_1_maj_135_U9 ( .A(ref_1_n46), .B(ref_1_maj_135_n24), .Z(
        ref_1_maj_135_n26) );
  XOR2_X1 ref_1_maj_135_U8 ( .A(ref_1_n54), .B(ref_1_maj_135_n25), .Z(
        ref_1_maj_135_n27) );
  XOR2_X1 ref_1_maj_135_U7 ( .A(ref_1_n39), .B(ref_1_n43), .Z(
        ref_1_maj_135_n24) );
  XOR2_X1 ref_1_maj_135_U6 ( .A(ref_1_n48), .B(ref_1_n52), .Z(
        ref_1_maj_135_n25) );
  OR2_X1 ref_1_maj_135_U5 ( .A1(ref_1_maj_135_n23), .A2(ref_1_maj_135_n22), 
        .ZN(ref_1_maj_135_n32) );
  NAND2_X1 ref_1_maj_135_U4 ( .A1(ref_1_maj_135_n22), .A2(ref_1_maj_135_n23), 
        .ZN(ref_1_maj_135_n34) );
  NAND2_X1 ref_1_maj_135_U3 ( .A1(ref_1_maj_135_n32), .A2(ref_1_maj_135_n31), 
        .ZN(ref_1_maj_135_n33) );
  NAND2_X1 ref_1_maj_135_U2 ( .A1(ref_1_maj_135_n34), .A2(ref_1_maj_135_n33), 
        .ZN(ref_1_maj_135_port_o) );
  OR2_X1 ref_1_maj_136_U19 ( .A1(ref_1_maj_136_n27), .A2(ref_1_maj_136_n26), 
        .ZN(ref_1_maj_136_n28) );
  NAND2_X1 ref_1_maj_136_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_136_n28), .ZN(
        ref_1_maj_136_n29) );
  NAND2_X1 ref_1_maj_136_U17 ( .A1(ref_1_maj_136_n26), .A2(ref_1_maj_136_n27), 
        .ZN(ref_1_maj_136_n30) );
  NAND2_X1 ref_1_maj_136_U16 ( .A1(ref_1_maj_136_n30), .A2(ref_1_maj_136_n29), 
        .ZN(ref_1_maj_136_n31) );
  NAND2_X1 ref_1_maj_136_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_136_n25), .ZN(
        ref_1_maj_136_n18) );
  NAND2_X1 ref_1_maj_136_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_136_n19) );
  NAND2_X1 ref_1_maj_136_U13 ( .A1(ref_1_maj_136_n19), .A2(ref_1_maj_136_n18), 
        .ZN(ref_1_maj_136_n22) );
  NAND2_X1 ref_1_maj_136_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_136_n24), .ZN(
        ref_1_maj_136_n20) );
  NAND2_X1 ref_1_maj_136_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_136_n21) );
  NAND2_X1 ref_1_maj_136_U10 ( .A1(ref_1_maj_136_n21), .A2(ref_1_maj_136_n20), 
        .ZN(ref_1_maj_136_n23) );
  XOR2_X1 ref_1_maj_136_U9 ( .A(ref_1_n26), .B(ref_1_maj_136_n24), .Z(
        ref_1_maj_136_n26) );
  XOR2_X1 ref_1_maj_136_U8 ( .A(ref_1_n35), .B(ref_1_maj_136_n25), .Z(
        ref_1_maj_136_n27) );
  XOR2_X1 ref_1_maj_136_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_136_n24) );
  XOR2_X1 ref_1_maj_136_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_136_n25) );
  OR2_X1 ref_1_maj_136_U5 ( .A1(ref_1_maj_136_n23), .A2(ref_1_maj_136_n22), 
        .ZN(ref_1_maj_136_n32) );
  NAND2_X1 ref_1_maj_136_U4 ( .A1(ref_1_maj_136_n22), .A2(ref_1_maj_136_n23), 
        .ZN(ref_1_maj_136_n34) );
  NAND2_X1 ref_1_maj_136_U3 ( .A1(ref_1_maj_136_n32), .A2(ref_1_maj_136_n31), 
        .ZN(ref_1_maj_136_n33) );
  NAND2_X1 ref_1_maj_136_U2 ( .A1(ref_1_maj_136_n34), .A2(ref_1_maj_136_n33), 
        .ZN(ref_1_maj_136_port_o) );
  OR2_X1 ref_1_maj_137_U19 ( .A1(ref_1_maj_137_n27), .A2(ref_1_maj_137_n26), 
        .ZN(ref_1_maj_137_n28) );
  NAND2_X1 ref_1_maj_137_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_137_n28), .ZN(
        ref_1_maj_137_n29) );
  NAND2_X1 ref_1_maj_137_U17 ( .A1(ref_1_maj_137_n26), .A2(ref_1_maj_137_n27), 
        .ZN(ref_1_maj_137_n30) );
  NAND2_X1 ref_1_maj_137_U16 ( .A1(ref_1_maj_137_n30), .A2(ref_1_maj_137_n29), 
        .ZN(ref_1_maj_137_n31) );
  NAND2_X1 ref_1_maj_137_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_137_n25), .ZN(
        ref_1_maj_137_n18) );
  NAND2_X1 ref_1_maj_137_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_137_n19) );
  NAND2_X1 ref_1_maj_137_U13 ( .A1(ref_1_maj_137_n19), .A2(ref_1_maj_137_n18), 
        .ZN(ref_1_maj_137_n22) );
  NAND2_X1 ref_1_maj_137_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_137_n24), .ZN(
        ref_1_maj_137_n20) );
  NAND2_X1 ref_1_maj_137_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_137_n21) );
  NAND2_X1 ref_1_maj_137_U10 ( .A1(ref_1_maj_137_n21), .A2(ref_1_maj_137_n20), 
        .ZN(ref_1_maj_137_n23) );
  XOR2_X1 ref_1_maj_137_U9 ( .A(ref_1_n26), .B(ref_1_maj_137_n24), .Z(
        ref_1_maj_137_n26) );
  XOR2_X1 ref_1_maj_137_U8 ( .A(ref_1_n35), .B(ref_1_maj_137_n25), .Z(
        ref_1_maj_137_n27) );
  XOR2_X1 ref_1_maj_137_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_137_n24) );
  XOR2_X1 ref_1_maj_137_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_137_n25) );
  OR2_X1 ref_1_maj_137_U5 ( .A1(ref_1_maj_137_n23), .A2(ref_1_maj_137_n22), 
        .ZN(ref_1_maj_137_n32) );
  NAND2_X1 ref_1_maj_137_U4 ( .A1(ref_1_maj_137_n22), .A2(ref_1_maj_137_n23), 
        .ZN(ref_1_maj_137_n34) );
  NAND2_X1 ref_1_maj_137_U3 ( .A1(ref_1_maj_137_n32), .A2(ref_1_maj_137_n31), 
        .ZN(ref_1_maj_137_n33) );
  NAND2_X1 ref_1_maj_137_U2 ( .A1(ref_1_maj_137_n34), .A2(ref_1_maj_137_n33), 
        .ZN(ref_1_maj_137_port_o) );
  OR2_X1 ref_1_maj_138_U19 ( .A1(ref_1_maj_138_n27), .A2(ref_1_maj_138_n26), 
        .ZN(ref_1_maj_138_n28) );
  NAND2_X1 ref_1_maj_138_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_138_n28), .ZN(
        ref_1_maj_138_n29) );
  NAND2_X1 ref_1_maj_138_U17 ( .A1(ref_1_maj_138_n26), .A2(ref_1_maj_138_n27), 
        .ZN(ref_1_maj_138_n30) );
  NAND2_X1 ref_1_maj_138_U16 ( .A1(ref_1_maj_138_n30), .A2(ref_1_maj_138_n29), 
        .ZN(ref_1_maj_138_n31) );
  NAND2_X1 ref_1_maj_138_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_138_n25), .ZN(
        ref_1_maj_138_n18) );
  NAND2_X1 ref_1_maj_138_U14 ( .A1(ref_1_n29), .A2(ref_1_n32), .ZN(
        ref_1_maj_138_n19) );
  NAND2_X1 ref_1_maj_138_U13 ( .A1(ref_1_maj_138_n19), .A2(ref_1_maj_138_n18), 
        .ZN(ref_1_maj_138_n22) );
  NAND2_X1 ref_1_maj_138_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_138_n24), .ZN(
        ref_1_maj_138_n20) );
  NAND2_X1 ref_1_maj_138_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_138_n21) );
  NAND2_X1 ref_1_maj_138_U10 ( .A1(ref_1_maj_138_n21), .A2(ref_1_maj_138_n20), 
        .ZN(ref_1_maj_138_n23) );
  XOR2_X1 ref_1_maj_138_U9 ( .A(ref_1_n26), .B(ref_1_maj_138_n24), .Z(
        ref_1_maj_138_n26) );
  XOR2_X1 ref_1_maj_138_U8 ( .A(ref_1_n35), .B(ref_1_maj_138_n25), .Z(
        ref_1_maj_138_n27) );
  XOR2_X1 ref_1_maj_138_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_138_n24) );
  XOR2_X1 ref_1_maj_138_U6 ( .A(ref_1_n29), .B(ref_1_n32), .Z(
        ref_1_maj_138_n25) );
  OR2_X1 ref_1_maj_138_U5 ( .A1(ref_1_maj_138_n23), .A2(ref_1_maj_138_n22), 
        .ZN(ref_1_maj_138_n32) );
  NAND2_X1 ref_1_maj_138_U4 ( .A1(ref_1_maj_138_n22), .A2(ref_1_maj_138_n23), 
        .ZN(ref_1_maj_138_n34) );
  NAND2_X1 ref_1_maj_138_U3 ( .A1(ref_1_maj_138_n32), .A2(ref_1_maj_138_n31), 
        .ZN(ref_1_maj_138_n33) );
  NAND2_X1 ref_1_maj_138_U2 ( .A1(ref_1_maj_138_n34), .A2(ref_1_maj_138_n33), 
        .ZN(ref_1_maj_138_port_o) );
  OR2_X1 ref_1_maj_139_U19 ( .A1(ref_1_maj_139_n27), .A2(ref_1_maj_139_n26), 
        .ZN(ref_1_maj_139_n28) );
  NAND2_X1 ref_1_maj_139_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_139_n28), .ZN(
        ref_1_maj_139_n29) );
  NAND2_X1 ref_1_maj_139_U17 ( .A1(ref_1_maj_139_n26), .A2(ref_1_maj_139_n27), 
        .ZN(ref_1_maj_139_n30) );
  NAND2_X1 ref_1_maj_139_U16 ( .A1(ref_1_maj_139_n30), .A2(ref_1_maj_139_n29), 
        .ZN(ref_1_maj_139_n31) );
  NAND2_X1 ref_1_maj_139_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_139_n25), .ZN(
        ref_1_maj_139_n18) );
  NAND2_X1 ref_1_maj_139_U14 ( .A1(ref_1_n30), .A2(ref_1_n32), .ZN(
        ref_1_maj_139_n19) );
  NAND2_X1 ref_1_maj_139_U13 ( .A1(ref_1_maj_139_n19), .A2(ref_1_maj_139_n18), 
        .ZN(ref_1_maj_139_n22) );
  NAND2_X1 ref_1_maj_139_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_139_n24), .ZN(
        ref_1_maj_139_n20) );
  NAND2_X1 ref_1_maj_139_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_139_n21) );
  NAND2_X1 ref_1_maj_139_U10 ( .A1(ref_1_maj_139_n21), .A2(ref_1_maj_139_n20), 
        .ZN(ref_1_maj_139_n23) );
  XOR2_X1 ref_1_maj_139_U9 ( .A(ref_1_n27), .B(ref_1_maj_139_n24), .Z(
        ref_1_maj_139_n26) );
  XOR2_X1 ref_1_maj_139_U8 ( .A(ref_1_n36), .B(ref_1_maj_139_n25), .Z(
        ref_1_maj_139_n27) );
  XOR2_X1 ref_1_maj_139_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_139_n24) );
  XOR2_X1 ref_1_maj_139_U6 ( .A(ref_1_n30), .B(ref_1_n32), .Z(
        ref_1_maj_139_n25) );
  OR2_X1 ref_1_maj_139_U5 ( .A1(ref_1_maj_139_n23), .A2(ref_1_maj_139_n22), 
        .ZN(ref_1_maj_139_n32) );
  NAND2_X1 ref_1_maj_139_U4 ( .A1(ref_1_maj_139_n22), .A2(ref_1_maj_139_n23), 
        .ZN(ref_1_maj_139_n34) );
  NAND2_X1 ref_1_maj_139_U3 ( .A1(ref_1_maj_139_n32), .A2(ref_1_maj_139_n31), 
        .ZN(ref_1_maj_139_n33) );
  NAND2_X1 ref_1_maj_139_U2 ( .A1(ref_1_maj_139_n34), .A2(ref_1_maj_139_n33), 
        .ZN(ref_1_maj_139_port_o) );
  OR2_X1 ref_1_maj_140_U19 ( .A1(ref_1_maj_140_n27), .A2(ref_1_maj_140_n26), 
        .ZN(ref_1_maj_140_n28) );
  NAND2_X1 ref_1_maj_140_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_140_n28), .ZN(
        ref_1_maj_140_n29) );
  NAND2_X1 ref_1_maj_140_U17 ( .A1(ref_1_maj_140_n26), .A2(ref_1_maj_140_n27), 
        .ZN(ref_1_maj_140_n30) );
  NAND2_X1 ref_1_maj_140_U16 ( .A1(ref_1_maj_140_n30), .A2(ref_1_maj_140_n29), 
        .ZN(ref_1_maj_140_n31) );
  NAND2_X1 ref_1_maj_140_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_140_n25), .ZN(
        ref_1_maj_140_n18) );
  NAND2_X1 ref_1_maj_140_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_140_n19) );
  NAND2_X1 ref_1_maj_140_U13 ( .A1(ref_1_maj_140_n19), .A2(ref_1_maj_140_n18), 
        .ZN(ref_1_maj_140_n22) );
  NAND2_X1 ref_1_maj_140_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_140_n24), .ZN(
        ref_1_maj_140_n20) );
  NAND2_X1 ref_1_maj_140_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_140_n21) );
  NAND2_X1 ref_1_maj_140_U10 ( .A1(ref_1_maj_140_n21), .A2(ref_1_maj_140_n20), 
        .ZN(ref_1_maj_140_n23) );
  XOR2_X1 ref_1_maj_140_U9 ( .A(ref_1_n7), .B(ref_1_maj_140_n24), .Z(
        ref_1_maj_140_n26) );
  XOR2_X1 ref_1_maj_140_U8 ( .A(ref_1_n16), .B(ref_1_maj_140_n25), .Z(
        ref_1_maj_140_n27) );
  XOR2_X1 ref_1_maj_140_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_140_n24)
         );
  XOR2_X1 ref_1_maj_140_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_140_n25) );
  OR2_X1 ref_1_maj_140_U5 ( .A1(ref_1_maj_140_n23), .A2(ref_1_maj_140_n22), 
        .ZN(ref_1_maj_140_n32) );
  NAND2_X1 ref_1_maj_140_U4 ( .A1(ref_1_maj_140_n22), .A2(ref_1_maj_140_n23), 
        .ZN(ref_1_maj_140_n34) );
  NAND2_X1 ref_1_maj_140_U3 ( .A1(ref_1_maj_140_n32), .A2(ref_1_maj_140_n31), 
        .ZN(ref_1_maj_140_n33) );
  NAND2_X1 ref_1_maj_140_U2 ( .A1(ref_1_maj_140_n34), .A2(ref_1_maj_140_n33), 
        .ZN(ref_1_maj_140_port_o) );
  OR2_X1 ref_1_maj_141_U19 ( .A1(ref_1_maj_141_n27), .A2(ref_1_maj_141_n26), 
        .ZN(ref_1_maj_141_n28) );
  NAND2_X1 ref_1_maj_141_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_141_n28), .ZN(
        ref_1_maj_141_n29) );
  NAND2_X1 ref_1_maj_141_U17 ( .A1(ref_1_maj_141_n26), .A2(ref_1_maj_141_n27), 
        .ZN(ref_1_maj_141_n30) );
  NAND2_X1 ref_1_maj_141_U16 ( .A1(ref_1_maj_141_n30), .A2(ref_1_maj_141_n29), 
        .ZN(ref_1_maj_141_n31) );
  NAND2_X1 ref_1_maj_141_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_141_n25), .ZN(
        ref_1_maj_141_n18) );
  NAND2_X1 ref_1_maj_141_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_141_n19) );
  NAND2_X1 ref_1_maj_141_U13 ( .A1(ref_1_maj_141_n19), .A2(ref_1_maj_141_n18), 
        .ZN(ref_1_maj_141_n22) );
  NAND2_X1 ref_1_maj_141_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_141_n24), .ZN(
        ref_1_maj_141_n20) );
  NAND2_X1 ref_1_maj_141_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_141_n21) );
  NAND2_X1 ref_1_maj_141_U10 ( .A1(ref_1_maj_141_n21), .A2(ref_1_maj_141_n20), 
        .ZN(ref_1_maj_141_n23) );
  XOR2_X1 ref_1_maj_141_U9 ( .A(ref_1_n7), .B(ref_1_maj_141_n24), .Z(
        ref_1_maj_141_n26) );
  XOR2_X1 ref_1_maj_141_U8 ( .A(ref_1_n16), .B(ref_1_maj_141_n25), .Z(
        ref_1_maj_141_n27) );
  XOR2_X1 ref_1_maj_141_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_141_n24)
         );
  XOR2_X1 ref_1_maj_141_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_141_n25) );
  OR2_X1 ref_1_maj_141_U5 ( .A1(ref_1_maj_141_n23), .A2(ref_1_maj_141_n22), 
        .ZN(ref_1_maj_141_n32) );
  NAND2_X1 ref_1_maj_141_U4 ( .A1(ref_1_maj_141_n22), .A2(ref_1_maj_141_n23), 
        .ZN(ref_1_maj_141_n34) );
  NAND2_X1 ref_1_maj_141_U3 ( .A1(ref_1_maj_141_n32), .A2(ref_1_maj_141_n31), 
        .ZN(ref_1_maj_141_n33) );
  NAND2_X1 ref_1_maj_141_U2 ( .A1(ref_1_maj_141_n34), .A2(ref_1_maj_141_n33), 
        .ZN(ref_1_maj_141_port_o) );
  OR2_X1 ref_1_maj_142_U19 ( .A1(ref_1_maj_142_n27), .A2(ref_1_maj_142_n26), 
        .ZN(ref_1_maj_142_n28) );
  NAND2_X1 ref_1_maj_142_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_142_n28), .ZN(
        ref_1_maj_142_n29) );
  NAND2_X1 ref_1_maj_142_U17 ( .A1(ref_1_maj_142_n26), .A2(ref_1_maj_142_n27), 
        .ZN(ref_1_maj_142_n30) );
  NAND2_X1 ref_1_maj_142_U16 ( .A1(ref_1_maj_142_n30), .A2(ref_1_maj_142_n29), 
        .ZN(ref_1_maj_142_n31) );
  NAND2_X1 ref_1_maj_142_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_142_n25), .ZN(
        ref_1_maj_142_n18) );
  NAND2_X1 ref_1_maj_142_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_142_n19) );
  NAND2_X1 ref_1_maj_142_U13 ( .A1(ref_1_maj_142_n19), .A2(ref_1_maj_142_n18), 
        .ZN(ref_1_maj_142_n22) );
  NAND2_X1 ref_1_maj_142_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_142_n24), .ZN(
        ref_1_maj_142_n20) );
  NAND2_X1 ref_1_maj_142_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_142_n21) );
  NAND2_X1 ref_1_maj_142_U10 ( .A1(ref_1_maj_142_n21), .A2(ref_1_maj_142_n20), 
        .ZN(ref_1_maj_142_n23) );
  XOR2_X1 ref_1_maj_142_U9 ( .A(ref_1_n7), .B(ref_1_maj_142_n24), .Z(
        ref_1_maj_142_n26) );
  XOR2_X1 ref_1_maj_142_U8 ( .A(ref_1_n16), .B(ref_1_maj_142_n25), .Z(
        ref_1_maj_142_n27) );
  XOR2_X1 ref_1_maj_142_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_142_n24)
         );
  XOR2_X1 ref_1_maj_142_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_142_n25) );
  OR2_X1 ref_1_maj_142_U5 ( .A1(ref_1_maj_142_n23), .A2(ref_1_maj_142_n22), 
        .ZN(ref_1_maj_142_n32) );
  NAND2_X1 ref_1_maj_142_U4 ( .A1(ref_1_maj_142_n22), .A2(ref_1_maj_142_n23), 
        .ZN(ref_1_maj_142_n34) );
  NAND2_X1 ref_1_maj_142_U3 ( .A1(ref_1_maj_142_n32), .A2(ref_1_maj_142_n31), 
        .ZN(ref_1_maj_142_n33) );
  NAND2_X1 ref_1_maj_142_U2 ( .A1(ref_1_maj_142_n34), .A2(ref_1_maj_142_n33), 
        .ZN(ref_1_maj_142_port_o) );
  OR2_X1 ref_1_maj_143_U19 ( .A1(ref_1_maj_143_n27), .A2(ref_1_maj_143_n26), 
        .ZN(ref_1_maj_143_n28) );
  NAND2_X1 ref_1_maj_143_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_143_n28), .ZN(
        ref_1_maj_143_n29) );
  NAND2_X1 ref_1_maj_143_U17 ( .A1(ref_1_maj_143_n26), .A2(ref_1_maj_143_n27), 
        .ZN(ref_1_maj_143_n30) );
  NAND2_X1 ref_1_maj_143_U16 ( .A1(ref_1_maj_143_n30), .A2(ref_1_maj_143_n29), 
        .ZN(ref_1_maj_143_n31) );
  NAND2_X1 ref_1_maj_143_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_143_n25), .ZN(
        ref_1_maj_143_n18) );
  NAND2_X1 ref_1_maj_143_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_143_n19) );
  NAND2_X1 ref_1_maj_143_U13 ( .A1(ref_1_maj_143_n19), .A2(ref_1_maj_143_n18), 
        .ZN(ref_1_maj_143_n22) );
  NAND2_X1 ref_1_maj_143_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_143_n24), .ZN(
        ref_1_maj_143_n20) );
  NAND2_X1 ref_1_maj_143_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_143_n21) );
  NAND2_X1 ref_1_maj_143_U10 ( .A1(ref_1_maj_143_n21), .A2(ref_1_maj_143_n20), 
        .ZN(ref_1_maj_143_n23) );
  XOR2_X1 ref_1_maj_143_U9 ( .A(ref_1_n8), .B(ref_1_maj_143_n24), .Z(
        ref_1_maj_143_n26) );
  XOR2_X1 ref_1_maj_143_U8 ( .A(ref_1_n17), .B(ref_1_maj_143_n25), .Z(
        ref_1_maj_143_n27) );
  XOR2_X1 ref_1_maj_143_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_143_n24)
         );
  XOR2_X1 ref_1_maj_143_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_143_n25) );
  OR2_X1 ref_1_maj_143_U5 ( .A1(ref_1_maj_143_n23), .A2(ref_1_maj_143_n22), 
        .ZN(ref_1_maj_143_n32) );
  NAND2_X1 ref_1_maj_143_U4 ( .A1(ref_1_maj_143_n22), .A2(ref_1_maj_143_n23), 
        .ZN(ref_1_maj_143_n34) );
  NAND2_X1 ref_1_maj_143_U3 ( .A1(ref_1_maj_143_n32), .A2(ref_1_maj_143_n31), 
        .ZN(ref_1_maj_143_n33) );
  NAND2_X1 ref_1_maj_143_U2 ( .A1(ref_1_maj_143_n34), .A2(ref_1_maj_143_n33), 
        .ZN(ref_1_maj_143_port_o) );
  OR2_X1 ref_1_maj_144_U19 ( .A1(ref_1_maj_144_n27), .A2(ref_1_maj_144_n26), 
        .ZN(ref_1_maj_144_n28) );
  NAND2_X1 ref_1_maj_144_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_144_n28), .ZN(
        ref_1_maj_144_n29) );
  NAND2_X1 ref_1_maj_144_U17 ( .A1(ref_1_maj_144_n26), .A2(ref_1_maj_144_n27), 
        .ZN(ref_1_maj_144_n30) );
  NAND2_X1 ref_1_maj_144_U16 ( .A1(ref_1_maj_144_n30), .A2(ref_1_maj_144_n29), 
        .ZN(ref_1_maj_144_n31) );
  NAND2_X1 ref_1_maj_144_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_144_n25), .ZN(
        ref_1_maj_144_n18) );
  NAND2_X1 ref_1_maj_144_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_144_n19) );
  NAND2_X1 ref_1_maj_144_U13 ( .A1(ref_1_maj_144_n19), .A2(ref_1_maj_144_n18), 
        .ZN(ref_1_maj_144_n22) );
  NAND2_X1 ref_1_maj_144_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_144_n24), .ZN(
        ref_1_maj_144_n20) );
  NAND2_X1 ref_1_maj_144_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_144_n21) );
  NAND2_X1 ref_1_maj_144_U10 ( .A1(ref_1_maj_144_n21), .A2(ref_1_maj_144_n20), 
        .ZN(ref_1_maj_144_n23) );
  XOR2_X1 ref_1_maj_144_U9 ( .A(ref_1_n65), .B(ref_1_maj_144_n24), .Z(
        ref_1_maj_144_n26) );
  XOR2_X1 ref_1_maj_144_U8 ( .A(ref_1_n73), .B(ref_1_maj_144_n25), .Z(
        ref_1_maj_144_n27) );
  XOR2_X1 ref_1_maj_144_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_144_n24) );
  XOR2_X1 ref_1_maj_144_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_144_n25) );
  OR2_X1 ref_1_maj_144_U5 ( .A1(ref_1_maj_144_n23), .A2(ref_1_maj_144_n22), 
        .ZN(ref_1_maj_144_n32) );
  NAND2_X1 ref_1_maj_144_U4 ( .A1(ref_1_maj_144_n22), .A2(ref_1_maj_144_n23), 
        .ZN(ref_1_maj_144_n34) );
  NAND2_X1 ref_1_maj_144_U3 ( .A1(ref_1_maj_144_n32), .A2(ref_1_maj_144_n31), 
        .ZN(ref_1_maj_144_n33) );
  NAND2_X1 ref_1_maj_144_U2 ( .A1(ref_1_maj_144_n34), .A2(ref_1_maj_144_n33), 
        .ZN(ref_1_maj_144_port_o) );
  OR2_X1 ref_1_maj_145_U19 ( .A1(ref_1_maj_145_n27), .A2(ref_1_maj_145_n26), 
        .ZN(ref_1_maj_145_n28) );
  NAND2_X1 ref_1_maj_145_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_145_n28), .ZN(
        ref_1_maj_145_n29) );
  NAND2_X1 ref_1_maj_145_U17 ( .A1(ref_1_maj_145_n26), .A2(ref_1_maj_145_n27), 
        .ZN(ref_1_maj_145_n30) );
  NAND2_X1 ref_1_maj_145_U16 ( .A1(ref_1_maj_145_n30), .A2(ref_1_maj_145_n29), 
        .ZN(ref_1_maj_145_n31) );
  NAND2_X1 ref_1_maj_145_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_145_n25), .ZN(
        ref_1_maj_145_n18) );
  NAND2_X1 ref_1_maj_145_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_145_n19) );
  NAND2_X1 ref_1_maj_145_U13 ( .A1(ref_1_maj_145_n19), .A2(ref_1_maj_145_n18), 
        .ZN(ref_1_maj_145_n22) );
  NAND2_X1 ref_1_maj_145_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_145_n24), .ZN(
        ref_1_maj_145_n20) );
  NAND2_X1 ref_1_maj_145_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_145_n21) );
  NAND2_X1 ref_1_maj_145_U10 ( .A1(ref_1_maj_145_n21), .A2(ref_1_maj_145_n20), 
        .ZN(ref_1_maj_145_n23) );
  XOR2_X1 ref_1_maj_145_U9 ( .A(ref_1_n65), .B(ref_1_maj_145_n24), .Z(
        ref_1_maj_145_n26) );
  XOR2_X1 ref_1_maj_145_U8 ( .A(ref_1_n75), .B(ref_1_maj_145_n25), .Z(
        ref_1_maj_145_n27) );
  XOR2_X1 ref_1_maj_145_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_145_n24) );
  XOR2_X1 ref_1_maj_145_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_145_n25) );
  OR2_X1 ref_1_maj_145_U5 ( .A1(ref_1_maj_145_n23), .A2(ref_1_maj_145_n22), 
        .ZN(ref_1_maj_145_n32) );
  NAND2_X1 ref_1_maj_145_U4 ( .A1(ref_1_maj_145_n22), .A2(ref_1_maj_145_n23), 
        .ZN(ref_1_maj_145_n34) );
  NAND2_X1 ref_1_maj_145_U3 ( .A1(ref_1_maj_145_n32), .A2(ref_1_maj_145_n31), 
        .ZN(ref_1_maj_145_n33) );
  NAND2_X1 ref_1_maj_145_U2 ( .A1(ref_1_maj_145_n34), .A2(ref_1_maj_145_n33), 
        .ZN(ref_1_maj_145_port_o) );
  OR2_X1 ref_1_maj_146_U19 ( .A1(ref_1_maj_146_n27), .A2(ref_1_maj_146_n26), 
        .ZN(ref_1_maj_146_n28) );
  NAND2_X1 ref_1_maj_146_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_146_n28), .ZN(
        ref_1_maj_146_n29) );
  NAND2_X1 ref_1_maj_146_U17 ( .A1(ref_1_maj_146_n26), .A2(ref_1_maj_146_n27), 
        .ZN(ref_1_maj_146_n30) );
  NAND2_X1 ref_1_maj_146_U16 ( .A1(ref_1_maj_146_n30), .A2(ref_1_maj_146_n29), 
        .ZN(ref_1_maj_146_n31) );
  NAND2_X1 ref_1_maj_146_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_146_n25), .ZN(
        ref_1_maj_146_n18) );
  NAND2_X1 ref_1_maj_146_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_146_n19) );
  NAND2_X1 ref_1_maj_146_U13 ( .A1(ref_1_maj_146_n19), .A2(ref_1_maj_146_n18), 
        .ZN(ref_1_maj_146_n22) );
  NAND2_X1 ref_1_maj_146_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_146_n24), .ZN(
        ref_1_maj_146_n20) );
  NAND2_X1 ref_1_maj_146_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_146_n21) );
  NAND2_X1 ref_1_maj_146_U10 ( .A1(ref_1_maj_146_n21), .A2(ref_1_maj_146_n20), 
        .ZN(ref_1_maj_146_n23) );
  XOR2_X1 ref_1_maj_146_U9 ( .A(ref_1_n65), .B(ref_1_maj_146_n24), .Z(
        ref_1_maj_146_n26) );
  XOR2_X1 ref_1_maj_146_U8 ( .A(ref_1_n74), .B(ref_1_maj_146_n25), .Z(
        ref_1_maj_146_n27) );
  XOR2_X1 ref_1_maj_146_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_146_n24) );
  XOR2_X1 ref_1_maj_146_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_146_n25) );
  OR2_X1 ref_1_maj_146_U5 ( .A1(ref_1_maj_146_n23), .A2(ref_1_maj_146_n22), 
        .ZN(ref_1_maj_146_n32) );
  NAND2_X1 ref_1_maj_146_U4 ( .A1(ref_1_maj_146_n22), .A2(ref_1_maj_146_n23), 
        .ZN(ref_1_maj_146_n34) );
  NAND2_X1 ref_1_maj_146_U3 ( .A1(ref_1_maj_146_n32), .A2(ref_1_maj_146_n31), 
        .ZN(ref_1_maj_146_n33) );
  NAND2_X1 ref_1_maj_146_U2 ( .A1(ref_1_maj_146_n34), .A2(ref_1_maj_146_n33), 
        .ZN(ref_1_maj_146_port_o) );
  OR2_X1 ref_1_maj_147_U19 ( .A1(ref_1_maj_147_n27), .A2(ref_1_maj_147_n26), 
        .ZN(ref_1_maj_147_n28) );
  NAND2_X1 ref_1_maj_147_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_147_n28), .ZN(
        ref_1_maj_147_n29) );
  NAND2_X1 ref_1_maj_147_U17 ( .A1(ref_1_maj_147_n26), .A2(ref_1_maj_147_n27), 
        .ZN(ref_1_maj_147_n30) );
  NAND2_X1 ref_1_maj_147_U16 ( .A1(ref_1_maj_147_n30), .A2(ref_1_maj_147_n29), 
        .ZN(ref_1_maj_147_n31) );
  NAND2_X1 ref_1_maj_147_U15 ( .A1(ref_1_n73), .A2(ref_1_maj_147_n25), .ZN(
        ref_1_maj_147_n18) );
  NAND2_X1 ref_1_maj_147_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_147_n19) );
  NAND2_X1 ref_1_maj_147_U13 ( .A1(ref_1_maj_147_n19), .A2(ref_1_maj_147_n18), 
        .ZN(ref_1_maj_147_n22) );
  NAND2_X1 ref_1_maj_147_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_147_n24), .ZN(
        ref_1_maj_147_n20) );
  NAND2_X1 ref_1_maj_147_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_147_n21) );
  NAND2_X1 ref_1_maj_147_U10 ( .A1(ref_1_maj_147_n21), .A2(ref_1_maj_147_n20), 
        .ZN(ref_1_maj_147_n23) );
  XOR2_X1 ref_1_maj_147_U9 ( .A(ref_1_n65), .B(ref_1_maj_147_n24), .Z(
        ref_1_maj_147_n26) );
  XOR2_X1 ref_1_maj_147_U8 ( .A(ref_1_n73), .B(ref_1_maj_147_n25), .Z(
        ref_1_maj_147_n27) );
  XOR2_X1 ref_1_maj_147_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_147_n24) );
  XOR2_X1 ref_1_maj_147_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_147_n25) );
  OR2_X1 ref_1_maj_147_U5 ( .A1(ref_1_maj_147_n23), .A2(ref_1_maj_147_n22), 
        .ZN(ref_1_maj_147_n32) );
  NAND2_X1 ref_1_maj_147_U4 ( .A1(ref_1_maj_147_n22), .A2(ref_1_maj_147_n23), 
        .ZN(ref_1_maj_147_n34) );
  NAND2_X1 ref_1_maj_147_U3 ( .A1(ref_1_maj_147_n32), .A2(ref_1_maj_147_n31), 
        .ZN(ref_1_maj_147_n33) );
  NAND2_X1 ref_1_maj_147_U2 ( .A1(ref_1_maj_147_n34), .A2(ref_1_maj_147_n33), 
        .ZN(ref_1_maj_147_port_o) );
  OR2_X1 ref_1_maj_148_U19 ( .A1(ref_1_maj_148_n27), .A2(ref_1_maj_148_n26), 
        .ZN(ref_1_maj_148_n28) );
  NAND2_X1 ref_1_maj_148_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_148_n28), .ZN(
        ref_1_maj_148_n29) );
  NAND2_X1 ref_1_maj_148_U17 ( .A1(ref_1_maj_148_n26), .A2(ref_1_maj_148_n27), 
        .ZN(ref_1_maj_148_n30) );
  NAND2_X1 ref_1_maj_148_U16 ( .A1(ref_1_maj_148_n30), .A2(ref_1_maj_148_n29), 
        .ZN(ref_1_maj_148_n31) );
  NAND2_X1 ref_1_maj_148_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_148_n25), .ZN(
        ref_1_maj_148_n18) );
  NAND2_X1 ref_1_maj_148_U14 ( .A1(ref_1_n50), .A2(ref_1_n52), .ZN(
        ref_1_maj_148_n19) );
  NAND2_X1 ref_1_maj_148_U13 ( .A1(ref_1_maj_148_n19), .A2(ref_1_maj_148_n18), 
        .ZN(ref_1_maj_148_n22) );
  NAND2_X1 ref_1_maj_148_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_148_n24), .ZN(
        ref_1_maj_148_n20) );
  NAND2_X1 ref_1_maj_148_U11 ( .A1(ref_1_n41), .A2(ref_1_n43), .ZN(
        ref_1_maj_148_n21) );
  NAND2_X1 ref_1_maj_148_U10 ( .A1(ref_1_maj_148_n21), .A2(ref_1_maj_148_n20), 
        .ZN(ref_1_maj_148_n23) );
  XOR2_X1 ref_1_maj_148_U9 ( .A(ref_1_n46), .B(ref_1_maj_148_n24), .Z(
        ref_1_maj_148_n26) );
  XOR2_X1 ref_1_maj_148_U8 ( .A(ref_1_n56), .B(ref_1_maj_148_n25), .Z(
        ref_1_maj_148_n27) );
  XOR2_X1 ref_1_maj_148_U7 ( .A(ref_1_n41), .B(ref_1_n43), .Z(
        ref_1_maj_148_n24) );
  XOR2_X1 ref_1_maj_148_U6 ( .A(ref_1_n50), .B(ref_1_n52), .Z(
        ref_1_maj_148_n25) );
  OR2_X1 ref_1_maj_148_U5 ( .A1(ref_1_maj_148_n23), .A2(ref_1_maj_148_n22), 
        .ZN(ref_1_maj_148_n32) );
  NAND2_X1 ref_1_maj_148_U4 ( .A1(ref_1_maj_148_n22), .A2(ref_1_maj_148_n23), 
        .ZN(ref_1_maj_148_n34) );
  NAND2_X1 ref_1_maj_148_U3 ( .A1(ref_1_maj_148_n32), .A2(ref_1_maj_148_n31), 
        .ZN(ref_1_maj_148_n33) );
  NAND2_X1 ref_1_maj_148_U2 ( .A1(ref_1_maj_148_n34), .A2(ref_1_maj_148_n33), 
        .ZN(ref_1_maj_148_port_o) );
  OR2_X1 ref_1_maj_149_U19 ( .A1(ref_1_maj_149_n27), .A2(ref_1_maj_149_n26), 
        .ZN(ref_1_maj_149_n28) );
  NAND2_X1 ref_1_maj_149_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_149_n28), .ZN(
        ref_1_maj_149_n29) );
  NAND2_X1 ref_1_maj_149_U17 ( .A1(ref_1_maj_149_n26), .A2(ref_1_maj_149_n27), 
        .ZN(ref_1_maj_149_n30) );
  NAND2_X1 ref_1_maj_149_U16 ( .A1(ref_1_maj_149_n30), .A2(ref_1_maj_149_n29), 
        .ZN(ref_1_maj_149_n31) );
  NAND2_X1 ref_1_maj_149_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_149_n25), .ZN(
        ref_1_maj_149_n18) );
  NAND2_X1 ref_1_maj_149_U14 ( .A1(ref_1_n49), .A2(ref_1_n52), .ZN(
        ref_1_maj_149_n19) );
  NAND2_X1 ref_1_maj_149_U13 ( .A1(ref_1_maj_149_n19), .A2(ref_1_maj_149_n18), 
        .ZN(ref_1_maj_149_n22) );
  NAND2_X1 ref_1_maj_149_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_149_n24), .ZN(
        ref_1_maj_149_n20) );
  NAND2_X1 ref_1_maj_149_U11 ( .A1(ref_1_n40), .A2(ref_1_n43), .ZN(
        ref_1_maj_149_n21) );
  NAND2_X1 ref_1_maj_149_U10 ( .A1(ref_1_maj_149_n21), .A2(ref_1_maj_149_n20), 
        .ZN(ref_1_maj_149_n23) );
  XOR2_X1 ref_1_maj_149_U9 ( .A(ref_1_n46), .B(ref_1_maj_149_n24), .Z(
        ref_1_maj_149_n26) );
  XOR2_X1 ref_1_maj_149_U8 ( .A(ref_1_n55), .B(ref_1_maj_149_n25), .Z(
        ref_1_maj_149_n27) );
  XOR2_X1 ref_1_maj_149_U7 ( .A(ref_1_n40), .B(ref_1_n43), .Z(
        ref_1_maj_149_n24) );
  XOR2_X1 ref_1_maj_149_U6 ( .A(ref_1_n49), .B(ref_1_n52), .Z(
        ref_1_maj_149_n25) );
  OR2_X1 ref_1_maj_149_U5 ( .A1(ref_1_maj_149_n23), .A2(ref_1_maj_149_n22), 
        .ZN(ref_1_maj_149_n32) );
  NAND2_X1 ref_1_maj_149_U4 ( .A1(ref_1_maj_149_n22), .A2(ref_1_maj_149_n23), 
        .ZN(ref_1_maj_149_n34) );
  NAND2_X1 ref_1_maj_149_U3 ( .A1(ref_1_maj_149_n32), .A2(ref_1_maj_149_n31), 
        .ZN(ref_1_maj_149_n33) );
  NAND2_X1 ref_1_maj_149_U2 ( .A1(ref_1_maj_149_n34), .A2(ref_1_maj_149_n33), 
        .ZN(ref_1_maj_149_port_o) );
  OR2_X1 ref_1_maj_150_U19 ( .A1(ref_1_maj_150_n27), .A2(ref_1_maj_150_n26), 
        .ZN(ref_1_maj_150_n28) );
  NAND2_X1 ref_1_maj_150_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_150_n28), .ZN(
        ref_1_maj_150_n29) );
  NAND2_X1 ref_1_maj_150_U17 ( .A1(ref_1_maj_150_n26), .A2(ref_1_maj_150_n27), 
        .ZN(ref_1_maj_150_n30) );
  NAND2_X1 ref_1_maj_150_U16 ( .A1(ref_1_maj_150_n30), .A2(ref_1_maj_150_n29), 
        .ZN(ref_1_maj_150_n31) );
  NAND2_X1 ref_1_maj_150_U15 ( .A1(ref_1_n54), .A2(ref_1_maj_150_n25), .ZN(
        ref_1_maj_150_n18) );
  NAND2_X1 ref_1_maj_150_U14 ( .A1(ref_1_n48), .A2(ref_1_n52), .ZN(
        ref_1_maj_150_n19) );
  NAND2_X1 ref_1_maj_150_U13 ( .A1(ref_1_maj_150_n19), .A2(ref_1_maj_150_n18), 
        .ZN(ref_1_maj_150_n22) );
  NAND2_X1 ref_1_maj_150_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_150_n24), .ZN(
        ref_1_maj_150_n20) );
  NAND2_X1 ref_1_maj_150_U11 ( .A1(ref_1_n39), .A2(ref_1_n43), .ZN(
        ref_1_maj_150_n21) );
  NAND2_X1 ref_1_maj_150_U10 ( .A1(ref_1_maj_150_n21), .A2(ref_1_maj_150_n20), 
        .ZN(ref_1_maj_150_n23) );
  XOR2_X1 ref_1_maj_150_U9 ( .A(ref_1_n46), .B(ref_1_maj_150_n24), .Z(
        ref_1_maj_150_n26) );
  XOR2_X1 ref_1_maj_150_U8 ( .A(ref_1_n54), .B(ref_1_maj_150_n25), .Z(
        ref_1_maj_150_n27) );
  XOR2_X1 ref_1_maj_150_U7 ( .A(ref_1_n39), .B(ref_1_n43), .Z(
        ref_1_maj_150_n24) );
  XOR2_X1 ref_1_maj_150_U6 ( .A(ref_1_n48), .B(ref_1_n52), .Z(
        ref_1_maj_150_n25) );
  OR2_X1 ref_1_maj_150_U5 ( .A1(ref_1_maj_150_n23), .A2(ref_1_maj_150_n22), 
        .ZN(ref_1_maj_150_n32) );
  NAND2_X1 ref_1_maj_150_U4 ( .A1(ref_1_maj_150_n22), .A2(ref_1_maj_150_n23), 
        .ZN(ref_1_maj_150_n34) );
  NAND2_X1 ref_1_maj_150_U3 ( .A1(ref_1_maj_150_n32), .A2(ref_1_maj_150_n31), 
        .ZN(ref_1_maj_150_n33) );
  NAND2_X1 ref_1_maj_150_U2 ( .A1(ref_1_maj_150_n34), .A2(ref_1_maj_150_n33), 
        .ZN(ref_1_maj_150_port_o) );
  OR2_X1 ref_1_maj_151_U19 ( .A1(ref_1_maj_151_n27), .A2(ref_1_maj_151_n26), 
        .ZN(ref_1_maj_151_n28) );
  NAND2_X1 ref_1_maj_151_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_151_n28), .ZN(
        ref_1_maj_151_n29) );
  NAND2_X1 ref_1_maj_151_U17 ( .A1(ref_1_maj_151_n26), .A2(ref_1_maj_151_n27), 
        .ZN(ref_1_maj_151_n30) );
  NAND2_X1 ref_1_maj_151_U16 ( .A1(ref_1_maj_151_n30), .A2(ref_1_maj_151_n29), 
        .ZN(ref_1_maj_151_n31) );
  NAND2_X1 ref_1_maj_151_U15 ( .A1(ref_1_refreshed_1_5_), .A2(
        ref_1_maj_151_n25), .ZN(ref_1_maj_151_n18) );
  NAND2_X1 ref_1_maj_151_U14 ( .A1(ref_1_refreshed_1_3_), .A2(ref_1_n52), .ZN(
        ref_1_maj_151_n19) );
  NAND2_X1 ref_1_maj_151_U13 ( .A1(ref_1_maj_151_n19), .A2(ref_1_maj_151_n18), 
        .ZN(ref_1_maj_151_n22) );
  NAND2_X1 ref_1_maj_151_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_151_n24), .ZN(
        ref_1_maj_151_n20) );
  NAND2_X1 ref_1_maj_151_U11 ( .A1(ref_1_refreshed_1_0_), .A2(ref_1_n43), .ZN(
        ref_1_maj_151_n21) );
  NAND2_X1 ref_1_maj_151_U10 ( .A1(ref_1_maj_151_n21), .A2(ref_1_maj_151_n20), 
        .ZN(ref_1_maj_151_n23) );
  XOR2_X1 ref_1_maj_151_U9 ( .A(ref_1_n46), .B(ref_1_maj_151_n24), .Z(
        ref_1_maj_151_n26) );
  XOR2_X1 ref_1_maj_151_U8 ( .A(ref_1_refreshed_1_5_), .B(ref_1_maj_151_n25), 
        .Z(ref_1_maj_151_n27) );
  XOR2_X1 ref_1_maj_151_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_n43), .Z(
        ref_1_maj_151_n24) );
  XOR2_X1 ref_1_maj_151_U6 ( .A(ref_1_refreshed_1_3_), .B(ref_1_n52), .Z(
        ref_1_maj_151_n25) );
  OR2_X1 ref_1_maj_151_U5 ( .A1(ref_1_maj_151_n23), .A2(ref_1_maj_151_n22), 
        .ZN(ref_1_maj_151_n32) );
  NAND2_X1 ref_1_maj_151_U4 ( .A1(ref_1_maj_151_n22), .A2(ref_1_maj_151_n23), 
        .ZN(ref_1_maj_151_n34) );
  NAND2_X1 ref_1_maj_151_U3 ( .A1(ref_1_maj_151_n32), .A2(ref_1_maj_151_n31), 
        .ZN(ref_1_maj_151_n33) );
  NAND2_X1 ref_1_maj_151_U2 ( .A1(ref_1_maj_151_n34), .A2(ref_1_maj_151_n33), 
        .ZN(ref_1_maj_151_port_o) );
  OR2_X1 ref_1_maj_152_U19 ( .A1(ref_1_maj_152_n27), .A2(ref_1_maj_152_n26), 
        .ZN(ref_1_maj_152_n28) );
  NAND2_X1 ref_1_maj_152_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_152_n28), .ZN(
        ref_1_maj_152_n29) );
  NAND2_X1 ref_1_maj_152_U17 ( .A1(ref_1_maj_152_n26), .A2(ref_1_maj_152_n27), 
        .ZN(ref_1_maj_152_n30) );
  NAND2_X1 ref_1_maj_152_U16 ( .A1(ref_1_maj_152_n30), .A2(ref_1_maj_152_n29), 
        .ZN(ref_1_maj_152_n31) );
  NAND2_X1 ref_1_maj_152_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_152_n25), .ZN(
        ref_1_maj_152_n18) );
  NAND2_X1 ref_1_maj_152_U14 ( .A1(ref_1_n30), .A2(ref_1_n34), .ZN(
        ref_1_maj_152_n19) );
  NAND2_X1 ref_1_maj_152_U13 ( .A1(ref_1_maj_152_n19), .A2(ref_1_maj_152_n18), 
        .ZN(ref_1_maj_152_n22) );
  NAND2_X1 ref_1_maj_152_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_152_n24), .ZN(
        ref_1_maj_152_n20) );
  NAND2_X1 ref_1_maj_152_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_152_n21) );
  NAND2_X1 ref_1_maj_152_U10 ( .A1(ref_1_maj_152_n21), .A2(ref_1_maj_152_n20), 
        .ZN(ref_1_maj_152_n23) );
  XOR2_X1 ref_1_maj_152_U9 ( .A(ref_1_n27), .B(ref_1_maj_152_n24), .Z(
        ref_1_maj_152_n26) );
  XOR2_X1 ref_1_maj_152_U8 ( .A(ref_1_n36), .B(ref_1_maj_152_n25), .Z(
        ref_1_maj_152_n27) );
  XOR2_X1 ref_1_maj_152_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_152_n24) );
  XOR2_X1 ref_1_maj_152_U6 ( .A(ref_1_n30), .B(ref_1_n34), .Z(
        ref_1_maj_152_n25) );
  OR2_X1 ref_1_maj_152_U5 ( .A1(ref_1_maj_152_n23), .A2(ref_1_maj_152_n22), 
        .ZN(ref_1_maj_152_n32) );
  NAND2_X1 ref_1_maj_152_U4 ( .A1(ref_1_maj_152_n22), .A2(ref_1_maj_152_n23), 
        .ZN(ref_1_maj_152_n34) );
  NAND2_X1 ref_1_maj_152_U3 ( .A1(ref_1_maj_152_n32), .A2(ref_1_maj_152_n31), 
        .ZN(ref_1_maj_152_n33) );
  NAND2_X1 ref_1_maj_152_U2 ( .A1(ref_1_maj_152_n34), .A2(ref_1_maj_152_n33), 
        .ZN(ref_1_maj_152_port_o) );
  OR2_X1 ref_1_maj_153_U19 ( .A1(ref_1_maj_153_n27), .A2(ref_1_maj_153_n26), 
        .ZN(ref_1_maj_153_n28) );
  NAND2_X1 ref_1_maj_153_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_153_n28), .ZN(
        ref_1_maj_153_n29) );
  NAND2_X1 ref_1_maj_153_U17 ( .A1(ref_1_maj_153_n26), .A2(ref_1_maj_153_n27), 
        .ZN(ref_1_maj_153_n30) );
  NAND2_X1 ref_1_maj_153_U16 ( .A1(ref_1_maj_153_n30), .A2(ref_1_maj_153_n29), 
        .ZN(ref_1_maj_153_n31) );
  NAND2_X1 ref_1_maj_153_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_153_n25), .ZN(
        ref_1_maj_153_n18) );
  NAND2_X1 ref_1_maj_153_U14 ( .A1(ref_1_n30), .A2(ref_1_n33), .ZN(
        ref_1_maj_153_n19) );
  NAND2_X1 ref_1_maj_153_U13 ( .A1(ref_1_maj_153_n19), .A2(ref_1_maj_153_n18), 
        .ZN(ref_1_maj_153_n22) );
  NAND2_X1 ref_1_maj_153_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_153_n24), .ZN(
        ref_1_maj_153_n20) );
  NAND2_X1 ref_1_maj_153_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_153_n21) );
  NAND2_X1 ref_1_maj_153_U10 ( .A1(ref_1_maj_153_n21), .A2(ref_1_maj_153_n20), 
        .ZN(ref_1_maj_153_n23) );
  XOR2_X1 ref_1_maj_153_U9 ( .A(ref_1_n27), .B(ref_1_maj_153_n24), .Z(
        ref_1_maj_153_n26) );
  XOR2_X1 ref_1_maj_153_U8 ( .A(ref_1_n36), .B(ref_1_maj_153_n25), .Z(
        ref_1_maj_153_n27) );
  XOR2_X1 ref_1_maj_153_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_153_n24) );
  XOR2_X1 ref_1_maj_153_U6 ( .A(ref_1_n30), .B(ref_1_n33), .Z(
        ref_1_maj_153_n25) );
  OR2_X1 ref_1_maj_153_U5 ( .A1(ref_1_maj_153_n23), .A2(ref_1_maj_153_n22), 
        .ZN(ref_1_maj_153_n32) );
  NAND2_X1 ref_1_maj_153_U4 ( .A1(ref_1_maj_153_n22), .A2(ref_1_maj_153_n23), 
        .ZN(ref_1_maj_153_n34) );
  NAND2_X1 ref_1_maj_153_U3 ( .A1(ref_1_maj_153_n32), .A2(ref_1_maj_153_n31), 
        .ZN(ref_1_maj_153_n33) );
  NAND2_X1 ref_1_maj_153_U2 ( .A1(ref_1_maj_153_n34), .A2(ref_1_maj_153_n33), 
        .ZN(ref_1_maj_153_port_o) );
  OR2_X1 ref_1_maj_154_U19 ( .A1(ref_1_maj_154_n27), .A2(ref_1_maj_154_n26), 
        .ZN(ref_1_maj_154_n28) );
  NAND2_X1 ref_1_maj_154_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_154_n28), .ZN(
        ref_1_maj_154_n29) );
  NAND2_X1 ref_1_maj_154_U17 ( .A1(ref_1_maj_154_n26), .A2(ref_1_maj_154_n27), 
        .ZN(ref_1_maj_154_n30) );
  NAND2_X1 ref_1_maj_154_U16 ( .A1(ref_1_maj_154_n30), .A2(ref_1_maj_154_n29), 
        .ZN(ref_1_maj_154_n31) );
  NAND2_X1 ref_1_maj_154_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_154_n25), .ZN(
        ref_1_maj_154_n18) );
  NAND2_X1 ref_1_maj_154_U14 ( .A1(ref_1_n30), .A2(ref_1_n32), .ZN(
        ref_1_maj_154_n19) );
  NAND2_X1 ref_1_maj_154_U13 ( .A1(ref_1_maj_154_n19), .A2(ref_1_maj_154_n18), 
        .ZN(ref_1_maj_154_n22) );
  NAND2_X1 ref_1_maj_154_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_154_n24), .ZN(
        ref_1_maj_154_n20) );
  NAND2_X1 ref_1_maj_154_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_154_n21) );
  NAND2_X1 ref_1_maj_154_U10 ( .A1(ref_1_maj_154_n21), .A2(ref_1_maj_154_n20), 
        .ZN(ref_1_maj_154_n23) );
  XOR2_X1 ref_1_maj_154_U9 ( .A(ref_1_n27), .B(ref_1_maj_154_n24), .Z(
        ref_1_maj_154_n26) );
  XOR2_X1 ref_1_maj_154_U8 ( .A(ref_1_n36), .B(ref_1_maj_154_n25), .Z(
        ref_1_maj_154_n27) );
  XOR2_X1 ref_1_maj_154_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_154_n24) );
  XOR2_X1 ref_1_maj_154_U6 ( .A(ref_1_n30), .B(ref_1_n32), .Z(
        ref_1_maj_154_n25) );
  OR2_X1 ref_1_maj_154_U5 ( .A1(ref_1_maj_154_n23), .A2(ref_1_maj_154_n22), 
        .ZN(ref_1_maj_154_n32) );
  NAND2_X1 ref_1_maj_154_U4 ( .A1(ref_1_maj_154_n22), .A2(ref_1_maj_154_n23), 
        .ZN(ref_1_maj_154_n34) );
  NAND2_X1 ref_1_maj_154_U3 ( .A1(ref_1_maj_154_n32), .A2(ref_1_maj_154_n31), 
        .ZN(ref_1_maj_154_n33) );
  NAND2_X1 ref_1_maj_154_U2 ( .A1(ref_1_maj_154_n34), .A2(ref_1_maj_154_n33), 
        .ZN(ref_1_maj_154_port_o) );
  OR2_X1 ref_1_maj_155_U19 ( .A1(ref_1_maj_155_n27), .A2(ref_1_maj_155_n26), 
        .ZN(ref_1_maj_155_n28) );
  NAND2_X1 ref_1_maj_155_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_155_n28), .ZN(
        ref_1_maj_155_n29) );
  NAND2_X1 ref_1_maj_155_U17 ( .A1(ref_1_maj_155_n26), .A2(ref_1_maj_155_n27), 
        .ZN(ref_1_maj_155_n30) );
  NAND2_X1 ref_1_maj_155_U16 ( .A1(ref_1_maj_155_n30), .A2(ref_1_maj_155_n29), 
        .ZN(ref_1_maj_155_n31) );
  NAND2_X1 ref_1_maj_155_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_155_n25), .ZN(
        ref_1_maj_155_n18) );
  NAND2_X1 ref_1_maj_155_U14 ( .A1(ref_1_n30), .A2(ref_1_refreshed_2_4_), .ZN(
        ref_1_maj_155_n19) );
  NAND2_X1 ref_1_maj_155_U13 ( .A1(ref_1_maj_155_n19), .A2(ref_1_maj_155_n18), 
        .ZN(ref_1_maj_155_n22) );
  NAND2_X1 ref_1_maj_155_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_155_n24), .ZN(
        ref_1_maj_155_n20) );
  NAND2_X1 ref_1_maj_155_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_155_n21) );
  NAND2_X1 ref_1_maj_155_U10 ( .A1(ref_1_maj_155_n21), .A2(ref_1_maj_155_n20), 
        .ZN(ref_1_maj_155_n23) );
  XOR2_X1 ref_1_maj_155_U9 ( .A(ref_1_n27), .B(ref_1_maj_155_n24), .Z(
        ref_1_maj_155_n26) );
  XOR2_X1 ref_1_maj_155_U8 ( .A(ref_1_n36), .B(ref_1_maj_155_n25), .Z(
        ref_1_maj_155_n27) );
  XOR2_X1 ref_1_maj_155_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_155_n24) );
  XOR2_X1 ref_1_maj_155_U6 ( .A(ref_1_n30), .B(ref_1_refreshed_2_4_), .Z(
        ref_1_maj_155_n25) );
  OR2_X1 ref_1_maj_155_U5 ( .A1(ref_1_maj_155_n23), .A2(ref_1_maj_155_n22), 
        .ZN(ref_1_maj_155_n32) );
  NAND2_X1 ref_1_maj_155_U4 ( .A1(ref_1_maj_155_n22), .A2(ref_1_maj_155_n23), 
        .ZN(ref_1_maj_155_n34) );
  NAND2_X1 ref_1_maj_155_U3 ( .A1(ref_1_maj_155_n32), .A2(ref_1_maj_155_n31), 
        .ZN(ref_1_maj_155_n33) );
  NAND2_X1 ref_1_maj_155_U2 ( .A1(ref_1_maj_155_n34), .A2(ref_1_maj_155_n33), 
        .ZN(ref_1_maj_155_port_o) );
  OR2_X1 ref_1_maj_156_U19 ( .A1(ref_1_maj_156_n27), .A2(ref_1_maj_156_n26), 
        .ZN(ref_1_maj_156_n28) );
  NAND2_X1 ref_1_maj_156_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_156_n28), .ZN(
        ref_1_maj_156_n29) );
  NAND2_X1 ref_1_maj_156_U17 ( .A1(ref_1_maj_156_n26), .A2(ref_1_maj_156_n27), 
        .ZN(ref_1_maj_156_n30) );
  NAND2_X1 ref_1_maj_156_U16 ( .A1(ref_1_maj_156_n30), .A2(ref_1_maj_156_n29), 
        .ZN(ref_1_maj_156_n31) );
  NAND2_X1 ref_1_maj_156_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_156_n25), .ZN(
        ref_1_maj_156_n18) );
  NAND2_X1 ref_1_maj_156_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_156_n19) );
  NAND2_X1 ref_1_maj_156_U13 ( .A1(ref_1_maj_156_n19), .A2(ref_1_maj_156_n18), 
        .ZN(ref_1_maj_156_n22) );
  NAND2_X1 ref_1_maj_156_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_156_n24), .ZN(
        ref_1_maj_156_n20) );
  NAND2_X1 ref_1_maj_156_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_156_n21) );
  NAND2_X1 ref_1_maj_156_U10 ( .A1(ref_1_maj_156_n21), .A2(ref_1_maj_156_n20), 
        .ZN(ref_1_maj_156_n23) );
  XOR2_X1 ref_1_maj_156_U9 ( .A(ref_1_n8), .B(ref_1_maj_156_n24), .Z(
        ref_1_maj_156_n26) );
  XOR2_X1 ref_1_maj_156_U8 ( .A(ref_1_n17), .B(ref_1_maj_156_n25), .Z(
        ref_1_maj_156_n27) );
  XOR2_X1 ref_1_maj_156_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_156_n24)
         );
  XOR2_X1 ref_1_maj_156_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_156_n25) );
  OR2_X1 ref_1_maj_156_U5 ( .A1(ref_1_maj_156_n23), .A2(ref_1_maj_156_n22), 
        .ZN(ref_1_maj_156_n32) );
  NAND2_X1 ref_1_maj_156_U4 ( .A1(ref_1_maj_156_n22), .A2(ref_1_maj_156_n23), 
        .ZN(ref_1_maj_156_n34) );
  NAND2_X1 ref_1_maj_156_U3 ( .A1(ref_1_maj_156_n32), .A2(ref_1_maj_156_n31), 
        .ZN(ref_1_maj_156_n33) );
  NAND2_X1 ref_1_maj_156_U2 ( .A1(ref_1_maj_156_n34), .A2(ref_1_maj_156_n33), 
        .ZN(ref_1_maj_156_port_o) );
  OR2_X1 ref_1_maj_157_U19 ( .A1(ref_1_maj_157_n27), .A2(ref_1_maj_157_n26), 
        .ZN(ref_1_maj_157_n28) );
  NAND2_X1 ref_1_maj_157_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_157_n28), .ZN(
        ref_1_maj_157_n29) );
  NAND2_X1 ref_1_maj_157_U17 ( .A1(ref_1_maj_157_n26), .A2(ref_1_maj_157_n27), 
        .ZN(ref_1_maj_157_n30) );
  NAND2_X1 ref_1_maj_157_U16 ( .A1(ref_1_maj_157_n30), .A2(ref_1_maj_157_n29), 
        .ZN(ref_1_maj_157_n31) );
  NAND2_X1 ref_1_maj_157_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_157_n25), .ZN(
        ref_1_maj_157_n18) );
  NAND2_X1 ref_1_maj_157_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_157_n19) );
  NAND2_X1 ref_1_maj_157_U13 ( .A1(ref_1_maj_157_n19), .A2(ref_1_maj_157_n18), 
        .ZN(ref_1_maj_157_n22) );
  NAND2_X1 ref_1_maj_157_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_157_n24), .ZN(
        ref_1_maj_157_n20) );
  NAND2_X1 ref_1_maj_157_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_157_n21) );
  NAND2_X1 ref_1_maj_157_U10 ( .A1(ref_1_maj_157_n21), .A2(ref_1_maj_157_n20), 
        .ZN(ref_1_maj_157_n23) );
  XOR2_X1 ref_1_maj_157_U9 ( .A(ref_1_n8), .B(ref_1_maj_157_n24), .Z(
        ref_1_maj_157_n26) );
  XOR2_X1 ref_1_maj_157_U8 ( .A(ref_1_n17), .B(ref_1_maj_157_n25), .Z(
        ref_1_maj_157_n27) );
  XOR2_X1 ref_1_maj_157_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_157_n24)
         );
  XOR2_X1 ref_1_maj_157_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_157_n25) );
  OR2_X1 ref_1_maj_157_U5 ( .A1(ref_1_maj_157_n23), .A2(ref_1_maj_157_n22), 
        .ZN(ref_1_maj_157_n32) );
  NAND2_X1 ref_1_maj_157_U4 ( .A1(ref_1_maj_157_n22), .A2(ref_1_maj_157_n23), 
        .ZN(ref_1_maj_157_n34) );
  NAND2_X1 ref_1_maj_157_U3 ( .A1(ref_1_maj_157_n32), .A2(ref_1_maj_157_n31), 
        .ZN(ref_1_maj_157_n33) );
  NAND2_X1 ref_1_maj_157_U2 ( .A1(ref_1_maj_157_n34), .A2(ref_1_maj_157_n33), 
        .ZN(ref_1_maj_157_port_o) );
  OR2_X1 ref_1_maj_158_U19 ( .A1(ref_1_maj_158_n27), .A2(ref_1_maj_158_n26), 
        .ZN(ref_1_maj_158_n28) );
  NAND2_X1 ref_1_maj_158_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_158_n28), .ZN(
        ref_1_maj_158_n29) );
  NAND2_X1 ref_1_maj_158_U17 ( .A1(ref_1_maj_158_n26), .A2(ref_1_maj_158_n27), 
        .ZN(ref_1_maj_158_n30) );
  NAND2_X1 ref_1_maj_158_U16 ( .A1(ref_1_maj_158_n30), .A2(ref_1_maj_158_n29), 
        .ZN(ref_1_maj_158_n31) );
  NAND2_X1 ref_1_maj_158_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_158_n25), .ZN(
        ref_1_maj_158_n18) );
  NAND2_X1 ref_1_maj_158_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_158_n19) );
  NAND2_X1 ref_1_maj_158_U13 ( .A1(ref_1_maj_158_n19), .A2(ref_1_maj_158_n18), 
        .ZN(ref_1_maj_158_n22) );
  NAND2_X1 ref_1_maj_158_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_158_n24), .ZN(
        ref_1_maj_158_n20) );
  NAND2_X1 ref_1_maj_158_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_158_n21) );
  NAND2_X1 ref_1_maj_158_U10 ( .A1(ref_1_maj_158_n21), .A2(ref_1_maj_158_n20), 
        .ZN(ref_1_maj_158_n23) );
  XOR2_X1 ref_1_maj_158_U9 ( .A(ref_1_n8), .B(ref_1_maj_158_n24), .Z(
        ref_1_maj_158_n26) );
  XOR2_X1 ref_1_maj_158_U8 ( .A(ref_1_n17), .B(ref_1_maj_158_n25), .Z(
        ref_1_maj_158_n27) );
  XOR2_X1 ref_1_maj_158_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_158_n24)
         );
  XOR2_X1 ref_1_maj_158_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_158_n25) );
  OR2_X1 ref_1_maj_158_U5 ( .A1(ref_1_maj_158_n23), .A2(ref_1_maj_158_n22), 
        .ZN(ref_1_maj_158_n32) );
  NAND2_X1 ref_1_maj_158_U4 ( .A1(ref_1_maj_158_n22), .A2(ref_1_maj_158_n23), 
        .ZN(ref_1_maj_158_n34) );
  NAND2_X1 ref_1_maj_158_U3 ( .A1(ref_1_maj_158_n32), .A2(ref_1_maj_158_n31), 
        .ZN(ref_1_maj_158_n33) );
  NAND2_X1 ref_1_maj_158_U2 ( .A1(ref_1_maj_158_n34), .A2(ref_1_maj_158_n33), 
        .ZN(ref_1_maj_158_port_o) );
  OR2_X1 ref_1_maj_159_U19 ( .A1(ref_1_maj_159_n27), .A2(ref_1_maj_159_n26), 
        .ZN(ref_1_maj_159_n28) );
  NAND2_X1 ref_1_maj_159_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_159_n28), .ZN(
        ref_1_maj_159_n29) );
  NAND2_X1 ref_1_maj_159_U17 ( .A1(ref_1_maj_159_n26), .A2(ref_1_maj_159_n27), 
        .ZN(ref_1_maj_159_n30) );
  NAND2_X1 ref_1_maj_159_U16 ( .A1(ref_1_maj_159_n30), .A2(ref_1_maj_159_n29), 
        .ZN(ref_1_maj_159_n31) );
  NAND2_X1 ref_1_maj_159_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_159_n25), .ZN(
        ref_1_maj_159_n18) );
  NAND2_X1 ref_1_maj_159_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_159_n19) );
  NAND2_X1 ref_1_maj_159_U13 ( .A1(ref_1_maj_159_n19), .A2(ref_1_maj_159_n18), 
        .ZN(ref_1_maj_159_n22) );
  NAND2_X1 ref_1_maj_159_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_159_n24), .ZN(
        ref_1_maj_159_n20) );
  NAND2_X1 ref_1_maj_159_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_159_n21) );
  NAND2_X1 ref_1_maj_159_U10 ( .A1(ref_1_maj_159_n21), .A2(ref_1_maj_159_n20), 
        .ZN(ref_1_maj_159_n23) );
  XOR2_X1 ref_1_maj_159_U9 ( .A(ref_1_n8), .B(ref_1_maj_159_n24), .Z(
        ref_1_maj_159_n26) );
  XOR2_X1 ref_1_maj_159_U8 ( .A(ref_1_n17), .B(ref_1_maj_159_n25), .Z(
        ref_1_maj_159_n27) );
  XOR2_X1 ref_1_maj_159_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_159_n24)
         );
  XOR2_X1 ref_1_maj_159_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_159_n25) );
  OR2_X1 ref_1_maj_159_U5 ( .A1(ref_1_maj_159_n23), .A2(ref_1_maj_159_n22), 
        .ZN(ref_1_maj_159_n32) );
  NAND2_X1 ref_1_maj_159_U4 ( .A1(ref_1_maj_159_n22), .A2(ref_1_maj_159_n23), 
        .ZN(ref_1_maj_159_n34) );
  NAND2_X1 ref_1_maj_159_U3 ( .A1(ref_1_maj_159_n32), .A2(ref_1_maj_159_n31), 
        .ZN(ref_1_maj_159_n33) );
  NAND2_X1 ref_1_maj_159_U2 ( .A1(ref_1_maj_159_n34), .A2(ref_1_maj_159_n33), 
        .ZN(ref_1_maj_159_port_o) );
  OR2_X1 ref_1_maj_160_U19 ( .A1(ref_1_maj_160_n27), .A2(ref_1_maj_160_n26), 
        .ZN(ref_1_maj_160_n28) );
  NAND2_X1 ref_1_maj_160_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_160_n28), .ZN(
        ref_1_maj_160_n29) );
  NAND2_X1 ref_1_maj_160_U17 ( .A1(ref_1_maj_160_n26), .A2(ref_1_maj_160_n27), 
        .ZN(ref_1_maj_160_n30) );
  NAND2_X1 ref_1_maj_160_U16 ( .A1(ref_1_maj_160_n30), .A2(ref_1_maj_160_n29), 
        .ZN(ref_1_maj_160_n31) );
  NAND2_X1 ref_1_maj_160_U15 ( .A1(ref_1_refreshed_0_5_), .A2(
        ref_1_maj_160_n25), .ZN(ref_1_maj_160_n18) );
  NAND2_X1 ref_1_maj_160_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_160_n19) );
  NAND2_X1 ref_1_maj_160_U13 ( .A1(ref_1_maj_160_n19), .A2(ref_1_maj_160_n18), 
        .ZN(ref_1_maj_160_n22) );
  NAND2_X1 ref_1_maj_160_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_160_n24), .ZN(
        ref_1_maj_160_n20) );
  NAND2_X1 ref_1_maj_160_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_160_n21) );
  NAND2_X1 ref_1_maj_160_U10 ( .A1(ref_1_maj_160_n21), .A2(ref_1_maj_160_n20), 
        .ZN(ref_1_maj_160_n23) );
  XOR2_X1 ref_1_maj_160_U9 ( .A(ref_1_n65), .B(ref_1_maj_160_n24), .Z(
        ref_1_maj_160_n26) );
  XOR2_X1 ref_1_maj_160_U8 ( .A(ref_1_refreshed_0_5_), .B(ref_1_maj_160_n25), 
        .Z(ref_1_maj_160_n27) );
  XOR2_X1 ref_1_maj_160_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_160_n24) );
  XOR2_X1 ref_1_maj_160_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_160_n25) );
  OR2_X1 ref_1_maj_160_U5 ( .A1(ref_1_maj_160_n23), .A2(ref_1_maj_160_n22), 
        .ZN(ref_1_maj_160_n32) );
  NAND2_X1 ref_1_maj_160_U4 ( .A1(ref_1_maj_160_n22), .A2(ref_1_maj_160_n23), 
        .ZN(ref_1_maj_160_n34) );
  NAND2_X1 ref_1_maj_160_U3 ( .A1(ref_1_maj_160_n32), .A2(ref_1_maj_160_n31), 
        .ZN(ref_1_maj_160_n33) );
  NAND2_X1 ref_1_maj_160_U2 ( .A1(ref_1_maj_160_n34), .A2(ref_1_maj_160_n33), 
        .ZN(ref_1_maj_160_port_o) );
  OR2_X1 ref_1_maj_161_U19 ( .A1(ref_1_maj_161_n27), .A2(ref_1_maj_161_n26), 
        .ZN(ref_1_maj_161_n28) );
  NAND2_X1 ref_1_maj_161_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_161_n28), .ZN(
        ref_1_maj_161_n29) );
  NAND2_X1 ref_1_maj_161_U17 ( .A1(ref_1_maj_161_n26), .A2(ref_1_maj_161_n27), 
        .ZN(ref_1_maj_161_n30) );
  NAND2_X1 ref_1_maj_161_U16 ( .A1(ref_1_maj_161_n30), .A2(ref_1_maj_161_n29), 
        .ZN(ref_1_maj_161_n31) );
  NAND2_X1 ref_1_maj_161_U15 ( .A1(ref_1_refreshed_0_5_), .A2(
        ref_1_maj_161_n25), .ZN(ref_1_maj_161_n18) );
  NAND2_X1 ref_1_maj_161_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_161_n19) );
  NAND2_X1 ref_1_maj_161_U13 ( .A1(ref_1_maj_161_n19), .A2(ref_1_maj_161_n18), 
        .ZN(ref_1_maj_161_n22) );
  NAND2_X1 ref_1_maj_161_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_161_n24), .ZN(
        ref_1_maj_161_n20) );
  NAND2_X1 ref_1_maj_161_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_161_n21) );
  NAND2_X1 ref_1_maj_161_U10 ( .A1(ref_1_maj_161_n21), .A2(ref_1_maj_161_n20), 
        .ZN(ref_1_maj_161_n23) );
  XOR2_X1 ref_1_maj_161_U9 ( .A(ref_1_n65), .B(ref_1_maj_161_n24), .Z(
        ref_1_maj_161_n26) );
  XOR2_X1 ref_1_maj_161_U8 ( .A(ref_1_refreshed_0_5_), .B(ref_1_maj_161_n25), 
        .Z(ref_1_maj_161_n27) );
  XOR2_X1 ref_1_maj_161_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_161_n24) );
  XOR2_X1 ref_1_maj_161_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_161_n25) );
  OR2_X1 ref_1_maj_161_U5 ( .A1(ref_1_maj_161_n23), .A2(ref_1_maj_161_n22), 
        .ZN(ref_1_maj_161_n32) );
  NAND2_X1 ref_1_maj_161_U4 ( .A1(ref_1_maj_161_n22), .A2(ref_1_maj_161_n23), 
        .ZN(ref_1_maj_161_n34) );
  NAND2_X1 ref_1_maj_161_U3 ( .A1(ref_1_maj_161_n32), .A2(ref_1_maj_161_n31), 
        .ZN(ref_1_maj_161_n33) );
  NAND2_X1 ref_1_maj_161_U2 ( .A1(ref_1_maj_161_n34), .A2(ref_1_maj_161_n33), 
        .ZN(ref_1_maj_161_port_o) );
  OR2_X1 ref_1_maj_162_U19 ( .A1(ref_1_maj_162_n27), .A2(ref_1_maj_162_n26), 
        .ZN(ref_1_maj_162_n28) );
  NAND2_X1 ref_1_maj_162_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_162_n28), .ZN(
        ref_1_maj_162_n29) );
  NAND2_X1 ref_1_maj_162_U17 ( .A1(ref_1_maj_162_n26), .A2(ref_1_maj_162_n27), 
        .ZN(ref_1_maj_162_n30) );
  NAND2_X1 ref_1_maj_162_U16 ( .A1(ref_1_maj_162_n30), .A2(ref_1_maj_162_n29), 
        .ZN(ref_1_maj_162_n31) );
  NAND2_X1 ref_1_maj_162_U15 ( .A1(ref_1_refreshed_0_5_), .A2(
        ref_1_maj_162_n25), .ZN(ref_1_maj_162_n18) );
  NAND2_X1 ref_1_maj_162_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_162_n19) );
  NAND2_X1 ref_1_maj_162_U13 ( .A1(ref_1_maj_162_n19), .A2(ref_1_maj_162_n18), 
        .ZN(ref_1_maj_162_n22) );
  NAND2_X1 ref_1_maj_162_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_162_n24), .ZN(
        ref_1_maj_162_n20) );
  NAND2_X1 ref_1_maj_162_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_162_n21) );
  NAND2_X1 ref_1_maj_162_U10 ( .A1(ref_1_maj_162_n21), .A2(ref_1_maj_162_n20), 
        .ZN(ref_1_maj_162_n23) );
  XOR2_X1 ref_1_maj_162_U9 ( .A(ref_1_n65), .B(ref_1_maj_162_n24), .Z(
        ref_1_maj_162_n26) );
  XOR2_X1 ref_1_maj_162_U8 ( .A(ref_1_refreshed_0_5_), .B(ref_1_maj_162_n25), 
        .Z(ref_1_maj_162_n27) );
  XOR2_X1 ref_1_maj_162_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_162_n24) );
  XOR2_X1 ref_1_maj_162_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_162_n25) );
  OR2_X1 ref_1_maj_162_U5 ( .A1(ref_1_maj_162_n23), .A2(ref_1_maj_162_n22), 
        .ZN(ref_1_maj_162_n32) );
  NAND2_X1 ref_1_maj_162_U4 ( .A1(ref_1_maj_162_n22), .A2(ref_1_maj_162_n23), 
        .ZN(ref_1_maj_162_n34) );
  NAND2_X1 ref_1_maj_162_U3 ( .A1(ref_1_maj_162_n32), .A2(ref_1_maj_162_n31), 
        .ZN(ref_1_maj_162_n33) );
  NAND2_X1 ref_1_maj_162_U2 ( .A1(ref_1_maj_162_n34), .A2(ref_1_maj_162_n33), 
        .ZN(ref_1_maj_162_port_o) );
  OR2_X1 ref_1_maj_163_U19 ( .A1(ref_1_maj_163_n27), .A2(ref_1_maj_163_n26), 
        .ZN(ref_1_maj_163_n28) );
  NAND2_X1 ref_1_maj_163_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_163_n28), .ZN(
        ref_1_maj_163_n29) );
  NAND2_X1 ref_1_maj_163_U17 ( .A1(ref_1_maj_163_n26), .A2(ref_1_maj_163_n27), 
        .ZN(ref_1_maj_163_n30) );
  NAND2_X1 ref_1_maj_163_U16 ( .A1(ref_1_maj_163_n30), .A2(ref_1_maj_163_n29), 
        .ZN(ref_1_maj_163_n31) );
  NAND2_X1 ref_1_maj_163_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_163_n25), .ZN(
        ref_1_maj_163_n18) );
  NAND2_X1 ref_1_maj_163_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_163_n19) );
  NAND2_X1 ref_1_maj_163_U13 ( .A1(ref_1_maj_163_n19), .A2(ref_1_maj_163_n18), 
        .ZN(ref_1_maj_163_n22) );
  NAND2_X1 ref_1_maj_163_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_163_n24), .ZN(
        ref_1_maj_163_n20) );
  NAND2_X1 ref_1_maj_163_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_163_n21) );
  NAND2_X1 ref_1_maj_163_U10 ( .A1(ref_1_maj_163_n21), .A2(ref_1_maj_163_n20), 
        .ZN(ref_1_maj_163_n23) );
  XOR2_X1 ref_1_maj_163_U9 ( .A(ref_1_n66), .B(ref_1_maj_163_n24), .Z(
        ref_1_maj_163_n26) );
  XOR2_X1 ref_1_maj_163_U8 ( .A(ref_1_n74), .B(ref_1_maj_163_n25), .Z(
        ref_1_maj_163_n27) );
  XOR2_X1 ref_1_maj_163_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_163_n24) );
  XOR2_X1 ref_1_maj_163_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_163_n25) );
  OR2_X1 ref_1_maj_163_U5 ( .A1(ref_1_maj_163_n23), .A2(ref_1_maj_163_n22), 
        .ZN(ref_1_maj_163_n32) );
  NAND2_X1 ref_1_maj_163_U4 ( .A1(ref_1_maj_163_n22), .A2(ref_1_maj_163_n23), 
        .ZN(ref_1_maj_163_n34) );
  NAND2_X1 ref_1_maj_163_U3 ( .A1(ref_1_maj_163_n32), .A2(ref_1_maj_163_n31), 
        .ZN(ref_1_maj_163_n33) );
  NAND2_X1 ref_1_maj_163_U2 ( .A1(ref_1_maj_163_n34), .A2(ref_1_maj_163_n33), 
        .ZN(ref_1_maj_163_port_o) );
  OR2_X1 ref_1_maj_164_U19 ( .A1(ref_1_maj_164_n27), .A2(ref_1_maj_164_n26), 
        .ZN(ref_1_maj_164_n28) );
  NAND2_X1 ref_1_maj_164_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_164_n28), .ZN(
        ref_1_maj_164_n29) );
  NAND2_X1 ref_1_maj_164_U17 ( .A1(ref_1_maj_164_n26), .A2(ref_1_maj_164_n27), 
        .ZN(ref_1_maj_164_n30) );
  NAND2_X1 ref_1_maj_164_U16 ( .A1(ref_1_maj_164_n30), .A2(ref_1_maj_164_n29), 
        .ZN(ref_1_maj_164_n31) );
  NAND2_X1 ref_1_maj_164_U15 ( .A1(ref_1_refreshed_1_5_), .A2(
        ref_1_maj_164_n25), .ZN(ref_1_maj_164_n18) );
  NAND2_X1 ref_1_maj_164_U14 ( .A1(ref_1_refreshed_1_3_), .A2(ref_1_n52), .ZN(
        ref_1_maj_164_n19) );
  NAND2_X1 ref_1_maj_164_U13 ( .A1(ref_1_maj_164_n19), .A2(ref_1_maj_164_n18), 
        .ZN(ref_1_maj_164_n22) );
  NAND2_X1 ref_1_maj_164_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_164_n24), .ZN(
        ref_1_maj_164_n20) );
  NAND2_X1 ref_1_maj_164_U11 ( .A1(ref_1_refreshed_1_0_), .A2(ref_1_n43), .ZN(
        ref_1_maj_164_n21) );
  NAND2_X1 ref_1_maj_164_U10 ( .A1(ref_1_maj_164_n21), .A2(ref_1_maj_164_n20), 
        .ZN(ref_1_maj_164_n23) );
  XOR2_X1 ref_1_maj_164_U9 ( .A(ref_1_n46), .B(ref_1_maj_164_n24), .Z(
        ref_1_maj_164_n26) );
  XOR2_X1 ref_1_maj_164_U8 ( .A(ref_1_refreshed_1_5_), .B(ref_1_maj_164_n25), 
        .Z(ref_1_maj_164_n27) );
  XOR2_X1 ref_1_maj_164_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_n43), .Z(
        ref_1_maj_164_n24) );
  XOR2_X1 ref_1_maj_164_U6 ( .A(ref_1_refreshed_1_3_), .B(ref_1_n52), .Z(
        ref_1_maj_164_n25) );
  OR2_X1 ref_1_maj_164_U5 ( .A1(ref_1_maj_164_n23), .A2(ref_1_maj_164_n22), 
        .ZN(ref_1_maj_164_n32) );
  NAND2_X1 ref_1_maj_164_U4 ( .A1(ref_1_maj_164_n22), .A2(ref_1_maj_164_n23), 
        .ZN(ref_1_maj_164_n34) );
  NAND2_X1 ref_1_maj_164_U3 ( .A1(ref_1_maj_164_n32), .A2(ref_1_maj_164_n31), 
        .ZN(ref_1_maj_164_n33) );
  NAND2_X1 ref_1_maj_164_U2 ( .A1(ref_1_maj_164_n34), .A2(ref_1_maj_164_n33), 
        .ZN(ref_1_maj_164_port_o) );
  OR2_X1 ref_1_maj_165_U19 ( .A1(ref_1_maj_165_n27), .A2(ref_1_maj_165_n26), 
        .ZN(ref_1_maj_165_n28) );
  NAND2_X1 ref_1_maj_165_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_165_n28), .ZN(
        ref_1_maj_165_n29) );
  NAND2_X1 ref_1_maj_165_U17 ( .A1(ref_1_maj_165_n26), .A2(ref_1_maj_165_n27), 
        .ZN(ref_1_maj_165_n30) );
  NAND2_X1 ref_1_maj_165_U16 ( .A1(ref_1_maj_165_n30), .A2(ref_1_maj_165_n29), 
        .ZN(ref_1_maj_165_n31) );
  NAND2_X1 ref_1_maj_165_U15 ( .A1(ref_1_refreshed_1_5_), .A2(
        ref_1_maj_165_n25), .ZN(ref_1_maj_165_n18) );
  NAND2_X1 ref_1_maj_165_U14 ( .A1(ref_1_refreshed_1_3_), .A2(ref_1_n52), .ZN(
        ref_1_maj_165_n19) );
  NAND2_X1 ref_1_maj_165_U13 ( .A1(ref_1_maj_165_n19), .A2(ref_1_maj_165_n18), 
        .ZN(ref_1_maj_165_n22) );
  NAND2_X1 ref_1_maj_165_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_165_n24), .ZN(
        ref_1_maj_165_n20) );
  NAND2_X1 ref_1_maj_165_U11 ( .A1(ref_1_refreshed_1_0_), .A2(ref_1_n43), .ZN(
        ref_1_maj_165_n21) );
  NAND2_X1 ref_1_maj_165_U10 ( .A1(ref_1_maj_165_n21), .A2(ref_1_maj_165_n20), 
        .ZN(ref_1_maj_165_n23) );
  XOR2_X1 ref_1_maj_165_U9 ( .A(ref_1_n46), .B(ref_1_maj_165_n24), .Z(
        ref_1_maj_165_n26) );
  XOR2_X1 ref_1_maj_165_U8 ( .A(ref_1_refreshed_1_5_), .B(ref_1_maj_165_n25), 
        .Z(ref_1_maj_165_n27) );
  XOR2_X1 ref_1_maj_165_U7 ( .A(ref_1_refreshed_1_0_), .B(ref_1_n43), .Z(
        ref_1_maj_165_n24) );
  XOR2_X1 ref_1_maj_165_U6 ( .A(ref_1_refreshed_1_3_), .B(ref_1_n52), .Z(
        ref_1_maj_165_n25) );
  OR2_X1 ref_1_maj_165_U5 ( .A1(ref_1_maj_165_n23), .A2(ref_1_maj_165_n22), 
        .ZN(ref_1_maj_165_n32) );
  NAND2_X1 ref_1_maj_165_U4 ( .A1(ref_1_maj_165_n22), .A2(ref_1_maj_165_n23), 
        .ZN(ref_1_maj_165_n34) );
  NAND2_X1 ref_1_maj_165_U3 ( .A1(ref_1_maj_165_n32), .A2(ref_1_maj_165_n31), 
        .ZN(ref_1_maj_165_n33) );
  NAND2_X1 ref_1_maj_165_U2 ( .A1(ref_1_maj_165_n34), .A2(ref_1_maj_165_n33), 
        .ZN(ref_1_maj_165_port_o) );
  OR2_X1 ref_1_maj_166_U19 ( .A1(ref_1_maj_166_n27), .A2(ref_1_maj_166_n26), 
        .ZN(ref_1_maj_166_n28) );
  NAND2_X1 ref_1_maj_166_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_166_n28), .ZN(
        ref_1_maj_166_n29) );
  NAND2_X1 ref_1_maj_166_U17 ( .A1(ref_1_maj_166_n26), .A2(ref_1_maj_166_n27), 
        .ZN(ref_1_maj_166_n30) );
  NAND2_X1 ref_1_maj_166_U16 ( .A1(ref_1_maj_166_n30), .A2(ref_1_maj_166_n29), 
        .ZN(ref_1_maj_166_n31) );
  NAND2_X1 ref_1_maj_166_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_166_n25), .ZN(
        ref_1_maj_166_n18) );
  NAND2_X1 ref_1_maj_166_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_166_n19) );
  NAND2_X1 ref_1_maj_166_U13 ( .A1(ref_1_maj_166_n19), .A2(ref_1_maj_166_n18), 
        .ZN(ref_1_maj_166_n22) );
  NAND2_X1 ref_1_maj_166_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_166_n24), .ZN(
        ref_1_maj_166_n20) );
  NAND2_X1 ref_1_maj_166_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_166_n21) );
  NAND2_X1 ref_1_maj_166_U10 ( .A1(ref_1_maj_166_n21), .A2(ref_1_maj_166_n20), 
        .ZN(ref_1_maj_166_n23) );
  XOR2_X1 ref_1_maj_166_U9 ( .A(ref_1_n47), .B(ref_1_maj_166_n24), .Z(
        ref_1_maj_166_n26) );
  XOR2_X1 ref_1_maj_166_U8 ( .A(ref_1_n55), .B(ref_1_maj_166_n25), .Z(
        ref_1_maj_166_n27) );
  XOR2_X1 ref_1_maj_166_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_166_n24) );
  XOR2_X1 ref_1_maj_166_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_166_n25) );
  OR2_X1 ref_1_maj_166_U5 ( .A1(ref_1_maj_166_n23), .A2(ref_1_maj_166_n22), 
        .ZN(ref_1_maj_166_n32) );
  NAND2_X1 ref_1_maj_166_U4 ( .A1(ref_1_maj_166_n22), .A2(ref_1_maj_166_n23), 
        .ZN(ref_1_maj_166_n34) );
  NAND2_X1 ref_1_maj_166_U3 ( .A1(ref_1_maj_166_n32), .A2(ref_1_maj_166_n31), 
        .ZN(ref_1_maj_166_n33) );
  NAND2_X1 ref_1_maj_166_U2 ( .A1(ref_1_maj_166_n34), .A2(ref_1_maj_166_n33), 
        .ZN(ref_1_maj_166_port_o) );
  OR2_X1 ref_1_maj_167_U19 ( .A1(ref_1_maj_167_n27), .A2(ref_1_maj_167_n26), 
        .ZN(ref_1_maj_167_n28) );
  NAND2_X1 ref_1_maj_167_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_167_n28), .ZN(
        ref_1_maj_167_n29) );
  NAND2_X1 ref_1_maj_167_U17 ( .A1(ref_1_maj_167_n26), .A2(ref_1_maj_167_n27), 
        .ZN(ref_1_maj_167_n30) );
  NAND2_X1 ref_1_maj_167_U16 ( .A1(ref_1_maj_167_n30), .A2(ref_1_maj_167_n29), 
        .ZN(ref_1_maj_167_n31) );
  NAND2_X1 ref_1_maj_167_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_167_n25), .ZN(
        ref_1_maj_167_n18) );
  NAND2_X1 ref_1_maj_167_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_167_n19) );
  NAND2_X1 ref_1_maj_167_U13 ( .A1(ref_1_maj_167_n19), .A2(ref_1_maj_167_n18), 
        .ZN(ref_1_maj_167_n22) );
  NAND2_X1 ref_1_maj_167_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_167_n24), .ZN(
        ref_1_maj_167_n20) );
  NAND2_X1 ref_1_maj_167_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_167_n21) );
  NAND2_X1 ref_1_maj_167_U10 ( .A1(ref_1_maj_167_n21), .A2(ref_1_maj_167_n20), 
        .ZN(ref_1_maj_167_n23) );
  XOR2_X1 ref_1_maj_167_U9 ( .A(ref_1_n47), .B(ref_1_maj_167_n24), .Z(
        ref_1_maj_167_n26) );
  XOR2_X1 ref_1_maj_167_U8 ( .A(ref_1_n55), .B(ref_1_maj_167_n25), .Z(
        ref_1_maj_167_n27) );
  XOR2_X1 ref_1_maj_167_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_167_n24) );
  XOR2_X1 ref_1_maj_167_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_167_n25) );
  OR2_X1 ref_1_maj_167_U5 ( .A1(ref_1_maj_167_n23), .A2(ref_1_maj_167_n22), 
        .ZN(ref_1_maj_167_n32) );
  NAND2_X1 ref_1_maj_167_U4 ( .A1(ref_1_maj_167_n22), .A2(ref_1_maj_167_n23), 
        .ZN(ref_1_maj_167_n34) );
  NAND2_X1 ref_1_maj_167_U3 ( .A1(ref_1_maj_167_n32), .A2(ref_1_maj_167_n31), 
        .ZN(ref_1_maj_167_n33) );
  NAND2_X1 ref_1_maj_167_U2 ( .A1(ref_1_maj_167_n34), .A2(ref_1_maj_167_n33), 
        .ZN(ref_1_maj_167_port_o) );
  OR2_X1 ref_1_maj_168_U19 ( .A1(ref_1_maj_168_n27), .A2(ref_1_maj_168_n26), 
        .ZN(ref_1_maj_168_n28) );
  NAND2_X1 ref_1_maj_168_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_168_n28), .ZN(
        ref_1_maj_168_n29) );
  NAND2_X1 ref_1_maj_168_U17 ( .A1(ref_1_maj_168_n26), .A2(ref_1_maj_168_n27), 
        .ZN(ref_1_maj_168_n30) );
  NAND2_X1 ref_1_maj_168_U16 ( .A1(ref_1_maj_168_n30), .A2(ref_1_maj_168_n29), 
        .ZN(ref_1_maj_168_n31) );
  NAND2_X1 ref_1_maj_168_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_168_n25), .ZN(
        ref_1_maj_168_n18) );
  NAND2_X1 ref_1_maj_168_U14 ( .A1(ref_1_n30), .A2(ref_1_refreshed_2_4_), .ZN(
        ref_1_maj_168_n19) );
  NAND2_X1 ref_1_maj_168_U13 ( .A1(ref_1_maj_168_n19), .A2(ref_1_maj_168_n18), 
        .ZN(ref_1_maj_168_n22) );
  NAND2_X1 ref_1_maj_168_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_168_n24), .ZN(
        ref_1_maj_168_n20) );
  NAND2_X1 ref_1_maj_168_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_168_n21) );
  NAND2_X1 ref_1_maj_168_U10 ( .A1(ref_1_maj_168_n21), .A2(ref_1_maj_168_n20), 
        .ZN(ref_1_maj_168_n23) );
  XOR2_X1 ref_1_maj_168_U9 ( .A(ref_1_n27), .B(ref_1_maj_168_n24), .Z(
        ref_1_maj_168_n26) );
  XOR2_X1 ref_1_maj_168_U8 ( .A(ref_1_n36), .B(ref_1_maj_168_n25), .Z(
        ref_1_maj_168_n27) );
  XOR2_X1 ref_1_maj_168_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_168_n24) );
  XOR2_X1 ref_1_maj_168_U6 ( .A(ref_1_n30), .B(ref_1_refreshed_2_4_), .Z(
        ref_1_maj_168_n25) );
  OR2_X1 ref_1_maj_168_U5 ( .A1(ref_1_maj_168_n23), .A2(ref_1_maj_168_n22), 
        .ZN(ref_1_maj_168_n32) );
  NAND2_X1 ref_1_maj_168_U4 ( .A1(ref_1_maj_168_n22), .A2(ref_1_maj_168_n23), 
        .ZN(ref_1_maj_168_n34) );
  NAND2_X1 ref_1_maj_168_U3 ( .A1(ref_1_maj_168_n32), .A2(ref_1_maj_168_n31), 
        .ZN(ref_1_maj_168_n33) );
  NAND2_X1 ref_1_maj_168_U2 ( .A1(ref_1_maj_168_n34), .A2(ref_1_maj_168_n33), 
        .ZN(ref_1_maj_168_port_o) );
  OR2_X1 ref_1_maj_169_U19 ( .A1(ref_1_maj_169_n27), .A2(ref_1_maj_169_n26), 
        .ZN(ref_1_maj_169_n28) );
  NAND2_X1 ref_1_maj_169_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_169_n28), .ZN(
        ref_1_maj_169_n29) );
  NAND2_X1 ref_1_maj_169_U17 ( .A1(ref_1_maj_169_n26), .A2(ref_1_maj_169_n27), 
        .ZN(ref_1_maj_169_n30) );
  NAND2_X1 ref_1_maj_169_U16 ( .A1(ref_1_maj_169_n30), .A2(ref_1_maj_169_n29), 
        .ZN(ref_1_maj_169_n31) );
  NAND2_X1 ref_1_maj_169_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_169_n25), .ZN(
        ref_1_maj_169_n18) );
  NAND2_X1 ref_1_maj_169_U14 ( .A1(ref_1_n30), .A2(ref_1_refreshed_2_4_), .ZN(
        ref_1_maj_169_n19) );
  NAND2_X1 ref_1_maj_169_U13 ( .A1(ref_1_maj_169_n19), .A2(ref_1_maj_169_n18), 
        .ZN(ref_1_maj_169_n22) );
  NAND2_X1 ref_1_maj_169_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_169_n24), .ZN(
        ref_1_maj_169_n20) );
  NAND2_X1 ref_1_maj_169_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_169_n21) );
  NAND2_X1 ref_1_maj_169_U10 ( .A1(ref_1_maj_169_n21), .A2(ref_1_maj_169_n20), 
        .ZN(ref_1_maj_169_n23) );
  XOR2_X1 ref_1_maj_169_U9 ( .A(ref_1_n27), .B(ref_1_maj_169_n24), .Z(
        ref_1_maj_169_n26) );
  XOR2_X1 ref_1_maj_169_U8 ( .A(ref_1_n36), .B(ref_1_maj_169_n25), .Z(
        ref_1_maj_169_n27) );
  XOR2_X1 ref_1_maj_169_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_169_n24) );
  XOR2_X1 ref_1_maj_169_U6 ( .A(ref_1_n30), .B(ref_1_refreshed_2_4_), .Z(
        ref_1_maj_169_n25) );
  OR2_X1 ref_1_maj_169_U5 ( .A1(ref_1_maj_169_n23), .A2(ref_1_maj_169_n22), 
        .ZN(ref_1_maj_169_n32) );
  NAND2_X1 ref_1_maj_169_U4 ( .A1(ref_1_maj_169_n22), .A2(ref_1_maj_169_n23), 
        .ZN(ref_1_maj_169_n34) );
  NAND2_X1 ref_1_maj_169_U3 ( .A1(ref_1_maj_169_n32), .A2(ref_1_maj_169_n31), 
        .ZN(ref_1_maj_169_n33) );
  NAND2_X1 ref_1_maj_169_U2 ( .A1(ref_1_maj_169_n34), .A2(ref_1_maj_169_n33), 
        .ZN(ref_1_maj_169_port_o) );
  OR2_X1 ref_1_maj_170_U19 ( .A1(ref_1_maj_170_n27), .A2(ref_1_maj_170_n26), 
        .ZN(ref_1_maj_170_n28) );
  NAND2_X1 ref_1_maj_170_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_170_n28), .ZN(
        ref_1_maj_170_n29) );
  NAND2_X1 ref_1_maj_170_U17 ( .A1(ref_1_maj_170_n26), .A2(ref_1_maj_170_n27), 
        .ZN(ref_1_maj_170_n30) );
  NAND2_X1 ref_1_maj_170_U16 ( .A1(ref_1_maj_170_n30), .A2(ref_1_maj_170_n29), 
        .ZN(ref_1_maj_170_n31) );
  NAND2_X1 ref_1_maj_170_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_170_n25), .ZN(
        ref_1_maj_170_n18) );
  NAND2_X1 ref_1_maj_170_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_170_n19) );
  NAND2_X1 ref_1_maj_170_U13 ( .A1(ref_1_maj_170_n19), .A2(ref_1_maj_170_n18), 
        .ZN(ref_1_maj_170_n22) );
  NAND2_X1 ref_1_maj_170_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_170_n24), .ZN(
        ref_1_maj_170_n20) );
  NAND2_X1 ref_1_maj_170_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_170_n21) );
  NAND2_X1 ref_1_maj_170_U10 ( .A1(ref_1_maj_170_n21), .A2(ref_1_maj_170_n20), 
        .ZN(ref_1_maj_170_n23) );
  XOR2_X1 ref_1_maj_170_U9 ( .A(ref_1_n28), .B(ref_1_maj_170_n24), .Z(
        ref_1_maj_170_n26) );
  XOR2_X1 ref_1_maj_170_U8 ( .A(ref_1_n37), .B(ref_1_maj_170_n25), .Z(
        ref_1_maj_170_n27) );
  XOR2_X1 ref_1_maj_170_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_170_n24) );
  XOR2_X1 ref_1_maj_170_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_170_n25) );
  OR2_X1 ref_1_maj_170_U5 ( .A1(ref_1_maj_170_n23), .A2(ref_1_maj_170_n22), 
        .ZN(ref_1_maj_170_n32) );
  NAND2_X1 ref_1_maj_170_U4 ( .A1(ref_1_maj_170_n22), .A2(ref_1_maj_170_n23), 
        .ZN(ref_1_maj_170_n34) );
  NAND2_X1 ref_1_maj_170_U3 ( .A1(ref_1_maj_170_n32), .A2(ref_1_maj_170_n31), 
        .ZN(ref_1_maj_170_n33) );
  NAND2_X1 ref_1_maj_170_U2 ( .A1(ref_1_maj_170_n34), .A2(ref_1_maj_170_n33), 
        .ZN(ref_1_maj_170_port_o) );
  OR2_X1 ref_1_maj_171_U19 ( .A1(ref_1_maj_171_n27), .A2(ref_1_maj_171_n26), 
        .ZN(ref_1_maj_171_n28) );
  NAND2_X1 ref_1_maj_171_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_171_n28), .ZN(
        ref_1_maj_171_n29) );
  NAND2_X1 ref_1_maj_171_U17 ( .A1(ref_1_maj_171_n26), .A2(ref_1_maj_171_n27), 
        .ZN(ref_1_maj_171_n30) );
  NAND2_X1 ref_1_maj_171_U16 ( .A1(ref_1_maj_171_n30), .A2(ref_1_maj_171_n29), 
        .ZN(ref_1_maj_171_n31) );
  NAND2_X1 ref_1_maj_171_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_171_n25), .ZN(
        ref_1_maj_171_n18) );
  NAND2_X1 ref_1_maj_171_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_171_n19) );
  NAND2_X1 ref_1_maj_171_U13 ( .A1(ref_1_maj_171_n19), .A2(ref_1_maj_171_n18), 
        .ZN(ref_1_maj_171_n22) );
  NAND2_X1 ref_1_maj_171_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_171_n24), .ZN(
        ref_1_maj_171_n20) );
  NAND2_X1 ref_1_maj_171_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_171_n21) );
  NAND2_X1 ref_1_maj_171_U10 ( .A1(ref_1_maj_171_n21), .A2(ref_1_maj_171_n20), 
        .ZN(ref_1_maj_171_n23) );
  XOR2_X1 ref_1_maj_171_U9 ( .A(ref_1_n28), .B(ref_1_maj_171_n24), .Z(
        ref_1_maj_171_n26) );
  XOR2_X1 ref_1_maj_171_U8 ( .A(ref_1_n37), .B(ref_1_maj_171_n25), .Z(
        ref_1_maj_171_n27) );
  XOR2_X1 ref_1_maj_171_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_171_n24) );
  XOR2_X1 ref_1_maj_171_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_171_n25) );
  OR2_X1 ref_1_maj_171_U5 ( .A1(ref_1_maj_171_n23), .A2(ref_1_maj_171_n22), 
        .ZN(ref_1_maj_171_n32) );
  NAND2_X1 ref_1_maj_171_U4 ( .A1(ref_1_maj_171_n22), .A2(ref_1_maj_171_n23), 
        .ZN(ref_1_maj_171_n34) );
  NAND2_X1 ref_1_maj_171_U3 ( .A1(ref_1_maj_171_n32), .A2(ref_1_maj_171_n31), 
        .ZN(ref_1_maj_171_n33) );
  NAND2_X1 ref_1_maj_171_U2 ( .A1(ref_1_maj_171_n34), .A2(ref_1_maj_171_n33), 
        .ZN(ref_1_maj_171_port_o) );
  OR2_X1 ref_1_maj_172_U19 ( .A1(ref_1_maj_172_n27), .A2(ref_1_maj_172_n26), 
        .ZN(ref_1_maj_172_n28) );
  NAND2_X1 ref_1_maj_172_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_172_n28), .ZN(
        ref_1_maj_172_n29) );
  NAND2_X1 ref_1_maj_172_U17 ( .A1(ref_1_maj_172_n26), .A2(ref_1_maj_172_n27), 
        .ZN(ref_1_maj_172_n30) );
  NAND2_X1 ref_1_maj_172_U16 ( .A1(ref_1_maj_172_n30), .A2(ref_1_maj_172_n29), 
        .ZN(ref_1_maj_172_n31) );
  NAND2_X1 ref_1_maj_172_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_172_n25), .ZN(
        ref_1_maj_172_n18) );
  NAND2_X1 ref_1_maj_172_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_172_n19) );
  NAND2_X1 ref_1_maj_172_U13 ( .A1(ref_1_maj_172_n19), .A2(ref_1_maj_172_n18), 
        .ZN(ref_1_maj_172_n22) );
  NAND2_X1 ref_1_maj_172_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_172_n24), .ZN(
        ref_1_maj_172_n20) );
  NAND2_X1 ref_1_maj_172_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_172_n21) );
  NAND2_X1 ref_1_maj_172_U10 ( .A1(ref_1_maj_172_n21), .A2(ref_1_maj_172_n20), 
        .ZN(ref_1_maj_172_n23) );
  XOR2_X1 ref_1_maj_172_U9 ( .A(ref_1_n8), .B(ref_1_maj_172_n24), .Z(
        ref_1_maj_172_n26) );
  XOR2_X1 ref_1_maj_172_U8 ( .A(ref_1_n17), .B(ref_1_maj_172_n25), .Z(
        ref_1_maj_172_n27) );
  XOR2_X1 ref_1_maj_172_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_172_n24)
         );
  XOR2_X1 ref_1_maj_172_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_172_n25) );
  OR2_X1 ref_1_maj_172_U5 ( .A1(ref_1_maj_172_n23), .A2(ref_1_maj_172_n22), 
        .ZN(ref_1_maj_172_n32) );
  NAND2_X1 ref_1_maj_172_U4 ( .A1(ref_1_maj_172_n22), .A2(ref_1_maj_172_n23), 
        .ZN(ref_1_maj_172_n34) );
  NAND2_X1 ref_1_maj_172_U3 ( .A1(ref_1_maj_172_n32), .A2(ref_1_maj_172_n31), 
        .ZN(ref_1_maj_172_n33) );
  NAND2_X1 ref_1_maj_172_U2 ( .A1(ref_1_maj_172_n34), .A2(ref_1_maj_172_n33), 
        .ZN(ref_1_maj_172_port_o) );
  OR2_X1 ref_1_maj_173_U19 ( .A1(ref_1_maj_173_n27), .A2(ref_1_maj_173_n26), 
        .ZN(ref_1_maj_173_n28) );
  NAND2_X1 ref_1_maj_173_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_173_n28), .ZN(
        ref_1_maj_173_n29) );
  NAND2_X1 ref_1_maj_173_U17 ( .A1(ref_1_maj_173_n26), .A2(ref_1_maj_173_n27), 
        .ZN(ref_1_maj_173_n30) );
  NAND2_X1 ref_1_maj_173_U16 ( .A1(ref_1_maj_173_n30), .A2(ref_1_maj_173_n29), 
        .ZN(ref_1_maj_173_n31) );
  NAND2_X1 ref_1_maj_173_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_173_n25), .ZN(
        ref_1_maj_173_n18) );
  NAND2_X1 ref_1_maj_173_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_173_n19) );
  NAND2_X1 ref_1_maj_173_U13 ( .A1(ref_1_maj_173_n19), .A2(ref_1_maj_173_n18), 
        .ZN(ref_1_maj_173_n22) );
  NAND2_X1 ref_1_maj_173_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_173_n24), .ZN(
        ref_1_maj_173_n20) );
  NAND2_X1 ref_1_maj_173_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_173_n21) );
  NAND2_X1 ref_1_maj_173_U10 ( .A1(ref_1_maj_173_n21), .A2(ref_1_maj_173_n20), 
        .ZN(ref_1_maj_173_n23) );
  XOR2_X1 ref_1_maj_173_U9 ( .A(ref_1_n8), .B(ref_1_maj_173_n24), .Z(
        ref_1_maj_173_n26) );
  XOR2_X1 ref_1_maj_173_U8 ( .A(ref_1_n17), .B(ref_1_maj_173_n25), .Z(
        ref_1_maj_173_n27) );
  XOR2_X1 ref_1_maj_173_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_173_n24)
         );
  XOR2_X1 ref_1_maj_173_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_173_n25) );
  OR2_X1 ref_1_maj_173_U5 ( .A1(ref_1_maj_173_n23), .A2(ref_1_maj_173_n22), 
        .ZN(ref_1_maj_173_n32) );
  NAND2_X1 ref_1_maj_173_U4 ( .A1(ref_1_maj_173_n22), .A2(ref_1_maj_173_n23), 
        .ZN(ref_1_maj_173_n34) );
  NAND2_X1 ref_1_maj_173_U3 ( .A1(ref_1_maj_173_n32), .A2(ref_1_maj_173_n31), 
        .ZN(ref_1_maj_173_n33) );
  NAND2_X1 ref_1_maj_173_U2 ( .A1(ref_1_maj_173_n34), .A2(ref_1_maj_173_n33), 
        .ZN(ref_1_maj_173_port_o) );
  OR2_X1 ref_1_maj_174_U19 ( .A1(ref_1_maj_174_n27), .A2(ref_1_maj_174_n26), 
        .ZN(ref_1_maj_174_n28) );
  NAND2_X1 ref_1_maj_174_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_174_n28), .ZN(
        ref_1_maj_174_n29) );
  NAND2_X1 ref_1_maj_174_U17 ( .A1(ref_1_maj_174_n26), .A2(ref_1_maj_174_n27), 
        .ZN(ref_1_maj_174_n30) );
  NAND2_X1 ref_1_maj_174_U16 ( .A1(ref_1_maj_174_n30), .A2(ref_1_maj_174_n29), 
        .ZN(ref_1_maj_174_n31) );
  NAND2_X1 ref_1_maj_174_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_174_n25), .ZN(
        ref_1_maj_174_n18) );
  NAND2_X1 ref_1_maj_174_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_174_n19) );
  NAND2_X1 ref_1_maj_174_U13 ( .A1(ref_1_maj_174_n19), .A2(ref_1_maj_174_n18), 
        .ZN(ref_1_maj_174_n22) );
  NAND2_X1 ref_1_maj_174_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_174_n24), .ZN(
        ref_1_maj_174_n20) );
  NAND2_X1 ref_1_maj_174_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_174_n21) );
  NAND2_X1 ref_1_maj_174_U10 ( .A1(ref_1_maj_174_n21), .A2(ref_1_maj_174_n20), 
        .ZN(ref_1_maj_174_n23) );
  XOR2_X1 ref_1_maj_174_U9 ( .A(ref_1_n9), .B(ref_1_maj_174_n24), .Z(
        ref_1_maj_174_n26) );
  XOR2_X1 ref_1_maj_174_U8 ( .A(ref_1_n18), .B(ref_1_maj_174_n25), .Z(
        ref_1_maj_174_n27) );
  XOR2_X1 ref_1_maj_174_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_174_n24)
         );
  XOR2_X1 ref_1_maj_174_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_174_n25) );
  OR2_X1 ref_1_maj_174_U5 ( .A1(ref_1_maj_174_n23), .A2(ref_1_maj_174_n22), 
        .ZN(ref_1_maj_174_n32) );
  NAND2_X1 ref_1_maj_174_U4 ( .A1(ref_1_maj_174_n22), .A2(ref_1_maj_174_n23), 
        .ZN(ref_1_maj_174_n34) );
  NAND2_X1 ref_1_maj_174_U3 ( .A1(ref_1_maj_174_n32), .A2(ref_1_maj_174_n31), 
        .ZN(ref_1_maj_174_n33) );
  NAND2_X1 ref_1_maj_174_U2 ( .A1(ref_1_maj_174_n34), .A2(ref_1_maj_174_n33), 
        .ZN(ref_1_maj_174_port_o) );
  OR2_X1 ref_1_maj_175_U19 ( .A1(ref_1_maj_175_n27), .A2(ref_1_maj_175_n26), 
        .ZN(ref_1_maj_175_n28) );
  NAND2_X1 ref_1_maj_175_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_175_n28), .ZN(
        ref_1_maj_175_n29) );
  NAND2_X1 ref_1_maj_175_U17 ( .A1(ref_1_maj_175_n26), .A2(ref_1_maj_175_n27), 
        .ZN(ref_1_maj_175_n30) );
  NAND2_X1 ref_1_maj_175_U16 ( .A1(ref_1_maj_175_n30), .A2(ref_1_maj_175_n29), 
        .ZN(ref_1_maj_175_n31) );
  NAND2_X1 ref_1_maj_175_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_175_n25), .ZN(
        ref_1_maj_175_n18) );
  NAND2_X1 ref_1_maj_175_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_175_n19) );
  NAND2_X1 ref_1_maj_175_U13 ( .A1(ref_1_maj_175_n19), .A2(ref_1_maj_175_n18), 
        .ZN(ref_1_maj_175_n22) );
  NAND2_X1 ref_1_maj_175_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_175_n24), .ZN(
        ref_1_maj_175_n20) );
  NAND2_X1 ref_1_maj_175_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_175_n21) );
  NAND2_X1 ref_1_maj_175_U10 ( .A1(ref_1_maj_175_n21), .A2(ref_1_maj_175_n20), 
        .ZN(ref_1_maj_175_n23) );
  XOR2_X1 ref_1_maj_175_U9 ( .A(ref_1_n9), .B(ref_1_maj_175_n24), .Z(
        ref_1_maj_175_n26) );
  XOR2_X1 ref_1_maj_175_U8 ( .A(ref_1_n18), .B(ref_1_maj_175_n25), .Z(
        ref_1_maj_175_n27) );
  XOR2_X1 ref_1_maj_175_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_175_n24)
         );
  XOR2_X1 ref_1_maj_175_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_175_n25) );
  OR2_X1 ref_1_maj_175_U5 ( .A1(ref_1_maj_175_n23), .A2(ref_1_maj_175_n22), 
        .ZN(ref_1_maj_175_n32) );
  NAND2_X1 ref_1_maj_175_U4 ( .A1(ref_1_maj_175_n22), .A2(ref_1_maj_175_n23), 
        .ZN(ref_1_maj_175_n34) );
  NAND2_X1 ref_1_maj_175_U3 ( .A1(ref_1_maj_175_n32), .A2(ref_1_maj_175_n31), 
        .ZN(ref_1_maj_175_n33) );
  NAND2_X1 ref_1_maj_175_U2 ( .A1(ref_1_maj_175_n34), .A2(ref_1_maj_175_n33), 
        .ZN(ref_1_maj_175_port_o) );
  OR2_X1 ref_1_maj_176_U19 ( .A1(ref_1_maj_176_n27), .A2(ref_1_maj_176_n26), 
        .ZN(ref_1_maj_176_n28) );
  NAND2_X1 ref_1_maj_176_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_176_n28), .ZN(
        ref_1_maj_176_n29) );
  NAND2_X1 ref_1_maj_176_U17 ( .A1(ref_1_maj_176_n26), .A2(ref_1_maj_176_n27), 
        .ZN(ref_1_maj_176_n30) );
  NAND2_X1 ref_1_maj_176_U16 ( .A1(ref_1_maj_176_n30), .A2(ref_1_maj_176_n29), 
        .ZN(ref_1_maj_176_n31) );
  NAND2_X1 ref_1_maj_176_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_176_n25), .ZN(
        ref_1_maj_176_n18) );
  NAND2_X1 ref_1_maj_176_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_176_n19) );
  NAND2_X1 ref_1_maj_176_U13 ( .A1(ref_1_maj_176_n19), .A2(ref_1_maj_176_n18), 
        .ZN(ref_1_maj_176_n22) );
  NAND2_X1 ref_1_maj_176_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_176_n24), .ZN(
        ref_1_maj_176_n20) );
  NAND2_X1 ref_1_maj_176_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_176_n21) );
  NAND2_X1 ref_1_maj_176_U10 ( .A1(ref_1_maj_176_n21), .A2(ref_1_maj_176_n20), 
        .ZN(ref_1_maj_176_n23) );
  XOR2_X1 ref_1_maj_176_U9 ( .A(ref_1_n66), .B(ref_1_maj_176_n24), .Z(
        ref_1_maj_176_n26) );
  XOR2_X1 ref_1_maj_176_U8 ( .A(ref_1_n74), .B(ref_1_maj_176_n25), .Z(
        ref_1_maj_176_n27) );
  XOR2_X1 ref_1_maj_176_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_176_n24) );
  XOR2_X1 ref_1_maj_176_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_176_n25) );
  OR2_X1 ref_1_maj_176_U5 ( .A1(ref_1_maj_176_n23), .A2(ref_1_maj_176_n22), 
        .ZN(ref_1_maj_176_n32) );
  NAND2_X1 ref_1_maj_176_U4 ( .A1(ref_1_maj_176_n22), .A2(ref_1_maj_176_n23), 
        .ZN(ref_1_maj_176_n34) );
  NAND2_X1 ref_1_maj_176_U3 ( .A1(ref_1_maj_176_n32), .A2(ref_1_maj_176_n31), 
        .ZN(ref_1_maj_176_n33) );
  NAND2_X1 ref_1_maj_176_U2 ( .A1(ref_1_maj_176_n34), .A2(ref_1_maj_176_n33), 
        .ZN(ref_1_maj_176_port_o) );
  OR2_X1 ref_1_maj_177_U19 ( .A1(ref_1_maj_177_n27), .A2(ref_1_maj_177_n26), 
        .ZN(ref_1_maj_177_n28) );
  NAND2_X1 ref_1_maj_177_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_177_n28), .ZN(
        ref_1_maj_177_n29) );
  NAND2_X1 ref_1_maj_177_U17 ( .A1(ref_1_maj_177_n26), .A2(ref_1_maj_177_n27), 
        .ZN(ref_1_maj_177_n30) );
  NAND2_X1 ref_1_maj_177_U16 ( .A1(ref_1_maj_177_n30), .A2(ref_1_maj_177_n29), 
        .ZN(ref_1_maj_177_n31) );
  NAND2_X1 ref_1_maj_177_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_177_n25), .ZN(
        ref_1_maj_177_n18) );
  NAND2_X1 ref_1_maj_177_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_177_n19) );
  NAND2_X1 ref_1_maj_177_U13 ( .A1(ref_1_maj_177_n19), .A2(ref_1_maj_177_n18), 
        .ZN(ref_1_maj_177_n22) );
  NAND2_X1 ref_1_maj_177_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_177_n24), .ZN(
        ref_1_maj_177_n20) );
  NAND2_X1 ref_1_maj_177_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_177_n21) );
  NAND2_X1 ref_1_maj_177_U10 ( .A1(ref_1_maj_177_n21), .A2(ref_1_maj_177_n20), 
        .ZN(ref_1_maj_177_n23) );
  XOR2_X1 ref_1_maj_177_U9 ( .A(ref_1_n66), .B(ref_1_maj_177_n24), .Z(
        ref_1_maj_177_n26) );
  XOR2_X1 ref_1_maj_177_U8 ( .A(ref_1_n74), .B(ref_1_maj_177_n25), .Z(
        ref_1_maj_177_n27) );
  XOR2_X1 ref_1_maj_177_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_177_n24) );
  XOR2_X1 ref_1_maj_177_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_177_n25) );
  OR2_X1 ref_1_maj_177_U5 ( .A1(ref_1_maj_177_n23), .A2(ref_1_maj_177_n22), 
        .ZN(ref_1_maj_177_n32) );
  NAND2_X1 ref_1_maj_177_U4 ( .A1(ref_1_maj_177_n22), .A2(ref_1_maj_177_n23), 
        .ZN(ref_1_maj_177_n34) );
  NAND2_X1 ref_1_maj_177_U3 ( .A1(ref_1_maj_177_n32), .A2(ref_1_maj_177_n31), 
        .ZN(ref_1_maj_177_n33) );
  NAND2_X1 ref_1_maj_177_U2 ( .A1(ref_1_maj_177_n34), .A2(ref_1_maj_177_n33), 
        .ZN(ref_1_maj_177_port_o) );
  OR2_X1 ref_1_maj_178_U19 ( .A1(ref_1_maj_178_n27), .A2(ref_1_maj_178_n26), 
        .ZN(ref_1_maj_178_n28) );
  NAND2_X1 ref_1_maj_178_U18 ( .A1(ref_1_n76), .A2(ref_1_maj_178_n28), .ZN(
        ref_1_maj_178_n29) );
  NAND2_X1 ref_1_maj_178_U17 ( .A1(ref_1_maj_178_n26), .A2(ref_1_maj_178_n27), 
        .ZN(ref_1_maj_178_n30) );
  NAND2_X1 ref_1_maj_178_U16 ( .A1(ref_1_maj_178_n30), .A2(ref_1_maj_178_n29), 
        .ZN(ref_1_maj_178_n31) );
  NAND2_X1 ref_1_maj_178_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_178_n25), .ZN(
        ref_1_maj_178_n18) );
  NAND2_X1 ref_1_maj_178_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_178_n19) );
  NAND2_X1 ref_1_maj_178_U13 ( .A1(ref_1_maj_178_n19), .A2(ref_1_maj_178_n18), 
        .ZN(ref_1_maj_178_n22) );
  NAND2_X1 ref_1_maj_178_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_178_n24), .ZN(
        ref_1_maj_178_n20) );
  NAND2_X1 ref_1_maj_178_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_178_n21) );
  NAND2_X1 ref_1_maj_178_U10 ( .A1(ref_1_maj_178_n21), .A2(ref_1_maj_178_n20), 
        .ZN(ref_1_maj_178_n23) );
  XOR2_X1 ref_1_maj_178_U9 ( .A(ref_1_n66), .B(ref_1_maj_178_n24), .Z(
        ref_1_maj_178_n26) );
  XOR2_X1 ref_1_maj_178_U8 ( .A(ref_1_n74), .B(ref_1_maj_178_n25), .Z(
        ref_1_maj_178_n27) );
  XOR2_X1 ref_1_maj_178_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_178_n24) );
  XOR2_X1 ref_1_maj_178_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_178_n25) );
  OR2_X1 ref_1_maj_178_U5 ( .A1(ref_1_maj_178_n23), .A2(ref_1_maj_178_n22), 
        .ZN(ref_1_maj_178_n32) );
  NAND2_X1 ref_1_maj_178_U4 ( .A1(ref_1_maj_178_n22), .A2(ref_1_maj_178_n23), 
        .ZN(ref_1_maj_178_n34) );
  NAND2_X1 ref_1_maj_178_U3 ( .A1(ref_1_maj_178_n32), .A2(ref_1_maj_178_n31), 
        .ZN(ref_1_maj_178_n33) );
  NAND2_X1 ref_1_maj_178_U2 ( .A1(ref_1_maj_178_n34), .A2(ref_1_maj_178_n33), 
        .ZN(ref_1_maj_178_port_o) );
  OR2_X1 ref_1_maj_179_U19 ( .A1(ref_1_maj_179_n27), .A2(ref_1_maj_179_n26), 
        .ZN(ref_1_maj_179_n28) );
  NAND2_X1 ref_1_maj_179_U18 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_179_n28), .ZN(ref_1_maj_179_n29) );
  NAND2_X1 ref_1_maj_179_U17 ( .A1(ref_1_maj_179_n26), .A2(ref_1_maj_179_n27), 
        .ZN(ref_1_maj_179_n30) );
  NAND2_X1 ref_1_maj_179_U16 ( .A1(ref_1_maj_179_n30), .A2(ref_1_maj_179_n29), 
        .ZN(ref_1_maj_179_n31) );
  NAND2_X1 ref_1_maj_179_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_179_n25), .ZN(
        ref_1_maj_179_n18) );
  NAND2_X1 ref_1_maj_179_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_179_n19) );
  NAND2_X1 ref_1_maj_179_U13 ( .A1(ref_1_maj_179_n19), .A2(ref_1_maj_179_n18), 
        .ZN(ref_1_maj_179_n22) );
  NAND2_X1 ref_1_maj_179_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_179_n24), .ZN(
        ref_1_maj_179_n20) );
  NAND2_X1 ref_1_maj_179_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_179_n21) );
  NAND2_X1 ref_1_maj_179_U10 ( .A1(ref_1_maj_179_n21), .A2(ref_1_maj_179_n20), 
        .ZN(ref_1_maj_179_n23) );
  XOR2_X1 ref_1_maj_179_U9 ( .A(ref_1_n66), .B(ref_1_maj_179_n24), .Z(
        ref_1_maj_179_n26) );
  XOR2_X1 ref_1_maj_179_U8 ( .A(ref_1_n74), .B(ref_1_maj_179_n25), .Z(
        ref_1_maj_179_n27) );
  XOR2_X1 ref_1_maj_179_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_179_n24) );
  XOR2_X1 ref_1_maj_179_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_179_n25) );
  OR2_X1 ref_1_maj_179_U5 ( .A1(ref_1_maj_179_n23), .A2(ref_1_maj_179_n22), 
        .ZN(ref_1_maj_179_n32) );
  NAND2_X1 ref_1_maj_179_U4 ( .A1(ref_1_maj_179_n22), .A2(ref_1_maj_179_n23), 
        .ZN(ref_1_maj_179_n34) );
  NAND2_X1 ref_1_maj_179_U3 ( .A1(ref_1_maj_179_n32), .A2(ref_1_maj_179_n31), 
        .ZN(ref_1_maj_179_n33) );
  NAND2_X1 ref_1_maj_179_U2 ( .A1(ref_1_maj_179_n34), .A2(ref_1_maj_179_n33), 
        .ZN(ref_1_maj_179_port_o) );
  OR2_X1 ref_1_maj_180_U19 ( .A1(ref_1_maj_180_n27), .A2(ref_1_maj_180_n26), 
        .ZN(ref_1_maj_180_n28) );
  NAND2_X1 ref_1_maj_180_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_180_n28), .ZN(
        ref_1_maj_180_n29) );
  NAND2_X1 ref_1_maj_180_U17 ( .A1(ref_1_maj_180_n26), .A2(ref_1_maj_180_n27), 
        .ZN(ref_1_maj_180_n30) );
  NAND2_X1 ref_1_maj_180_U16 ( .A1(ref_1_maj_180_n30), .A2(ref_1_maj_180_n29), 
        .ZN(ref_1_maj_180_n31) );
  NAND2_X1 ref_1_maj_180_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_180_n25), .ZN(
        ref_1_maj_180_n18) );
  NAND2_X1 ref_1_maj_180_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_180_n19) );
  NAND2_X1 ref_1_maj_180_U13 ( .A1(ref_1_maj_180_n19), .A2(ref_1_maj_180_n18), 
        .ZN(ref_1_maj_180_n22) );
  NAND2_X1 ref_1_maj_180_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_180_n24), .ZN(
        ref_1_maj_180_n20) );
  NAND2_X1 ref_1_maj_180_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_180_n21) );
  NAND2_X1 ref_1_maj_180_U10 ( .A1(ref_1_maj_180_n21), .A2(ref_1_maj_180_n20), 
        .ZN(ref_1_maj_180_n23) );
  XOR2_X1 ref_1_maj_180_U9 ( .A(ref_1_n47), .B(ref_1_maj_180_n24), .Z(
        ref_1_maj_180_n26) );
  XOR2_X1 ref_1_maj_180_U8 ( .A(ref_1_n55), .B(ref_1_maj_180_n25), .Z(
        ref_1_maj_180_n27) );
  XOR2_X1 ref_1_maj_180_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_180_n24) );
  XOR2_X1 ref_1_maj_180_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_180_n25) );
  OR2_X1 ref_1_maj_180_U5 ( .A1(ref_1_maj_180_n23), .A2(ref_1_maj_180_n22), 
        .ZN(ref_1_maj_180_n32) );
  NAND2_X1 ref_1_maj_180_U4 ( .A1(ref_1_maj_180_n22), .A2(ref_1_maj_180_n23), 
        .ZN(ref_1_maj_180_n34) );
  NAND2_X1 ref_1_maj_180_U3 ( .A1(ref_1_maj_180_n32), .A2(ref_1_maj_180_n31), 
        .ZN(ref_1_maj_180_n33) );
  NAND2_X1 ref_1_maj_180_U2 ( .A1(ref_1_maj_180_n34), .A2(ref_1_maj_180_n33), 
        .ZN(ref_1_maj_180_port_o) );
  OR2_X1 ref_1_maj_181_U19 ( .A1(ref_1_maj_181_n27), .A2(ref_1_maj_181_n26), 
        .ZN(ref_1_maj_181_n28) );
  NAND2_X1 ref_1_maj_181_U18 ( .A1(ref_1_n57), .A2(ref_1_maj_181_n28), .ZN(
        ref_1_maj_181_n29) );
  NAND2_X1 ref_1_maj_181_U17 ( .A1(ref_1_maj_181_n26), .A2(ref_1_maj_181_n27), 
        .ZN(ref_1_maj_181_n30) );
  NAND2_X1 ref_1_maj_181_U16 ( .A1(ref_1_maj_181_n30), .A2(ref_1_maj_181_n29), 
        .ZN(ref_1_maj_181_n31) );
  NAND2_X1 ref_1_maj_181_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_181_n25), .ZN(
        ref_1_maj_181_n18) );
  NAND2_X1 ref_1_maj_181_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_181_n19) );
  NAND2_X1 ref_1_maj_181_U13 ( .A1(ref_1_maj_181_n19), .A2(ref_1_maj_181_n18), 
        .ZN(ref_1_maj_181_n22) );
  NAND2_X1 ref_1_maj_181_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_181_n24), .ZN(
        ref_1_maj_181_n20) );
  NAND2_X1 ref_1_maj_181_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_181_n21) );
  NAND2_X1 ref_1_maj_181_U10 ( .A1(ref_1_maj_181_n21), .A2(ref_1_maj_181_n20), 
        .ZN(ref_1_maj_181_n23) );
  XOR2_X1 ref_1_maj_181_U9 ( .A(ref_1_n47), .B(ref_1_maj_181_n24), .Z(
        ref_1_maj_181_n26) );
  XOR2_X1 ref_1_maj_181_U8 ( .A(ref_1_n55), .B(ref_1_maj_181_n25), .Z(
        ref_1_maj_181_n27) );
  XOR2_X1 ref_1_maj_181_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_181_n24) );
  XOR2_X1 ref_1_maj_181_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_181_n25) );
  OR2_X1 ref_1_maj_181_U5 ( .A1(ref_1_maj_181_n23), .A2(ref_1_maj_181_n22), 
        .ZN(ref_1_maj_181_n32) );
  NAND2_X1 ref_1_maj_181_U4 ( .A1(ref_1_maj_181_n22), .A2(ref_1_maj_181_n23), 
        .ZN(ref_1_maj_181_n34) );
  NAND2_X1 ref_1_maj_181_U3 ( .A1(ref_1_maj_181_n32), .A2(ref_1_maj_181_n31), 
        .ZN(ref_1_maj_181_n33) );
  NAND2_X1 ref_1_maj_181_U2 ( .A1(ref_1_maj_181_n34), .A2(ref_1_maj_181_n33), 
        .ZN(ref_1_maj_181_port_o) );
  OR2_X1 ref_1_maj_182_U19 ( .A1(ref_1_maj_182_n27), .A2(ref_1_maj_182_n26), 
        .ZN(ref_1_maj_182_n28) );
  NAND2_X1 ref_1_maj_182_U18 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_182_n28), .ZN(ref_1_maj_182_n29) );
  NAND2_X1 ref_1_maj_182_U17 ( .A1(ref_1_maj_182_n26), .A2(ref_1_maj_182_n27), 
        .ZN(ref_1_maj_182_n30) );
  NAND2_X1 ref_1_maj_182_U16 ( .A1(ref_1_maj_182_n30), .A2(ref_1_maj_182_n29), 
        .ZN(ref_1_maj_182_n31) );
  NAND2_X1 ref_1_maj_182_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_182_n25), .ZN(
        ref_1_maj_182_n18) );
  NAND2_X1 ref_1_maj_182_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_182_n19) );
  NAND2_X1 ref_1_maj_182_U13 ( .A1(ref_1_maj_182_n19), .A2(ref_1_maj_182_n18), 
        .ZN(ref_1_maj_182_n22) );
  NAND2_X1 ref_1_maj_182_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_182_n24), .ZN(
        ref_1_maj_182_n20) );
  NAND2_X1 ref_1_maj_182_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_182_n21) );
  NAND2_X1 ref_1_maj_182_U10 ( .A1(ref_1_maj_182_n21), .A2(ref_1_maj_182_n20), 
        .ZN(ref_1_maj_182_n23) );
  XOR2_X1 ref_1_maj_182_U9 ( .A(ref_1_n47), .B(ref_1_maj_182_n24), .Z(
        ref_1_maj_182_n26) );
  XOR2_X1 ref_1_maj_182_U8 ( .A(ref_1_n55), .B(ref_1_maj_182_n25), .Z(
        ref_1_maj_182_n27) );
  XOR2_X1 ref_1_maj_182_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_182_n24) );
  XOR2_X1 ref_1_maj_182_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_182_n25) );
  OR2_X1 ref_1_maj_182_U5 ( .A1(ref_1_maj_182_n23), .A2(ref_1_maj_182_n22), 
        .ZN(ref_1_maj_182_n32) );
  NAND2_X1 ref_1_maj_182_U4 ( .A1(ref_1_maj_182_n22), .A2(ref_1_maj_182_n23), 
        .ZN(ref_1_maj_182_n34) );
  NAND2_X1 ref_1_maj_182_U3 ( .A1(ref_1_maj_182_n32), .A2(ref_1_maj_182_n31), 
        .ZN(ref_1_maj_182_n33) );
  NAND2_X1 ref_1_maj_182_U2 ( .A1(ref_1_maj_182_n34), .A2(ref_1_maj_182_n33), 
        .ZN(ref_1_maj_182_port_o) );
  OR2_X1 ref_1_maj_183_U19 ( .A1(ref_1_maj_183_n27), .A2(ref_1_maj_183_n26), 
        .ZN(ref_1_maj_183_n28) );
  NAND2_X1 ref_1_maj_183_U18 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_183_n28), .ZN(ref_1_maj_183_n29) );
  NAND2_X1 ref_1_maj_183_U17 ( .A1(ref_1_maj_183_n26), .A2(ref_1_maj_183_n27), 
        .ZN(ref_1_maj_183_n30) );
  NAND2_X1 ref_1_maj_183_U16 ( .A1(ref_1_maj_183_n30), .A2(ref_1_maj_183_n29), 
        .ZN(ref_1_maj_183_n31) );
  NAND2_X1 ref_1_maj_183_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_183_n25), .ZN(
        ref_1_maj_183_n18) );
  NAND2_X1 ref_1_maj_183_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_183_n19) );
  NAND2_X1 ref_1_maj_183_U13 ( .A1(ref_1_maj_183_n19), .A2(ref_1_maj_183_n18), 
        .ZN(ref_1_maj_183_n22) );
  NAND2_X1 ref_1_maj_183_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_183_n24), .ZN(
        ref_1_maj_183_n20) );
  NAND2_X1 ref_1_maj_183_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_183_n21) );
  NAND2_X1 ref_1_maj_183_U10 ( .A1(ref_1_maj_183_n21), .A2(ref_1_maj_183_n20), 
        .ZN(ref_1_maj_183_n23) );
  XOR2_X1 ref_1_maj_183_U9 ( .A(ref_1_n47), .B(ref_1_maj_183_n24), .Z(
        ref_1_maj_183_n26) );
  XOR2_X1 ref_1_maj_183_U8 ( .A(ref_1_n55), .B(ref_1_maj_183_n25), .Z(
        ref_1_maj_183_n27) );
  XOR2_X1 ref_1_maj_183_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_183_n24) );
  XOR2_X1 ref_1_maj_183_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_183_n25) );
  OR2_X1 ref_1_maj_183_U5 ( .A1(ref_1_maj_183_n23), .A2(ref_1_maj_183_n22), 
        .ZN(ref_1_maj_183_n32) );
  NAND2_X1 ref_1_maj_183_U4 ( .A1(ref_1_maj_183_n22), .A2(ref_1_maj_183_n23), 
        .ZN(ref_1_maj_183_n34) );
  NAND2_X1 ref_1_maj_183_U3 ( .A1(ref_1_maj_183_n32), .A2(ref_1_maj_183_n31), 
        .ZN(ref_1_maj_183_n33) );
  NAND2_X1 ref_1_maj_183_U2 ( .A1(ref_1_maj_183_n34), .A2(ref_1_maj_183_n33), 
        .ZN(ref_1_maj_183_port_o) );
  OR2_X1 ref_1_maj_184_U19 ( .A1(ref_1_maj_184_n27), .A2(ref_1_maj_184_n26), 
        .ZN(ref_1_maj_184_n28) );
  NAND2_X1 ref_1_maj_184_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_184_n28), .ZN(
        ref_1_maj_184_n29) );
  NAND2_X1 ref_1_maj_184_U17 ( .A1(ref_1_maj_184_n26), .A2(ref_1_maj_184_n27), 
        .ZN(ref_1_maj_184_n30) );
  NAND2_X1 ref_1_maj_184_U16 ( .A1(ref_1_maj_184_n30), .A2(ref_1_maj_184_n29), 
        .ZN(ref_1_maj_184_n31) );
  NAND2_X1 ref_1_maj_184_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_184_n25), .ZN(
        ref_1_maj_184_n18) );
  NAND2_X1 ref_1_maj_184_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_184_n19) );
  NAND2_X1 ref_1_maj_184_U13 ( .A1(ref_1_maj_184_n19), .A2(ref_1_maj_184_n18), 
        .ZN(ref_1_maj_184_n22) );
  NAND2_X1 ref_1_maj_184_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_184_n24), .ZN(
        ref_1_maj_184_n20) );
  NAND2_X1 ref_1_maj_184_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_184_n21) );
  NAND2_X1 ref_1_maj_184_U10 ( .A1(ref_1_maj_184_n21), .A2(ref_1_maj_184_n20), 
        .ZN(ref_1_maj_184_n23) );
  XOR2_X1 ref_1_maj_184_U9 ( .A(ref_1_n28), .B(ref_1_maj_184_n24), .Z(
        ref_1_maj_184_n26) );
  XOR2_X1 ref_1_maj_184_U8 ( .A(ref_1_n37), .B(ref_1_maj_184_n25), .Z(
        ref_1_maj_184_n27) );
  XOR2_X1 ref_1_maj_184_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_184_n24) );
  XOR2_X1 ref_1_maj_184_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_184_n25) );
  OR2_X1 ref_1_maj_184_U5 ( .A1(ref_1_maj_184_n23), .A2(ref_1_maj_184_n22), 
        .ZN(ref_1_maj_184_n32) );
  NAND2_X1 ref_1_maj_184_U4 ( .A1(ref_1_maj_184_n22), .A2(ref_1_maj_184_n23), 
        .ZN(ref_1_maj_184_n34) );
  NAND2_X1 ref_1_maj_184_U3 ( .A1(ref_1_maj_184_n32), .A2(ref_1_maj_184_n31), 
        .ZN(ref_1_maj_184_n33) );
  NAND2_X1 ref_1_maj_184_U2 ( .A1(ref_1_maj_184_n34), .A2(ref_1_maj_184_n33), 
        .ZN(ref_1_maj_184_port_o) );
  OR2_X1 ref_1_maj_185_U19 ( .A1(ref_1_maj_185_n27), .A2(ref_1_maj_185_n26), 
        .ZN(ref_1_maj_185_n28) );
  NAND2_X1 ref_1_maj_185_U18 ( .A1(ref_1_n38), .A2(ref_1_maj_185_n28), .ZN(
        ref_1_maj_185_n29) );
  NAND2_X1 ref_1_maj_185_U17 ( .A1(ref_1_maj_185_n26), .A2(ref_1_maj_185_n27), 
        .ZN(ref_1_maj_185_n30) );
  NAND2_X1 ref_1_maj_185_U16 ( .A1(ref_1_maj_185_n30), .A2(ref_1_maj_185_n29), 
        .ZN(ref_1_maj_185_n31) );
  NAND2_X1 ref_1_maj_185_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_185_n25), .ZN(
        ref_1_maj_185_n18) );
  NAND2_X1 ref_1_maj_185_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_185_n19) );
  NAND2_X1 ref_1_maj_185_U13 ( .A1(ref_1_maj_185_n19), .A2(ref_1_maj_185_n18), 
        .ZN(ref_1_maj_185_n22) );
  NAND2_X1 ref_1_maj_185_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_185_n24), .ZN(
        ref_1_maj_185_n20) );
  NAND2_X1 ref_1_maj_185_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_185_n21) );
  NAND2_X1 ref_1_maj_185_U10 ( .A1(ref_1_maj_185_n21), .A2(ref_1_maj_185_n20), 
        .ZN(ref_1_maj_185_n23) );
  XOR2_X1 ref_1_maj_185_U9 ( .A(ref_1_n28), .B(ref_1_maj_185_n24), .Z(
        ref_1_maj_185_n26) );
  XOR2_X1 ref_1_maj_185_U8 ( .A(ref_1_n37), .B(ref_1_maj_185_n25), .Z(
        ref_1_maj_185_n27) );
  XOR2_X1 ref_1_maj_185_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_185_n24) );
  XOR2_X1 ref_1_maj_185_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_185_n25) );
  OR2_X1 ref_1_maj_185_U5 ( .A1(ref_1_maj_185_n23), .A2(ref_1_maj_185_n22), 
        .ZN(ref_1_maj_185_n32) );
  NAND2_X1 ref_1_maj_185_U4 ( .A1(ref_1_maj_185_n22), .A2(ref_1_maj_185_n23), 
        .ZN(ref_1_maj_185_n34) );
  NAND2_X1 ref_1_maj_185_U3 ( .A1(ref_1_maj_185_n32), .A2(ref_1_maj_185_n31), 
        .ZN(ref_1_maj_185_n33) );
  NAND2_X1 ref_1_maj_185_U2 ( .A1(ref_1_maj_185_n34), .A2(ref_1_maj_185_n33), 
        .ZN(ref_1_maj_185_port_o) );
  OR2_X1 ref_1_maj_186_U19 ( .A1(ref_1_maj_186_n27), .A2(ref_1_maj_186_n26), 
        .ZN(ref_1_maj_186_n28) );
  NAND2_X1 ref_1_maj_186_U18 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_186_n28), .ZN(ref_1_maj_186_n29) );
  NAND2_X1 ref_1_maj_186_U17 ( .A1(ref_1_maj_186_n26), .A2(ref_1_maj_186_n27), 
        .ZN(ref_1_maj_186_n30) );
  NAND2_X1 ref_1_maj_186_U16 ( .A1(ref_1_maj_186_n30), .A2(ref_1_maj_186_n29), 
        .ZN(ref_1_maj_186_n31) );
  NAND2_X1 ref_1_maj_186_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_186_n25), .ZN(
        ref_1_maj_186_n18) );
  NAND2_X1 ref_1_maj_186_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_186_n19) );
  NAND2_X1 ref_1_maj_186_U13 ( .A1(ref_1_maj_186_n19), .A2(ref_1_maj_186_n18), 
        .ZN(ref_1_maj_186_n22) );
  NAND2_X1 ref_1_maj_186_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_186_n24), .ZN(
        ref_1_maj_186_n20) );
  NAND2_X1 ref_1_maj_186_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_186_n21) );
  NAND2_X1 ref_1_maj_186_U10 ( .A1(ref_1_maj_186_n21), .A2(ref_1_maj_186_n20), 
        .ZN(ref_1_maj_186_n23) );
  XOR2_X1 ref_1_maj_186_U9 ( .A(ref_1_n28), .B(ref_1_maj_186_n24), .Z(
        ref_1_maj_186_n26) );
  XOR2_X1 ref_1_maj_186_U8 ( .A(ref_1_n37), .B(ref_1_maj_186_n25), .Z(
        ref_1_maj_186_n27) );
  XOR2_X1 ref_1_maj_186_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_186_n24) );
  XOR2_X1 ref_1_maj_186_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_186_n25) );
  OR2_X1 ref_1_maj_186_U5 ( .A1(ref_1_maj_186_n23), .A2(ref_1_maj_186_n22), 
        .ZN(ref_1_maj_186_n32) );
  NAND2_X1 ref_1_maj_186_U4 ( .A1(ref_1_maj_186_n22), .A2(ref_1_maj_186_n23), 
        .ZN(ref_1_maj_186_n34) );
  NAND2_X1 ref_1_maj_186_U3 ( .A1(ref_1_maj_186_n32), .A2(ref_1_maj_186_n31), 
        .ZN(ref_1_maj_186_n33) );
  NAND2_X1 ref_1_maj_186_U2 ( .A1(ref_1_maj_186_n34), .A2(ref_1_maj_186_n33), 
        .ZN(ref_1_maj_186_port_o) );
  OR2_X1 ref_1_maj_187_U19 ( .A1(ref_1_maj_187_n27), .A2(ref_1_maj_187_n26), 
        .ZN(ref_1_maj_187_n28) );
  NAND2_X1 ref_1_maj_187_U18 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_187_n28), .ZN(ref_1_maj_187_n29) );
  NAND2_X1 ref_1_maj_187_U17 ( .A1(ref_1_maj_187_n26), .A2(ref_1_maj_187_n27), 
        .ZN(ref_1_maj_187_n30) );
  NAND2_X1 ref_1_maj_187_U16 ( .A1(ref_1_maj_187_n30), .A2(ref_1_maj_187_n29), 
        .ZN(ref_1_maj_187_n31) );
  NAND2_X1 ref_1_maj_187_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_187_n25), .ZN(
        ref_1_maj_187_n18) );
  NAND2_X1 ref_1_maj_187_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_187_n19) );
  NAND2_X1 ref_1_maj_187_U13 ( .A1(ref_1_maj_187_n19), .A2(ref_1_maj_187_n18), 
        .ZN(ref_1_maj_187_n22) );
  NAND2_X1 ref_1_maj_187_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_187_n24), .ZN(
        ref_1_maj_187_n20) );
  NAND2_X1 ref_1_maj_187_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_187_n21) );
  NAND2_X1 ref_1_maj_187_U10 ( .A1(ref_1_maj_187_n21), .A2(ref_1_maj_187_n20), 
        .ZN(ref_1_maj_187_n23) );
  XOR2_X1 ref_1_maj_187_U9 ( .A(ref_1_n28), .B(ref_1_maj_187_n24), .Z(
        ref_1_maj_187_n26) );
  XOR2_X1 ref_1_maj_187_U8 ( .A(ref_1_n37), .B(ref_1_maj_187_n25), .Z(
        ref_1_maj_187_n27) );
  XOR2_X1 ref_1_maj_187_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_187_n24) );
  XOR2_X1 ref_1_maj_187_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_187_n25) );
  OR2_X1 ref_1_maj_187_U5 ( .A1(ref_1_maj_187_n23), .A2(ref_1_maj_187_n22), 
        .ZN(ref_1_maj_187_n32) );
  NAND2_X1 ref_1_maj_187_U4 ( .A1(ref_1_maj_187_n22), .A2(ref_1_maj_187_n23), 
        .ZN(ref_1_maj_187_n34) );
  NAND2_X1 ref_1_maj_187_U3 ( .A1(ref_1_maj_187_n32), .A2(ref_1_maj_187_n31), 
        .ZN(ref_1_maj_187_n33) );
  NAND2_X1 ref_1_maj_187_U2 ( .A1(ref_1_maj_187_n34), .A2(ref_1_maj_187_n33), 
        .ZN(ref_1_maj_187_port_o) );
  OR2_X1 ref_1_maj_188_U19 ( .A1(ref_1_maj_188_n27), .A2(ref_1_maj_188_n26), 
        .ZN(ref_1_maj_188_n28) );
  NAND2_X1 ref_1_maj_188_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_188_n28), .ZN(
        ref_1_maj_188_n29) );
  NAND2_X1 ref_1_maj_188_U17 ( .A1(ref_1_maj_188_n26), .A2(ref_1_maj_188_n27), 
        .ZN(ref_1_maj_188_n30) );
  NAND2_X1 ref_1_maj_188_U16 ( .A1(ref_1_maj_188_n30), .A2(ref_1_maj_188_n29), 
        .ZN(ref_1_maj_188_n31) );
  NAND2_X1 ref_1_maj_188_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_188_n25), .ZN(
        ref_1_maj_188_n18) );
  NAND2_X1 ref_1_maj_188_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_188_n19) );
  NAND2_X1 ref_1_maj_188_U13 ( .A1(ref_1_maj_188_n19), .A2(ref_1_maj_188_n18), 
        .ZN(ref_1_maj_188_n22) );
  NAND2_X1 ref_1_maj_188_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_188_n24), .ZN(
        ref_1_maj_188_n20) );
  NAND2_X1 ref_1_maj_188_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_188_n21) );
  NAND2_X1 ref_1_maj_188_U10 ( .A1(ref_1_maj_188_n21), .A2(ref_1_maj_188_n20), 
        .ZN(ref_1_maj_188_n23) );
  XOR2_X1 ref_1_maj_188_U9 ( .A(ref_1_n9), .B(ref_1_maj_188_n24), .Z(
        ref_1_maj_188_n26) );
  XOR2_X1 ref_1_maj_188_U8 ( .A(ref_1_n18), .B(ref_1_maj_188_n25), .Z(
        ref_1_maj_188_n27) );
  XOR2_X1 ref_1_maj_188_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_188_n24)
         );
  XOR2_X1 ref_1_maj_188_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_188_n25) );
  OR2_X1 ref_1_maj_188_U5 ( .A1(ref_1_maj_188_n23), .A2(ref_1_maj_188_n22), 
        .ZN(ref_1_maj_188_n32) );
  NAND2_X1 ref_1_maj_188_U4 ( .A1(ref_1_maj_188_n22), .A2(ref_1_maj_188_n23), 
        .ZN(ref_1_maj_188_n34) );
  NAND2_X1 ref_1_maj_188_U3 ( .A1(ref_1_maj_188_n32), .A2(ref_1_maj_188_n31), 
        .ZN(ref_1_maj_188_n33) );
  NAND2_X1 ref_1_maj_188_U2 ( .A1(ref_1_maj_188_n34), .A2(ref_1_maj_188_n33), 
        .ZN(ref_1_maj_188_port_o) );
  OR2_X1 ref_1_maj_189_U19 ( .A1(ref_1_maj_189_n27), .A2(ref_1_maj_189_n26), 
        .ZN(ref_1_maj_189_n28) );
  NAND2_X1 ref_1_maj_189_U18 ( .A1(ref_1_n19), .A2(ref_1_maj_189_n28), .ZN(
        ref_1_maj_189_n29) );
  NAND2_X1 ref_1_maj_189_U17 ( .A1(ref_1_maj_189_n26), .A2(ref_1_maj_189_n27), 
        .ZN(ref_1_maj_189_n30) );
  NAND2_X1 ref_1_maj_189_U16 ( .A1(ref_1_maj_189_n30), .A2(ref_1_maj_189_n29), 
        .ZN(ref_1_maj_189_n31) );
  NAND2_X1 ref_1_maj_189_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_189_n25), .ZN(
        ref_1_maj_189_n18) );
  NAND2_X1 ref_1_maj_189_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_189_n19) );
  NAND2_X1 ref_1_maj_189_U13 ( .A1(ref_1_maj_189_n19), .A2(ref_1_maj_189_n18), 
        .ZN(ref_1_maj_189_n22) );
  NAND2_X1 ref_1_maj_189_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_189_n24), .ZN(
        ref_1_maj_189_n20) );
  NAND2_X1 ref_1_maj_189_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_189_n21) );
  NAND2_X1 ref_1_maj_189_U10 ( .A1(ref_1_maj_189_n21), .A2(ref_1_maj_189_n20), 
        .ZN(ref_1_maj_189_n23) );
  XOR2_X1 ref_1_maj_189_U9 ( .A(ref_1_n9), .B(ref_1_maj_189_n24), .Z(
        ref_1_maj_189_n26) );
  XOR2_X1 ref_1_maj_189_U8 ( .A(ref_1_n18), .B(ref_1_maj_189_n25), .Z(
        ref_1_maj_189_n27) );
  XOR2_X1 ref_1_maj_189_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_189_n24)
         );
  XOR2_X1 ref_1_maj_189_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_189_n25) );
  OR2_X1 ref_1_maj_189_U5 ( .A1(ref_1_maj_189_n23), .A2(ref_1_maj_189_n22), 
        .ZN(ref_1_maj_189_n32) );
  NAND2_X1 ref_1_maj_189_U4 ( .A1(ref_1_maj_189_n22), .A2(ref_1_maj_189_n23), 
        .ZN(ref_1_maj_189_n34) );
  NAND2_X1 ref_1_maj_189_U3 ( .A1(ref_1_maj_189_n32), .A2(ref_1_maj_189_n31), 
        .ZN(ref_1_maj_189_n33) );
  NAND2_X1 ref_1_maj_189_U2 ( .A1(ref_1_maj_189_n34), .A2(ref_1_maj_189_n33), 
        .ZN(ref_1_maj_189_port_o) );
  OR2_X1 ref_1_maj_190_U19 ( .A1(ref_1_maj_190_n27), .A2(ref_1_maj_190_n26), 
        .ZN(ref_1_maj_190_n28) );
  NAND2_X1 ref_1_maj_190_U18 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_190_n28), .ZN(ref_1_maj_190_n29) );
  NAND2_X1 ref_1_maj_190_U17 ( .A1(ref_1_maj_190_n26), .A2(ref_1_maj_190_n27), 
        .ZN(ref_1_maj_190_n30) );
  NAND2_X1 ref_1_maj_190_U16 ( .A1(ref_1_maj_190_n30), .A2(ref_1_maj_190_n29), 
        .ZN(ref_1_maj_190_n31) );
  NAND2_X1 ref_1_maj_190_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_190_n25), .ZN(
        ref_1_maj_190_n18) );
  NAND2_X1 ref_1_maj_190_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_190_n19) );
  NAND2_X1 ref_1_maj_190_U13 ( .A1(ref_1_maj_190_n19), .A2(ref_1_maj_190_n18), 
        .ZN(ref_1_maj_190_n22) );
  NAND2_X1 ref_1_maj_190_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_190_n24), .ZN(
        ref_1_maj_190_n20) );
  NAND2_X1 ref_1_maj_190_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_190_n21) );
  NAND2_X1 ref_1_maj_190_U10 ( .A1(ref_1_maj_190_n21), .A2(ref_1_maj_190_n20), 
        .ZN(ref_1_maj_190_n23) );
  XOR2_X1 ref_1_maj_190_U9 ( .A(ref_1_n9), .B(ref_1_maj_190_n24), .Z(
        ref_1_maj_190_n26) );
  XOR2_X1 ref_1_maj_190_U8 ( .A(ref_1_n18), .B(ref_1_maj_190_n25), .Z(
        ref_1_maj_190_n27) );
  XOR2_X1 ref_1_maj_190_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_190_n24)
         );
  XOR2_X1 ref_1_maj_190_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_190_n25) );
  OR2_X1 ref_1_maj_190_U5 ( .A1(ref_1_maj_190_n23), .A2(ref_1_maj_190_n22), 
        .ZN(ref_1_maj_190_n32) );
  NAND2_X1 ref_1_maj_190_U4 ( .A1(ref_1_maj_190_n22), .A2(ref_1_maj_190_n23), 
        .ZN(ref_1_maj_190_n34) );
  NAND2_X1 ref_1_maj_190_U3 ( .A1(ref_1_maj_190_n32), .A2(ref_1_maj_190_n31), 
        .ZN(ref_1_maj_190_n33) );
  NAND2_X1 ref_1_maj_190_U2 ( .A1(ref_1_maj_190_n34), .A2(ref_1_maj_190_n33), 
        .ZN(ref_1_maj_190_port_o) );
  OR2_X1 ref_1_maj_191_U19 ( .A1(ref_1_maj_191_n27), .A2(ref_1_maj_191_n26), 
        .ZN(ref_1_maj_191_n28) );
  NAND2_X1 ref_1_maj_191_U18 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_191_n28), .ZN(ref_1_maj_191_n29) );
  NAND2_X1 ref_1_maj_191_U17 ( .A1(ref_1_maj_191_n26), .A2(ref_1_maj_191_n27), 
        .ZN(ref_1_maj_191_n30) );
  NAND2_X1 ref_1_maj_191_U16 ( .A1(ref_1_maj_191_n30), .A2(ref_1_maj_191_n29), 
        .ZN(ref_1_maj_191_n31) );
  NAND2_X1 ref_1_maj_191_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_191_n25), .ZN(
        ref_1_maj_191_n18) );
  NAND2_X1 ref_1_maj_191_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_191_n19) );
  NAND2_X1 ref_1_maj_191_U13 ( .A1(ref_1_maj_191_n19), .A2(ref_1_maj_191_n18), 
        .ZN(ref_1_maj_191_n22) );
  NAND2_X1 ref_1_maj_191_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_191_n24), .ZN(
        ref_1_maj_191_n20) );
  NAND2_X1 ref_1_maj_191_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_191_n21) );
  NAND2_X1 ref_1_maj_191_U10 ( .A1(ref_1_maj_191_n21), .A2(ref_1_maj_191_n20), 
        .ZN(ref_1_maj_191_n23) );
  XOR2_X1 ref_1_maj_191_U9 ( .A(ref_1_n9), .B(ref_1_maj_191_n24), .Z(
        ref_1_maj_191_n26) );
  XOR2_X1 ref_1_maj_191_U8 ( .A(ref_1_n18), .B(ref_1_maj_191_n25), .Z(
        ref_1_maj_191_n27) );
  XOR2_X1 ref_1_maj_191_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_191_n24)
         );
  XOR2_X1 ref_1_maj_191_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_191_n25) );
  OR2_X1 ref_1_maj_191_U5 ( .A1(ref_1_maj_191_n23), .A2(ref_1_maj_191_n22), 
        .ZN(ref_1_maj_191_n32) );
  NAND2_X1 ref_1_maj_191_U4 ( .A1(ref_1_maj_191_n22), .A2(ref_1_maj_191_n23), 
        .ZN(ref_1_maj_191_n34) );
  NAND2_X1 ref_1_maj_191_U3 ( .A1(ref_1_maj_191_n32), .A2(ref_1_maj_191_n31), 
        .ZN(ref_1_maj_191_n33) );
  NAND2_X1 ref_1_maj_191_U2 ( .A1(ref_1_maj_191_n34), .A2(ref_1_maj_191_n33), 
        .ZN(ref_1_maj_191_port_o) );
  OR2_X1 ref_1_maj_192_U19 ( .A1(ref_1_maj_192_n27), .A2(ref_1_maj_192_n26), 
        .ZN(ref_1_maj_192_n28) );
  NAND2_X1 ref_1_maj_192_U18 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_192_n28), .ZN(ref_1_maj_192_n29) );
  NAND2_X1 ref_1_maj_192_U17 ( .A1(ref_1_maj_192_n26), .A2(ref_1_maj_192_n27), 
        .ZN(ref_1_maj_192_n30) );
  NAND2_X1 ref_1_maj_192_U16 ( .A1(ref_1_maj_192_n30), .A2(ref_1_maj_192_n29), 
        .ZN(ref_1_maj_192_n31) );
  NAND2_X1 ref_1_maj_192_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_192_n25), .ZN(
        ref_1_maj_192_n18) );
  NAND2_X1 ref_1_maj_192_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_192_n19) );
  NAND2_X1 ref_1_maj_192_U13 ( .A1(ref_1_maj_192_n19), .A2(ref_1_maj_192_n18), 
        .ZN(ref_1_maj_192_n22) );
  NAND2_X1 ref_1_maj_192_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_192_n24), .ZN(
        ref_1_maj_192_n20) );
  NAND2_X1 ref_1_maj_192_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_192_n21) );
  NAND2_X1 ref_1_maj_192_U10 ( .A1(ref_1_maj_192_n21), .A2(ref_1_maj_192_n20), 
        .ZN(ref_1_maj_192_n23) );
  XOR2_X1 ref_1_maj_192_U9 ( .A(ref_1_n66), .B(ref_1_maj_192_n24), .Z(
        ref_1_maj_192_n26) );
  XOR2_X1 ref_1_maj_192_U8 ( .A(ref_1_n74), .B(ref_1_maj_192_n25), .Z(
        ref_1_maj_192_n27) );
  XOR2_X1 ref_1_maj_192_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_192_n24) );
  XOR2_X1 ref_1_maj_192_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_192_n25) );
  OR2_X1 ref_1_maj_192_U5 ( .A1(ref_1_maj_192_n23), .A2(ref_1_maj_192_n22), 
        .ZN(ref_1_maj_192_n32) );
  NAND2_X1 ref_1_maj_192_U4 ( .A1(ref_1_maj_192_n22), .A2(ref_1_maj_192_n23), 
        .ZN(ref_1_maj_192_n34) );
  NAND2_X1 ref_1_maj_192_U3 ( .A1(ref_1_maj_192_n32), .A2(ref_1_maj_192_n31), 
        .ZN(ref_1_maj_192_n33) );
  NAND2_X1 ref_1_maj_192_U2 ( .A1(ref_1_maj_192_n34), .A2(ref_1_maj_192_n33), 
        .ZN(ref_1_maj_192_port_o) );
  OR2_X1 ref_1_maj_193_U19 ( .A1(ref_1_maj_193_n27), .A2(ref_1_maj_193_n26), 
        .ZN(ref_1_maj_193_n28) );
  NAND2_X1 ref_1_maj_193_U18 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_193_n28), .ZN(ref_1_maj_193_n29) );
  NAND2_X1 ref_1_maj_193_U17 ( .A1(ref_1_maj_193_n26), .A2(ref_1_maj_193_n27), 
        .ZN(ref_1_maj_193_n30) );
  NAND2_X1 ref_1_maj_193_U16 ( .A1(ref_1_maj_193_n30), .A2(ref_1_maj_193_n29), 
        .ZN(ref_1_maj_193_n31) );
  NAND2_X1 ref_1_maj_193_U15 ( .A1(ref_1_n74), .A2(ref_1_maj_193_n25), .ZN(
        ref_1_maj_193_n18) );
  NAND2_X1 ref_1_maj_193_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_193_n19) );
  NAND2_X1 ref_1_maj_193_U13 ( .A1(ref_1_maj_193_n19), .A2(ref_1_maj_193_n18), 
        .ZN(ref_1_maj_193_n22) );
  NAND2_X1 ref_1_maj_193_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_193_n24), .ZN(
        ref_1_maj_193_n20) );
  NAND2_X1 ref_1_maj_193_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_193_n21) );
  NAND2_X1 ref_1_maj_193_U10 ( .A1(ref_1_maj_193_n21), .A2(ref_1_maj_193_n20), 
        .ZN(ref_1_maj_193_n23) );
  XOR2_X1 ref_1_maj_193_U9 ( .A(ref_1_n66), .B(ref_1_maj_193_n24), .Z(
        ref_1_maj_193_n26) );
  XOR2_X1 ref_1_maj_193_U8 ( .A(ref_1_n74), .B(ref_1_maj_193_n25), .Z(
        ref_1_maj_193_n27) );
  XOR2_X1 ref_1_maj_193_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_193_n24) );
  XOR2_X1 ref_1_maj_193_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_193_n25) );
  OR2_X1 ref_1_maj_193_U5 ( .A1(ref_1_maj_193_n23), .A2(ref_1_maj_193_n22), 
        .ZN(ref_1_maj_193_n32) );
  NAND2_X1 ref_1_maj_193_U4 ( .A1(ref_1_maj_193_n22), .A2(ref_1_maj_193_n23), 
        .ZN(ref_1_maj_193_n34) );
  NAND2_X1 ref_1_maj_193_U3 ( .A1(ref_1_maj_193_n32), .A2(ref_1_maj_193_n31), 
        .ZN(ref_1_maj_193_n33) );
  NAND2_X1 ref_1_maj_193_U2 ( .A1(ref_1_maj_193_n34), .A2(ref_1_maj_193_n33), 
        .ZN(ref_1_maj_193_port_o) );
  OR2_X1 ref_1_maj_194_U19 ( .A1(ref_1_maj_194_n27), .A2(ref_1_maj_194_n26), 
        .ZN(ref_1_maj_194_n28) );
  NAND2_X1 ref_1_maj_194_U18 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_194_n28), .ZN(ref_1_maj_194_n29) );
  NAND2_X1 ref_1_maj_194_U17 ( .A1(ref_1_maj_194_n26), .A2(ref_1_maj_194_n27), 
        .ZN(ref_1_maj_194_n30) );
  NAND2_X1 ref_1_maj_194_U16 ( .A1(ref_1_maj_194_n30), .A2(ref_1_maj_194_n29), 
        .ZN(ref_1_maj_194_n31) );
  NAND2_X1 ref_1_maj_194_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_194_n25), .ZN(
        ref_1_maj_194_n18) );
  NAND2_X1 ref_1_maj_194_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_194_n19) );
  NAND2_X1 ref_1_maj_194_U13 ( .A1(ref_1_maj_194_n19), .A2(ref_1_maj_194_n18), 
        .ZN(ref_1_maj_194_n22) );
  NAND2_X1 ref_1_maj_194_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_194_n24), .ZN(
        ref_1_maj_194_n20) );
  NAND2_X1 ref_1_maj_194_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_194_n21) );
  NAND2_X1 ref_1_maj_194_U10 ( .A1(ref_1_maj_194_n21), .A2(ref_1_maj_194_n20), 
        .ZN(ref_1_maj_194_n23) );
  XOR2_X1 ref_1_maj_194_U9 ( .A(ref_1_n64), .B(ref_1_maj_194_n24), .Z(
        ref_1_maj_194_n26) );
  XOR2_X1 ref_1_maj_194_U8 ( .A(ref_1_n75), .B(ref_1_maj_194_n25), .Z(
        ref_1_maj_194_n27) );
  XOR2_X1 ref_1_maj_194_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_194_n24) );
  XOR2_X1 ref_1_maj_194_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_194_n25) );
  OR2_X1 ref_1_maj_194_U5 ( .A1(ref_1_maj_194_n23), .A2(ref_1_maj_194_n22), 
        .ZN(ref_1_maj_194_n32) );
  NAND2_X1 ref_1_maj_194_U4 ( .A1(ref_1_maj_194_n22), .A2(ref_1_maj_194_n23), 
        .ZN(ref_1_maj_194_n34) );
  NAND2_X1 ref_1_maj_194_U3 ( .A1(ref_1_maj_194_n32), .A2(ref_1_maj_194_n31), 
        .ZN(ref_1_maj_194_n33) );
  NAND2_X1 ref_1_maj_194_U2 ( .A1(ref_1_maj_194_n34), .A2(ref_1_maj_194_n33), 
        .ZN(ref_1_maj_194_port_o) );
  OR2_X1 ref_1_maj_195_U19 ( .A1(ref_1_maj_195_n27), .A2(ref_1_maj_195_n26), 
        .ZN(ref_1_maj_195_n28) );
  NAND2_X1 ref_1_maj_195_U18 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_195_n28), .ZN(ref_1_maj_195_n29) );
  NAND2_X1 ref_1_maj_195_U17 ( .A1(ref_1_maj_195_n26), .A2(ref_1_maj_195_n27), 
        .ZN(ref_1_maj_195_n30) );
  NAND2_X1 ref_1_maj_195_U16 ( .A1(ref_1_maj_195_n30), .A2(ref_1_maj_195_n29), 
        .ZN(ref_1_maj_195_n31) );
  NAND2_X1 ref_1_maj_195_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_195_n25), .ZN(
        ref_1_maj_195_n18) );
  NAND2_X1 ref_1_maj_195_U14 ( .A1(ref_1_n69), .A2(ref_1_n72), .ZN(
        ref_1_maj_195_n19) );
  NAND2_X1 ref_1_maj_195_U13 ( .A1(ref_1_maj_195_n19), .A2(ref_1_maj_195_n18), 
        .ZN(ref_1_maj_195_n22) );
  NAND2_X1 ref_1_maj_195_U12 ( .A1(ref_1_n66), .A2(ref_1_maj_195_n24), .ZN(
        ref_1_maj_195_n20) );
  NAND2_X1 ref_1_maj_195_U11 ( .A1(ref_1_n60), .A2(ref_1_n63), .ZN(
        ref_1_maj_195_n21) );
  NAND2_X1 ref_1_maj_195_U10 ( .A1(ref_1_maj_195_n21), .A2(ref_1_maj_195_n20), 
        .ZN(ref_1_maj_195_n23) );
  XOR2_X1 ref_1_maj_195_U9 ( .A(ref_1_n66), .B(ref_1_maj_195_n24), .Z(
        ref_1_maj_195_n26) );
  XOR2_X1 ref_1_maj_195_U8 ( .A(ref_1_n75), .B(ref_1_maj_195_n25), .Z(
        ref_1_maj_195_n27) );
  XOR2_X1 ref_1_maj_195_U7 ( .A(ref_1_n60), .B(ref_1_n63), .Z(
        ref_1_maj_195_n24) );
  XOR2_X1 ref_1_maj_195_U6 ( .A(ref_1_n69), .B(ref_1_n72), .Z(
        ref_1_maj_195_n25) );
  OR2_X1 ref_1_maj_195_U5 ( .A1(ref_1_maj_195_n23), .A2(ref_1_maj_195_n22), 
        .ZN(ref_1_maj_195_n32) );
  NAND2_X1 ref_1_maj_195_U4 ( .A1(ref_1_maj_195_n22), .A2(ref_1_maj_195_n23), 
        .ZN(ref_1_maj_195_n34) );
  NAND2_X1 ref_1_maj_195_U3 ( .A1(ref_1_maj_195_n32), .A2(ref_1_maj_195_n31), 
        .ZN(ref_1_maj_195_n33) );
  NAND2_X1 ref_1_maj_195_U2 ( .A1(ref_1_maj_195_n34), .A2(ref_1_maj_195_n33), 
        .ZN(ref_1_maj_195_port_o) );
  OR2_X1 ref_1_maj_196_U19 ( .A1(ref_1_maj_196_n27), .A2(ref_1_maj_196_n26), 
        .ZN(ref_1_maj_196_n28) );
  NAND2_X1 ref_1_maj_196_U18 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_196_n28), .ZN(ref_1_maj_196_n29) );
  NAND2_X1 ref_1_maj_196_U17 ( .A1(ref_1_maj_196_n26), .A2(ref_1_maj_196_n27), 
        .ZN(ref_1_maj_196_n30) );
  NAND2_X1 ref_1_maj_196_U16 ( .A1(ref_1_maj_196_n30), .A2(ref_1_maj_196_n29), 
        .ZN(ref_1_maj_196_n31) );
  NAND2_X1 ref_1_maj_196_U15 ( .A1(ref_1_n55), .A2(ref_1_maj_196_n25), .ZN(
        ref_1_maj_196_n18) );
  NAND2_X1 ref_1_maj_196_U14 ( .A1(ref_1_n49), .A2(ref_1_n53), .ZN(
        ref_1_maj_196_n19) );
  NAND2_X1 ref_1_maj_196_U13 ( .A1(ref_1_maj_196_n19), .A2(ref_1_maj_196_n18), 
        .ZN(ref_1_maj_196_n22) );
  NAND2_X1 ref_1_maj_196_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_196_n24), .ZN(
        ref_1_maj_196_n20) );
  NAND2_X1 ref_1_maj_196_U11 ( .A1(ref_1_n40), .A2(ref_1_n44), .ZN(
        ref_1_maj_196_n21) );
  NAND2_X1 ref_1_maj_196_U10 ( .A1(ref_1_maj_196_n21), .A2(ref_1_maj_196_n20), 
        .ZN(ref_1_maj_196_n23) );
  XOR2_X1 ref_1_maj_196_U9 ( .A(ref_1_n47), .B(ref_1_maj_196_n24), .Z(
        ref_1_maj_196_n26) );
  XOR2_X1 ref_1_maj_196_U8 ( .A(ref_1_n55), .B(ref_1_maj_196_n25), .Z(
        ref_1_maj_196_n27) );
  XOR2_X1 ref_1_maj_196_U7 ( .A(ref_1_n40), .B(ref_1_n44), .Z(
        ref_1_maj_196_n24) );
  XOR2_X1 ref_1_maj_196_U6 ( .A(ref_1_n49), .B(ref_1_n53), .Z(
        ref_1_maj_196_n25) );
  OR2_X1 ref_1_maj_196_U5 ( .A1(ref_1_maj_196_n23), .A2(ref_1_maj_196_n22), 
        .ZN(ref_1_maj_196_n32) );
  NAND2_X1 ref_1_maj_196_U4 ( .A1(ref_1_maj_196_n22), .A2(ref_1_maj_196_n23), 
        .ZN(ref_1_maj_196_n34) );
  NAND2_X1 ref_1_maj_196_U3 ( .A1(ref_1_maj_196_n32), .A2(ref_1_maj_196_n31), 
        .ZN(ref_1_maj_196_n33) );
  NAND2_X1 ref_1_maj_196_U2 ( .A1(ref_1_maj_196_n34), .A2(ref_1_maj_196_n33), 
        .ZN(ref_1_maj_196_port_o) );
  OR2_X1 ref_1_maj_197_U19 ( .A1(ref_1_maj_197_n27), .A2(ref_1_maj_197_n26), 
        .ZN(ref_1_maj_197_n28) );
  NAND2_X1 ref_1_maj_197_U18 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_197_n28), .ZN(ref_1_maj_197_n29) );
  NAND2_X1 ref_1_maj_197_U17 ( .A1(ref_1_maj_197_n26), .A2(ref_1_maj_197_n27), 
        .ZN(ref_1_maj_197_n30) );
  NAND2_X1 ref_1_maj_197_U16 ( .A1(ref_1_maj_197_n30), .A2(ref_1_maj_197_n29), 
        .ZN(ref_1_maj_197_n31) );
  NAND2_X1 ref_1_maj_197_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_197_n25), .ZN(
        ref_1_maj_197_n18) );
  NAND2_X1 ref_1_maj_197_U14 ( .A1(ref_1_n50), .A2(ref_1_n51), .ZN(
        ref_1_maj_197_n19) );
  NAND2_X1 ref_1_maj_197_U13 ( .A1(ref_1_maj_197_n19), .A2(ref_1_maj_197_n18), 
        .ZN(ref_1_maj_197_n22) );
  NAND2_X1 ref_1_maj_197_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_197_n24), .ZN(
        ref_1_maj_197_n20) );
  NAND2_X1 ref_1_maj_197_U11 ( .A1(ref_1_n41), .A2(ref_1_n42), .ZN(
        ref_1_maj_197_n21) );
  NAND2_X1 ref_1_maj_197_U10 ( .A1(ref_1_maj_197_n21), .A2(ref_1_maj_197_n20), 
        .ZN(ref_1_maj_197_n23) );
  XOR2_X1 ref_1_maj_197_U9 ( .A(ref_1_n45), .B(ref_1_maj_197_n24), .Z(
        ref_1_maj_197_n26) );
  XOR2_X1 ref_1_maj_197_U8 ( .A(ref_1_n56), .B(ref_1_maj_197_n25), .Z(
        ref_1_maj_197_n27) );
  XOR2_X1 ref_1_maj_197_U7 ( .A(ref_1_n41), .B(ref_1_n42), .Z(
        ref_1_maj_197_n24) );
  XOR2_X1 ref_1_maj_197_U6 ( .A(ref_1_n50), .B(ref_1_n51), .Z(
        ref_1_maj_197_n25) );
  OR2_X1 ref_1_maj_197_U5 ( .A1(ref_1_maj_197_n23), .A2(ref_1_maj_197_n22), 
        .ZN(ref_1_maj_197_n32) );
  NAND2_X1 ref_1_maj_197_U4 ( .A1(ref_1_maj_197_n22), .A2(ref_1_maj_197_n23), 
        .ZN(ref_1_maj_197_n34) );
  NAND2_X1 ref_1_maj_197_U3 ( .A1(ref_1_maj_197_n32), .A2(ref_1_maj_197_n31), 
        .ZN(ref_1_maj_197_n33) );
  NAND2_X1 ref_1_maj_197_U2 ( .A1(ref_1_maj_197_n34), .A2(ref_1_maj_197_n33), 
        .ZN(ref_1_maj_197_port_o) );
  OR2_X1 ref_1_maj_198_U19 ( .A1(ref_1_maj_198_n27), .A2(ref_1_maj_198_n26), 
        .ZN(ref_1_maj_198_n28) );
  NAND2_X1 ref_1_maj_198_U18 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_198_n28), .ZN(ref_1_maj_198_n29) );
  NAND2_X1 ref_1_maj_198_U17 ( .A1(ref_1_maj_198_n26), .A2(ref_1_maj_198_n27), 
        .ZN(ref_1_maj_198_n30) );
  NAND2_X1 ref_1_maj_198_U16 ( .A1(ref_1_maj_198_n30), .A2(ref_1_maj_198_n29), 
        .ZN(ref_1_maj_198_n31) );
  NAND2_X1 ref_1_maj_198_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_198_n25), .ZN(
        ref_1_maj_198_n18) );
  NAND2_X1 ref_1_maj_198_U14 ( .A1(ref_1_n50), .A2(ref_1_n53), .ZN(
        ref_1_maj_198_n19) );
  NAND2_X1 ref_1_maj_198_U13 ( .A1(ref_1_maj_198_n19), .A2(ref_1_maj_198_n18), 
        .ZN(ref_1_maj_198_n22) );
  NAND2_X1 ref_1_maj_198_U12 ( .A1(ref_1_n47), .A2(ref_1_maj_198_n24), .ZN(
        ref_1_maj_198_n20) );
  NAND2_X1 ref_1_maj_198_U11 ( .A1(ref_1_n41), .A2(ref_1_n44), .ZN(
        ref_1_maj_198_n21) );
  NAND2_X1 ref_1_maj_198_U10 ( .A1(ref_1_maj_198_n21), .A2(ref_1_maj_198_n20), 
        .ZN(ref_1_maj_198_n23) );
  XOR2_X1 ref_1_maj_198_U9 ( .A(ref_1_n47), .B(ref_1_maj_198_n24), .Z(
        ref_1_maj_198_n26) );
  XOR2_X1 ref_1_maj_198_U8 ( .A(ref_1_n56), .B(ref_1_maj_198_n25), .Z(
        ref_1_maj_198_n27) );
  XOR2_X1 ref_1_maj_198_U7 ( .A(ref_1_n41), .B(ref_1_n44), .Z(
        ref_1_maj_198_n24) );
  XOR2_X1 ref_1_maj_198_U6 ( .A(ref_1_n50), .B(ref_1_n53), .Z(
        ref_1_maj_198_n25) );
  OR2_X1 ref_1_maj_198_U5 ( .A1(ref_1_maj_198_n23), .A2(ref_1_maj_198_n22), 
        .ZN(ref_1_maj_198_n32) );
  NAND2_X1 ref_1_maj_198_U4 ( .A1(ref_1_maj_198_n22), .A2(ref_1_maj_198_n23), 
        .ZN(ref_1_maj_198_n34) );
  NAND2_X1 ref_1_maj_198_U3 ( .A1(ref_1_maj_198_n32), .A2(ref_1_maj_198_n31), 
        .ZN(ref_1_maj_198_n33) );
  NAND2_X1 ref_1_maj_198_U2 ( .A1(ref_1_maj_198_n34), .A2(ref_1_maj_198_n33), 
        .ZN(ref_1_maj_198_port_o) );
  OR2_X1 ref_1_maj_199_U19 ( .A1(ref_1_maj_199_n27), .A2(ref_1_maj_199_n26), 
        .ZN(ref_1_maj_199_n28) );
  NAND2_X1 ref_1_maj_199_U18 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_199_n28), .ZN(ref_1_maj_199_n29) );
  NAND2_X1 ref_1_maj_199_U17 ( .A1(ref_1_maj_199_n26), .A2(ref_1_maj_199_n27), 
        .ZN(ref_1_maj_199_n30) );
  NAND2_X1 ref_1_maj_199_U16 ( .A1(ref_1_maj_199_n30), .A2(ref_1_maj_199_n29), 
        .ZN(ref_1_maj_199_n31) );
  NAND2_X1 ref_1_maj_199_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_199_n25), .ZN(
        ref_1_maj_199_n18) );
  NAND2_X1 ref_1_maj_199_U14 ( .A1(ref_1_n50), .A2(ref_1_n52), .ZN(
        ref_1_maj_199_n19) );
  NAND2_X1 ref_1_maj_199_U13 ( .A1(ref_1_maj_199_n19), .A2(ref_1_maj_199_n18), 
        .ZN(ref_1_maj_199_n22) );
  NAND2_X1 ref_1_maj_199_U12 ( .A1(ref_1_n46), .A2(ref_1_maj_199_n24), .ZN(
        ref_1_maj_199_n20) );
  NAND2_X1 ref_1_maj_199_U11 ( .A1(ref_1_n41), .A2(ref_1_n43), .ZN(
        ref_1_maj_199_n21) );
  NAND2_X1 ref_1_maj_199_U10 ( .A1(ref_1_maj_199_n21), .A2(ref_1_maj_199_n20), 
        .ZN(ref_1_maj_199_n23) );
  XOR2_X1 ref_1_maj_199_U9 ( .A(ref_1_n46), .B(ref_1_maj_199_n24), .Z(
        ref_1_maj_199_n26) );
  XOR2_X1 ref_1_maj_199_U8 ( .A(ref_1_n56), .B(ref_1_maj_199_n25), .Z(
        ref_1_maj_199_n27) );
  XOR2_X1 ref_1_maj_199_U7 ( .A(ref_1_n41), .B(ref_1_n43), .Z(
        ref_1_maj_199_n24) );
  XOR2_X1 ref_1_maj_199_U6 ( .A(ref_1_n50), .B(ref_1_n52), .Z(
        ref_1_maj_199_n25) );
  OR2_X1 ref_1_maj_199_U5 ( .A1(ref_1_maj_199_n23), .A2(ref_1_maj_199_n22), 
        .ZN(ref_1_maj_199_n32) );
  NAND2_X1 ref_1_maj_199_U4 ( .A1(ref_1_maj_199_n22), .A2(ref_1_maj_199_n23), 
        .ZN(ref_1_maj_199_n34) );
  NAND2_X1 ref_1_maj_199_U3 ( .A1(ref_1_maj_199_n32), .A2(ref_1_maj_199_n31), 
        .ZN(ref_1_maj_199_n33) );
  NAND2_X1 ref_1_maj_199_U2 ( .A1(ref_1_maj_199_n34), .A2(ref_1_maj_199_n33), 
        .ZN(ref_1_maj_199_port_o) );
  OR2_X1 ref_1_maj_200_U19 ( .A1(ref_1_maj_200_n27), .A2(ref_1_maj_200_n26), 
        .ZN(ref_1_maj_200_n28) );
  NAND2_X1 ref_1_maj_200_U18 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_200_n28), .ZN(ref_1_maj_200_n29) );
  NAND2_X1 ref_1_maj_200_U17 ( .A1(ref_1_maj_200_n26), .A2(ref_1_maj_200_n27), 
        .ZN(ref_1_maj_200_n30) );
  NAND2_X1 ref_1_maj_200_U16 ( .A1(ref_1_maj_200_n30), .A2(ref_1_maj_200_n29), 
        .ZN(ref_1_maj_200_n31) );
  NAND2_X1 ref_1_maj_200_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_200_n25), .ZN(
        ref_1_maj_200_n18) );
  NAND2_X1 ref_1_maj_200_U14 ( .A1(ref_1_n31), .A2(ref_1_n33), .ZN(
        ref_1_maj_200_n19) );
  NAND2_X1 ref_1_maj_200_U13 ( .A1(ref_1_maj_200_n19), .A2(ref_1_maj_200_n18), 
        .ZN(ref_1_maj_200_n22) );
  NAND2_X1 ref_1_maj_200_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_200_n24), .ZN(
        ref_1_maj_200_n20) );
  NAND2_X1 ref_1_maj_200_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_200_n21) );
  NAND2_X1 ref_1_maj_200_U10 ( .A1(ref_1_maj_200_n21), .A2(ref_1_maj_200_n20), 
        .ZN(ref_1_maj_200_n23) );
  XOR2_X1 ref_1_maj_200_U9 ( .A(ref_1_n28), .B(ref_1_maj_200_n24), .Z(
        ref_1_maj_200_n26) );
  XOR2_X1 ref_1_maj_200_U8 ( .A(ref_1_n37), .B(ref_1_maj_200_n25), .Z(
        ref_1_maj_200_n27) );
  XOR2_X1 ref_1_maj_200_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_200_n24) );
  XOR2_X1 ref_1_maj_200_U6 ( .A(ref_1_n31), .B(ref_1_n33), .Z(
        ref_1_maj_200_n25) );
  OR2_X1 ref_1_maj_200_U5 ( .A1(ref_1_maj_200_n23), .A2(ref_1_maj_200_n22), 
        .ZN(ref_1_maj_200_n32) );
  NAND2_X1 ref_1_maj_200_U4 ( .A1(ref_1_maj_200_n22), .A2(ref_1_maj_200_n23), 
        .ZN(ref_1_maj_200_n34) );
  NAND2_X1 ref_1_maj_200_U3 ( .A1(ref_1_maj_200_n32), .A2(ref_1_maj_200_n31), 
        .ZN(ref_1_maj_200_n33) );
  NAND2_X1 ref_1_maj_200_U2 ( .A1(ref_1_maj_200_n34), .A2(ref_1_maj_200_n33), 
        .ZN(ref_1_maj_200_port_o) );
  OR2_X1 ref_1_maj_201_U19 ( .A1(ref_1_maj_201_n27), .A2(ref_1_maj_201_n26), 
        .ZN(ref_1_maj_201_n28) );
  NAND2_X1 ref_1_maj_201_U18 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_201_n28), .ZN(ref_1_maj_201_n29) );
  NAND2_X1 ref_1_maj_201_U17 ( .A1(ref_1_maj_201_n26), .A2(ref_1_maj_201_n27), 
        .ZN(ref_1_maj_201_n30) );
  NAND2_X1 ref_1_maj_201_U16 ( .A1(ref_1_maj_201_n30), .A2(ref_1_maj_201_n29), 
        .ZN(ref_1_maj_201_n31) );
  NAND2_X1 ref_1_maj_201_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_201_n25), .ZN(
        ref_1_maj_201_n18) );
  NAND2_X1 ref_1_maj_201_U14 ( .A1(ref_1_n29), .A2(ref_1_n34), .ZN(
        ref_1_maj_201_n19) );
  NAND2_X1 ref_1_maj_201_U13 ( .A1(ref_1_maj_201_n19), .A2(ref_1_maj_201_n18), 
        .ZN(ref_1_maj_201_n22) );
  NAND2_X1 ref_1_maj_201_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_201_n24), .ZN(
        ref_1_maj_201_n20) );
  NAND2_X1 ref_1_maj_201_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_201_n21) );
  NAND2_X1 ref_1_maj_201_U10 ( .A1(ref_1_maj_201_n21), .A2(ref_1_maj_201_n20), 
        .ZN(ref_1_maj_201_n23) );
  XOR2_X1 ref_1_maj_201_U9 ( .A(ref_1_n26), .B(ref_1_maj_201_n24), .Z(
        ref_1_maj_201_n26) );
  XOR2_X1 ref_1_maj_201_U8 ( .A(ref_1_n35), .B(ref_1_maj_201_n25), .Z(
        ref_1_maj_201_n27) );
  XOR2_X1 ref_1_maj_201_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_201_n24) );
  XOR2_X1 ref_1_maj_201_U6 ( .A(ref_1_n29), .B(ref_1_n34), .Z(
        ref_1_maj_201_n25) );
  OR2_X1 ref_1_maj_201_U5 ( .A1(ref_1_maj_201_n23), .A2(ref_1_maj_201_n22), 
        .ZN(ref_1_maj_201_n32) );
  NAND2_X1 ref_1_maj_201_U4 ( .A1(ref_1_maj_201_n22), .A2(ref_1_maj_201_n23), 
        .ZN(ref_1_maj_201_n34) );
  NAND2_X1 ref_1_maj_201_U3 ( .A1(ref_1_maj_201_n32), .A2(ref_1_maj_201_n31), 
        .ZN(ref_1_maj_201_n33) );
  NAND2_X1 ref_1_maj_201_U2 ( .A1(ref_1_maj_201_n34), .A2(ref_1_maj_201_n33), 
        .ZN(ref_1_maj_201_port_o) );
  OR2_X1 ref_1_maj_202_U19 ( .A1(ref_1_maj_202_n27), .A2(ref_1_maj_202_n26), 
        .ZN(ref_1_maj_202_n28) );
  NAND2_X1 ref_1_maj_202_U18 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_202_n28), .ZN(ref_1_maj_202_n29) );
  NAND2_X1 ref_1_maj_202_U17 ( .A1(ref_1_maj_202_n26), .A2(ref_1_maj_202_n27), 
        .ZN(ref_1_maj_202_n30) );
  NAND2_X1 ref_1_maj_202_U16 ( .A1(ref_1_maj_202_n30), .A2(ref_1_maj_202_n29), 
        .ZN(ref_1_maj_202_n31) );
  NAND2_X1 ref_1_maj_202_U15 ( .A1(ref_1_n37), .A2(ref_1_maj_202_n25), .ZN(
        ref_1_maj_202_n18) );
  NAND2_X1 ref_1_maj_202_U14 ( .A1(ref_1_n31), .A2(ref_1_n34), .ZN(
        ref_1_maj_202_n19) );
  NAND2_X1 ref_1_maj_202_U13 ( .A1(ref_1_maj_202_n19), .A2(ref_1_maj_202_n18), 
        .ZN(ref_1_maj_202_n22) );
  NAND2_X1 ref_1_maj_202_U12 ( .A1(ref_1_n28), .A2(ref_1_maj_202_n24), .ZN(
        ref_1_maj_202_n20) );
  NAND2_X1 ref_1_maj_202_U11 ( .A1(ref_1_n22), .A2(ref_1_n25), .ZN(
        ref_1_maj_202_n21) );
  NAND2_X1 ref_1_maj_202_U10 ( .A1(ref_1_maj_202_n21), .A2(ref_1_maj_202_n20), 
        .ZN(ref_1_maj_202_n23) );
  XOR2_X1 ref_1_maj_202_U9 ( .A(ref_1_n28), .B(ref_1_maj_202_n24), .Z(
        ref_1_maj_202_n26) );
  XOR2_X1 ref_1_maj_202_U8 ( .A(ref_1_n37), .B(ref_1_maj_202_n25), .Z(
        ref_1_maj_202_n27) );
  XOR2_X1 ref_1_maj_202_U7 ( .A(ref_1_n22), .B(ref_1_n25), .Z(
        ref_1_maj_202_n24) );
  XOR2_X1 ref_1_maj_202_U6 ( .A(ref_1_n31), .B(ref_1_n34), .Z(
        ref_1_maj_202_n25) );
  OR2_X1 ref_1_maj_202_U5 ( .A1(ref_1_maj_202_n23), .A2(ref_1_maj_202_n22), 
        .ZN(ref_1_maj_202_n32) );
  NAND2_X1 ref_1_maj_202_U4 ( .A1(ref_1_maj_202_n22), .A2(ref_1_maj_202_n23), 
        .ZN(ref_1_maj_202_n34) );
  NAND2_X1 ref_1_maj_202_U3 ( .A1(ref_1_maj_202_n32), .A2(ref_1_maj_202_n31), 
        .ZN(ref_1_maj_202_n33) );
  NAND2_X1 ref_1_maj_202_U2 ( .A1(ref_1_maj_202_n34), .A2(ref_1_maj_202_n33), 
        .ZN(ref_1_maj_202_port_o) );
  OR2_X1 ref_1_maj_203_U19 ( .A1(ref_1_maj_203_n27), .A2(ref_1_maj_203_n26), 
        .ZN(ref_1_maj_203_n28) );
  NAND2_X1 ref_1_maj_203_U18 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_203_n28), .ZN(ref_1_maj_203_n29) );
  NAND2_X1 ref_1_maj_203_U17 ( .A1(ref_1_maj_203_n26), .A2(ref_1_maj_203_n27), 
        .ZN(ref_1_maj_203_n30) );
  NAND2_X1 ref_1_maj_203_U16 ( .A1(ref_1_maj_203_n30), .A2(ref_1_maj_203_n29), 
        .ZN(ref_1_maj_203_n31) );
  NAND2_X1 ref_1_maj_203_U15 ( .A1(ref_1_n36), .A2(ref_1_maj_203_n25), .ZN(
        ref_1_maj_203_n18) );
  NAND2_X1 ref_1_maj_203_U14 ( .A1(ref_1_n30), .A2(ref_1_n34), .ZN(
        ref_1_maj_203_n19) );
  NAND2_X1 ref_1_maj_203_U13 ( .A1(ref_1_maj_203_n19), .A2(ref_1_maj_203_n18), 
        .ZN(ref_1_maj_203_n22) );
  NAND2_X1 ref_1_maj_203_U12 ( .A1(ref_1_n27), .A2(ref_1_maj_203_n24), .ZN(
        ref_1_maj_203_n20) );
  NAND2_X1 ref_1_maj_203_U11 ( .A1(ref_1_n21), .A2(ref_1_n24), .ZN(
        ref_1_maj_203_n21) );
  NAND2_X1 ref_1_maj_203_U10 ( .A1(ref_1_maj_203_n21), .A2(ref_1_maj_203_n20), 
        .ZN(ref_1_maj_203_n23) );
  XOR2_X1 ref_1_maj_203_U9 ( .A(ref_1_n27), .B(ref_1_maj_203_n24), .Z(
        ref_1_maj_203_n26) );
  XOR2_X1 ref_1_maj_203_U8 ( .A(ref_1_n36), .B(ref_1_maj_203_n25), .Z(
        ref_1_maj_203_n27) );
  XOR2_X1 ref_1_maj_203_U7 ( .A(ref_1_n21), .B(ref_1_n24), .Z(
        ref_1_maj_203_n24) );
  XOR2_X1 ref_1_maj_203_U6 ( .A(ref_1_n30), .B(ref_1_n34), .Z(
        ref_1_maj_203_n25) );
  OR2_X1 ref_1_maj_203_U5 ( .A1(ref_1_maj_203_n23), .A2(ref_1_maj_203_n22), 
        .ZN(ref_1_maj_203_n32) );
  NAND2_X1 ref_1_maj_203_U4 ( .A1(ref_1_maj_203_n22), .A2(ref_1_maj_203_n23), 
        .ZN(ref_1_maj_203_n34) );
  NAND2_X1 ref_1_maj_203_U3 ( .A1(ref_1_maj_203_n32), .A2(ref_1_maj_203_n31), 
        .ZN(ref_1_maj_203_n33) );
  NAND2_X1 ref_1_maj_203_U2 ( .A1(ref_1_maj_203_n34), .A2(ref_1_maj_203_n33), 
        .ZN(ref_1_maj_203_port_o) );
  OR2_X1 ref_1_maj_204_U19 ( .A1(ref_1_maj_204_n27), .A2(ref_1_maj_204_n26), 
        .ZN(ref_1_maj_204_n28) );
  NAND2_X1 ref_1_maj_204_U18 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_204_n28), .ZN(ref_1_maj_204_n29) );
  NAND2_X1 ref_1_maj_204_U17 ( .A1(ref_1_maj_204_n26), .A2(ref_1_maj_204_n27), 
        .ZN(ref_1_maj_204_n30) );
  NAND2_X1 ref_1_maj_204_U16 ( .A1(ref_1_maj_204_n30), .A2(ref_1_maj_204_n29), 
        .ZN(ref_1_maj_204_n31) );
  NAND2_X1 ref_1_maj_204_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_204_n25), .ZN(
        ref_1_maj_204_n18) );
  NAND2_X1 ref_1_maj_204_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_204_n19) );
  NAND2_X1 ref_1_maj_204_U13 ( .A1(ref_1_maj_204_n19), .A2(ref_1_maj_204_n18), 
        .ZN(ref_1_maj_204_n22) );
  NAND2_X1 ref_1_maj_204_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_204_n24), .ZN(
        ref_1_maj_204_n20) );
  NAND2_X1 ref_1_maj_204_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_204_n21) );
  NAND2_X1 ref_1_maj_204_U10 ( .A1(ref_1_maj_204_n21), .A2(ref_1_maj_204_n20), 
        .ZN(ref_1_maj_204_n23) );
  XOR2_X1 ref_1_maj_204_U9 ( .A(ref_1_n9), .B(ref_1_maj_204_n24), .Z(
        ref_1_maj_204_n26) );
  XOR2_X1 ref_1_maj_204_U8 ( .A(ref_1_n18), .B(ref_1_maj_204_n25), .Z(
        ref_1_maj_204_n27) );
  XOR2_X1 ref_1_maj_204_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_204_n24)
         );
  XOR2_X1 ref_1_maj_204_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_204_n25) );
  OR2_X1 ref_1_maj_204_U5 ( .A1(ref_1_maj_204_n23), .A2(ref_1_maj_204_n22), 
        .ZN(ref_1_maj_204_n32) );
  NAND2_X1 ref_1_maj_204_U4 ( .A1(ref_1_maj_204_n22), .A2(ref_1_maj_204_n23), 
        .ZN(ref_1_maj_204_n34) );
  NAND2_X1 ref_1_maj_204_U3 ( .A1(ref_1_maj_204_n32), .A2(ref_1_maj_204_n31), 
        .ZN(ref_1_maj_204_n33) );
  NAND2_X1 ref_1_maj_204_U2 ( .A1(ref_1_maj_204_n34), .A2(ref_1_maj_204_n33), 
        .ZN(ref_1_maj_204_port_o) );
  OR2_X1 ref_1_maj_205_U19 ( .A1(ref_1_maj_205_n27), .A2(ref_1_maj_205_n26), 
        .ZN(ref_1_maj_205_n28) );
  NAND2_X1 ref_1_maj_205_U18 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_205_n28), .ZN(ref_1_maj_205_n29) );
  NAND2_X1 ref_1_maj_205_U17 ( .A1(ref_1_maj_205_n26), .A2(ref_1_maj_205_n27), 
        .ZN(ref_1_maj_205_n30) );
  NAND2_X1 ref_1_maj_205_U16 ( .A1(ref_1_maj_205_n30), .A2(ref_1_maj_205_n29), 
        .ZN(ref_1_maj_205_n31) );
  NAND2_X1 ref_1_maj_205_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_205_n25), .ZN(
        ref_1_maj_205_n18) );
  NAND2_X1 ref_1_maj_205_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_205_n19) );
  NAND2_X1 ref_1_maj_205_U13 ( .A1(ref_1_maj_205_n19), .A2(ref_1_maj_205_n18), 
        .ZN(ref_1_maj_205_n22) );
  NAND2_X1 ref_1_maj_205_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_205_n24), .ZN(
        ref_1_maj_205_n20) );
  NAND2_X1 ref_1_maj_205_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_205_n21) );
  NAND2_X1 ref_1_maj_205_U10 ( .A1(ref_1_maj_205_n21), .A2(ref_1_maj_205_n20), 
        .ZN(ref_1_maj_205_n23) );
  XOR2_X1 ref_1_maj_205_U9 ( .A(ref_1_n7), .B(ref_1_maj_205_n24), .Z(
        ref_1_maj_205_n26) );
  XOR2_X1 ref_1_maj_205_U8 ( .A(ref_1_n16), .B(ref_1_maj_205_n25), .Z(
        ref_1_maj_205_n27) );
  XOR2_X1 ref_1_maj_205_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_205_n24)
         );
  XOR2_X1 ref_1_maj_205_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_205_n25) );
  OR2_X1 ref_1_maj_205_U5 ( .A1(ref_1_maj_205_n23), .A2(ref_1_maj_205_n22), 
        .ZN(ref_1_maj_205_n32) );
  NAND2_X1 ref_1_maj_205_U4 ( .A1(ref_1_maj_205_n22), .A2(ref_1_maj_205_n23), 
        .ZN(ref_1_maj_205_n34) );
  NAND2_X1 ref_1_maj_205_U3 ( .A1(ref_1_maj_205_n32), .A2(ref_1_maj_205_n31), 
        .ZN(ref_1_maj_205_n33) );
  NAND2_X1 ref_1_maj_205_U2 ( .A1(ref_1_maj_205_n34), .A2(ref_1_maj_205_n33), 
        .ZN(ref_1_maj_205_port_o) );
  OR2_X1 ref_1_maj_206_U19 ( .A1(ref_1_maj_206_n27), .A2(ref_1_maj_206_n26), 
        .ZN(ref_1_maj_206_n28) );
  NAND2_X1 ref_1_maj_206_U18 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_206_n28), .ZN(ref_1_maj_206_n29) );
  NAND2_X1 ref_1_maj_206_U17 ( .A1(ref_1_maj_206_n26), .A2(ref_1_maj_206_n27), 
        .ZN(ref_1_maj_206_n30) );
  NAND2_X1 ref_1_maj_206_U16 ( .A1(ref_1_maj_206_n30), .A2(ref_1_maj_206_n29), 
        .ZN(ref_1_maj_206_n31) );
  NAND2_X1 ref_1_maj_206_U15 ( .A1(ref_1_n18), .A2(ref_1_maj_206_n25), .ZN(
        ref_1_maj_206_n18) );
  NAND2_X1 ref_1_maj_206_U14 ( .A1(ref_1_n12), .A2(ref_1_n15), .ZN(
        ref_1_maj_206_n19) );
  NAND2_X1 ref_1_maj_206_U13 ( .A1(ref_1_maj_206_n19), .A2(ref_1_maj_206_n18), 
        .ZN(ref_1_maj_206_n22) );
  NAND2_X1 ref_1_maj_206_U12 ( .A1(ref_1_n9), .A2(ref_1_maj_206_n24), .ZN(
        ref_1_maj_206_n20) );
  NAND2_X1 ref_1_maj_206_U11 ( .A1(ref_1_n3), .A2(ref_1_n6), .ZN(
        ref_1_maj_206_n21) );
  NAND2_X1 ref_1_maj_206_U10 ( .A1(ref_1_maj_206_n21), .A2(ref_1_maj_206_n20), 
        .ZN(ref_1_maj_206_n23) );
  XOR2_X1 ref_1_maj_206_U9 ( .A(ref_1_n9), .B(ref_1_maj_206_n24), .Z(
        ref_1_maj_206_n26) );
  XOR2_X1 ref_1_maj_206_U8 ( .A(ref_1_n18), .B(ref_1_maj_206_n25), .Z(
        ref_1_maj_206_n27) );
  XOR2_X1 ref_1_maj_206_U7 ( .A(ref_1_n3), .B(ref_1_n6), .Z(ref_1_maj_206_n24)
         );
  XOR2_X1 ref_1_maj_206_U6 ( .A(ref_1_n12), .B(ref_1_n15), .Z(
        ref_1_maj_206_n25) );
  OR2_X1 ref_1_maj_206_U5 ( .A1(ref_1_maj_206_n23), .A2(ref_1_maj_206_n22), 
        .ZN(ref_1_maj_206_n32) );
  NAND2_X1 ref_1_maj_206_U4 ( .A1(ref_1_maj_206_n22), .A2(ref_1_maj_206_n23), 
        .ZN(ref_1_maj_206_n34) );
  NAND2_X1 ref_1_maj_206_U3 ( .A1(ref_1_maj_206_n32), .A2(ref_1_maj_206_n31), 
        .ZN(ref_1_maj_206_n33) );
  NAND2_X1 ref_1_maj_206_U2 ( .A1(ref_1_maj_206_n34), .A2(ref_1_maj_206_n33), 
        .ZN(ref_1_maj_206_port_o) );
  OR2_X1 ref_1_maj_207_U19 ( .A1(ref_1_maj_207_n27), .A2(ref_1_maj_207_n26), 
        .ZN(ref_1_maj_207_n28) );
  NAND2_X1 ref_1_maj_207_U18 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_207_n28), .ZN(ref_1_maj_207_n29) );
  NAND2_X1 ref_1_maj_207_U17 ( .A1(ref_1_maj_207_n26), .A2(ref_1_maj_207_n27), 
        .ZN(ref_1_maj_207_n30) );
  NAND2_X1 ref_1_maj_207_U16 ( .A1(ref_1_maj_207_n30), .A2(ref_1_maj_207_n29), 
        .ZN(ref_1_maj_207_n31) );
  NAND2_X1 ref_1_maj_207_U15 ( .A1(ref_1_n17), .A2(ref_1_maj_207_n25), .ZN(
        ref_1_maj_207_n18) );
  NAND2_X1 ref_1_maj_207_U14 ( .A1(ref_1_n11), .A2(ref_1_n14), .ZN(
        ref_1_maj_207_n19) );
  NAND2_X1 ref_1_maj_207_U13 ( .A1(ref_1_maj_207_n19), .A2(ref_1_maj_207_n18), 
        .ZN(ref_1_maj_207_n22) );
  NAND2_X1 ref_1_maj_207_U12 ( .A1(ref_1_n8), .A2(ref_1_maj_207_n24), .ZN(
        ref_1_maj_207_n20) );
  NAND2_X1 ref_1_maj_207_U11 ( .A1(ref_1_n2), .A2(ref_1_n5), .ZN(
        ref_1_maj_207_n21) );
  NAND2_X1 ref_1_maj_207_U10 ( .A1(ref_1_maj_207_n21), .A2(ref_1_maj_207_n20), 
        .ZN(ref_1_maj_207_n23) );
  XOR2_X1 ref_1_maj_207_U9 ( .A(ref_1_n8), .B(ref_1_maj_207_n24), .Z(
        ref_1_maj_207_n26) );
  XOR2_X1 ref_1_maj_207_U8 ( .A(ref_1_n17), .B(ref_1_maj_207_n25), .Z(
        ref_1_maj_207_n27) );
  XOR2_X1 ref_1_maj_207_U7 ( .A(ref_1_n2), .B(ref_1_n5), .Z(ref_1_maj_207_n24)
         );
  XOR2_X1 ref_1_maj_207_U6 ( .A(ref_1_n11), .B(ref_1_n14), .Z(
        ref_1_maj_207_n25) );
  OR2_X1 ref_1_maj_207_U5 ( .A1(ref_1_maj_207_n23), .A2(ref_1_maj_207_n22), 
        .ZN(ref_1_maj_207_n32) );
  NAND2_X1 ref_1_maj_207_U4 ( .A1(ref_1_maj_207_n22), .A2(ref_1_maj_207_n23), 
        .ZN(ref_1_maj_207_n34) );
  NAND2_X1 ref_1_maj_207_U3 ( .A1(ref_1_maj_207_n32), .A2(ref_1_maj_207_n31), 
        .ZN(ref_1_maj_207_n33) );
  NAND2_X1 ref_1_maj_207_U2 ( .A1(ref_1_maj_207_n34), .A2(ref_1_maj_207_n33), 
        .ZN(ref_1_maj_207_port_o) );
  OR2_X1 ref_1_maj_208_U19 ( .A1(ref_1_maj_208_n27), .A2(ref_1_maj_208_n26), 
        .ZN(ref_1_maj_208_n28) );
  NAND2_X1 ref_1_maj_208_U18 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_208_n28), .ZN(ref_1_maj_208_n29) );
  NAND2_X1 ref_1_maj_208_U17 ( .A1(ref_1_maj_208_n26), .A2(ref_1_maj_208_n27), 
        .ZN(ref_1_maj_208_n30) );
  NAND2_X1 ref_1_maj_208_U16 ( .A1(ref_1_maj_208_n30), .A2(ref_1_maj_208_n29), 
        .ZN(ref_1_maj_208_n31) );
  NAND2_X1 ref_1_maj_208_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_208_n25), .ZN(
        ref_1_maj_208_n18) );
  NAND2_X1 ref_1_maj_208_U14 ( .A1(ref_1_n68), .A2(ref_1_n71), .ZN(
        ref_1_maj_208_n19) );
  NAND2_X1 ref_1_maj_208_U13 ( .A1(ref_1_maj_208_n19), .A2(ref_1_maj_208_n18), 
        .ZN(ref_1_maj_208_n22) );
  NAND2_X1 ref_1_maj_208_U12 ( .A1(ref_1_n65), .A2(ref_1_maj_208_n24), .ZN(
        ref_1_maj_208_n20) );
  NAND2_X1 ref_1_maj_208_U11 ( .A1(ref_1_n59), .A2(ref_1_n62), .ZN(
        ref_1_maj_208_n21) );
  NAND2_X1 ref_1_maj_208_U10 ( .A1(ref_1_maj_208_n21), .A2(ref_1_maj_208_n20), 
        .ZN(ref_1_maj_208_n23) );
  XOR2_X1 ref_1_maj_208_U9 ( .A(ref_1_n65), .B(ref_1_maj_208_n24), .Z(
        ref_1_maj_208_n26) );
  XOR2_X1 ref_1_maj_208_U8 ( .A(ref_1_n75), .B(ref_1_maj_208_n25), .Z(
        ref_1_maj_208_n27) );
  XOR2_X1 ref_1_maj_208_U7 ( .A(ref_1_n59), .B(ref_1_n62), .Z(
        ref_1_maj_208_n24) );
  XOR2_X1 ref_1_maj_208_U6 ( .A(ref_1_n68), .B(ref_1_n71), .Z(
        ref_1_maj_208_n25) );
  OR2_X1 ref_1_maj_208_U5 ( .A1(ref_1_maj_208_n23), .A2(ref_1_maj_208_n22), 
        .ZN(ref_1_maj_208_n32) );
  NAND2_X1 ref_1_maj_208_U4 ( .A1(ref_1_maj_208_n22), .A2(ref_1_maj_208_n23), 
        .ZN(ref_1_maj_208_n34) );
  NAND2_X1 ref_1_maj_208_U3 ( .A1(ref_1_maj_208_n32), .A2(ref_1_maj_208_n31), 
        .ZN(ref_1_maj_208_n33) );
  NAND2_X1 ref_1_maj_208_U2 ( .A1(ref_1_maj_208_n34), .A2(ref_1_maj_208_n33), 
        .ZN(ref_1_maj_208_port_o) );
  OR2_X1 ref_1_maj_209_U19 ( .A1(ref_1_maj_209_n27), .A2(ref_1_maj_209_n26), 
        .ZN(ref_1_maj_209_n28) );
  NAND2_X1 ref_1_maj_209_U18 ( .A1(ref_1_maj_209_n26), .A2(ref_1_maj_209_n27), 
        .ZN(ref_1_maj_209_n30) );
  NAND2_X1 ref_1_maj_209_U17 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_209_n28), .ZN(ref_1_maj_209_n29) );
  NAND2_X1 ref_1_maj_209_U16 ( .A1(ref_1_maj_209_n30), .A2(ref_1_maj_209_n29), 
        .ZN(ref_1_maj_209_n31) );
  NAND2_X1 ref_1_maj_209_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_209_n25), .ZN(
        ref_1_maj_209_n18) );
  NAND2_X1 ref_1_maj_209_U14 ( .A1(ref_1_n67), .A2(ref_1_n70), .ZN(
        ref_1_maj_209_n19) );
  NAND2_X1 ref_1_maj_209_U13 ( .A1(ref_1_maj_209_n19), .A2(ref_1_maj_209_n18), 
        .ZN(ref_1_maj_209_n22) );
  NAND2_X1 ref_1_maj_209_U12 ( .A1(ref_1_n64), .A2(ref_1_maj_209_n24), .ZN(
        ref_1_maj_209_n20) );
  NAND2_X1 ref_1_maj_209_U11 ( .A1(ref_1_n58), .A2(ref_1_n61), .ZN(
        ref_1_maj_209_n21) );
  NAND2_X1 ref_1_maj_209_U10 ( .A1(ref_1_maj_209_n21), .A2(ref_1_maj_209_n20), 
        .ZN(ref_1_maj_209_n23) );
  XOR2_X1 ref_1_maj_209_U9 ( .A(ref_1_n64), .B(ref_1_maj_209_n24), .Z(
        ref_1_maj_209_n26) );
  XOR2_X1 ref_1_maj_209_U8 ( .A(ref_1_n75), .B(ref_1_maj_209_n25), .Z(
        ref_1_maj_209_n27) );
  XOR2_X1 ref_1_maj_209_U7 ( .A(ref_1_n58), .B(ref_1_n61), .Z(
        ref_1_maj_209_n24) );
  XOR2_X1 ref_1_maj_209_U6 ( .A(ref_1_n67), .B(ref_1_n70), .Z(
        ref_1_maj_209_n25) );
  OR2_X1 ref_1_maj_209_U5 ( .A1(ref_1_maj_209_n23), .A2(ref_1_maj_209_n22), 
        .ZN(ref_1_maj_209_n32) );
  NAND2_X1 ref_1_maj_209_U4 ( .A1(ref_1_maj_209_n22), .A2(ref_1_maj_209_n23), 
        .ZN(ref_1_maj_209_n34) );
  NAND2_X1 ref_1_maj_209_U3 ( .A1(ref_1_maj_209_n32), .A2(ref_1_maj_209_n31), 
        .ZN(ref_1_maj_209_n33) );
  NAND2_X1 ref_1_maj_209_U2 ( .A1(ref_1_maj_209_n34), .A2(ref_1_maj_209_n33), 
        .ZN(ref_1_maj_209_port_o) );
  OR2_X1 ref_1_maj_210_U19 ( .A1(ref_1_maj_210_n27), .A2(ref_1_maj_210_n26), 
        .ZN(ref_1_maj_210_n28) );
  NAND2_X1 ref_1_maj_210_U18 ( .A1(ref_1_maj_210_n26), .A2(ref_1_maj_210_n27), 
        .ZN(ref_1_maj_210_n30) );
  NAND2_X1 ref_1_maj_210_U17 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_210_n28), .ZN(ref_1_maj_210_n29) );
  NAND2_X1 ref_1_maj_210_U16 ( .A1(ref_1_maj_210_n30), .A2(ref_1_maj_210_n29), 
        .ZN(ref_1_maj_210_n31) );
  NAND2_X1 ref_1_maj_210_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_210_n25), .ZN(
        ref_1_maj_210_n18) );
  NAND2_X1 ref_1_maj_210_U14 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_210_n19) );
  NAND2_X1 ref_1_maj_210_U13 ( .A1(ref_1_maj_210_n19), .A2(ref_1_maj_210_n18), 
        .ZN(ref_1_maj_210_n22) );
  NAND2_X1 ref_1_maj_210_U12 ( .A1(ref_1_refreshed_0_2_), .A2(
        ref_1_maj_210_n24), .ZN(ref_1_maj_210_n20) );
  NAND2_X1 ref_1_maj_210_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_210_n21) );
  NAND2_X1 ref_1_maj_210_U10 ( .A1(ref_1_maj_210_n21), .A2(ref_1_maj_210_n20), 
        .ZN(ref_1_maj_210_n23) );
  XOR2_X1 ref_1_maj_210_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_210_n24), 
        .Z(ref_1_maj_210_n26) );
  XOR2_X1 ref_1_maj_210_U8 ( .A(ref_1_n75), .B(ref_1_maj_210_n25), .Z(
        ref_1_maj_210_n27) );
  XOR2_X1 ref_1_maj_210_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), .Z(ref_1_maj_210_n24) );
  XOR2_X1 ref_1_maj_210_U6 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), .Z(ref_1_maj_210_n25) );
  OR2_X1 ref_1_maj_210_U5 ( .A1(ref_1_maj_210_n23), .A2(ref_1_maj_210_n22), 
        .ZN(ref_1_maj_210_n32) );
  NAND2_X1 ref_1_maj_210_U4 ( .A1(ref_1_maj_210_n22), .A2(ref_1_maj_210_n23), 
        .ZN(ref_1_maj_210_n34) );
  NAND2_X1 ref_1_maj_210_U3 ( .A1(ref_1_maj_210_n32), .A2(ref_1_maj_210_n31), 
        .ZN(ref_1_maj_210_n33) );
  NAND2_X1 ref_1_maj_210_U2 ( .A1(ref_1_maj_210_n34), .A2(ref_1_maj_210_n33), 
        .ZN(ref_1_maj_210_port_o) );
  OR2_X1 ref_1_maj_211_U19 ( .A1(ref_1_maj_211_n27), .A2(ref_1_maj_211_n26), 
        .ZN(ref_1_maj_211_n28) );
  NAND2_X1 ref_1_maj_211_U18 ( .A1(ref_1_maj_211_n26), .A2(ref_1_maj_211_n27), 
        .ZN(ref_1_maj_211_n30) );
  NAND2_X1 ref_1_maj_211_U17 ( .A1(ref_1_refreshed_0_6_), .A2(
        ref_1_maj_211_n28), .ZN(ref_1_maj_211_n29) );
  NAND2_X1 ref_1_maj_211_U16 ( .A1(ref_1_maj_211_n30), .A2(ref_1_maj_211_n29), 
        .ZN(ref_1_maj_211_n31) );
  NAND2_X1 ref_1_maj_211_U15 ( .A1(ref_1_n75), .A2(ref_1_maj_211_n25), .ZN(
        ref_1_maj_211_n18) );
  NAND2_X1 ref_1_maj_211_U14 ( .A1(ref_1_refreshed_0_3_), .A2(
        ref_1_refreshed_0_4_), .ZN(ref_1_maj_211_n19) );
  NAND2_X1 ref_1_maj_211_U13 ( .A1(ref_1_maj_211_n19), .A2(ref_1_maj_211_n18), 
        .ZN(ref_1_maj_211_n22) );
  NAND2_X1 ref_1_maj_211_U12 ( .A1(ref_1_refreshed_0_2_), .A2(
        ref_1_maj_211_n24), .ZN(ref_1_maj_211_n20) );
  NAND2_X1 ref_1_maj_211_U11 ( .A1(ref_1_refreshed_0_0_), .A2(
        ref_1_refreshed_0_1_), .ZN(ref_1_maj_211_n21) );
  NAND2_X1 ref_1_maj_211_U10 ( .A1(ref_1_maj_211_n21), .A2(ref_1_maj_211_n20), 
        .ZN(ref_1_maj_211_n23) );
  XOR2_X1 ref_1_maj_211_U9 ( .A(ref_1_refreshed_0_2_), .B(ref_1_maj_211_n24), 
        .Z(ref_1_maj_211_n26) );
  XOR2_X1 ref_1_maj_211_U8 ( .A(ref_1_n75), .B(ref_1_maj_211_n25), .Z(
        ref_1_maj_211_n27) );
  XOR2_X1 ref_1_maj_211_U7 ( .A(ref_1_refreshed_0_0_), .B(ref_1_refreshed_0_1_), .Z(ref_1_maj_211_n24) );
  XOR2_X1 ref_1_maj_211_U6 ( .A(ref_1_refreshed_0_3_), .B(ref_1_refreshed_0_4_), .Z(ref_1_maj_211_n25) );
  OR2_X1 ref_1_maj_211_U5 ( .A1(ref_1_maj_211_n23), .A2(ref_1_maj_211_n22), 
        .ZN(ref_1_maj_211_n32) );
  NAND2_X1 ref_1_maj_211_U4 ( .A1(ref_1_maj_211_n22), .A2(ref_1_maj_211_n23), 
        .ZN(ref_1_maj_211_n34) );
  NAND2_X1 ref_1_maj_211_U3 ( .A1(ref_1_maj_211_n32), .A2(ref_1_maj_211_n31), 
        .ZN(ref_1_maj_211_n33) );
  NAND2_X1 ref_1_maj_211_U2 ( .A1(ref_1_maj_211_n34), .A2(ref_1_maj_211_n33), 
        .ZN(ref_1_maj_211_port_o) );
  OR2_X1 ref_1_maj_212_U19 ( .A1(ref_1_maj_212_n27), .A2(ref_1_maj_212_n26), 
        .ZN(ref_1_maj_212_n28) );
  NAND2_X1 ref_1_maj_212_U18 ( .A1(ref_1_maj_212_n26), .A2(ref_1_maj_212_n27), 
        .ZN(ref_1_maj_212_n30) );
  NAND2_X1 ref_1_maj_212_U17 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_212_n28), .ZN(ref_1_maj_212_n29) );
  NAND2_X1 ref_1_maj_212_U16 ( .A1(ref_1_maj_212_n30), .A2(ref_1_maj_212_n29), 
        .ZN(ref_1_maj_212_n31) );
  NAND2_X1 ref_1_maj_212_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_212_n25), .ZN(
        ref_1_maj_212_n18) );
  NAND2_X1 ref_1_maj_212_U14 ( .A1(ref_1_n50), .A2(ref_1_n51), .ZN(
        ref_1_maj_212_n19) );
  NAND2_X1 ref_1_maj_212_U13 ( .A1(ref_1_maj_212_n19), .A2(ref_1_maj_212_n18), 
        .ZN(ref_1_maj_212_n22) );
  NAND2_X1 ref_1_maj_212_U12 ( .A1(ref_1_n45), .A2(ref_1_maj_212_n24), .ZN(
        ref_1_maj_212_n20) );
  NAND2_X1 ref_1_maj_212_U11 ( .A1(ref_1_n41), .A2(ref_1_n42), .ZN(
        ref_1_maj_212_n21) );
  NAND2_X1 ref_1_maj_212_U10 ( .A1(ref_1_maj_212_n21), .A2(ref_1_maj_212_n20), 
        .ZN(ref_1_maj_212_n23) );
  XOR2_X1 ref_1_maj_212_U9 ( .A(ref_1_n45), .B(ref_1_maj_212_n24), .Z(
        ref_1_maj_212_n26) );
  XOR2_X1 ref_1_maj_212_U8 ( .A(ref_1_n56), .B(ref_1_maj_212_n25), .Z(
        ref_1_maj_212_n27) );
  XOR2_X1 ref_1_maj_212_U7 ( .A(ref_1_n41), .B(ref_1_n42), .Z(
        ref_1_maj_212_n24) );
  XOR2_X1 ref_1_maj_212_U6 ( .A(ref_1_n50), .B(ref_1_n51), .Z(
        ref_1_maj_212_n25) );
  OR2_X1 ref_1_maj_212_U5 ( .A1(ref_1_maj_212_n23), .A2(ref_1_maj_212_n22), 
        .ZN(ref_1_maj_212_n32) );
  NAND2_X1 ref_1_maj_212_U4 ( .A1(ref_1_maj_212_n22), .A2(ref_1_maj_212_n23), 
        .ZN(ref_1_maj_212_n34) );
  NAND2_X1 ref_1_maj_212_U3 ( .A1(ref_1_maj_212_n32), .A2(ref_1_maj_212_n31), 
        .ZN(ref_1_maj_212_n33) );
  NAND2_X1 ref_1_maj_212_U2 ( .A1(ref_1_maj_212_n34), .A2(ref_1_maj_212_n33), 
        .ZN(ref_1_maj_212_port_o) );
  OR2_X1 ref_1_maj_213_U19 ( .A1(ref_1_maj_213_n27), .A2(ref_1_maj_213_n26), 
        .ZN(ref_1_maj_213_n28) );
  NAND2_X1 ref_1_maj_213_U18 ( .A1(ref_1_maj_213_n26), .A2(ref_1_maj_213_n27), 
        .ZN(ref_1_maj_213_n30) );
  NAND2_X1 ref_1_maj_213_U17 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_213_n28), .ZN(ref_1_maj_213_n29) );
  NAND2_X1 ref_1_maj_213_U16 ( .A1(ref_1_maj_213_n30), .A2(ref_1_maj_213_n29), 
        .ZN(ref_1_maj_213_n31) );
  NAND2_X1 ref_1_maj_213_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_213_n25), .ZN(
        ref_1_maj_213_n18) );
  NAND2_X1 ref_1_maj_213_U14 ( .A1(ref_1_n50), .A2(ref_1_refreshed_1_4_), .ZN(
        ref_1_maj_213_n19) );
  NAND2_X1 ref_1_maj_213_U13 ( .A1(ref_1_maj_213_n19), .A2(ref_1_maj_213_n18), 
        .ZN(ref_1_maj_213_n22) );
  NAND2_X1 ref_1_maj_213_U12 ( .A1(ref_1_refreshed_1_2_), .A2(
        ref_1_maj_213_n24), .ZN(ref_1_maj_213_n20) );
  NAND2_X1 ref_1_maj_213_U11 ( .A1(ref_1_n41), .A2(ref_1_refreshed_1_1_), .ZN(
        ref_1_maj_213_n21) );
  NAND2_X1 ref_1_maj_213_U10 ( .A1(ref_1_maj_213_n21), .A2(ref_1_maj_213_n20), 
        .ZN(ref_1_maj_213_n23) );
  XOR2_X1 ref_1_maj_213_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_213_n24), 
        .Z(ref_1_maj_213_n26) );
  XOR2_X1 ref_1_maj_213_U8 ( .A(ref_1_n56), .B(ref_1_maj_213_n25), .Z(
        ref_1_maj_213_n27) );
  XOR2_X1 ref_1_maj_213_U7 ( .A(ref_1_n41), .B(ref_1_refreshed_1_1_), .Z(
        ref_1_maj_213_n24) );
  XOR2_X1 ref_1_maj_213_U6 ( .A(ref_1_n50), .B(ref_1_refreshed_1_4_), .Z(
        ref_1_maj_213_n25) );
  OR2_X1 ref_1_maj_213_U5 ( .A1(ref_1_maj_213_n23), .A2(ref_1_maj_213_n22), 
        .ZN(ref_1_maj_213_n32) );
  NAND2_X1 ref_1_maj_213_U4 ( .A1(ref_1_maj_213_n22), .A2(ref_1_maj_213_n23), 
        .ZN(ref_1_maj_213_n34) );
  NAND2_X1 ref_1_maj_213_U3 ( .A1(ref_1_maj_213_n32), .A2(ref_1_maj_213_n31), 
        .ZN(ref_1_maj_213_n33) );
  NAND2_X1 ref_1_maj_213_U2 ( .A1(ref_1_maj_213_n34), .A2(ref_1_maj_213_n33), 
        .ZN(ref_1_maj_213_port_o) );
  OR2_X1 ref_1_maj_214_U19 ( .A1(ref_1_maj_214_n27), .A2(ref_1_maj_214_n26), 
        .ZN(ref_1_maj_214_n28) );
  NAND2_X1 ref_1_maj_214_U18 ( .A1(ref_1_maj_214_n26), .A2(ref_1_maj_214_n27), 
        .ZN(ref_1_maj_214_n30) );
  NAND2_X1 ref_1_maj_214_U17 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_214_n28), .ZN(ref_1_maj_214_n29) );
  NAND2_X1 ref_1_maj_214_U16 ( .A1(ref_1_maj_214_n30), .A2(ref_1_maj_214_n29), 
        .ZN(ref_1_maj_214_n31) );
  NAND2_X1 ref_1_maj_214_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_214_n25), .ZN(
        ref_1_maj_214_n18) );
  NAND2_X1 ref_1_maj_214_U14 ( .A1(ref_1_n50), .A2(ref_1_refreshed_1_4_), .ZN(
        ref_1_maj_214_n19) );
  NAND2_X1 ref_1_maj_214_U13 ( .A1(ref_1_maj_214_n19), .A2(ref_1_maj_214_n18), 
        .ZN(ref_1_maj_214_n22) );
  NAND2_X1 ref_1_maj_214_U12 ( .A1(ref_1_refreshed_1_2_), .A2(
        ref_1_maj_214_n24), .ZN(ref_1_maj_214_n20) );
  NAND2_X1 ref_1_maj_214_U11 ( .A1(ref_1_n41), .A2(ref_1_refreshed_1_1_), .ZN(
        ref_1_maj_214_n21) );
  NAND2_X1 ref_1_maj_214_U10 ( .A1(ref_1_maj_214_n21), .A2(ref_1_maj_214_n20), 
        .ZN(ref_1_maj_214_n23) );
  XOR2_X1 ref_1_maj_214_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_214_n24), 
        .Z(ref_1_maj_214_n26) );
  XOR2_X1 ref_1_maj_214_U8 ( .A(ref_1_n56), .B(ref_1_maj_214_n25), .Z(
        ref_1_maj_214_n27) );
  XOR2_X1 ref_1_maj_214_U7 ( .A(ref_1_n41), .B(ref_1_refreshed_1_1_), .Z(
        ref_1_maj_214_n24) );
  XOR2_X1 ref_1_maj_214_U6 ( .A(ref_1_n50), .B(ref_1_refreshed_1_4_), .Z(
        ref_1_maj_214_n25) );
  OR2_X1 ref_1_maj_214_U5 ( .A1(ref_1_maj_214_n23), .A2(ref_1_maj_214_n22), 
        .ZN(ref_1_maj_214_n32) );
  NAND2_X1 ref_1_maj_214_U4 ( .A1(ref_1_maj_214_n22), .A2(ref_1_maj_214_n23), 
        .ZN(ref_1_maj_214_n34) );
  NAND2_X1 ref_1_maj_214_U3 ( .A1(ref_1_maj_214_n32), .A2(ref_1_maj_214_n31), 
        .ZN(ref_1_maj_214_n33) );
  NAND2_X1 ref_1_maj_214_U2 ( .A1(ref_1_maj_214_n34), .A2(ref_1_maj_214_n33), 
        .ZN(ref_1_maj_214_port_o) );
  OR2_X1 ref_1_maj_215_U19 ( .A1(ref_1_maj_215_n27), .A2(ref_1_maj_215_n26), 
        .ZN(ref_1_maj_215_n28) );
  NAND2_X1 ref_1_maj_215_U18 ( .A1(ref_1_maj_215_n26), .A2(ref_1_maj_215_n27), 
        .ZN(ref_1_maj_215_n30) );
  NAND2_X1 ref_1_maj_215_U17 ( .A1(ref_1_refreshed_1_6_), .A2(
        ref_1_maj_215_n28), .ZN(ref_1_maj_215_n29) );
  NAND2_X1 ref_1_maj_215_U16 ( .A1(ref_1_maj_215_n30), .A2(ref_1_maj_215_n29), 
        .ZN(ref_1_maj_215_n31) );
  NAND2_X1 ref_1_maj_215_U15 ( .A1(ref_1_n56), .A2(ref_1_maj_215_n25), .ZN(
        ref_1_maj_215_n18) );
  NAND2_X1 ref_1_maj_215_U14 ( .A1(ref_1_n50), .A2(ref_1_refreshed_1_4_), .ZN(
        ref_1_maj_215_n19) );
  NAND2_X1 ref_1_maj_215_U13 ( .A1(ref_1_maj_215_n19), .A2(ref_1_maj_215_n18), 
        .ZN(ref_1_maj_215_n22) );
  NAND2_X1 ref_1_maj_215_U12 ( .A1(ref_1_refreshed_1_2_), .A2(
        ref_1_maj_215_n24), .ZN(ref_1_maj_215_n20) );
  NAND2_X1 ref_1_maj_215_U11 ( .A1(ref_1_n41), .A2(ref_1_refreshed_1_1_), .ZN(
        ref_1_maj_215_n21) );
  NAND2_X1 ref_1_maj_215_U10 ( .A1(ref_1_maj_215_n21), .A2(ref_1_maj_215_n20), 
        .ZN(ref_1_maj_215_n23) );
  XOR2_X1 ref_1_maj_215_U9 ( .A(ref_1_refreshed_1_2_), .B(ref_1_maj_215_n24), 
        .Z(ref_1_maj_215_n26) );
  XOR2_X1 ref_1_maj_215_U8 ( .A(ref_1_n56), .B(ref_1_maj_215_n25), .Z(
        ref_1_maj_215_n27) );
  XOR2_X1 ref_1_maj_215_U7 ( .A(ref_1_n41), .B(ref_1_refreshed_1_1_), .Z(
        ref_1_maj_215_n24) );
  XOR2_X1 ref_1_maj_215_U6 ( .A(ref_1_n50), .B(ref_1_refreshed_1_4_), .Z(
        ref_1_maj_215_n25) );
  OR2_X1 ref_1_maj_215_U5 ( .A1(ref_1_maj_215_n23), .A2(ref_1_maj_215_n22), 
        .ZN(ref_1_maj_215_n32) );
  NAND2_X1 ref_1_maj_215_U4 ( .A1(ref_1_maj_215_n22), .A2(ref_1_maj_215_n23), 
        .ZN(ref_1_maj_215_n34) );
  NAND2_X1 ref_1_maj_215_U3 ( .A1(ref_1_maj_215_n32), .A2(ref_1_maj_215_n31), 
        .ZN(ref_1_maj_215_n33) );
  NAND2_X1 ref_1_maj_215_U2 ( .A1(ref_1_maj_215_n34), .A2(ref_1_maj_215_n33), 
        .ZN(ref_1_maj_215_port_o) );
  OR2_X1 ref_1_maj_216_U19 ( .A1(ref_1_maj_216_n27), .A2(ref_1_maj_216_n26), 
        .ZN(ref_1_maj_216_n28) );
  NAND2_X1 ref_1_maj_216_U18 ( .A1(ref_1_maj_216_n26), .A2(ref_1_maj_216_n27), 
        .ZN(ref_1_maj_216_n30) );
  NAND2_X1 ref_1_maj_216_U17 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_216_n28), .ZN(ref_1_maj_216_n29) );
  NAND2_X1 ref_1_maj_216_U16 ( .A1(ref_1_maj_216_n30), .A2(ref_1_maj_216_n29), 
        .ZN(ref_1_maj_216_n31) );
  NAND2_X1 ref_1_maj_216_U15 ( .A1(ref_1_n35), .A2(ref_1_maj_216_n25), .ZN(
        ref_1_maj_216_n18) );
  NAND2_X1 ref_1_maj_216_U14 ( .A1(ref_1_n29), .A2(ref_1_n34), .ZN(
        ref_1_maj_216_n19) );
  NAND2_X1 ref_1_maj_216_U13 ( .A1(ref_1_maj_216_n19), .A2(ref_1_maj_216_n18), 
        .ZN(ref_1_maj_216_n22) );
  NAND2_X1 ref_1_maj_216_U12 ( .A1(ref_1_n26), .A2(ref_1_maj_216_n24), .ZN(
        ref_1_maj_216_n20) );
  NAND2_X1 ref_1_maj_216_U11 ( .A1(ref_1_n20), .A2(ref_1_n23), .ZN(
        ref_1_maj_216_n21) );
  NAND2_X1 ref_1_maj_216_U10 ( .A1(ref_1_maj_216_n21), .A2(ref_1_maj_216_n20), 
        .ZN(ref_1_maj_216_n23) );
  XOR2_X1 ref_1_maj_216_U9 ( .A(ref_1_n26), .B(ref_1_maj_216_n24), .Z(
        ref_1_maj_216_n26) );
  XOR2_X1 ref_1_maj_216_U8 ( .A(ref_1_n35), .B(ref_1_maj_216_n25), .Z(
        ref_1_maj_216_n27) );
  XOR2_X1 ref_1_maj_216_U7 ( .A(ref_1_n20), .B(ref_1_n23), .Z(
        ref_1_maj_216_n24) );
  XOR2_X1 ref_1_maj_216_U6 ( .A(ref_1_n29), .B(ref_1_n34), .Z(
        ref_1_maj_216_n25) );
  OR2_X1 ref_1_maj_216_U5 ( .A1(ref_1_maj_216_n23), .A2(ref_1_maj_216_n22), 
        .ZN(ref_1_maj_216_n32) );
  NAND2_X1 ref_1_maj_216_U4 ( .A1(ref_1_maj_216_n22), .A2(ref_1_maj_216_n23), 
        .ZN(ref_1_maj_216_n34) );
  NAND2_X1 ref_1_maj_216_U3 ( .A1(ref_1_maj_216_n32), .A2(ref_1_maj_216_n31), 
        .ZN(ref_1_maj_216_n33) );
  NAND2_X1 ref_1_maj_216_U2 ( .A1(ref_1_maj_216_n34), .A2(ref_1_maj_216_n33), 
        .ZN(ref_1_maj_216_port_o) );
  OR2_X1 ref_1_maj_217_U19 ( .A1(ref_1_maj_217_n27), .A2(ref_1_maj_217_n26), 
        .ZN(ref_1_maj_217_n28) );
  NAND2_X1 ref_1_maj_217_U18 ( .A1(ref_1_maj_217_n26), .A2(ref_1_maj_217_n27), 
        .ZN(ref_1_maj_217_n30) );
  NAND2_X1 ref_1_maj_217_U17 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_217_n28), .ZN(ref_1_maj_217_n29) );
  NAND2_X1 ref_1_maj_217_U16 ( .A1(ref_1_maj_217_n30), .A2(ref_1_maj_217_n29), 
        .ZN(ref_1_maj_217_n31) );
  NAND2_X1 ref_1_maj_217_U15 ( .A1(ref_1_refreshed_2_5_), .A2(
        ref_1_maj_217_n25), .ZN(ref_1_maj_217_n18) );
  NAND2_X1 ref_1_maj_217_U14 ( .A1(ref_1_refreshed_2_3_), .A2(ref_1_n34), .ZN(
        ref_1_maj_217_n19) );
  NAND2_X1 ref_1_maj_217_U13 ( .A1(ref_1_maj_217_n19), .A2(ref_1_maj_217_n18), 
        .ZN(ref_1_maj_217_n22) );
  NAND2_X1 ref_1_maj_217_U12 ( .A1(ref_1_refreshed_2_2_), .A2(
        ref_1_maj_217_n24), .ZN(ref_1_maj_217_n20) );
  NAND2_X1 ref_1_maj_217_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_217_n21) );
  NAND2_X1 ref_1_maj_217_U10 ( .A1(ref_1_maj_217_n21), .A2(ref_1_maj_217_n20), 
        .ZN(ref_1_maj_217_n23) );
  XOR2_X1 ref_1_maj_217_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_217_n24), 
        .Z(ref_1_maj_217_n26) );
  XOR2_X1 ref_1_maj_217_U8 ( .A(ref_1_refreshed_2_5_), .B(ref_1_maj_217_n25), 
        .Z(ref_1_maj_217_n27) );
  XOR2_X1 ref_1_maj_217_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), .Z(ref_1_maj_217_n24) );
  XOR2_X1 ref_1_maj_217_U6 ( .A(ref_1_refreshed_2_3_), .B(ref_1_n34), .Z(
        ref_1_maj_217_n25) );
  OR2_X1 ref_1_maj_217_U5 ( .A1(ref_1_maj_217_n23), .A2(ref_1_maj_217_n22), 
        .ZN(ref_1_maj_217_n32) );
  NAND2_X1 ref_1_maj_217_U4 ( .A1(ref_1_maj_217_n22), .A2(ref_1_maj_217_n23), 
        .ZN(ref_1_maj_217_n34) );
  NAND2_X1 ref_1_maj_217_U3 ( .A1(ref_1_maj_217_n32), .A2(ref_1_maj_217_n31), 
        .ZN(ref_1_maj_217_n33) );
  NAND2_X1 ref_1_maj_217_U2 ( .A1(ref_1_maj_217_n34), .A2(ref_1_maj_217_n33), 
        .ZN(ref_1_maj_217_port_o) );
  OR2_X1 ref_1_maj_218_U19 ( .A1(ref_1_maj_218_n27), .A2(ref_1_maj_218_n26), 
        .ZN(ref_1_maj_218_n28) );
  NAND2_X1 ref_1_maj_218_U18 ( .A1(ref_1_maj_218_n26), .A2(ref_1_maj_218_n27), 
        .ZN(ref_1_maj_218_n30) );
  NAND2_X1 ref_1_maj_218_U17 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_218_n28), .ZN(ref_1_maj_218_n29) );
  NAND2_X1 ref_1_maj_218_U16 ( .A1(ref_1_maj_218_n30), .A2(ref_1_maj_218_n29), 
        .ZN(ref_1_maj_218_n31) );
  NAND2_X1 ref_1_maj_218_U15 ( .A1(ref_1_refreshed_2_5_), .A2(
        ref_1_maj_218_n25), .ZN(ref_1_maj_218_n18) );
  NAND2_X1 ref_1_maj_218_U14 ( .A1(ref_1_refreshed_2_3_), .A2(ref_1_n34), .ZN(
        ref_1_maj_218_n19) );
  NAND2_X1 ref_1_maj_218_U13 ( .A1(ref_1_maj_218_n19), .A2(ref_1_maj_218_n18), 
        .ZN(ref_1_maj_218_n22) );
  NAND2_X1 ref_1_maj_218_U12 ( .A1(ref_1_refreshed_2_2_), .A2(
        ref_1_maj_218_n24), .ZN(ref_1_maj_218_n20) );
  NAND2_X1 ref_1_maj_218_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_218_n21) );
  NAND2_X1 ref_1_maj_218_U10 ( .A1(ref_1_maj_218_n21), .A2(ref_1_maj_218_n20), 
        .ZN(ref_1_maj_218_n23) );
  XOR2_X1 ref_1_maj_218_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_218_n24), 
        .Z(ref_1_maj_218_n26) );
  XOR2_X1 ref_1_maj_218_U8 ( .A(ref_1_refreshed_2_5_), .B(ref_1_maj_218_n25), 
        .Z(ref_1_maj_218_n27) );
  XOR2_X1 ref_1_maj_218_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), .Z(ref_1_maj_218_n24) );
  XOR2_X1 ref_1_maj_218_U6 ( .A(ref_1_refreshed_2_3_), .B(ref_1_n34), .Z(
        ref_1_maj_218_n25) );
  OR2_X1 ref_1_maj_218_U5 ( .A1(ref_1_maj_218_n23), .A2(ref_1_maj_218_n22), 
        .ZN(ref_1_maj_218_n32) );
  NAND2_X1 ref_1_maj_218_U4 ( .A1(ref_1_maj_218_n22), .A2(ref_1_maj_218_n23), 
        .ZN(ref_1_maj_218_n34) );
  NAND2_X1 ref_1_maj_218_U3 ( .A1(ref_1_maj_218_n32), .A2(ref_1_maj_218_n31), 
        .ZN(ref_1_maj_218_n33) );
  NAND2_X1 ref_1_maj_218_U2 ( .A1(ref_1_maj_218_n34), .A2(ref_1_maj_218_n33), 
        .ZN(ref_1_maj_218_port_o) );
  OR2_X1 ref_1_maj_219_U19 ( .A1(ref_1_maj_219_n27), .A2(ref_1_maj_219_n26), 
        .ZN(ref_1_maj_219_n28) );
  NAND2_X1 ref_1_maj_219_U18 ( .A1(ref_1_maj_219_n26), .A2(ref_1_maj_219_n27), 
        .ZN(ref_1_maj_219_n30) );
  NAND2_X1 ref_1_maj_219_U17 ( .A1(ref_1_refreshed_2_6_), .A2(
        ref_1_maj_219_n28), .ZN(ref_1_maj_219_n29) );
  NAND2_X1 ref_1_maj_219_U16 ( .A1(ref_1_maj_219_n30), .A2(ref_1_maj_219_n29), 
        .ZN(ref_1_maj_219_n31) );
  NAND2_X1 ref_1_maj_219_U15 ( .A1(ref_1_refreshed_2_5_), .A2(
        ref_1_maj_219_n25), .ZN(ref_1_maj_219_n18) );
  NAND2_X1 ref_1_maj_219_U14 ( .A1(ref_1_refreshed_2_3_), .A2(ref_1_n34), .ZN(
        ref_1_maj_219_n19) );
  NAND2_X1 ref_1_maj_219_U13 ( .A1(ref_1_maj_219_n19), .A2(ref_1_maj_219_n18), 
        .ZN(ref_1_maj_219_n22) );
  NAND2_X1 ref_1_maj_219_U12 ( .A1(ref_1_refreshed_2_2_), .A2(
        ref_1_maj_219_n24), .ZN(ref_1_maj_219_n20) );
  NAND2_X1 ref_1_maj_219_U11 ( .A1(ref_1_refreshed_2_0_), .A2(
        ref_1_refreshed_2_1_), .ZN(ref_1_maj_219_n21) );
  NAND2_X1 ref_1_maj_219_U10 ( .A1(ref_1_maj_219_n21), .A2(ref_1_maj_219_n20), 
        .ZN(ref_1_maj_219_n23) );
  XOR2_X1 ref_1_maj_219_U9 ( .A(ref_1_refreshed_2_2_), .B(ref_1_maj_219_n24), 
        .Z(ref_1_maj_219_n26) );
  XOR2_X1 ref_1_maj_219_U8 ( .A(ref_1_refreshed_2_5_), .B(ref_1_maj_219_n25), 
        .Z(ref_1_maj_219_n27) );
  XOR2_X1 ref_1_maj_219_U7 ( .A(ref_1_refreshed_2_0_), .B(ref_1_refreshed_2_1_), .Z(ref_1_maj_219_n24) );
  XOR2_X1 ref_1_maj_219_U6 ( .A(ref_1_refreshed_2_3_), .B(ref_1_n34), .Z(
        ref_1_maj_219_n25) );
  OR2_X1 ref_1_maj_219_U5 ( .A1(ref_1_maj_219_n23), .A2(ref_1_maj_219_n22), 
        .ZN(ref_1_maj_219_n32) );
  NAND2_X1 ref_1_maj_219_U4 ( .A1(ref_1_maj_219_n22), .A2(ref_1_maj_219_n23), 
        .ZN(ref_1_maj_219_n34) );
  NAND2_X1 ref_1_maj_219_U3 ( .A1(ref_1_maj_219_n32), .A2(ref_1_maj_219_n31), 
        .ZN(ref_1_maj_219_n33) );
  NAND2_X1 ref_1_maj_219_U2 ( .A1(ref_1_maj_219_n34), .A2(ref_1_maj_219_n33), 
        .ZN(ref_1_maj_219_port_o) );
  OR2_X1 ref_1_maj_220_U19 ( .A1(ref_1_maj_220_n27), .A2(ref_1_maj_220_n26), 
        .ZN(ref_1_maj_220_n28) );
  NAND2_X1 ref_1_maj_220_U18 ( .A1(ref_1_maj_220_n26), .A2(ref_1_maj_220_n27), 
        .ZN(ref_1_maj_220_n30) );
  NAND2_X1 ref_1_maj_220_U17 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_220_n28), .ZN(ref_1_maj_220_n29) );
  NAND2_X1 ref_1_maj_220_U16 ( .A1(ref_1_maj_220_n30), .A2(ref_1_maj_220_n29), 
        .ZN(ref_1_maj_220_n31) );
  NAND2_X1 ref_1_maj_220_U15 ( .A1(ref_1_n16), .A2(ref_1_maj_220_n25), .ZN(
        ref_1_maj_220_n18) );
  NAND2_X1 ref_1_maj_220_U14 ( .A1(ref_1_n10), .A2(ref_1_n13), .ZN(
        ref_1_maj_220_n19) );
  NAND2_X1 ref_1_maj_220_U13 ( .A1(ref_1_maj_220_n19), .A2(ref_1_maj_220_n18), 
        .ZN(ref_1_maj_220_n22) );
  NAND2_X1 ref_1_maj_220_U12 ( .A1(ref_1_n7), .A2(ref_1_maj_220_n24), .ZN(
        ref_1_maj_220_n20) );
  NAND2_X1 ref_1_maj_220_U11 ( .A1(ref_1_n1), .A2(ref_1_n4), .ZN(
        ref_1_maj_220_n21) );
  NAND2_X1 ref_1_maj_220_U10 ( .A1(ref_1_maj_220_n21), .A2(ref_1_maj_220_n20), 
        .ZN(ref_1_maj_220_n23) );
  XOR2_X1 ref_1_maj_220_U9 ( .A(ref_1_n7), .B(ref_1_maj_220_n24), .Z(
        ref_1_maj_220_n26) );
  XOR2_X1 ref_1_maj_220_U8 ( .A(ref_1_n16), .B(ref_1_maj_220_n25), .Z(
        ref_1_maj_220_n27) );
  XOR2_X1 ref_1_maj_220_U7 ( .A(ref_1_n1), .B(ref_1_n4), .Z(ref_1_maj_220_n24)
         );
  XOR2_X1 ref_1_maj_220_U6 ( .A(ref_1_n10), .B(ref_1_n13), .Z(
        ref_1_maj_220_n25) );
  OR2_X1 ref_1_maj_220_U5 ( .A1(ref_1_maj_220_n23), .A2(ref_1_maj_220_n22), 
        .ZN(ref_1_maj_220_n32) );
  NAND2_X1 ref_1_maj_220_U4 ( .A1(ref_1_maj_220_n22), .A2(ref_1_maj_220_n23), 
        .ZN(ref_1_maj_220_n34) );
  NAND2_X1 ref_1_maj_220_U3 ( .A1(ref_1_maj_220_n32), .A2(ref_1_maj_220_n31), 
        .ZN(ref_1_maj_220_n33) );
  NAND2_X1 ref_1_maj_220_U2 ( .A1(ref_1_maj_220_n34), .A2(ref_1_maj_220_n33), 
        .ZN(ref_1_maj_220_port_o) );
  OR2_X1 ref_1_maj_221_U19 ( .A1(ref_1_maj_221_n27), .A2(ref_1_maj_221_n26), 
        .ZN(ref_1_maj_221_n28) );
  NAND2_X1 ref_1_maj_221_U18 ( .A1(ref_1_maj_221_n26), .A2(ref_1_maj_221_n27), 
        .ZN(ref_1_maj_221_n30) );
  NAND2_X1 ref_1_maj_221_U17 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_221_n28), .ZN(ref_1_maj_221_n29) );
  NAND2_X1 ref_1_maj_221_U16 ( .A1(ref_1_maj_221_n30), .A2(ref_1_maj_221_n29), 
        .ZN(ref_1_maj_221_n31) );
  NAND2_X1 ref_1_maj_221_U15 ( .A1(ref_1_refreshed_3_5_), .A2(
        ref_1_maj_221_n25), .ZN(ref_1_maj_221_n18) );
  NAND2_X1 ref_1_maj_221_U14 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_221_n19) );
  NAND2_X1 ref_1_maj_221_U13 ( .A1(ref_1_maj_221_n19), .A2(ref_1_maj_221_n18), 
        .ZN(ref_1_maj_221_n22) );
  NAND2_X1 ref_1_maj_221_U12 ( .A1(ref_1_refreshed_3_2_), .A2(
        ref_1_maj_221_n24), .ZN(ref_1_maj_221_n20) );
  NAND2_X1 ref_1_maj_221_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_221_n21) );
  NAND2_X1 ref_1_maj_221_U10 ( .A1(ref_1_maj_221_n21), .A2(ref_1_maj_221_n20), 
        .ZN(ref_1_maj_221_n23) );
  XOR2_X1 ref_1_maj_221_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_221_n24), 
        .Z(ref_1_maj_221_n26) );
  XOR2_X1 ref_1_maj_221_U8 ( .A(ref_1_refreshed_3_5_), .B(ref_1_maj_221_n25), 
        .Z(ref_1_maj_221_n27) );
  XOR2_X1 ref_1_maj_221_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), .Z(ref_1_maj_221_n24) );
  XOR2_X1 ref_1_maj_221_U6 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), .Z(ref_1_maj_221_n25) );
  OR2_X1 ref_1_maj_221_U5 ( .A1(ref_1_maj_221_n23), .A2(ref_1_maj_221_n22), 
        .ZN(ref_1_maj_221_n32) );
  NAND2_X1 ref_1_maj_221_U4 ( .A1(ref_1_maj_221_n22), .A2(ref_1_maj_221_n23), 
        .ZN(ref_1_maj_221_n34) );
  NAND2_X1 ref_1_maj_221_U3 ( .A1(ref_1_maj_221_n32), .A2(ref_1_maj_221_n31), 
        .ZN(ref_1_maj_221_n33) );
  NAND2_X1 ref_1_maj_221_U2 ( .A1(ref_1_maj_221_n34), .A2(ref_1_maj_221_n33), 
        .ZN(ref_1_maj_221_port_o) );
  OR2_X1 ref_1_maj_222_U19 ( .A1(ref_1_maj_222_n27), .A2(ref_1_maj_222_n26), 
        .ZN(ref_1_maj_222_n28) );
  NAND2_X1 ref_1_maj_222_U18 ( .A1(ref_1_maj_222_n26), .A2(ref_1_maj_222_n27), 
        .ZN(ref_1_maj_222_n30) );
  NAND2_X1 ref_1_maj_222_U17 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_222_n28), .ZN(ref_1_maj_222_n29) );
  NAND2_X1 ref_1_maj_222_U16 ( .A1(ref_1_maj_222_n30), .A2(ref_1_maj_222_n29), 
        .ZN(ref_1_maj_222_n31) );
  NAND2_X1 ref_1_maj_222_U15 ( .A1(ref_1_refreshed_3_5_), .A2(
        ref_1_maj_222_n25), .ZN(ref_1_maj_222_n18) );
  NAND2_X1 ref_1_maj_222_U14 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_222_n19) );
  NAND2_X1 ref_1_maj_222_U13 ( .A1(ref_1_maj_222_n19), .A2(ref_1_maj_222_n18), 
        .ZN(ref_1_maj_222_n22) );
  NAND2_X1 ref_1_maj_222_U12 ( .A1(ref_1_refreshed_3_2_), .A2(
        ref_1_maj_222_n24), .ZN(ref_1_maj_222_n20) );
  NAND2_X1 ref_1_maj_222_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_222_n21) );
  NAND2_X1 ref_1_maj_222_U10 ( .A1(ref_1_maj_222_n21), .A2(ref_1_maj_222_n20), 
        .ZN(ref_1_maj_222_n23) );
  XOR2_X1 ref_1_maj_222_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_222_n24), 
        .Z(ref_1_maj_222_n26) );
  XOR2_X1 ref_1_maj_222_U8 ( .A(ref_1_refreshed_3_5_), .B(ref_1_maj_222_n25), 
        .Z(ref_1_maj_222_n27) );
  XOR2_X1 ref_1_maj_222_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), .Z(ref_1_maj_222_n24) );
  XOR2_X1 ref_1_maj_222_U6 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), .Z(ref_1_maj_222_n25) );
  OR2_X1 ref_1_maj_222_U5 ( .A1(ref_1_maj_222_n23), .A2(ref_1_maj_222_n22), 
        .ZN(ref_1_maj_222_n32) );
  NAND2_X1 ref_1_maj_222_U4 ( .A1(ref_1_maj_222_n22), .A2(ref_1_maj_222_n23), 
        .ZN(ref_1_maj_222_n34) );
  NAND2_X1 ref_1_maj_222_U3 ( .A1(ref_1_maj_222_n32), .A2(ref_1_maj_222_n31), 
        .ZN(ref_1_maj_222_n33) );
  NAND2_X1 ref_1_maj_222_U2 ( .A1(ref_1_maj_222_n34), .A2(ref_1_maj_222_n33), 
        .ZN(ref_1_maj_222_port_o) );
  OR2_X1 ref_1_maj_223_U19 ( .A1(ref_1_maj_223_n27), .A2(ref_1_maj_223_n26), 
        .ZN(ref_1_maj_223_n28) );
  NAND2_X1 ref_1_maj_223_U18 ( .A1(ref_1_maj_223_n26), .A2(ref_1_maj_223_n27), 
        .ZN(ref_1_maj_223_n30) );
  NAND2_X1 ref_1_maj_223_U17 ( .A1(ref_1_refreshed_3_6_), .A2(
        ref_1_maj_223_n28), .ZN(ref_1_maj_223_n29) );
  NAND2_X1 ref_1_maj_223_U16 ( .A1(ref_1_maj_223_n30), .A2(ref_1_maj_223_n29), 
        .ZN(ref_1_maj_223_n31) );
  NAND2_X1 ref_1_maj_223_U15 ( .A1(ref_1_refreshed_3_5_), .A2(
        ref_1_maj_223_n25), .ZN(ref_1_maj_223_n18) );
  NAND2_X1 ref_1_maj_223_U14 ( .A1(ref_1_refreshed_3_3_), .A2(
        ref_1_refreshed_3_4_), .ZN(ref_1_maj_223_n19) );
  NAND2_X1 ref_1_maj_223_U13 ( .A1(ref_1_maj_223_n19), .A2(ref_1_maj_223_n18), 
        .ZN(ref_1_maj_223_n22) );
  NAND2_X1 ref_1_maj_223_U12 ( .A1(ref_1_refreshed_3_2_), .A2(
        ref_1_maj_223_n24), .ZN(ref_1_maj_223_n20) );
  NAND2_X1 ref_1_maj_223_U11 ( .A1(ref_1_refreshed_3_0_), .A2(
        ref_1_refreshed_3_1_), .ZN(ref_1_maj_223_n21) );
  NAND2_X1 ref_1_maj_223_U10 ( .A1(ref_1_maj_223_n21), .A2(ref_1_maj_223_n20), 
        .ZN(ref_1_maj_223_n23) );
  XOR2_X1 ref_1_maj_223_U9 ( .A(ref_1_refreshed_3_2_), .B(ref_1_maj_223_n24), 
        .Z(ref_1_maj_223_n26) );
  XOR2_X1 ref_1_maj_223_U8 ( .A(ref_1_refreshed_3_5_), .B(ref_1_maj_223_n25), 
        .Z(ref_1_maj_223_n27) );
  XOR2_X1 ref_1_maj_223_U7 ( .A(ref_1_refreshed_3_0_), .B(ref_1_refreshed_3_1_), .Z(ref_1_maj_223_n24) );
  XOR2_X1 ref_1_maj_223_U6 ( .A(ref_1_refreshed_3_3_), .B(ref_1_refreshed_3_4_), .Z(ref_1_maj_223_n25) );
  OR2_X1 ref_1_maj_223_U5 ( .A1(ref_1_maj_223_n23), .A2(ref_1_maj_223_n22), 
        .ZN(ref_1_maj_223_n32) );
  NAND2_X1 ref_1_maj_223_U4 ( .A1(ref_1_maj_223_n22), .A2(ref_1_maj_223_n23), 
        .ZN(ref_1_maj_223_n34) );
  NAND2_X1 ref_1_maj_223_U3 ( .A1(ref_1_maj_223_n32), .A2(ref_1_maj_223_n31), 
        .ZN(ref_1_maj_223_n33) );
  NAND2_X1 ref_1_maj_223_U2 ( .A1(ref_1_maj_223_n34), .A2(ref_1_maj_223_n33), 
        .ZN(ref_1_maj_223_port_o) );
endmodule

