
module CINI_HPC3 ( port_a_0, port_a_1, port_a_2, port_b_0, port_b_1, port_b_2, 
        port_c_0, port_c_1, port_c_2, port_rand_ref, port_rand_mul, clk, reset
 );
  input [6:0] port_a_0;
  input [6:0] port_a_1;
  input [6:0] port_a_2;
  input [6:0] port_b_0;
  input [6:0] port_b_1;
  input [6:0] port_b_2;
  output [6:0] port_c_0;
  output [6:0] port_c_1;
  output [6:0] port_c_2;
  input [2:0] port_rand_ref;
  input [2:0] port_rand_mul;
  input clk, reset;
  wire   simpleAnd_42_port_z, simpleAnd_43_port_z, simpleAnd_44_port_z,
         simpleAnd_45_port_z, simpleAnd_46_port_z, simpleAnd_47_port_z,
         simpleAnd_48_port_z, simpleAnd_49_port_z, simpleAnd_50_port_z,
         simpleAnd_51_port_z, simpleAnd_52_port_z, simpleAnd_53_port_z,
         simpleAnd_54_port_z, simpleAnd_55_port_z, simpleAnd_56_port_z,
         simpleAnd_57_port_z, simpleAnd_58_port_z, simpleAnd_59_port_z,
         simpleAnd_60_port_z, simpleAnd_61_port_z, simpleAnd_62_port_z,
         simpleAnd_63_port_z, simpleAnd_64_port_z, simpleAnd_65_port_z,
         simpleAnd_66_port_z, simpleAnd_67_port_z, simpleAnd_68_port_z,
         simpleAnd_69_port_z, simpleAnd_70_port_z, simpleAnd_71_port_z,
         simpleAnd_72_port_z, simpleAnd_73_port_z, simpleAnd_74_port_z,
         simpleAnd_75_port_z, simpleAnd_76_port_z, simpleAnd_77_port_z,
         simpleAnd_78_port_z, simpleAnd_79_port_z, simpleAnd_80_port_z,
         simpleAnd_81_port_z, simpleAnd_82_port_z, simpleAnd_83_port_z,
         maj_84_port_o, maj_85_port_o, maj_86_port_o, maj_87_port_o,
         maj_88_port_o, maj_89_port_o, maj_90_port_o, maj_91_port_o,
         maj_92_port_o, maj_93_port_o, maj_94_port_o, maj_95_port_o,
         maj_96_port_o, maj_97_port_o, maj_98_port_o, maj_99_port_o,
         maj_100_port_o, maj_101_port_o, maj_102_port_o, maj_103_port_o,
         maj_104_port_o, maj_105_port_o, maj_106_port_o, maj_107_port_o,
         maj_108_port_o, maj_109_port_o, maj_110_port_o, maj_111_port_o,
         maj_112_port_o, maj_113_port_o, maj_114_port_o, maj_115_port_o,
         maj_116_port_o, maj_117_port_o, maj_118_port_o, maj_119_port_o,
         maj_120_port_o, maj_121_port_o, maj_122_port_o, maj_123_port_o,
         maj_124_port_o, maj_125_port_o, maj_126_port_o, maj_127_port_o,
         maj_128_port_o, maj_129_port_o, maj_130_port_o, maj_131_port_o,
         maj_132_port_o, maj_133_port_o, maj_134_port_o, maj_135_port_o,
         maj_136_port_o, maj_137_port_o, maj_138_port_o, maj_139_port_o,
         maj_140_port_o, maj_141_port_o, maj_142_port_o, maj_143_port_o,
         maj_144_port_o, maj_145_port_o, maj_146_port_o, maj_147_port_o,
         maj_148_port_o, maj_149_port_o, maj_150_port_o, maj_151_port_o,
         maj_152_port_o, maj_153_port_o, maj_154_port_o, maj_155_port_o,
         maj_156_port_o, maj_157_port_o, maj_158_port_o, maj_159_port_o,
         maj_160_port_o, maj_161_port_o, maj_162_port_o, maj_163_port_o,
         maj_164_port_o, maj_165_port_o, maj_166_port_o, maj_167_port_o, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, maj_84_n17, maj_84_n16,
         maj_84_n15, maj_84_n14, maj_84_n13, maj_84_n12, maj_84_n11,
         maj_84_n10, maj_84_n9, maj_84_n8, maj_84_n7, maj_84_n6, maj_84_n5,
         maj_84_n4, maj_84_n3, maj_84_n2, maj_84_n1, maj_85_n34, maj_85_n33,
         maj_85_n32, maj_85_n31, maj_85_n30, maj_85_n29, maj_85_n28,
         maj_85_n27, maj_85_n26, maj_85_n25, maj_85_n24, maj_85_n23,
         maj_85_n22, maj_85_n21, maj_85_n20, maj_85_n19, maj_85_n18,
         maj_86_n34, maj_86_n33, maj_86_n32, maj_86_n31, maj_86_n30,
         maj_86_n29, maj_86_n28, maj_86_n27, maj_86_n26, maj_86_n25,
         maj_86_n24, maj_86_n23, maj_86_n22, maj_86_n21, maj_86_n20,
         maj_86_n19, maj_86_n18, maj_87_n34, maj_87_n33, maj_87_n32,
         maj_87_n31, maj_87_n30, maj_87_n29, maj_87_n28, maj_87_n27,
         maj_87_n26, maj_87_n25, maj_87_n24, maj_87_n23, maj_87_n22,
         maj_87_n21, maj_87_n20, maj_87_n19, maj_87_n18, maj_88_n34,
         maj_88_n33, maj_88_n32, maj_88_n31, maj_88_n30, maj_88_n29,
         maj_88_n28, maj_88_n27, maj_88_n26, maj_88_n25, maj_88_n24,
         maj_88_n23, maj_88_n22, maj_88_n21, maj_88_n20, maj_88_n19,
         maj_88_n18, maj_89_n34, maj_89_n33, maj_89_n32, maj_89_n31,
         maj_89_n30, maj_89_n29, maj_89_n28, maj_89_n27, maj_89_n26,
         maj_89_n25, maj_89_n24, maj_89_n23, maj_89_n22, maj_89_n21,
         maj_89_n20, maj_89_n19, maj_89_n18, maj_90_n34, maj_90_n33,
         maj_90_n32, maj_90_n31, maj_90_n30, maj_90_n29, maj_90_n28,
         maj_90_n27, maj_90_n26, maj_90_n25, maj_90_n24, maj_90_n23,
         maj_90_n22, maj_90_n21, maj_90_n20, maj_90_n19, maj_90_n18,
         maj_91_n34, maj_91_n33, maj_91_n32, maj_91_n31, maj_91_n30,
         maj_91_n29, maj_91_n28, maj_91_n27, maj_91_n26, maj_91_n25,
         maj_91_n24, maj_91_n23, maj_91_n22, maj_91_n21, maj_91_n20,
         maj_91_n19, maj_91_n18, maj_92_n34, maj_92_n33, maj_92_n32,
         maj_92_n31, maj_92_n30, maj_92_n29, maj_92_n28, maj_92_n27,
         maj_92_n26, maj_92_n25, maj_92_n24, maj_92_n23, maj_92_n22,
         maj_92_n21, maj_92_n20, maj_92_n19, maj_92_n18, maj_93_n34,
         maj_93_n33, maj_93_n32, maj_93_n31, maj_93_n30, maj_93_n29,
         maj_93_n28, maj_93_n27, maj_93_n26, maj_93_n25, maj_93_n24,
         maj_93_n23, maj_93_n22, maj_93_n21, maj_93_n20, maj_93_n19,
         maj_93_n18, maj_94_n34, maj_94_n33, maj_94_n32, maj_94_n31,
         maj_94_n30, maj_94_n29, maj_94_n28, maj_94_n27, maj_94_n26,
         maj_94_n25, maj_94_n24, maj_94_n23, maj_94_n22, maj_94_n21,
         maj_94_n20, maj_94_n19, maj_94_n18, maj_95_n34, maj_95_n33,
         maj_95_n32, maj_95_n31, maj_95_n30, maj_95_n29, maj_95_n28,
         maj_95_n27, maj_95_n26, maj_95_n25, maj_95_n24, maj_95_n23,
         maj_95_n22, maj_95_n21, maj_95_n20, maj_95_n19, maj_95_n18,
         maj_96_n34, maj_96_n33, maj_96_n32, maj_96_n31, maj_96_n30,
         maj_96_n29, maj_96_n28, maj_96_n27, maj_96_n26, maj_96_n25,
         maj_96_n24, maj_96_n23, maj_96_n22, maj_96_n21, maj_96_n20,
         maj_96_n19, maj_96_n18, maj_97_n34, maj_97_n33, maj_97_n32,
         maj_97_n31, maj_97_n30, maj_97_n29, maj_97_n28, maj_97_n27,
         maj_97_n26, maj_97_n25, maj_97_n24, maj_97_n23, maj_97_n22,
         maj_97_n21, maj_97_n20, maj_97_n19, maj_97_n18, maj_98_n34,
         maj_98_n33, maj_98_n32, maj_98_n31, maj_98_n30, maj_98_n29,
         maj_98_n28, maj_98_n27, maj_98_n26, maj_98_n25, maj_98_n24,
         maj_98_n23, maj_98_n22, maj_98_n21, maj_98_n20, maj_98_n19,
         maj_98_n18, maj_99_n34, maj_99_n33, maj_99_n32, maj_99_n31,
         maj_99_n30, maj_99_n29, maj_99_n28, maj_99_n27, maj_99_n26,
         maj_99_n25, maj_99_n24, maj_99_n23, maj_99_n22, maj_99_n21,
         maj_99_n20, maj_99_n19, maj_99_n18, maj_100_n34, maj_100_n33,
         maj_100_n32, maj_100_n31, maj_100_n30, maj_100_n29, maj_100_n28,
         maj_100_n27, maj_100_n26, maj_100_n25, maj_100_n24, maj_100_n23,
         maj_100_n22, maj_100_n21, maj_100_n20, maj_100_n19, maj_100_n18,
         maj_101_n34, maj_101_n33, maj_101_n32, maj_101_n31, maj_101_n30,
         maj_101_n29, maj_101_n28, maj_101_n27, maj_101_n26, maj_101_n25,
         maj_101_n24, maj_101_n23, maj_101_n22, maj_101_n21, maj_101_n20,
         maj_101_n19, maj_101_n18, maj_102_n34, maj_102_n33, maj_102_n32,
         maj_102_n31, maj_102_n30, maj_102_n29, maj_102_n28, maj_102_n27,
         maj_102_n26, maj_102_n25, maj_102_n24, maj_102_n23, maj_102_n22,
         maj_102_n21, maj_102_n20, maj_102_n19, maj_102_n18, maj_103_n34,
         maj_103_n33, maj_103_n32, maj_103_n31, maj_103_n30, maj_103_n29,
         maj_103_n28, maj_103_n27, maj_103_n26, maj_103_n25, maj_103_n24,
         maj_103_n23, maj_103_n22, maj_103_n21, maj_103_n20, maj_103_n19,
         maj_103_n18, maj_104_n34, maj_104_n33, maj_104_n32, maj_104_n31,
         maj_104_n30, maj_104_n29, maj_104_n28, maj_104_n27, maj_104_n26,
         maj_104_n25, maj_104_n24, maj_104_n23, maj_104_n22, maj_104_n21,
         maj_104_n20, maj_104_n19, maj_104_n18, maj_105_n34, maj_105_n33,
         maj_105_n32, maj_105_n31, maj_105_n30, maj_105_n29, maj_105_n28,
         maj_105_n27, maj_105_n26, maj_105_n25, maj_105_n24, maj_105_n23,
         maj_105_n22, maj_105_n21, maj_105_n20, maj_105_n19, maj_105_n18,
         maj_106_n34, maj_106_n33, maj_106_n32, maj_106_n31, maj_106_n30,
         maj_106_n29, maj_106_n28, maj_106_n27, maj_106_n26, maj_106_n25,
         maj_106_n24, maj_106_n23, maj_106_n22, maj_106_n21, maj_106_n20,
         maj_106_n19, maj_106_n18, maj_107_n34, maj_107_n33, maj_107_n32,
         maj_107_n31, maj_107_n30, maj_107_n29, maj_107_n28, maj_107_n27,
         maj_107_n26, maj_107_n25, maj_107_n24, maj_107_n23, maj_107_n22,
         maj_107_n21, maj_107_n20, maj_107_n19, maj_107_n18, maj_108_n34,
         maj_108_n33, maj_108_n32, maj_108_n31, maj_108_n30, maj_108_n29,
         maj_108_n28, maj_108_n27, maj_108_n26, maj_108_n25, maj_108_n24,
         maj_108_n23, maj_108_n22, maj_108_n21, maj_108_n20, maj_108_n19,
         maj_108_n18, maj_109_n34, maj_109_n33, maj_109_n32, maj_109_n31,
         maj_109_n30, maj_109_n29, maj_109_n28, maj_109_n27, maj_109_n26,
         maj_109_n25, maj_109_n24, maj_109_n23, maj_109_n22, maj_109_n21,
         maj_109_n20, maj_109_n19, maj_109_n18, maj_110_n34, maj_110_n33,
         maj_110_n32, maj_110_n31, maj_110_n30, maj_110_n29, maj_110_n28,
         maj_110_n27, maj_110_n26, maj_110_n25, maj_110_n24, maj_110_n23,
         maj_110_n22, maj_110_n21, maj_110_n20, maj_110_n19, maj_110_n18,
         maj_111_n34, maj_111_n33, maj_111_n32, maj_111_n31, maj_111_n30,
         maj_111_n29, maj_111_n28, maj_111_n27, maj_111_n26, maj_111_n25,
         maj_111_n24, maj_111_n23, maj_111_n22, maj_111_n21, maj_111_n20,
         maj_111_n19, maj_111_n18, maj_112_n34, maj_112_n33, maj_112_n32,
         maj_112_n31, maj_112_n30, maj_112_n29, maj_112_n28, maj_112_n27,
         maj_112_n26, maj_112_n25, maj_112_n24, maj_112_n23, maj_112_n22,
         maj_112_n21, maj_112_n20, maj_112_n19, maj_112_n18, maj_113_n34,
         maj_113_n33, maj_113_n32, maj_113_n31, maj_113_n30, maj_113_n29,
         maj_113_n28, maj_113_n27, maj_113_n26, maj_113_n25, maj_113_n24,
         maj_113_n23, maj_113_n22, maj_113_n21, maj_113_n20, maj_113_n19,
         maj_113_n18, maj_114_n34, maj_114_n33, maj_114_n32, maj_114_n31,
         maj_114_n30, maj_114_n29, maj_114_n28, maj_114_n27, maj_114_n26,
         maj_114_n25, maj_114_n24, maj_114_n23, maj_114_n22, maj_114_n21,
         maj_114_n20, maj_114_n19, maj_114_n18, maj_115_n34, maj_115_n33,
         maj_115_n32, maj_115_n31, maj_115_n30, maj_115_n29, maj_115_n28,
         maj_115_n27, maj_115_n26, maj_115_n25, maj_115_n24, maj_115_n23,
         maj_115_n22, maj_115_n21, maj_115_n20, maj_115_n19, maj_115_n18,
         maj_116_n34, maj_116_n33, maj_116_n32, maj_116_n31, maj_116_n30,
         maj_116_n29, maj_116_n28, maj_116_n27, maj_116_n26, maj_116_n25,
         maj_116_n24, maj_116_n23, maj_116_n22, maj_116_n21, maj_116_n20,
         maj_116_n19, maj_116_n18, maj_117_n34, maj_117_n33, maj_117_n32,
         maj_117_n31, maj_117_n30, maj_117_n29, maj_117_n28, maj_117_n27,
         maj_117_n26, maj_117_n25, maj_117_n24, maj_117_n23, maj_117_n22,
         maj_117_n21, maj_117_n20, maj_117_n19, maj_117_n18, maj_118_n34,
         maj_118_n33, maj_118_n32, maj_118_n31, maj_118_n30, maj_118_n29,
         maj_118_n28, maj_118_n27, maj_118_n26, maj_118_n25, maj_118_n24,
         maj_118_n23, maj_118_n22, maj_118_n21, maj_118_n20, maj_118_n19,
         maj_118_n18, maj_119_n34, maj_119_n33, maj_119_n32, maj_119_n31,
         maj_119_n30, maj_119_n29, maj_119_n28, maj_119_n27, maj_119_n26,
         maj_119_n25, maj_119_n24, maj_119_n23, maj_119_n22, maj_119_n21,
         maj_119_n20, maj_119_n19, maj_119_n18, maj_120_n34, maj_120_n33,
         maj_120_n32, maj_120_n31, maj_120_n30, maj_120_n29, maj_120_n28,
         maj_120_n27, maj_120_n26, maj_120_n25, maj_120_n24, maj_120_n23,
         maj_120_n22, maj_120_n21, maj_120_n20, maj_120_n19, maj_120_n18,
         maj_121_n34, maj_121_n33, maj_121_n32, maj_121_n31, maj_121_n30,
         maj_121_n29, maj_121_n28, maj_121_n27, maj_121_n26, maj_121_n25,
         maj_121_n24, maj_121_n23, maj_121_n22, maj_121_n21, maj_121_n20,
         maj_121_n19, maj_121_n18, maj_122_n34, maj_122_n33, maj_122_n32,
         maj_122_n31, maj_122_n30, maj_122_n29, maj_122_n28, maj_122_n27,
         maj_122_n26, maj_122_n25, maj_122_n24, maj_122_n23, maj_122_n22,
         maj_122_n21, maj_122_n20, maj_122_n19, maj_122_n18, maj_123_n34,
         maj_123_n33, maj_123_n32, maj_123_n31, maj_123_n30, maj_123_n29,
         maj_123_n28, maj_123_n27, maj_123_n26, maj_123_n25, maj_123_n24,
         maj_123_n23, maj_123_n22, maj_123_n21, maj_123_n20, maj_123_n19,
         maj_123_n18, maj_124_n34, maj_124_n33, maj_124_n32, maj_124_n31,
         maj_124_n30, maj_124_n29, maj_124_n28, maj_124_n27, maj_124_n26,
         maj_124_n25, maj_124_n24, maj_124_n23, maj_124_n22, maj_124_n21,
         maj_124_n20, maj_124_n19, maj_124_n18, maj_125_n34, maj_125_n33,
         maj_125_n32, maj_125_n31, maj_125_n30, maj_125_n29, maj_125_n28,
         maj_125_n27, maj_125_n26, maj_125_n25, maj_125_n24, maj_125_n23,
         maj_125_n22, maj_125_n21, maj_125_n20, maj_125_n19, maj_125_n18,
         maj_126_n34, maj_126_n33, maj_126_n32, maj_126_n31, maj_126_n30,
         maj_126_n29, maj_126_n28, maj_126_n27, maj_126_n26, maj_126_n25,
         maj_126_n24, maj_126_n23, maj_126_n22, maj_126_n21, maj_126_n20,
         maj_126_n19, maj_126_n18, maj_127_n34, maj_127_n33, maj_127_n32,
         maj_127_n31, maj_127_n30, maj_127_n29, maj_127_n28, maj_127_n27,
         maj_127_n26, maj_127_n25, maj_127_n24, maj_127_n23, maj_127_n22,
         maj_127_n21, maj_127_n20, maj_127_n19, maj_127_n18, maj_128_n34,
         maj_128_n33, maj_128_n32, maj_128_n31, maj_128_n30, maj_128_n29,
         maj_128_n28, maj_128_n27, maj_128_n26, maj_128_n25, maj_128_n24,
         maj_128_n23, maj_128_n22, maj_128_n21, maj_128_n20, maj_128_n19,
         maj_128_n18, maj_129_n34, maj_129_n33, maj_129_n32, maj_129_n31,
         maj_129_n30, maj_129_n29, maj_129_n28, maj_129_n27, maj_129_n26,
         maj_129_n25, maj_129_n24, maj_129_n23, maj_129_n22, maj_129_n21,
         maj_129_n20, maj_129_n19, maj_129_n18, maj_130_n34, maj_130_n33,
         maj_130_n32, maj_130_n31, maj_130_n30, maj_130_n29, maj_130_n28,
         maj_130_n27, maj_130_n26, maj_130_n25, maj_130_n24, maj_130_n23,
         maj_130_n22, maj_130_n21, maj_130_n20, maj_130_n19, maj_130_n18,
         maj_131_n34, maj_131_n33, maj_131_n32, maj_131_n31, maj_131_n30,
         maj_131_n29, maj_131_n28, maj_131_n27, maj_131_n26, maj_131_n25,
         maj_131_n24, maj_131_n23, maj_131_n22, maj_131_n21, maj_131_n20,
         maj_131_n19, maj_131_n18, maj_132_n34, maj_132_n33, maj_132_n32,
         maj_132_n31, maj_132_n30, maj_132_n29, maj_132_n28, maj_132_n27,
         maj_132_n26, maj_132_n25, maj_132_n24, maj_132_n23, maj_132_n22,
         maj_132_n21, maj_132_n20, maj_132_n19, maj_132_n18, maj_133_n34,
         maj_133_n33, maj_133_n32, maj_133_n31, maj_133_n30, maj_133_n29,
         maj_133_n28, maj_133_n27, maj_133_n26, maj_133_n25, maj_133_n24,
         maj_133_n23, maj_133_n22, maj_133_n21, maj_133_n20, maj_133_n19,
         maj_133_n18, maj_134_n34, maj_134_n33, maj_134_n32, maj_134_n31,
         maj_134_n30, maj_134_n29, maj_134_n28, maj_134_n27, maj_134_n26,
         maj_134_n25, maj_134_n24, maj_134_n23, maj_134_n22, maj_134_n21,
         maj_134_n20, maj_134_n19, maj_134_n18, maj_135_n34, maj_135_n33,
         maj_135_n32, maj_135_n31, maj_135_n30, maj_135_n29, maj_135_n28,
         maj_135_n27, maj_135_n26, maj_135_n25, maj_135_n24, maj_135_n23,
         maj_135_n22, maj_135_n21, maj_135_n20, maj_135_n19, maj_135_n18,
         maj_136_n34, maj_136_n33, maj_136_n32, maj_136_n31, maj_136_n30,
         maj_136_n29, maj_136_n28, maj_136_n27, maj_136_n26, maj_136_n25,
         maj_136_n24, maj_136_n23, maj_136_n22, maj_136_n21, maj_136_n20,
         maj_136_n19, maj_136_n18, maj_137_n34, maj_137_n33, maj_137_n32,
         maj_137_n31, maj_137_n30, maj_137_n29, maj_137_n28, maj_137_n27,
         maj_137_n26, maj_137_n25, maj_137_n24, maj_137_n23, maj_137_n22,
         maj_137_n21, maj_137_n20, maj_137_n19, maj_137_n18, maj_138_n34,
         maj_138_n33, maj_138_n32, maj_138_n31, maj_138_n30, maj_138_n29,
         maj_138_n28, maj_138_n27, maj_138_n26, maj_138_n25, maj_138_n24,
         maj_138_n23, maj_138_n22, maj_138_n21, maj_138_n20, maj_138_n19,
         maj_138_n18, maj_139_n34, maj_139_n33, maj_139_n32, maj_139_n31,
         maj_139_n30, maj_139_n29, maj_139_n28, maj_139_n27, maj_139_n26,
         maj_139_n25, maj_139_n24, maj_139_n23, maj_139_n22, maj_139_n21,
         maj_139_n20, maj_139_n19, maj_139_n18, maj_140_n34, maj_140_n33,
         maj_140_n32, maj_140_n31, maj_140_n30, maj_140_n29, maj_140_n28,
         maj_140_n27, maj_140_n26, maj_140_n25, maj_140_n24, maj_140_n23,
         maj_140_n22, maj_140_n21, maj_140_n20, maj_140_n19, maj_140_n18,
         maj_141_n34, maj_141_n33, maj_141_n32, maj_141_n31, maj_141_n30,
         maj_141_n29, maj_141_n28, maj_141_n27, maj_141_n26, maj_141_n25,
         maj_141_n24, maj_141_n23, maj_141_n22, maj_141_n21, maj_141_n20,
         maj_141_n19, maj_141_n18, maj_142_n34, maj_142_n33, maj_142_n32,
         maj_142_n31, maj_142_n30, maj_142_n29, maj_142_n28, maj_142_n27,
         maj_142_n26, maj_142_n25, maj_142_n24, maj_142_n23, maj_142_n22,
         maj_142_n21, maj_142_n20, maj_142_n19, maj_142_n18, maj_143_n34,
         maj_143_n33, maj_143_n32, maj_143_n31, maj_143_n30, maj_143_n29,
         maj_143_n28, maj_143_n27, maj_143_n26, maj_143_n25, maj_143_n24,
         maj_143_n23, maj_143_n22, maj_143_n21, maj_143_n20, maj_143_n19,
         maj_143_n18, maj_144_n34, maj_144_n33, maj_144_n32, maj_144_n31,
         maj_144_n30, maj_144_n29, maj_144_n28, maj_144_n27, maj_144_n26,
         maj_144_n25, maj_144_n24, maj_144_n23, maj_144_n22, maj_144_n21,
         maj_144_n20, maj_144_n19, maj_144_n18, maj_145_n34, maj_145_n33,
         maj_145_n32, maj_145_n31, maj_145_n30, maj_145_n29, maj_145_n28,
         maj_145_n27, maj_145_n26, maj_145_n25, maj_145_n24, maj_145_n23,
         maj_145_n22, maj_145_n21, maj_145_n20, maj_145_n19, maj_145_n18,
         maj_146_n34, maj_146_n33, maj_146_n32, maj_146_n31, maj_146_n30,
         maj_146_n29, maj_146_n28, maj_146_n27, maj_146_n26, maj_146_n25,
         maj_146_n24, maj_146_n23, maj_146_n22, maj_146_n21, maj_146_n20,
         maj_146_n19, maj_146_n18, maj_147_n34, maj_147_n33, maj_147_n32,
         maj_147_n31, maj_147_n30, maj_147_n29, maj_147_n28, maj_147_n27,
         maj_147_n26, maj_147_n25, maj_147_n24, maj_147_n23, maj_147_n22,
         maj_147_n21, maj_147_n20, maj_147_n19, maj_147_n18, maj_148_n34,
         maj_148_n33, maj_148_n32, maj_148_n31, maj_148_n30, maj_148_n29,
         maj_148_n28, maj_148_n27, maj_148_n26, maj_148_n25, maj_148_n24,
         maj_148_n23, maj_148_n22, maj_148_n21, maj_148_n20, maj_148_n19,
         maj_148_n18, maj_149_n34, maj_149_n33, maj_149_n32, maj_149_n31,
         maj_149_n30, maj_149_n29, maj_149_n28, maj_149_n27, maj_149_n26,
         maj_149_n25, maj_149_n24, maj_149_n23, maj_149_n22, maj_149_n21,
         maj_149_n20, maj_149_n19, maj_149_n18, maj_150_n34, maj_150_n33,
         maj_150_n32, maj_150_n31, maj_150_n30, maj_150_n29, maj_150_n28,
         maj_150_n27, maj_150_n26, maj_150_n25, maj_150_n24, maj_150_n23,
         maj_150_n22, maj_150_n21, maj_150_n20, maj_150_n19, maj_150_n18,
         maj_151_n34, maj_151_n33, maj_151_n32, maj_151_n31, maj_151_n30,
         maj_151_n29, maj_151_n28, maj_151_n27, maj_151_n26, maj_151_n25,
         maj_151_n24, maj_151_n23, maj_151_n22, maj_151_n21, maj_151_n20,
         maj_151_n19, maj_151_n18, maj_152_n34, maj_152_n33, maj_152_n32,
         maj_152_n31, maj_152_n30, maj_152_n29, maj_152_n28, maj_152_n27,
         maj_152_n26, maj_152_n25, maj_152_n24, maj_152_n23, maj_152_n22,
         maj_152_n21, maj_152_n20, maj_152_n19, maj_152_n18, maj_153_n34,
         maj_153_n33, maj_153_n32, maj_153_n31, maj_153_n30, maj_153_n29,
         maj_153_n28, maj_153_n27, maj_153_n26, maj_153_n25, maj_153_n24,
         maj_153_n23, maj_153_n22, maj_153_n21, maj_153_n20, maj_153_n19,
         maj_153_n18, maj_154_n34, maj_154_n33, maj_154_n32, maj_154_n31,
         maj_154_n30, maj_154_n29, maj_154_n28, maj_154_n27, maj_154_n26,
         maj_154_n25, maj_154_n24, maj_154_n23, maj_154_n22, maj_154_n21,
         maj_154_n20, maj_154_n19, maj_154_n18, maj_155_n34, maj_155_n33,
         maj_155_n32, maj_155_n31, maj_155_n30, maj_155_n29, maj_155_n28,
         maj_155_n27, maj_155_n26, maj_155_n25, maj_155_n24, maj_155_n23,
         maj_155_n22, maj_155_n21, maj_155_n20, maj_155_n19, maj_155_n18,
         maj_156_n34, maj_156_n33, maj_156_n32, maj_156_n31, maj_156_n30,
         maj_156_n29, maj_156_n28, maj_156_n27, maj_156_n26, maj_156_n25,
         maj_156_n24, maj_156_n23, maj_156_n22, maj_156_n21, maj_156_n20,
         maj_156_n19, maj_156_n18, maj_157_n34, maj_157_n33, maj_157_n32,
         maj_157_n31, maj_157_n30, maj_157_n29, maj_157_n28, maj_157_n27,
         maj_157_n26, maj_157_n25, maj_157_n24, maj_157_n23, maj_157_n22,
         maj_157_n21, maj_157_n20, maj_157_n19, maj_157_n18, maj_158_n34,
         maj_158_n33, maj_158_n32, maj_158_n31, maj_158_n30, maj_158_n29,
         maj_158_n28, maj_158_n27, maj_158_n26, maj_158_n25, maj_158_n24,
         maj_158_n23, maj_158_n22, maj_158_n21, maj_158_n20, maj_158_n19,
         maj_158_n18, maj_159_n34, maj_159_n33, maj_159_n32, maj_159_n31,
         maj_159_n30, maj_159_n29, maj_159_n28, maj_159_n27, maj_159_n26,
         maj_159_n25, maj_159_n24, maj_159_n23, maj_159_n22, maj_159_n21,
         maj_159_n20, maj_159_n19, maj_159_n18, maj_160_n34, maj_160_n33,
         maj_160_n32, maj_160_n31, maj_160_n30, maj_160_n29, maj_160_n28,
         maj_160_n27, maj_160_n26, maj_160_n25, maj_160_n24, maj_160_n23,
         maj_160_n22, maj_160_n21, maj_160_n20, maj_160_n19, maj_160_n18,
         maj_161_n34, maj_161_n33, maj_161_n32, maj_161_n31, maj_161_n30,
         maj_161_n29, maj_161_n28, maj_161_n27, maj_161_n26, maj_161_n25,
         maj_161_n24, maj_161_n23, maj_161_n22, maj_161_n21, maj_161_n20,
         maj_161_n19, maj_161_n18, maj_162_n34, maj_162_n33, maj_162_n32,
         maj_162_n31, maj_162_n30, maj_162_n29, maj_162_n28, maj_162_n27,
         maj_162_n26, maj_162_n25, maj_162_n24, maj_162_n23, maj_162_n22,
         maj_162_n21, maj_162_n20, maj_162_n19, maj_162_n18, maj_163_n34,
         maj_163_n33, maj_163_n32, maj_163_n31, maj_163_n30, maj_163_n29,
         maj_163_n28, maj_163_n27, maj_163_n26, maj_163_n25, maj_163_n24,
         maj_163_n23, maj_163_n22, maj_163_n21, maj_163_n20, maj_163_n19,
         maj_163_n18, maj_164_n34, maj_164_n33, maj_164_n32, maj_164_n31,
         maj_164_n30, maj_164_n29, maj_164_n28, maj_164_n27, maj_164_n26,
         maj_164_n25, maj_164_n24, maj_164_n23, maj_164_n22, maj_164_n21,
         maj_164_n20, maj_164_n19, maj_164_n18, maj_165_n34, maj_165_n33,
         maj_165_n32, maj_165_n31, maj_165_n30, maj_165_n29, maj_165_n28,
         maj_165_n27, maj_165_n26, maj_165_n25, maj_165_n24, maj_165_n23,
         maj_165_n22, maj_165_n21, maj_165_n20, maj_165_n19, maj_165_n18,
         maj_166_n34, maj_166_n33, maj_166_n32, maj_166_n31, maj_166_n30,
         maj_166_n29, maj_166_n28, maj_166_n27, maj_166_n26, maj_166_n25,
         maj_166_n24, maj_166_n23, maj_166_n22, maj_166_n21, maj_166_n20,
         maj_166_n19, maj_166_n18, maj_167_n34, maj_167_n33, maj_167_n32,
         maj_167_n31, maj_167_n30, maj_167_n29, maj_167_n28, maj_167_n27,
         maj_167_n26, maj_167_n25, maj_167_n24, maj_167_n23, maj_167_n22,
         maj_167_n21, maj_167_n20, maj_167_n19, maj_167_n18;
  wire   [6:0] u_0_0;
  wire   [6:0] v_0_0;
  wire   [6:0] u_0_1;
  wire   [6:0] v_0_1;
  wire   [6:0] u_1_0;
  wire   [6:0] v_1_0;
  wire   [6:0] u_1_1;
  wire   [6:0] v_1_1;
  wire   [6:0] u_2_0;
  wire   [6:0] v_2_0;
  wire   [6:0] u_2_1;
  wire   [6:0] v_2_1;
  wire   [6:0] temp_0_0;
  wire   [6:0] a_reg_0;
  wire   [6:0] v_reg_0_0;
  wire   [6:0] u_reg_0_0;
  wire   [6:0] v_reg_0_1;
  wire   [6:0] u_reg_0_1;
  wire   [6:0] temp_0_1;
  wire   [6:0] a_reg_1;
  wire   [6:0] v_reg_1_0;
  wire   [6:0] u_reg_1_0;
  wire   [6:0] v_reg_1_1;
  wire   [6:0] u_reg_1_1;
  wire   [6:0] temp_0_2;
  wire   [6:0] a_reg_2;
  wire   [6:0] v_reg_2_0;
  wire   [6:0] u_reg_2_0;
  wire   [6:0] v_reg_2_1;
  wire   [6:0] u_reg_2_1;

  DFF_X1 v_reg_1_0_reg_6_ ( .D(maj_161_port_o), .CK(clk), .Q(v_reg_1_0[6]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_5_ ( .D(maj_149_port_o), .CK(clk), .Q(v_reg_1_0[5]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_4_ ( .D(maj_137_port_o), .CK(clk), .Q(v_reg_1_0[4]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_3_ ( .D(maj_125_port_o), .CK(clk), .Q(v_reg_1_0[3]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_2_ ( .D(maj_113_port_o), .CK(clk), .Q(v_reg_1_0[2]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_1_ ( .D(maj_101_port_o), .CK(clk), .Q(v_reg_1_0[1]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_0_ ( .D(maj_89_port_o), .CK(clk), .Q(v_reg_1_0[0]), 
        .QN() );
  DFF_X1 a_reg_2_reg_6_ ( .D(port_a_2[6]), .CK(clk), .Q(a_reg_2[6]), .QN() );
  DFF_X1 a_reg_2_reg_5_ ( .D(port_a_2[5]), .CK(clk), .Q(a_reg_2[5]), .QN() );
  DFF_X1 a_reg_2_reg_4_ ( .D(port_a_2[4]), .CK(clk), .Q(a_reg_2[4]), .QN() );
  DFF_X1 a_reg_2_reg_3_ ( .D(port_a_2[3]), .CK(clk), .Q(a_reg_2[3]), .QN() );
  DFF_X1 a_reg_2_reg_2_ ( .D(port_a_2[2]), .CK(clk), .Q(a_reg_2[2]), .QN() );
  DFF_X1 a_reg_2_reg_1_ ( .D(port_a_2[1]), .CK(clk), .Q(a_reg_2[1]), .QN() );
  DFF_X1 a_reg_2_reg_0_ ( .D(port_a_2[0]), .CK(clk), .Q(a_reg_2[0]), .QN() );
  DFF_X1 u_reg_0_0_reg_6_ ( .D(maj_156_port_o), .CK(clk), .Q(u_reg_0_0[6]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_5_ ( .D(maj_144_port_o), .CK(clk), .Q(u_reg_0_0[5]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_4_ ( .D(maj_132_port_o), .CK(clk), .Q(u_reg_0_0[4]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_3_ ( .D(maj_120_port_o), .CK(clk), .Q(u_reg_0_0[3]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_2_ ( .D(maj_108_port_o), .CK(clk), .Q(u_reg_0_0[2]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_1_ ( .D(maj_96_port_o), .CK(clk), .Q(u_reg_0_0[1]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_0_ ( .D(maj_84_port_o), .CK(clk), .Q(u_reg_0_0[0]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_6_ ( .D(maj_159_port_o), .CK(clk), .Q(v_reg_0_1[6]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_5_ ( .D(maj_147_port_o), .CK(clk), .Q(v_reg_0_1[5]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_4_ ( .D(maj_135_port_o), .CK(clk), .Q(v_reg_0_1[4]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_3_ ( .D(maj_123_port_o), .CK(clk), .Q(v_reg_0_1[3]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_2_ ( .D(maj_111_port_o), .CK(clk), .Q(v_reg_0_1[2]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_1_ ( .D(maj_99_port_o), .CK(clk), .Q(v_reg_0_1[1]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_0_ ( .D(maj_87_port_o), .CK(clk), .Q(v_reg_0_1[0]), 
        .QN() );
  DFF_X1 ab_reg_2_reg_6_ ( .D(N20), .CK(clk), .Q(temp_0_2[6]), .QN() );
  DFF_X1 ab_reg_2_reg_5_ ( .D(N17), .CK(clk), .Q(temp_0_2[5]), .QN() );
  DFF_X1 ab_reg_2_reg_4_ ( .D(N14), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 ab_reg_2_reg_3_ ( .D(N11), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 ab_reg_2_reg_2_ ( .D(N8), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 ab_reg_2_reg_1_ ( .D(N5), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 ab_reg_2_reg_0_ ( .D(N2), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 u_reg_0_1_reg_6_ ( .D(maj_158_port_o), .CK(clk), .Q(u_reg_0_1[6]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_5_ ( .D(maj_146_port_o), .CK(clk), .Q(u_reg_0_1[5]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_4_ ( .D(maj_134_port_o), .CK(clk), .Q(u_reg_0_1[4]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_3_ ( .D(maj_122_port_o), .CK(clk), .Q(u_reg_0_1[3]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_2_ ( .D(maj_110_port_o), .CK(clk), .Q(u_reg_0_1[2]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_1_ ( .D(maj_98_port_o), .CK(clk), .Q(u_reg_0_1[1]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_0_ ( .D(maj_86_port_o), .CK(clk), .Q(u_reg_0_1[0]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_6_ ( .D(maj_157_port_o), .CK(clk), .Q(v_reg_0_0[6]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_5_ ( .D(maj_145_port_o), .CK(clk), .Q(v_reg_0_0[5]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_4_ ( .D(maj_133_port_o), .CK(clk), .Q(v_reg_0_0[4]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_3_ ( .D(maj_121_port_o), .CK(clk), .Q(v_reg_0_0[3]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_2_ ( .D(maj_109_port_o), .CK(clk), .Q(v_reg_0_0[2]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_1_ ( .D(maj_97_port_o), .CK(clk), .Q(v_reg_0_0[1]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_0_ ( .D(maj_85_port_o), .CK(clk), .Q(v_reg_0_0[0]), 
        .QN() );
  DFF_X1 a_reg_1_reg_6_ ( .D(port_a_1[6]), .CK(clk), .Q(a_reg_1[6]), .QN() );
  DFF_X1 a_reg_1_reg_5_ ( .D(port_a_1[5]), .CK(clk), .Q(a_reg_1[5]), .QN() );
  DFF_X1 a_reg_1_reg_4_ ( .D(port_a_1[4]), .CK(clk), .Q(a_reg_1[4]), .QN() );
  DFF_X1 a_reg_1_reg_3_ ( .D(port_a_1[3]), .CK(clk), .Q(a_reg_1[3]), .QN() );
  DFF_X1 a_reg_1_reg_2_ ( .D(port_a_1[2]), .CK(clk), .Q(a_reg_1[2]), .QN() );
  DFF_X1 a_reg_1_reg_1_ ( .D(port_a_1[1]), .CK(clk), .Q(a_reg_1[1]), .QN() );
  DFF_X1 a_reg_1_reg_0_ ( .D(port_a_1[0]), .CK(clk), .Q(a_reg_1[0]), .QN() );
  DFF_X1 u_reg_1_0_reg_6_ ( .D(maj_160_port_o), .CK(clk), .Q(u_reg_1_0[6]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_5_ ( .D(maj_148_port_o), .CK(clk), .Q(u_reg_1_0[5]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_4_ ( .D(maj_136_port_o), .CK(clk), .Q(u_reg_1_0[4]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_3_ ( .D(maj_124_port_o), .CK(clk), .Q(u_reg_1_0[3]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_2_ ( .D(maj_112_port_o), .CK(clk), .Q(u_reg_1_0[2]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_1_ ( .D(maj_100_port_o), .CK(clk), .Q(u_reg_1_0[1]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_0_ ( .D(maj_88_port_o), .CK(clk), .Q(u_reg_1_0[0]), 
        .QN() );
  DFF_X1 ab_reg_1_reg_6_ ( .D(N19), .CK(clk), .Q(temp_0_1[6]), .QN() );
  DFF_X1 ab_reg_1_reg_5_ ( .D(N16), .CK(clk), .Q(temp_0_1[5]), .QN() );
  DFF_X1 ab_reg_1_reg_4_ ( .D(N13), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 ab_reg_1_reg_3_ ( .D(N10), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 ab_reg_1_reg_2_ ( .D(N7), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 ab_reg_1_reg_1_ ( .D(N4), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 ab_reg_1_reg_0_ ( .D(N1), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 a_reg_0_reg_6_ ( .D(port_a_0[6]), .CK(clk), .Q(a_reg_0[6]), .QN() );
  DFF_X1 a_reg_0_reg_5_ ( .D(port_a_0[5]), .CK(clk), .Q(a_reg_0[5]), .QN() );
  DFF_X1 a_reg_0_reg_4_ ( .D(port_a_0[4]), .CK(clk), .Q(a_reg_0[4]), .QN() );
  DFF_X1 a_reg_0_reg_3_ ( .D(port_a_0[3]), .CK(clk), .Q(a_reg_0[3]), .QN() );
  DFF_X1 a_reg_0_reg_2_ ( .D(port_a_0[2]), .CK(clk), .Q(a_reg_0[2]), .QN() );
  DFF_X1 a_reg_0_reg_1_ ( .D(port_a_0[1]), .CK(clk), .Q(a_reg_0[1]), .QN() );
  DFF_X1 a_reg_0_reg_0_ ( .D(port_a_0[0]), .CK(clk), .Q(a_reg_0[0]), .QN() );
  DFF_X1 ab_reg_0_reg_6_ ( .D(N18), .CK(clk), .Q(temp_0_0[6]), .QN() );
  DFF_X1 ab_reg_0_reg_5_ ( .D(N15), .CK(clk), .Q(temp_0_0[5]), .QN() );
  DFF_X1 ab_reg_0_reg_4_ ( .D(N12), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 ab_reg_0_reg_3_ ( .D(N9), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 ab_reg_0_reg_2_ ( .D(N6), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 ab_reg_0_reg_1_ ( .D(N3), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 ab_reg_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 v_reg_2_1_reg_6_ ( .D(maj_167_port_o), .CK(clk), .Q(v_reg_2_1[6]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_5_ ( .D(maj_155_port_o), .CK(clk), .Q(v_reg_2_1[5]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_4_ ( .D(maj_143_port_o), .CK(clk), .Q(v_reg_2_1[4]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_3_ ( .D(maj_131_port_o), .CK(clk), .Q(v_reg_2_1[3]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_2_ ( .D(maj_119_port_o), .CK(clk), .Q(v_reg_2_1[2]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_1_ ( .D(maj_107_port_o), .CK(clk), .Q(v_reg_2_1[1]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_0_ ( .D(maj_95_port_o), .CK(clk), .Q(v_reg_2_1[0]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_6_ ( .D(maj_166_port_o), .CK(clk), .Q(u_reg_2_1[6]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_5_ ( .D(maj_154_port_o), .CK(clk), .Q(u_reg_2_1[5]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_4_ ( .D(maj_142_port_o), .CK(clk), .Q(u_reg_2_1[4]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_3_ ( .D(maj_130_port_o), .CK(clk), .Q(u_reg_2_1[3]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_2_ ( .D(maj_118_port_o), .CK(clk), .Q(u_reg_2_1[2]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_1_ ( .D(maj_106_port_o), .CK(clk), .Q(u_reg_2_1[1]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_0_ ( .D(maj_94_port_o), .CK(clk), .Q(u_reg_2_1[0]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_6_ ( .D(maj_165_port_o), .CK(clk), .Q(v_reg_2_0[6]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_5_ ( .D(maj_153_port_o), .CK(clk), .Q(v_reg_2_0[5]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_4_ ( .D(maj_141_port_o), .CK(clk), .Q(v_reg_2_0[4]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_3_ ( .D(maj_129_port_o), .CK(clk), .Q(v_reg_2_0[3]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_2_ ( .D(maj_117_port_o), .CK(clk), .Q(v_reg_2_0[2]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_1_ ( .D(maj_105_port_o), .CK(clk), .Q(v_reg_2_0[1]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_0_ ( .D(maj_93_port_o), .CK(clk), .Q(v_reg_2_0[0]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_6_ ( .D(maj_164_port_o), .CK(clk), .Q(u_reg_2_0[6]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_5_ ( .D(maj_152_port_o), .CK(clk), .Q(u_reg_2_0[5]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_4_ ( .D(maj_140_port_o), .CK(clk), .Q(u_reg_2_0[4]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_3_ ( .D(maj_128_port_o), .CK(clk), .Q(u_reg_2_0[3]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_2_ ( .D(maj_116_port_o), .CK(clk), .Q(u_reg_2_0[2]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_1_ ( .D(maj_104_port_o), .CK(clk), .Q(u_reg_2_0[1]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_0_ ( .D(maj_92_port_o), .CK(clk), .Q(u_reg_2_0[0]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_6_ ( .D(maj_163_port_o), .CK(clk), .Q(v_reg_1_1[6]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_5_ ( .D(maj_151_port_o), .CK(clk), .Q(v_reg_1_1[5]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_4_ ( .D(maj_139_port_o), .CK(clk), .Q(v_reg_1_1[4]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_3_ ( .D(maj_127_port_o), .CK(clk), .Q(v_reg_1_1[3]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_2_ ( .D(maj_115_port_o), .CK(clk), .Q(v_reg_1_1[2]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_1_ ( .D(maj_103_port_o), .CK(clk), .Q(v_reg_1_1[1]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_0_ ( .D(maj_91_port_o), .CK(clk), .Q(v_reg_1_1[0]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_6_ ( .D(maj_162_port_o), .CK(clk), .Q(u_reg_1_1[6]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_5_ ( .D(maj_150_port_o), .CK(clk), .Q(u_reg_1_1[5]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_4_ ( .D(maj_138_port_o), .CK(clk), .Q(u_reg_1_1[4]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_3_ ( .D(maj_126_port_o), .CK(clk), .Q(u_reg_1_1[3]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_2_ ( .D(maj_114_port_o), .CK(clk), .Q(u_reg_1_1[2]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_1_ ( .D(maj_102_port_o), .CK(clk), .Q(u_reg_1_1[1]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_0_ ( .D(maj_90_port_o), .CK(clk), .Q(u_reg_1_1[0]), 
        .QN() );
  XNOR2_X1 U171 ( .A(u_reg_2_1[0]), .B(u_reg_2_0[0]), .ZN(n56) );
  XNOR2_X1 U172 ( .A(u_reg_2_1[1]), .B(u_reg_2_0[1]), .ZN(n51) );
  XNOR2_X1 U173 ( .A(u_reg_2_1[2]), .B(u_reg_2_0[2]), .ZN(n46) );
  XNOR2_X1 U174 ( .A(u_reg_2_1[3]), .B(u_reg_2_0[3]), .ZN(n41) );
  XNOR2_X1 U175 ( .A(u_reg_2_1[4]), .B(u_reg_2_0[4]), .ZN(n36) );
  XNOR2_X1 U176 ( .A(u_reg_2_1[5]), .B(u_reg_2_0[5]), .ZN(n31) );
  XNOR2_X1 U177 ( .A(u_reg_2_1[6]), .B(u_reg_2_0[6]), .ZN(n26) );
  XNOR2_X1 U178 ( .A(u_reg_1_1[0]), .B(u_reg_1_0[0]), .ZN(n91) );
  XNOR2_X1 U179 ( .A(u_reg_1_1[1]), .B(u_reg_1_0[1]), .ZN(n86) );
  XNOR2_X1 U180 ( .A(u_reg_1_1[2]), .B(u_reg_1_0[2]), .ZN(n81) );
  XNOR2_X1 U181 ( .A(u_reg_1_1[3]), .B(u_reg_1_0[3]), .ZN(n76) );
  XNOR2_X1 U182 ( .A(u_reg_1_1[4]), .B(u_reg_1_0[4]), .ZN(n71) );
  XNOR2_X1 U183 ( .A(u_reg_1_1[5]), .B(u_reg_1_0[5]), .ZN(n66) );
  XNOR2_X1 U184 ( .A(u_reg_1_1[6]), .B(u_reg_1_0[6]), .ZN(n61) );
  XNOR2_X1 U185 ( .A(u_reg_0_1[0]), .B(u_reg_0_0[0]), .ZN(n126) );
  XNOR2_X1 U186 ( .A(u_reg_0_1[1]), .B(u_reg_0_0[1]), .ZN(n121) );
  XNOR2_X1 U187 ( .A(u_reg_0_1[2]), .B(u_reg_0_0[2]), .ZN(n116) );
  XNOR2_X1 U188 ( .A(u_reg_0_1[3]), .B(u_reg_0_0[3]), .ZN(n111) );
  XNOR2_X1 U189 ( .A(u_reg_0_1[4]), .B(u_reg_0_0[4]), .ZN(n106) );
  XNOR2_X1 U190 ( .A(u_reg_0_1[5]), .B(u_reg_0_0[5]), .ZN(n101) );
  XNOR2_X1 U191 ( .A(u_reg_0_1[6]), .B(u_reg_0_0[6]), .ZN(n96) );
  XOR2_X1 U192 ( .A(n52), .B(n53), .Z(port_c_2[0]) );
  XNOR2_X1 U193 ( .A(n54), .B(n55), .ZN(n53) );
  XOR2_X1 U194 ( .A(n56), .B(temp_0_2[0]), .Z(n52) );
  NAND2_X1 U195 ( .A1(v_reg_2_1[0]), .A2(a_reg_2[0]), .ZN(n54) );
  XOR2_X1 U196 ( .A(n47), .B(n48), .Z(port_c_2[1]) );
  XNOR2_X1 U197 ( .A(n49), .B(n50), .ZN(n48) );
  XOR2_X1 U198 ( .A(n51), .B(temp_0_2[1]), .Z(n47) );
  NAND2_X1 U199 ( .A1(v_reg_2_1[1]), .A2(a_reg_2[1]), .ZN(n49) );
  XOR2_X1 U200 ( .A(n42), .B(n43), .Z(port_c_2[2]) );
  XNOR2_X1 U201 ( .A(n44), .B(n45), .ZN(n43) );
  XOR2_X1 U202 ( .A(n46), .B(temp_0_2[2]), .Z(n42) );
  NAND2_X1 U203 ( .A1(v_reg_2_1[2]), .A2(a_reg_2[2]), .ZN(n44) );
  XOR2_X1 U204 ( .A(n37), .B(n38), .Z(port_c_2[3]) );
  XNOR2_X1 U205 ( .A(n39), .B(n40), .ZN(n38) );
  XOR2_X1 U206 ( .A(n41), .B(temp_0_2[3]), .Z(n37) );
  NAND2_X1 U207 ( .A1(v_reg_2_1[3]), .A2(a_reg_2[3]), .ZN(n39) );
  XOR2_X1 U208 ( .A(n32), .B(n33), .Z(port_c_2[4]) );
  XNOR2_X1 U209 ( .A(n34), .B(n35), .ZN(n33) );
  XOR2_X1 U210 ( .A(n36), .B(temp_0_2[4]), .Z(n32) );
  NAND2_X1 U211 ( .A1(v_reg_2_1[4]), .A2(a_reg_2[4]), .ZN(n34) );
  XOR2_X1 U212 ( .A(n27), .B(n28), .Z(port_c_2[5]) );
  XNOR2_X1 U213 ( .A(n29), .B(n30), .ZN(n28) );
  XOR2_X1 U214 ( .A(n31), .B(temp_0_2[5]), .Z(n27) );
  NAND2_X1 U215 ( .A1(v_reg_2_1[5]), .A2(a_reg_2[5]), .ZN(n29) );
  XOR2_X1 U216 ( .A(n22), .B(n23), .Z(port_c_2[6]) );
  XNOR2_X1 U217 ( .A(n24), .B(n25), .ZN(n23) );
  XOR2_X1 U218 ( .A(n26), .B(temp_0_2[6]), .Z(n22) );
  NAND2_X1 U219 ( .A1(v_reg_2_1[6]), .A2(a_reg_2[6]), .ZN(n24) );
  XOR2_X1 U220 ( .A(n87), .B(n88), .Z(port_c_1[0]) );
  XNOR2_X1 U221 ( .A(n89), .B(n90), .ZN(n88) );
  XOR2_X1 U222 ( .A(n91), .B(temp_0_1[0]), .Z(n87) );
  NAND2_X1 U223 ( .A1(v_reg_1_1[0]), .A2(a_reg_1[0]), .ZN(n89) );
  XOR2_X1 U224 ( .A(n82), .B(n83), .Z(port_c_1[1]) );
  XNOR2_X1 U225 ( .A(n84), .B(n85), .ZN(n83) );
  XOR2_X1 U226 ( .A(n86), .B(temp_0_1[1]), .Z(n82) );
  NAND2_X1 U227 ( .A1(v_reg_1_1[1]), .A2(a_reg_1[1]), .ZN(n84) );
  XOR2_X1 U228 ( .A(n77), .B(n78), .Z(port_c_1[2]) );
  XNOR2_X1 U229 ( .A(n79), .B(n80), .ZN(n78) );
  XOR2_X1 U230 ( .A(n81), .B(temp_0_1[2]), .Z(n77) );
  NAND2_X1 U231 ( .A1(v_reg_1_1[2]), .A2(a_reg_1[2]), .ZN(n79) );
  XOR2_X1 U232 ( .A(n72), .B(n73), .Z(port_c_1[3]) );
  XNOR2_X1 U233 ( .A(n74), .B(n75), .ZN(n73) );
  XOR2_X1 U234 ( .A(n76), .B(temp_0_1[3]), .Z(n72) );
  NAND2_X1 U235 ( .A1(v_reg_1_1[3]), .A2(a_reg_1[3]), .ZN(n74) );
  XOR2_X1 U236 ( .A(n67), .B(n68), .Z(port_c_1[4]) );
  XNOR2_X1 U237 ( .A(n69), .B(n70), .ZN(n68) );
  XOR2_X1 U238 ( .A(n71), .B(temp_0_1[4]), .Z(n67) );
  NAND2_X1 U239 ( .A1(v_reg_1_1[4]), .A2(a_reg_1[4]), .ZN(n69) );
  XOR2_X1 U240 ( .A(n62), .B(n63), .Z(port_c_1[5]) );
  XNOR2_X1 U241 ( .A(n64), .B(n65), .ZN(n63) );
  XOR2_X1 U242 ( .A(n66), .B(temp_0_1[5]), .Z(n62) );
  NAND2_X1 U243 ( .A1(v_reg_1_1[5]), .A2(a_reg_1[5]), .ZN(n64) );
  XOR2_X1 U244 ( .A(n57), .B(n58), .Z(port_c_1[6]) );
  XNOR2_X1 U245 ( .A(n59), .B(n60), .ZN(n58) );
  XOR2_X1 U246 ( .A(n61), .B(temp_0_1[6]), .Z(n57) );
  NAND2_X1 U247 ( .A1(v_reg_1_1[6]), .A2(a_reg_1[6]), .ZN(n59) );
  XOR2_X1 U248 ( .A(n122), .B(n123), .Z(port_c_0[0]) );
  XNOR2_X1 U249 ( .A(n124), .B(n125), .ZN(n123) );
  XOR2_X1 U250 ( .A(n126), .B(temp_0_0[0]), .Z(n122) );
  NAND2_X1 U251 ( .A1(v_reg_0_1[0]), .A2(a_reg_0[0]), .ZN(n124) );
  XOR2_X1 U252 ( .A(n117), .B(n118), .Z(port_c_0[1]) );
  XNOR2_X1 U253 ( .A(n119), .B(n120), .ZN(n118) );
  XOR2_X1 U254 ( .A(n121), .B(temp_0_0[1]), .Z(n117) );
  NAND2_X1 U255 ( .A1(v_reg_0_1[1]), .A2(a_reg_0[1]), .ZN(n119) );
  XOR2_X1 U256 ( .A(n112), .B(n113), .Z(port_c_0[2]) );
  XNOR2_X1 U257 ( .A(n114), .B(n115), .ZN(n113) );
  XOR2_X1 U258 ( .A(n116), .B(temp_0_0[2]), .Z(n112) );
  NAND2_X1 U259 ( .A1(v_reg_0_1[2]), .A2(a_reg_0[2]), .ZN(n114) );
  XOR2_X1 U260 ( .A(n107), .B(n108), .Z(port_c_0[3]) );
  XNOR2_X1 U261 ( .A(n109), .B(n110), .ZN(n108) );
  XOR2_X1 U262 ( .A(n111), .B(temp_0_0[3]), .Z(n107) );
  NAND2_X1 U263 ( .A1(v_reg_0_1[3]), .A2(a_reg_0[3]), .ZN(n109) );
  XOR2_X1 U264 ( .A(n102), .B(n103), .Z(port_c_0[4]) );
  XNOR2_X1 U265 ( .A(n104), .B(n105), .ZN(n103) );
  XOR2_X1 U266 ( .A(n106), .B(temp_0_0[4]), .Z(n102) );
  NAND2_X1 U267 ( .A1(v_reg_0_1[4]), .A2(a_reg_0[4]), .ZN(n104) );
  XOR2_X1 U268 ( .A(n97), .B(n98), .Z(port_c_0[5]) );
  XNOR2_X1 U269 ( .A(n99), .B(n100), .ZN(n98) );
  XOR2_X1 U270 ( .A(n101), .B(temp_0_0[5]), .Z(n97) );
  NAND2_X1 U271 ( .A1(v_reg_0_1[5]), .A2(a_reg_0[5]), .ZN(n99) );
  XOR2_X1 U272 ( .A(n92), .B(n93), .Z(port_c_0[6]) );
  XNOR2_X1 U273 ( .A(n94), .B(n95), .ZN(n93) );
  XOR2_X1 U274 ( .A(n96), .B(temp_0_0[6]), .Z(n92) );
  NAND2_X1 U275 ( .A1(v_reg_0_1[6]), .A2(a_reg_0[6]), .ZN(n94) );
  NAND2_X1 U276 ( .A1(v_reg_2_0[0]), .A2(a_reg_2[0]), .ZN(n55) );
  NAND2_X1 U277 ( .A1(v_reg_2_0[1]), .A2(a_reg_2[1]), .ZN(n50) );
  NAND2_X1 U278 ( .A1(v_reg_2_0[2]), .A2(a_reg_2[2]), .ZN(n45) );
  NAND2_X1 U279 ( .A1(v_reg_2_0[3]), .A2(a_reg_2[3]), .ZN(n40) );
  NAND2_X1 U280 ( .A1(v_reg_2_0[4]), .A2(a_reg_2[4]), .ZN(n35) );
  NAND2_X1 U281 ( .A1(v_reg_2_0[5]), .A2(a_reg_2[5]), .ZN(n30) );
  NAND2_X1 U282 ( .A1(v_reg_2_0[6]), .A2(a_reg_2[6]), .ZN(n25) );
  NAND2_X1 U283 ( .A1(v_reg_1_0[0]), .A2(a_reg_1[0]), .ZN(n90) );
  NAND2_X1 U284 ( .A1(v_reg_1_0[1]), .A2(a_reg_1[1]), .ZN(n85) );
  NAND2_X1 U285 ( .A1(v_reg_1_0[2]), .A2(a_reg_1[2]), .ZN(n80) );
  NAND2_X1 U286 ( .A1(v_reg_1_0[3]), .A2(a_reg_1[3]), .ZN(n75) );
  NAND2_X1 U287 ( .A1(v_reg_1_0[4]), .A2(a_reg_1[4]), .ZN(n70) );
  NAND2_X1 U288 ( .A1(v_reg_1_0[5]), .A2(a_reg_1[5]), .ZN(n65) );
  NAND2_X1 U289 ( .A1(v_reg_1_0[6]), .A2(a_reg_1[6]), .ZN(n60) );
  NAND2_X1 U290 ( .A1(v_reg_0_0[0]), .A2(a_reg_0[0]), .ZN(n125) );
  NAND2_X1 U291 ( .A1(v_reg_0_0[1]), .A2(a_reg_0[1]), .ZN(n120) );
  NAND2_X1 U292 ( .A1(v_reg_0_0[2]), .A2(a_reg_0[2]), .ZN(n115) );
  NAND2_X1 U293 ( .A1(v_reg_0_0[3]), .A2(a_reg_0[3]), .ZN(n110) );
  NAND2_X1 U294 ( .A1(v_reg_0_0[4]), .A2(a_reg_0[4]), .ZN(n105) );
  NAND2_X1 U295 ( .A1(v_reg_0_0[5]), .A2(a_reg_0[5]), .ZN(n100) );
  NAND2_X1 U296 ( .A1(v_reg_0_0[6]), .A2(a_reg_0[6]), .ZN(n95) );
  INV_X1 U297 ( .A(port_a_2[2]), .ZN(n19) );
  INV_X1 U298 ( .A(port_a_2[1]), .ZN(n20) );
  INV_X1 U299 ( .A(port_a_2[0]), .ZN(n21) );
  INV_X1 U300 ( .A(port_a_2[5]), .ZN(n16) );
  INV_X1 U301 ( .A(port_a_2[4]), .ZN(n17) );
  INV_X1 U302 ( .A(port_a_2[3]), .ZN(n18) );
  INV_X1 U303 ( .A(port_a_2[6]), .ZN(n15) );
  INV_X1 U304 ( .A(port_a_1[2]), .ZN(n12) );
  INV_X1 U305 ( .A(port_a_1[1]), .ZN(n13) );
  INV_X1 U306 ( .A(port_a_1[0]), .ZN(n14) );
  INV_X1 U307 ( .A(port_a_1[5]), .ZN(n9) );
  INV_X1 U308 ( .A(port_a_1[4]), .ZN(n10) );
  INV_X1 U309 ( .A(port_a_1[3]), .ZN(n11) );
  INV_X1 U310 ( .A(port_a_1[6]), .ZN(n8) );
  INV_X1 U311 ( .A(port_a_0[2]), .ZN(n5) );
  INV_X1 U312 ( .A(port_a_0[1]), .ZN(n6) );
  INV_X1 U313 ( .A(port_a_0[0]), .ZN(n7) );
  INV_X1 U314 ( .A(port_a_0[5]), .ZN(n2) );
  INV_X1 U315 ( .A(port_a_0[4]), .ZN(n3) );
  INV_X1 U316 ( .A(port_a_0[3]), .ZN(n4) );
  INV_X1 U317 ( .A(port_a_0[6]), .ZN(n1) );
  AND2_X1 U318 ( .A1(port_b_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U319 ( .A1(port_b_0[1]), .A2(port_a_0[1]), .ZN(N3) );
  AND2_X1 U320 ( .A1(port_b_0[2]), .A2(port_a_0[2]), .ZN(N6) );
  AND2_X1 U321 ( .A1(port_b_0[3]), .A2(port_a_0[3]), .ZN(N9) );
  AND2_X1 U322 ( .A1(port_b_0[4]), .A2(port_a_0[4]), .ZN(N12) );
  AND2_X1 U323 ( .A1(port_b_0[5]), .A2(port_a_0[5]), .ZN(N15) );
  AND2_X1 U324 ( .A1(port_b_0[6]), .A2(port_a_0[6]), .ZN(N18) );
  AND2_X1 U325 ( .A1(port_b_1[0]), .A2(port_a_1[0]), .ZN(N1) );
  AND2_X1 U326 ( .A1(port_b_1[1]), .A2(port_a_1[1]), .ZN(N4) );
  AND2_X1 U327 ( .A1(port_b_1[2]), .A2(port_a_1[2]), .ZN(N7) );
  AND2_X1 U328 ( .A1(port_b_1[3]), .A2(port_a_1[3]), .ZN(N10) );
  AND2_X1 U329 ( .A1(port_b_1[4]), .A2(port_a_1[4]), .ZN(N13) );
  AND2_X1 U330 ( .A1(port_b_1[5]), .A2(port_a_1[5]), .ZN(N16) );
  AND2_X1 U331 ( .A1(port_b_1[6]), .A2(port_a_1[6]), .ZN(N19) );
  AND2_X1 U332 ( .A1(port_b_2[0]), .A2(port_a_2[0]), .ZN(N2) );
  AND2_X1 U333 ( .A1(port_b_2[1]), .A2(port_a_2[1]), .ZN(N5) );
  AND2_X1 U334 ( .A1(port_b_2[2]), .A2(port_a_2[2]), .ZN(N8) );
  AND2_X1 U335 ( .A1(port_b_2[3]), .A2(port_a_2[3]), .ZN(N11) );
  AND2_X1 U336 ( .A1(port_b_2[4]), .A2(port_a_2[4]), .ZN(N14) );
  AND2_X1 U337 ( .A1(port_b_2[5]), .A2(port_a_2[5]), .ZN(N17) );
  AND2_X1 U338 ( .A1(port_b_2[6]), .A2(port_a_2[6]), .ZN(N20) );
  AND2_X1 simpleAnd_42_U1 ( .A1(port_rand_mul[0]), .A2(n7), .ZN(
        simpleAnd_42_port_z) );
  XOR2_X2 simpleXor_84_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_42_port_z), .Z(
        u_0_0[0]) );
  XOR2_X2 simpleXor_85_U1 ( .A(port_rand_mul[0]), .B(port_b_1[0]), .Z(v_0_0[0]) );
  AND2_X1 simpleAnd_43_U1 ( .A1(port_rand_mul[1]), .A2(n7), .ZN(
        simpleAnd_43_port_z) );
  XOR2_X2 simpleXor_86_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_43_port_z), .Z(
        u_0_1[0]) );
  XOR2_X2 simpleXor_87_U1 ( .A(port_rand_mul[1]), .B(port_b_2[0]), .Z(v_0_1[0]) );
  AND2_X1 simpleAnd_44_U1 ( .A1(port_rand_mul[0]), .A2(n14), .ZN(
        simpleAnd_44_port_z) );
  XOR2_X2 simpleXor_88_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_44_port_z), .Z(
        u_1_0[0]) );
  XOR2_X2 simpleXor_89_U1 ( .A(port_rand_mul[0]), .B(port_b_0[0]), .Z(v_1_0[0]) );
  AND2_X1 simpleAnd_45_U1 ( .A1(port_rand_mul[2]), .A2(n14), .ZN(
        simpleAnd_45_port_z) );
  XOR2_X2 simpleXor_90_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_45_port_z), .Z(
        u_1_1[0]) );
  XOR2_X2 simpleXor_91_U1 ( .A(port_rand_mul[2]), .B(port_b_2[0]), .Z(v_1_1[0]) );
  AND2_X1 simpleAnd_46_U1 ( .A1(port_rand_mul[1]), .A2(n21), .ZN(
        simpleAnd_46_port_z) );
  XOR2_X2 simpleXor_92_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_46_port_z), .Z(
        u_2_0[0]) );
  XOR2_X2 simpleXor_93_U1 ( .A(port_rand_mul[1]), .B(port_b_0[0]), .Z(v_2_0[0]) );
  AND2_X1 simpleAnd_47_U1 ( .A1(port_rand_mul[2]), .A2(n21), .ZN(
        simpleAnd_47_port_z) );
  XOR2_X2 simpleXor_94_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_47_port_z), .Z(
        u_2_1[0]) );
  XOR2_X2 simpleXor_95_U1 ( .A(port_rand_mul[2]), .B(port_b_1[0]), .Z(v_2_1[0]) );
  AND2_X1 simpleAnd_48_U1 ( .A1(port_rand_mul[0]), .A2(n6), .ZN(
        simpleAnd_48_port_z) );
  XOR2_X2 simpleXor_96_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_48_port_z), .Z(
        u_0_0[1]) );
  XOR2_X2 simpleXor_97_U1 ( .A(port_rand_mul[0]), .B(port_b_1[1]), .Z(v_0_0[1]) );
  AND2_X1 simpleAnd_49_U1 ( .A1(port_rand_mul[1]), .A2(n6), .ZN(
        simpleAnd_49_port_z) );
  XOR2_X2 simpleXor_98_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_49_port_z), .Z(
        u_0_1[1]) );
  XOR2_X2 simpleXor_99_U1 ( .A(port_rand_mul[1]), .B(port_b_2[1]), .Z(v_0_1[1]) );
  AND2_X1 simpleAnd_50_U1 ( .A1(port_rand_mul[0]), .A2(n13), .ZN(
        simpleAnd_50_port_z) );
  XOR2_X2 simpleXor_100_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_50_port_z), 
        .Z(u_1_0[1]) );
  XOR2_X2 simpleXor_101_U1 ( .A(port_rand_mul[0]), .B(port_b_0[1]), .Z(
        v_1_0[1]) );
  AND2_X1 simpleAnd_51_U1 ( .A1(port_rand_mul[2]), .A2(n13), .ZN(
        simpleAnd_51_port_z) );
  XOR2_X2 simpleXor_102_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_51_port_z), 
        .Z(u_1_1[1]) );
  XOR2_X2 simpleXor_103_U1 ( .A(port_rand_mul[2]), .B(port_b_2[1]), .Z(
        v_1_1[1]) );
  AND2_X1 simpleAnd_52_U1 ( .A1(port_rand_mul[1]), .A2(n20), .ZN(
        simpleAnd_52_port_z) );
  XOR2_X2 simpleXor_104_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_52_port_z), 
        .Z(u_2_0[1]) );
  XOR2_X2 simpleXor_105_U1 ( .A(port_rand_mul[1]), .B(port_b_0[1]), .Z(
        v_2_0[1]) );
  AND2_X1 simpleAnd_53_U1 ( .A1(port_rand_mul[2]), .A2(n20), .ZN(
        simpleAnd_53_port_z) );
  XOR2_X2 simpleXor_106_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_53_port_z), 
        .Z(u_2_1[1]) );
  XOR2_X2 simpleXor_107_U1 ( .A(port_rand_mul[2]), .B(port_b_1[1]), .Z(
        v_2_1[1]) );
  AND2_X1 simpleAnd_54_U1 ( .A1(port_rand_mul[0]), .A2(n5), .ZN(
        simpleAnd_54_port_z) );
  XOR2_X2 simpleXor_108_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_54_port_z), 
        .Z(u_0_0[2]) );
  XOR2_X2 simpleXor_109_U1 ( .A(port_rand_mul[0]), .B(port_b_1[2]), .Z(
        v_0_0[2]) );
  AND2_X1 simpleAnd_55_U1 ( .A1(port_rand_mul[1]), .A2(n5), .ZN(
        simpleAnd_55_port_z) );
  XOR2_X2 simpleXor_110_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_55_port_z), 
        .Z(u_0_1[2]) );
  XOR2_X2 simpleXor_111_U1 ( .A(port_rand_mul[1]), .B(port_b_2[2]), .Z(
        v_0_1[2]) );
  AND2_X1 simpleAnd_56_U1 ( .A1(port_rand_mul[0]), .A2(n12), .ZN(
        simpleAnd_56_port_z) );
  XOR2_X2 simpleXor_112_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_56_port_z), 
        .Z(u_1_0[2]) );
  XOR2_X2 simpleXor_113_U1 ( .A(port_rand_mul[0]), .B(port_b_0[2]), .Z(
        v_1_0[2]) );
  AND2_X1 simpleAnd_57_U1 ( .A1(port_rand_mul[2]), .A2(n12), .ZN(
        simpleAnd_57_port_z) );
  XOR2_X2 simpleXor_114_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_57_port_z), 
        .Z(u_1_1[2]) );
  XOR2_X2 simpleXor_115_U1 ( .A(port_rand_mul[2]), .B(port_b_2[2]), .Z(
        v_1_1[2]) );
  AND2_X1 simpleAnd_58_U1 ( .A1(port_rand_mul[1]), .A2(n19), .ZN(
        simpleAnd_58_port_z) );
  XOR2_X2 simpleXor_116_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_58_port_z), 
        .Z(u_2_0[2]) );
  XOR2_X2 simpleXor_117_U1 ( .A(port_rand_mul[1]), .B(port_b_0[2]), .Z(
        v_2_0[2]) );
  AND2_X1 simpleAnd_59_U1 ( .A1(port_rand_mul[2]), .A2(n19), .ZN(
        simpleAnd_59_port_z) );
  XOR2_X2 simpleXor_118_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_59_port_z), 
        .Z(u_2_1[2]) );
  XOR2_X2 simpleXor_119_U1 ( .A(port_rand_mul[2]), .B(port_b_1[2]), .Z(
        v_2_1[2]) );
  AND2_X1 simpleAnd_60_U1 ( .A1(port_rand_mul[0]), .A2(n4), .ZN(
        simpleAnd_60_port_z) );
  XOR2_X2 simpleXor_120_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_60_port_z), 
        .Z(u_0_0[3]) );
  XOR2_X2 simpleXor_121_U1 ( .A(port_rand_mul[0]), .B(port_b_1[3]), .Z(
        v_0_0[3]) );
  AND2_X1 simpleAnd_61_U1 ( .A1(port_rand_mul[1]), .A2(n4), .ZN(
        simpleAnd_61_port_z) );
  XOR2_X2 simpleXor_122_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_61_port_z), 
        .Z(u_0_1[3]) );
  XOR2_X2 simpleXor_123_U1 ( .A(port_rand_mul[1]), .B(port_b_2[3]), .Z(
        v_0_1[3]) );
  AND2_X1 simpleAnd_62_U1 ( .A1(port_rand_mul[0]), .A2(n11), .ZN(
        simpleAnd_62_port_z) );
  XOR2_X2 simpleXor_124_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_62_port_z), 
        .Z(u_1_0[3]) );
  XOR2_X2 simpleXor_125_U1 ( .A(port_rand_mul[0]), .B(port_b_0[3]), .Z(
        v_1_0[3]) );
  AND2_X1 simpleAnd_63_U1 ( .A1(port_rand_mul[2]), .A2(n11), .ZN(
        simpleAnd_63_port_z) );
  XOR2_X2 simpleXor_126_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_63_port_z), 
        .Z(u_1_1[3]) );
  XOR2_X2 simpleXor_127_U1 ( .A(port_rand_mul[2]), .B(port_b_2[3]), .Z(
        v_1_1[3]) );
  AND2_X1 simpleAnd_64_U1 ( .A1(port_rand_mul[1]), .A2(n18), .ZN(
        simpleAnd_64_port_z) );
  XOR2_X2 simpleXor_128_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_64_port_z), 
        .Z(u_2_0[3]) );
  XOR2_X2 simpleXor_129_U1 ( .A(port_rand_mul[1]), .B(port_b_0[3]), .Z(
        v_2_0[3]) );
  AND2_X1 simpleAnd_65_U1 ( .A1(port_rand_mul[2]), .A2(n18), .ZN(
        simpleAnd_65_port_z) );
  XOR2_X2 simpleXor_130_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_65_port_z), 
        .Z(u_2_1[3]) );
  XOR2_X2 simpleXor_131_U1 ( .A(port_rand_mul[2]), .B(port_b_1[3]), .Z(
        v_2_1[3]) );
  AND2_X1 simpleAnd_66_U1 ( .A1(port_rand_mul[0]), .A2(n3), .ZN(
        simpleAnd_66_port_z) );
  XOR2_X2 simpleXor_132_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_66_port_z), 
        .Z(u_0_0[4]) );
  XOR2_X2 simpleXor_133_U1 ( .A(port_rand_mul[0]), .B(port_b_1[4]), .Z(
        v_0_0[4]) );
  AND2_X1 simpleAnd_67_U1 ( .A1(port_rand_mul[1]), .A2(n3), .ZN(
        simpleAnd_67_port_z) );
  XOR2_X2 simpleXor_134_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_67_port_z), 
        .Z(u_0_1[4]) );
  XOR2_X2 simpleXor_135_U1 ( .A(port_rand_mul[1]), .B(port_b_2[4]), .Z(
        v_0_1[4]) );
  AND2_X1 simpleAnd_68_U1 ( .A1(port_rand_mul[0]), .A2(n10), .ZN(
        simpleAnd_68_port_z) );
  XOR2_X2 simpleXor_136_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_68_port_z), 
        .Z(u_1_0[4]) );
  XOR2_X2 simpleXor_137_U1 ( .A(port_rand_mul[0]), .B(port_b_0[4]), .Z(
        v_1_0[4]) );
  AND2_X1 simpleAnd_69_U1 ( .A1(port_rand_mul[2]), .A2(n10), .ZN(
        simpleAnd_69_port_z) );
  XOR2_X2 simpleXor_138_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_69_port_z), 
        .Z(u_1_1[4]) );
  XOR2_X2 simpleXor_139_U1 ( .A(port_rand_mul[2]), .B(port_b_2[4]), .Z(
        v_1_1[4]) );
  AND2_X1 simpleAnd_70_U1 ( .A1(port_rand_mul[1]), .A2(n17), .ZN(
        simpleAnd_70_port_z) );
  XOR2_X2 simpleXor_140_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_70_port_z), 
        .Z(u_2_0[4]) );
  XOR2_X2 simpleXor_141_U1 ( .A(port_rand_mul[1]), .B(port_b_0[4]), .Z(
        v_2_0[4]) );
  AND2_X1 simpleAnd_71_U1 ( .A1(port_rand_mul[2]), .A2(n17), .ZN(
        simpleAnd_71_port_z) );
  XOR2_X2 simpleXor_142_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_71_port_z), 
        .Z(u_2_1[4]) );
  XOR2_X2 simpleXor_143_U1 ( .A(port_rand_mul[2]), .B(port_b_1[4]), .Z(
        v_2_1[4]) );
  AND2_X1 simpleAnd_72_U1 ( .A1(port_rand_mul[0]), .A2(n2), .ZN(
        simpleAnd_72_port_z) );
  XOR2_X2 simpleXor_144_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_72_port_z), 
        .Z(u_0_0[5]) );
  XOR2_X2 simpleXor_145_U1 ( .A(port_rand_mul[0]), .B(port_b_1[5]), .Z(
        v_0_0[5]) );
  AND2_X1 simpleAnd_73_U1 ( .A1(port_rand_mul[1]), .A2(n2), .ZN(
        simpleAnd_73_port_z) );
  XOR2_X2 simpleXor_146_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_73_port_z), 
        .Z(u_0_1[5]) );
  XOR2_X2 simpleXor_147_U1 ( .A(port_rand_mul[1]), .B(port_b_2[5]), .Z(
        v_0_1[5]) );
  AND2_X1 simpleAnd_74_U1 ( .A1(port_rand_mul[0]), .A2(n9), .ZN(
        simpleAnd_74_port_z) );
  XOR2_X2 simpleXor_148_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_74_port_z), 
        .Z(u_1_0[5]) );
  XOR2_X2 simpleXor_149_U1 ( .A(port_rand_mul[0]), .B(port_b_0[5]), .Z(
        v_1_0[5]) );
  AND2_X1 simpleAnd_75_U1 ( .A1(port_rand_mul[2]), .A2(n9), .ZN(
        simpleAnd_75_port_z) );
  XOR2_X2 simpleXor_150_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_75_port_z), 
        .Z(u_1_1[5]) );
  XOR2_X2 simpleXor_151_U1 ( .A(port_rand_mul[2]), .B(port_b_2[5]), .Z(
        v_1_1[5]) );
  AND2_X1 simpleAnd_76_U1 ( .A1(port_rand_mul[1]), .A2(n16), .ZN(
        simpleAnd_76_port_z) );
  XOR2_X2 simpleXor_152_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_76_port_z), 
        .Z(u_2_0[5]) );
  XOR2_X2 simpleXor_153_U1 ( .A(port_rand_mul[1]), .B(port_b_0[5]), .Z(
        v_2_0[5]) );
  AND2_X1 simpleAnd_77_U1 ( .A1(port_rand_mul[2]), .A2(n16), .ZN(
        simpleAnd_77_port_z) );
  XOR2_X2 simpleXor_154_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_77_port_z), 
        .Z(u_2_1[5]) );
  XOR2_X2 simpleXor_155_U1 ( .A(port_rand_mul[2]), .B(port_b_1[5]), .Z(
        v_2_1[5]) );
  AND2_X1 simpleAnd_78_U1 ( .A1(port_rand_mul[0]), .A2(n1), .ZN(
        simpleAnd_78_port_z) );
  XOR2_X1 simpleXor_156_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_78_port_z), 
        .Z(u_0_0[6]) );
  XOR2_X1 simpleXor_157_U1 ( .A(port_rand_mul[0]), .B(port_b_1[6]), .Z(
        v_0_0[6]) );
  AND2_X1 simpleAnd_79_U1 ( .A1(port_rand_mul[1]), .A2(n1), .ZN(
        simpleAnd_79_port_z) );
  XOR2_X1 simpleXor_158_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_79_port_z), 
        .Z(u_0_1[6]) );
  XOR2_X1 simpleXor_159_U1 ( .A(port_rand_mul[1]), .B(port_b_2[6]), .Z(
        v_0_1[6]) );
  AND2_X1 simpleAnd_80_U1 ( .A1(port_rand_mul[0]), .A2(n8), .ZN(
        simpleAnd_80_port_z) );
  XOR2_X1 simpleXor_160_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_80_port_z), 
        .Z(u_1_0[6]) );
  XOR2_X1 simpleXor_161_U1 ( .A(port_rand_mul[0]), .B(port_b_0[6]), .Z(
        v_1_0[6]) );
  AND2_X1 simpleAnd_81_U1 ( .A1(port_rand_mul[2]), .A2(n8), .ZN(
        simpleAnd_81_port_z) );
  XOR2_X1 simpleXor_162_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_81_port_z), 
        .Z(u_1_1[6]) );
  XOR2_X1 simpleXor_163_U1 ( .A(port_rand_mul[2]), .B(port_b_2[6]), .Z(
        v_1_1[6]) );
  AND2_X1 simpleAnd_82_U1 ( .A1(port_rand_mul[1]), .A2(n15), .ZN(
        simpleAnd_82_port_z) );
  XOR2_X1 simpleXor_164_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_82_port_z), 
        .Z(u_2_0[6]) );
  XOR2_X1 simpleXor_165_U1 ( .A(port_rand_mul[1]), .B(port_b_0[6]), .Z(
        v_2_0[6]) );
  AND2_X1 simpleAnd_83_U1 ( .A1(port_rand_mul[2]), .A2(n15), .ZN(
        simpleAnd_83_port_z) );
  XOR2_X1 simpleXor_166_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_83_port_z), 
        .Z(u_2_1[6]) );
  XOR2_X1 simpleXor_167_U1 ( .A(port_rand_mul[2]), .B(port_b_1[6]), .Z(
        v_2_1[6]) );
  OR2_X1 maj_84_U19 ( .A1(maj_84_n8), .A2(maj_84_n9), .ZN(maj_84_n7) );
  NAND2_X1 maj_84_U18 ( .A1(u_0_0[6]), .A2(maj_84_n7), .ZN(maj_84_n6) );
  NAND2_X1 maj_84_U17 ( .A1(maj_84_n9), .A2(maj_84_n8), .ZN(maj_84_n5) );
  NAND2_X1 maj_84_U16 ( .A1(maj_84_n5), .A2(maj_84_n6), .ZN(maj_84_n4) );
  NAND2_X1 maj_84_U15 ( .A1(u_0_0[5]), .A2(maj_84_n10), .ZN(maj_84_n17) );
  NAND2_X1 maj_84_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_84_n16) );
  NAND2_X1 maj_84_U13 ( .A1(maj_84_n16), .A2(maj_84_n17), .ZN(maj_84_n13) );
  NAND2_X1 maj_84_U12 ( .A1(u_0_0[2]), .A2(maj_84_n11), .ZN(maj_84_n15) );
  NAND2_X1 maj_84_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_84_n14) );
  NAND2_X1 maj_84_U10 ( .A1(maj_84_n14), .A2(maj_84_n15), .ZN(maj_84_n12) );
  XOR2_X1 maj_84_U9 ( .A(u_0_0[2]), .B(maj_84_n11), .Z(maj_84_n9) );
  XOR2_X1 maj_84_U8 ( .A(u_0_0[5]), .B(maj_84_n10), .Z(maj_84_n8) );
  XOR2_X1 maj_84_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_84_n11) );
  XOR2_X1 maj_84_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_84_n10) );
  OR2_X1 maj_84_U5 ( .A1(maj_84_n12), .A2(maj_84_n13), .ZN(maj_84_n3) );
  NAND2_X1 maj_84_U4 ( .A1(maj_84_n13), .A2(maj_84_n12), .ZN(maj_84_n1) );
  NAND2_X1 maj_84_U3 ( .A1(maj_84_n3), .A2(maj_84_n4), .ZN(maj_84_n2) );
  NAND2_X1 maj_84_U2 ( .A1(maj_84_n1), .A2(maj_84_n2), .ZN(maj_84_port_o) );
  OR2_X1 maj_85_U19 ( .A1(maj_85_n27), .A2(maj_85_n26), .ZN(maj_85_n28) );
  NAND2_X1 maj_85_U18 ( .A1(v_0_0[6]), .A2(maj_85_n28), .ZN(maj_85_n29) );
  NAND2_X1 maj_85_U17 ( .A1(maj_85_n26), .A2(maj_85_n27), .ZN(maj_85_n30) );
  NAND2_X1 maj_85_U16 ( .A1(maj_85_n30), .A2(maj_85_n29), .ZN(maj_85_n31) );
  NAND2_X1 maj_85_U15 ( .A1(v_0_0[5]), .A2(maj_85_n25), .ZN(maj_85_n18) );
  NAND2_X1 maj_85_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_85_n19) );
  NAND2_X1 maj_85_U13 ( .A1(maj_85_n19), .A2(maj_85_n18), .ZN(maj_85_n22) );
  NAND2_X1 maj_85_U12 ( .A1(v_0_0[2]), .A2(maj_85_n24), .ZN(maj_85_n20) );
  NAND2_X1 maj_85_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_85_n21) );
  NAND2_X1 maj_85_U10 ( .A1(maj_85_n21), .A2(maj_85_n20), .ZN(maj_85_n23) );
  XOR2_X1 maj_85_U9 ( .A(v_0_0[2]), .B(maj_85_n24), .Z(maj_85_n26) );
  XOR2_X1 maj_85_U8 ( .A(v_0_0[5]), .B(maj_85_n25), .Z(maj_85_n27) );
  XOR2_X1 maj_85_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_85_n24) );
  XOR2_X1 maj_85_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_85_n25) );
  OR2_X1 maj_85_U5 ( .A1(maj_85_n23), .A2(maj_85_n22), .ZN(maj_85_n32) );
  NAND2_X1 maj_85_U4 ( .A1(maj_85_n22), .A2(maj_85_n23), .ZN(maj_85_n34) );
  NAND2_X1 maj_85_U3 ( .A1(maj_85_n32), .A2(maj_85_n31), .ZN(maj_85_n33) );
  NAND2_X1 maj_85_U2 ( .A1(maj_85_n34), .A2(maj_85_n33), .ZN(maj_85_port_o) );
  OR2_X1 maj_86_U19 ( .A1(maj_86_n27), .A2(maj_86_n26), .ZN(maj_86_n28) );
  NAND2_X1 maj_86_U18 ( .A1(u_0_1[6]), .A2(maj_86_n28), .ZN(maj_86_n29) );
  NAND2_X1 maj_86_U17 ( .A1(maj_86_n26), .A2(maj_86_n27), .ZN(maj_86_n30) );
  NAND2_X1 maj_86_U16 ( .A1(maj_86_n30), .A2(maj_86_n29), .ZN(maj_86_n31) );
  NAND2_X1 maj_86_U15 ( .A1(u_0_1[5]), .A2(maj_86_n25), .ZN(maj_86_n18) );
  NAND2_X1 maj_86_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_86_n19) );
  NAND2_X1 maj_86_U13 ( .A1(maj_86_n19), .A2(maj_86_n18), .ZN(maj_86_n22) );
  NAND2_X1 maj_86_U12 ( .A1(u_0_1[2]), .A2(maj_86_n24), .ZN(maj_86_n20) );
  NAND2_X1 maj_86_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_86_n21) );
  NAND2_X1 maj_86_U10 ( .A1(maj_86_n21), .A2(maj_86_n20), .ZN(maj_86_n23) );
  XOR2_X1 maj_86_U9 ( .A(u_0_1[2]), .B(maj_86_n24), .Z(maj_86_n26) );
  XOR2_X1 maj_86_U8 ( .A(u_0_1[5]), .B(maj_86_n25), .Z(maj_86_n27) );
  XOR2_X1 maj_86_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_86_n24) );
  XOR2_X1 maj_86_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_86_n25) );
  OR2_X1 maj_86_U5 ( .A1(maj_86_n23), .A2(maj_86_n22), .ZN(maj_86_n32) );
  NAND2_X1 maj_86_U4 ( .A1(maj_86_n22), .A2(maj_86_n23), .ZN(maj_86_n34) );
  NAND2_X1 maj_86_U3 ( .A1(maj_86_n32), .A2(maj_86_n31), .ZN(maj_86_n33) );
  NAND2_X1 maj_86_U2 ( .A1(maj_86_n34), .A2(maj_86_n33), .ZN(maj_86_port_o) );
  OR2_X1 maj_87_U19 ( .A1(maj_87_n27), .A2(maj_87_n26), .ZN(maj_87_n28) );
  NAND2_X1 maj_87_U18 ( .A1(v_0_1[6]), .A2(maj_87_n28), .ZN(maj_87_n29) );
  NAND2_X1 maj_87_U17 ( .A1(maj_87_n26), .A2(maj_87_n27), .ZN(maj_87_n30) );
  NAND2_X1 maj_87_U16 ( .A1(maj_87_n30), .A2(maj_87_n29), .ZN(maj_87_n31) );
  NAND2_X1 maj_87_U15 ( .A1(v_0_1[5]), .A2(maj_87_n25), .ZN(maj_87_n18) );
  NAND2_X1 maj_87_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_87_n19) );
  NAND2_X1 maj_87_U13 ( .A1(maj_87_n19), .A2(maj_87_n18), .ZN(maj_87_n22) );
  NAND2_X1 maj_87_U12 ( .A1(v_0_1[2]), .A2(maj_87_n24), .ZN(maj_87_n20) );
  NAND2_X1 maj_87_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_87_n21) );
  NAND2_X1 maj_87_U10 ( .A1(maj_87_n21), .A2(maj_87_n20), .ZN(maj_87_n23) );
  XOR2_X1 maj_87_U9 ( .A(v_0_1[2]), .B(maj_87_n24), .Z(maj_87_n26) );
  XOR2_X1 maj_87_U8 ( .A(v_0_1[5]), .B(maj_87_n25), .Z(maj_87_n27) );
  XOR2_X1 maj_87_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_87_n24) );
  XOR2_X1 maj_87_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_87_n25) );
  OR2_X1 maj_87_U5 ( .A1(maj_87_n23), .A2(maj_87_n22), .ZN(maj_87_n32) );
  NAND2_X1 maj_87_U4 ( .A1(maj_87_n22), .A2(maj_87_n23), .ZN(maj_87_n34) );
  NAND2_X1 maj_87_U3 ( .A1(maj_87_n32), .A2(maj_87_n31), .ZN(maj_87_n33) );
  NAND2_X1 maj_87_U2 ( .A1(maj_87_n34), .A2(maj_87_n33), .ZN(maj_87_port_o) );
  OR2_X1 maj_88_U19 ( .A1(maj_88_n27), .A2(maj_88_n26), .ZN(maj_88_n28) );
  NAND2_X1 maj_88_U18 ( .A1(u_1_0[6]), .A2(maj_88_n28), .ZN(maj_88_n29) );
  NAND2_X1 maj_88_U17 ( .A1(maj_88_n26), .A2(maj_88_n27), .ZN(maj_88_n30) );
  NAND2_X1 maj_88_U16 ( .A1(maj_88_n30), .A2(maj_88_n29), .ZN(maj_88_n31) );
  NAND2_X1 maj_88_U15 ( .A1(u_1_0[5]), .A2(maj_88_n25), .ZN(maj_88_n18) );
  NAND2_X1 maj_88_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_88_n19) );
  NAND2_X1 maj_88_U13 ( .A1(maj_88_n19), .A2(maj_88_n18), .ZN(maj_88_n22) );
  NAND2_X1 maj_88_U12 ( .A1(u_1_0[2]), .A2(maj_88_n24), .ZN(maj_88_n20) );
  NAND2_X1 maj_88_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_88_n21) );
  NAND2_X1 maj_88_U10 ( .A1(maj_88_n21), .A2(maj_88_n20), .ZN(maj_88_n23) );
  XOR2_X1 maj_88_U9 ( .A(u_1_0[2]), .B(maj_88_n24), .Z(maj_88_n26) );
  XOR2_X1 maj_88_U8 ( .A(u_1_0[5]), .B(maj_88_n25), .Z(maj_88_n27) );
  XOR2_X1 maj_88_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_88_n24) );
  XOR2_X1 maj_88_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_88_n25) );
  OR2_X1 maj_88_U5 ( .A1(maj_88_n23), .A2(maj_88_n22), .ZN(maj_88_n32) );
  NAND2_X1 maj_88_U4 ( .A1(maj_88_n22), .A2(maj_88_n23), .ZN(maj_88_n34) );
  NAND2_X1 maj_88_U3 ( .A1(maj_88_n32), .A2(maj_88_n31), .ZN(maj_88_n33) );
  NAND2_X1 maj_88_U2 ( .A1(maj_88_n34), .A2(maj_88_n33), .ZN(maj_88_port_o) );
  OR2_X1 maj_89_U19 ( .A1(maj_89_n27), .A2(maj_89_n26), .ZN(maj_89_n28) );
  NAND2_X1 maj_89_U18 ( .A1(v_1_0[6]), .A2(maj_89_n28), .ZN(maj_89_n29) );
  NAND2_X1 maj_89_U17 ( .A1(maj_89_n26), .A2(maj_89_n27), .ZN(maj_89_n30) );
  NAND2_X1 maj_89_U16 ( .A1(maj_89_n30), .A2(maj_89_n29), .ZN(maj_89_n31) );
  NAND2_X1 maj_89_U15 ( .A1(v_1_0[5]), .A2(maj_89_n25), .ZN(maj_89_n18) );
  NAND2_X1 maj_89_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_89_n19) );
  NAND2_X1 maj_89_U13 ( .A1(maj_89_n19), .A2(maj_89_n18), .ZN(maj_89_n22) );
  NAND2_X1 maj_89_U12 ( .A1(v_1_0[2]), .A2(maj_89_n24), .ZN(maj_89_n20) );
  NAND2_X1 maj_89_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_89_n21) );
  NAND2_X1 maj_89_U10 ( .A1(maj_89_n21), .A2(maj_89_n20), .ZN(maj_89_n23) );
  XOR2_X1 maj_89_U9 ( .A(v_1_0[2]), .B(maj_89_n24), .Z(maj_89_n26) );
  XOR2_X1 maj_89_U8 ( .A(v_1_0[5]), .B(maj_89_n25), .Z(maj_89_n27) );
  XOR2_X1 maj_89_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_89_n24) );
  XOR2_X1 maj_89_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_89_n25) );
  OR2_X1 maj_89_U5 ( .A1(maj_89_n23), .A2(maj_89_n22), .ZN(maj_89_n32) );
  NAND2_X1 maj_89_U4 ( .A1(maj_89_n22), .A2(maj_89_n23), .ZN(maj_89_n34) );
  NAND2_X1 maj_89_U3 ( .A1(maj_89_n32), .A2(maj_89_n31), .ZN(maj_89_n33) );
  NAND2_X1 maj_89_U2 ( .A1(maj_89_n34), .A2(maj_89_n33), .ZN(maj_89_port_o) );
  OR2_X1 maj_90_U19 ( .A1(maj_90_n27), .A2(maj_90_n26), .ZN(maj_90_n28) );
  NAND2_X1 maj_90_U18 ( .A1(u_1_1[6]), .A2(maj_90_n28), .ZN(maj_90_n29) );
  NAND2_X1 maj_90_U17 ( .A1(maj_90_n26), .A2(maj_90_n27), .ZN(maj_90_n30) );
  NAND2_X1 maj_90_U16 ( .A1(maj_90_n30), .A2(maj_90_n29), .ZN(maj_90_n31) );
  NAND2_X1 maj_90_U15 ( .A1(u_1_1[5]), .A2(maj_90_n25), .ZN(maj_90_n18) );
  NAND2_X1 maj_90_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_90_n19) );
  NAND2_X1 maj_90_U13 ( .A1(maj_90_n19), .A2(maj_90_n18), .ZN(maj_90_n22) );
  NAND2_X1 maj_90_U12 ( .A1(u_1_1[2]), .A2(maj_90_n24), .ZN(maj_90_n20) );
  NAND2_X1 maj_90_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_90_n21) );
  NAND2_X1 maj_90_U10 ( .A1(maj_90_n21), .A2(maj_90_n20), .ZN(maj_90_n23) );
  XOR2_X1 maj_90_U9 ( .A(u_1_1[2]), .B(maj_90_n24), .Z(maj_90_n26) );
  XOR2_X1 maj_90_U8 ( .A(u_1_1[5]), .B(maj_90_n25), .Z(maj_90_n27) );
  XOR2_X1 maj_90_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_90_n24) );
  XOR2_X1 maj_90_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_90_n25) );
  OR2_X1 maj_90_U5 ( .A1(maj_90_n23), .A2(maj_90_n22), .ZN(maj_90_n32) );
  NAND2_X1 maj_90_U4 ( .A1(maj_90_n22), .A2(maj_90_n23), .ZN(maj_90_n34) );
  NAND2_X1 maj_90_U3 ( .A1(maj_90_n32), .A2(maj_90_n31), .ZN(maj_90_n33) );
  NAND2_X1 maj_90_U2 ( .A1(maj_90_n34), .A2(maj_90_n33), .ZN(maj_90_port_o) );
  OR2_X1 maj_91_U19 ( .A1(maj_91_n27), .A2(maj_91_n26), .ZN(maj_91_n28) );
  NAND2_X1 maj_91_U18 ( .A1(v_1_1[6]), .A2(maj_91_n28), .ZN(maj_91_n29) );
  NAND2_X1 maj_91_U17 ( .A1(maj_91_n26), .A2(maj_91_n27), .ZN(maj_91_n30) );
  NAND2_X1 maj_91_U16 ( .A1(maj_91_n30), .A2(maj_91_n29), .ZN(maj_91_n31) );
  NAND2_X1 maj_91_U15 ( .A1(v_1_1[5]), .A2(maj_91_n25), .ZN(maj_91_n18) );
  NAND2_X1 maj_91_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_91_n19) );
  NAND2_X1 maj_91_U13 ( .A1(maj_91_n19), .A2(maj_91_n18), .ZN(maj_91_n22) );
  NAND2_X1 maj_91_U12 ( .A1(v_1_1[2]), .A2(maj_91_n24), .ZN(maj_91_n20) );
  NAND2_X1 maj_91_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_91_n21) );
  NAND2_X1 maj_91_U10 ( .A1(maj_91_n21), .A2(maj_91_n20), .ZN(maj_91_n23) );
  XOR2_X1 maj_91_U9 ( .A(v_1_1[2]), .B(maj_91_n24), .Z(maj_91_n26) );
  XOR2_X1 maj_91_U8 ( .A(v_1_1[5]), .B(maj_91_n25), .Z(maj_91_n27) );
  XOR2_X1 maj_91_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_91_n24) );
  XOR2_X1 maj_91_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_91_n25) );
  OR2_X1 maj_91_U5 ( .A1(maj_91_n23), .A2(maj_91_n22), .ZN(maj_91_n32) );
  NAND2_X1 maj_91_U4 ( .A1(maj_91_n22), .A2(maj_91_n23), .ZN(maj_91_n34) );
  NAND2_X1 maj_91_U3 ( .A1(maj_91_n32), .A2(maj_91_n31), .ZN(maj_91_n33) );
  NAND2_X1 maj_91_U2 ( .A1(maj_91_n34), .A2(maj_91_n33), .ZN(maj_91_port_o) );
  OR2_X1 maj_92_U19 ( .A1(maj_92_n27), .A2(maj_92_n26), .ZN(maj_92_n28) );
  NAND2_X1 maj_92_U18 ( .A1(u_2_0[6]), .A2(maj_92_n28), .ZN(maj_92_n29) );
  NAND2_X1 maj_92_U17 ( .A1(maj_92_n26), .A2(maj_92_n27), .ZN(maj_92_n30) );
  NAND2_X1 maj_92_U16 ( .A1(maj_92_n30), .A2(maj_92_n29), .ZN(maj_92_n31) );
  NAND2_X1 maj_92_U15 ( .A1(u_2_0[5]), .A2(maj_92_n25), .ZN(maj_92_n18) );
  NAND2_X1 maj_92_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_92_n19) );
  NAND2_X1 maj_92_U13 ( .A1(maj_92_n19), .A2(maj_92_n18), .ZN(maj_92_n22) );
  NAND2_X1 maj_92_U12 ( .A1(u_2_0[2]), .A2(maj_92_n24), .ZN(maj_92_n20) );
  NAND2_X1 maj_92_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_92_n21) );
  NAND2_X1 maj_92_U10 ( .A1(maj_92_n21), .A2(maj_92_n20), .ZN(maj_92_n23) );
  XOR2_X1 maj_92_U9 ( .A(u_2_0[2]), .B(maj_92_n24), .Z(maj_92_n26) );
  XOR2_X1 maj_92_U8 ( .A(u_2_0[5]), .B(maj_92_n25), .Z(maj_92_n27) );
  XOR2_X1 maj_92_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_92_n24) );
  XOR2_X1 maj_92_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_92_n25) );
  OR2_X1 maj_92_U5 ( .A1(maj_92_n23), .A2(maj_92_n22), .ZN(maj_92_n32) );
  NAND2_X1 maj_92_U4 ( .A1(maj_92_n22), .A2(maj_92_n23), .ZN(maj_92_n34) );
  NAND2_X1 maj_92_U3 ( .A1(maj_92_n32), .A2(maj_92_n31), .ZN(maj_92_n33) );
  NAND2_X1 maj_92_U2 ( .A1(maj_92_n34), .A2(maj_92_n33), .ZN(maj_92_port_o) );
  OR2_X1 maj_93_U19 ( .A1(maj_93_n27), .A2(maj_93_n26), .ZN(maj_93_n28) );
  NAND2_X1 maj_93_U18 ( .A1(v_2_0[6]), .A2(maj_93_n28), .ZN(maj_93_n29) );
  NAND2_X1 maj_93_U17 ( .A1(maj_93_n26), .A2(maj_93_n27), .ZN(maj_93_n30) );
  NAND2_X1 maj_93_U16 ( .A1(maj_93_n30), .A2(maj_93_n29), .ZN(maj_93_n31) );
  NAND2_X1 maj_93_U15 ( .A1(v_2_0[5]), .A2(maj_93_n25), .ZN(maj_93_n18) );
  NAND2_X1 maj_93_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_93_n19) );
  NAND2_X1 maj_93_U13 ( .A1(maj_93_n19), .A2(maj_93_n18), .ZN(maj_93_n22) );
  NAND2_X1 maj_93_U12 ( .A1(v_2_0[2]), .A2(maj_93_n24), .ZN(maj_93_n20) );
  NAND2_X1 maj_93_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_93_n21) );
  NAND2_X1 maj_93_U10 ( .A1(maj_93_n21), .A2(maj_93_n20), .ZN(maj_93_n23) );
  XOR2_X1 maj_93_U9 ( .A(v_2_0[2]), .B(maj_93_n24), .Z(maj_93_n26) );
  XOR2_X1 maj_93_U8 ( .A(v_2_0[5]), .B(maj_93_n25), .Z(maj_93_n27) );
  XOR2_X1 maj_93_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_93_n24) );
  XOR2_X1 maj_93_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_93_n25) );
  OR2_X1 maj_93_U5 ( .A1(maj_93_n23), .A2(maj_93_n22), .ZN(maj_93_n32) );
  NAND2_X1 maj_93_U4 ( .A1(maj_93_n22), .A2(maj_93_n23), .ZN(maj_93_n34) );
  NAND2_X1 maj_93_U3 ( .A1(maj_93_n32), .A2(maj_93_n31), .ZN(maj_93_n33) );
  NAND2_X1 maj_93_U2 ( .A1(maj_93_n34), .A2(maj_93_n33), .ZN(maj_93_port_o) );
  OR2_X1 maj_94_U19 ( .A1(maj_94_n27), .A2(maj_94_n26), .ZN(maj_94_n28) );
  NAND2_X1 maj_94_U18 ( .A1(u_2_1[6]), .A2(maj_94_n28), .ZN(maj_94_n29) );
  NAND2_X1 maj_94_U17 ( .A1(maj_94_n26), .A2(maj_94_n27), .ZN(maj_94_n30) );
  NAND2_X1 maj_94_U16 ( .A1(maj_94_n30), .A2(maj_94_n29), .ZN(maj_94_n31) );
  NAND2_X1 maj_94_U15 ( .A1(u_2_1[5]), .A2(maj_94_n25), .ZN(maj_94_n18) );
  NAND2_X1 maj_94_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_94_n19) );
  NAND2_X1 maj_94_U13 ( .A1(maj_94_n19), .A2(maj_94_n18), .ZN(maj_94_n22) );
  NAND2_X1 maj_94_U12 ( .A1(u_2_1[2]), .A2(maj_94_n24), .ZN(maj_94_n20) );
  NAND2_X1 maj_94_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_94_n21) );
  NAND2_X1 maj_94_U10 ( .A1(maj_94_n21), .A2(maj_94_n20), .ZN(maj_94_n23) );
  XOR2_X1 maj_94_U9 ( .A(u_2_1[2]), .B(maj_94_n24), .Z(maj_94_n26) );
  XOR2_X1 maj_94_U8 ( .A(u_2_1[5]), .B(maj_94_n25), .Z(maj_94_n27) );
  XOR2_X1 maj_94_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_94_n24) );
  XOR2_X1 maj_94_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_94_n25) );
  OR2_X1 maj_94_U5 ( .A1(maj_94_n23), .A2(maj_94_n22), .ZN(maj_94_n32) );
  NAND2_X1 maj_94_U4 ( .A1(maj_94_n22), .A2(maj_94_n23), .ZN(maj_94_n34) );
  NAND2_X1 maj_94_U3 ( .A1(maj_94_n32), .A2(maj_94_n31), .ZN(maj_94_n33) );
  NAND2_X1 maj_94_U2 ( .A1(maj_94_n34), .A2(maj_94_n33), .ZN(maj_94_port_o) );
  OR2_X1 maj_95_U19 ( .A1(maj_95_n27), .A2(maj_95_n26), .ZN(maj_95_n28) );
  NAND2_X1 maj_95_U18 ( .A1(v_2_1[6]), .A2(maj_95_n28), .ZN(maj_95_n29) );
  NAND2_X1 maj_95_U17 ( .A1(maj_95_n26), .A2(maj_95_n27), .ZN(maj_95_n30) );
  NAND2_X1 maj_95_U16 ( .A1(maj_95_n30), .A2(maj_95_n29), .ZN(maj_95_n31) );
  NAND2_X1 maj_95_U15 ( .A1(v_2_1[5]), .A2(maj_95_n25), .ZN(maj_95_n18) );
  NAND2_X1 maj_95_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_95_n19) );
  NAND2_X1 maj_95_U13 ( .A1(maj_95_n19), .A2(maj_95_n18), .ZN(maj_95_n22) );
  NAND2_X1 maj_95_U12 ( .A1(v_2_1[2]), .A2(maj_95_n24), .ZN(maj_95_n20) );
  NAND2_X1 maj_95_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_95_n21) );
  NAND2_X1 maj_95_U10 ( .A1(maj_95_n21), .A2(maj_95_n20), .ZN(maj_95_n23) );
  XOR2_X1 maj_95_U9 ( .A(v_2_1[2]), .B(maj_95_n24), .Z(maj_95_n26) );
  XOR2_X1 maj_95_U8 ( .A(v_2_1[5]), .B(maj_95_n25), .Z(maj_95_n27) );
  XOR2_X1 maj_95_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_95_n24) );
  XOR2_X1 maj_95_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_95_n25) );
  OR2_X1 maj_95_U5 ( .A1(maj_95_n23), .A2(maj_95_n22), .ZN(maj_95_n32) );
  NAND2_X1 maj_95_U4 ( .A1(maj_95_n22), .A2(maj_95_n23), .ZN(maj_95_n34) );
  NAND2_X1 maj_95_U3 ( .A1(maj_95_n32), .A2(maj_95_n31), .ZN(maj_95_n33) );
  NAND2_X1 maj_95_U2 ( .A1(maj_95_n34), .A2(maj_95_n33), .ZN(maj_95_port_o) );
  OR2_X1 maj_96_U19 ( .A1(maj_96_n27), .A2(maj_96_n26), .ZN(maj_96_n28) );
  NAND2_X1 maj_96_U18 ( .A1(u_0_0[6]), .A2(maj_96_n28), .ZN(maj_96_n29) );
  NAND2_X1 maj_96_U17 ( .A1(maj_96_n26), .A2(maj_96_n27), .ZN(maj_96_n30) );
  NAND2_X1 maj_96_U16 ( .A1(maj_96_n30), .A2(maj_96_n29), .ZN(maj_96_n31) );
  NAND2_X1 maj_96_U15 ( .A1(u_0_0[5]), .A2(maj_96_n25), .ZN(maj_96_n18) );
  NAND2_X1 maj_96_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_96_n19) );
  NAND2_X1 maj_96_U13 ( .A1(maj_96_n19), .A2(maj_96_n18), .ZN(maj_96_n22) );
  NAND2_X1 maj_96_U12 ( .A1(u_0_0[2]), .A2(maj_96_n24), .ZN(maj_96_n20) );
  NAND2_X1 maj_96_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_96_n21) );
  NAND2_X1 maj_96_U10 ( .A1(maj_96_n21), .A2(maj_96_n20), .ZN(maj_96_n23) );
  XOR2_X1 maj_96_U9 ( .A(u_0_0[2]), .B(maj_96_n24), .Z(maj_96_n26) );
  XOR2_X1 maj_96_U8 ( .A(u_0_0[5]), .B(maj_96_n25), .Z(maj_96_n27) );
  XOR2_X1 maj_96_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_96_n24) );
  XOR2_X1 maj_96_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_96_n25) );
  OR2_X1 maj_96_U5 ( .A1(maj_96_n23), .A2(maj_96_n22), .ZN(maj_96_n32) );
  NAND2_X1 maj_96_U4 ( .A1(maj_96_n22), .A2(maj_96_n23), .ZN(maj_96_n34) );
  NAND2_X1 maj_96_U3 ( .A1(maj_96_n32), .A2(maj_96_n31), .ZN(maj_96_n33) );
  NAND2_X1 maj_96_U2 ( .A1(maj_96_n34), .A2(maj_96_n33), .ZN(maj_96_port_o) );
  OR2_X1 maj_97_U19 ( .A1(maj_97_n27), .A2(maj_97_n26), .ZN(maj_97_n28) );
  NAND2_X1 maj_97_U18 ( .A1(v_0_0[6]), .A2(maj_97_n28), .ZN(maj_97_n29) );
  NAND2_X1 maj_97_U17 ( .A1(maj_97_n26), .A2(maj_97_n27), .ZN(maj_97_n30) );
  NAND2_X1 maj_97_U16 ( .A1(maj_97_n30), .A2(maj_97_n29), .ZN(maj_97_n31) );
  NAND2_X1 maj_97_U15 ( .A1(v_0_0[5]), .A2(maj_97_n25), .ZN(maj_97_n18) );
  NAND2_X1 maj_97_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_97_n19) );
  NAND2_X1 maj_97_U13 ( .A1(maj_97_n19), .A2(maj_97_n18), .ZN(maj_97_n22) );
  NAND2_X1 maj_97_U12 ( .A1(v_0_0[2]), .A2(maj_97_n24), .ZN(maj_97_n20) );
  NAND2_X1 maj_97_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_97_n21) );
  NAND2_X1 maj_97_U10 ( .A1(maj_97_n21), .A2(maj_97_n20), .ZN(maj_97_n23) );
  XOR2_X1 maj_97_U9 ( .A(v_0_0[2]), .B(maj_97_n24), .Z(maj_97_n26) );
  XOR2_X1 maj_97_U8 ( .A(v_0_0[5]), .B(maj_97_n25), .Z(maj_97_n27) );
  XOR2_X1 maj_97_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_97_n24) );
  XOR2_X1 maj_97_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_97_n25) );
  OR2_X1 maj_97_U5 ( .A1(maj_97_n23), .A2(maj_97_n22), .ZN(maj_97_n32) );
  NAND2_X1 maj_97_U4 ( .A1(maj_97_n22), .A2(maj_97_n23), .ZN(maj_97_n34) );
  NAND2_X1 maj_97_U3 ( .A1(maj_97_n32), .A2(maj_97_n31), .ZN(maj_97_n33) );
  NAND2_X1 maj_97_U2 ( .A1(maj_97_n34), .A2(maj_97_n33), .ZN(maj_97_port_o) );
  OR2_X1 maj_98_U19 ( .A1(maj_98_n27), .A2(maj_98_n26), .ZN(maj_98_n28) );
  NAND2_X1 maj_98_U18 ( .A1(u_0_1[6]), .A2(maj_98_n28), .ZN(maj_98_n29) );
  NAND2_X1 maj_98_U17 ( .A1(maj_98_n26), .A2(maj_98_n27), .ZN(maj_98_n30) );
  NAND2_X1 maj_98_U16 ( .A1(maj_98_n30), .A2(maj_98_n29), .ZN(maj_98_n31) );
  NAND2_X1 maj_98_U15 ( .A1(u_0_1[5]), .A2(maj_98_n25), .ZN(maj_98_n18) );
  NAND2_X1 maj_98_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_98_n19) );
  NAND2_X1 maj_98_U13 ( .A1(maj_98_n19), .A2(maj_98_n18), .ZN(maj_98_n22) );
  NAND2_X1 maj_98_U12 ( .A1(u_0_1[2]), .A2(maj_98_n24), .ZN(maj_98_n20) );
  NAND2_X1 maj_98_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_98_n21) );
  NAND2_X1 maj_98_U10 ( .A1(maj_98_n21), .A2(maj_98_n20), .ZN(maj_98_n23) );
  XOR2_X1 maj_98_U9 ( .A(u_0_1[2]), .B(maj_98_n24), .Z(maj_98_n26) );
  XOR2_X1 maj_98_U8 ( .A(u_0_1[5]), .B(maj_98_n25), .Z(maj_98_n27) );
  XOR2_X1 maj_98_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_98_n24) );
  XOR2_X1 maj_98_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_98_n25) );
  OR2_X1 maj_98_U5 ( .A1(maj_98_n23), .A2(maj_98_n22), .ZN(maj_98_n32) );
  NAND2_X1 maj_98_U4 ( .A1(maj_98_n22), .A2(maj_98_n23), .ZN(maj_98_n34) );
  NAND2_X1 maj_98_U3 ( .A1(maj_98_n32), .A2(maj_98_n31), .ZN(maj_98_n33) );
  NAND2_X1 maj_98_U2 ( .A1(maj_98_n34), .A2(maj_98_n33), .ZN(maj_98_port_o) );
  OR2_X1 maj_99_U19 ( .A1(maj_99_n27), .A2(maj_99_n26), .ZN(maj_99_n28) );
  NAND2_X1 maj_99_U18 ( .A1(v_0_1[6]), .A2(maj_99_n28), .ZN(maj_99_n29) );
  NAND2_X1 maj_99_U17 ( .A1(maj_99_n26), .A2(maj_99_n27), .ZN(maj_99_n30) );
  NAND2_X1 maj_99_U16 ( .A1(maj_99_n30), .A2(maj_99_n29), .ZN(maj_99_n31) );
  NAND2_X1 maj_99_U15 ( .A1(v_0_1[5]), .A2(maj_99_n25), .ZN(maj_99_n18) );
  NAND2_X1 maj_99_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_99_n19) );
  NAND2_X1 maj_99_U13 ( .A1(maj_99_n19), .A2(maj_99_n18), .ZN(maj_99_n22) );
  NAND2_X1 maj_99_U12 ( .A1(v_0_1[2]), .A2(maj_99_n24), .ZN(maj_99_n20) );
  NAND2_X1 maj_99_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_99_n21) );
  NAND2_X1 maj_99_U10 ( .A1(maj_99_n21), .A2(maj_99_n20), .ZN(maj_99_n23) );
  XOR2_X1 maj_99_U9 ( .A(v_0_1[2]), .B(maj_99_n24), .Z(maj_99_n26) );
  XOR2_X1 maj_99_U8 ( .A(v_0_1[5]), .B(maj_99_n25), .Z(maj_99_n27) );
  XOR2_X1 maj_99_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_99_n24) );
  XOR2_X1 maj_99_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_99_n25) );
  OR2_X1 maj_99_U5 ( .A1(maj_99_n23), .A2(maj_99_n22), .ZN(maj_99_n32) );
  NAND2_X1 maj_99_U4 ( .A1(maj_99_n22), .A2(maj_99_n23), .ZN(maj_99_n34) );
  NAND2_X1 maj_99_U3 ( .A1(maj_99_n32), .A2(maj_99_n31), .ZN(maj_99_n33) );
  NAND2_X1 maj_99_U2 ( .A1(maj_99_n34), .A2(maj_99_n33), .ZN(maj_99_port_o) );
  OR2_X1 maj_100_U19 ( .A1(maj_100_n27), .A2(maj_100_n26), .ZN(maj_100_n28) );
  NAND2_X1 maj_100_U18 ( .A1(u_1_0[6]), .A2(maj_100_n28), .ZN(maj_100_n29) );
  NAND2_X1 maj_100_U17 ( .A1(maj_100_n26), .A2(maj_100_n27), .ZN(maj_100_n30)
         );
  NAND2_X1 maj_100_U16 ( .A1(maj_100_n30), .A2(maj_100_n29), .ZN(maj_100_n31)
         );
  NAND2_X1 maj_100_U15 ( .A1(u_1_0[5]), .A2(maj_100_n25), .ZN(maj_100_n18) );
  NAND2_X1 maj_100_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_100_n19) );
  NAND2_X1 maj_100_U13 ( .A1(maj_100_n19), .A2(maj_100_n18), .ZN(maj_100_n22)
         );
  NAND2_X1 maj_100_U12 ( .A1(u_1_0[2]), .A2(maj_100_n24), .ZN(maj_100_n20) );
  NAND2_X1 maj_100_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_100_n21) );
  NAND2_X1 maj_100_U10 ( .A1(maj_100_n21), .A2(maj_100_n20), .ZN(maj_100_n23)
         );
  XOR2_X1 maj_100_U9 ( .A(u_1_0[2]), .B(maj_100_n24), .Z(maj_100_n26) );
  XOR2_X1 maj_100_U8 ( .A(u_1_0[5]), .B(maj_100_n25), .Z(maj_100_n27) );
  XOR2_X1 maj_100_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_100_n24) );
  XOR2_X1 maj_100_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_100_n25) );
  OR2_X1 maj_100_U5 ( .A1(maj_100_n23), .A2(maj_100_n22), .ZN(maj_100_n32) );
  NAND2_X1 maj_100_U4 ( .A1(maj_100_n22), .A2(maj_100_n23), .ZN(maj_100_n34)
         );
  NAND2_X1 maj_100_U3 ( .A1(maj_100_n32), .A2(maj_100_n31), .ZN(maj_100_n33)
         );
  NAND2_X1 maj_100_U2 ( .A1(maj_100_n34), .A2(maj_100_n33), .ZN(maj_100_port_o) );
  OR2_X1 maj_101_U19 ( .A1(maj_101_n27), .A2(maj_101_n26), .ZN(maj_101_n28) );
  NAND2_X1 maj_101_U18 ( .A1(v_1_0[6]), .A2(maj_101_n28), .ZN(maj_101_n29) );
  NAND2_X1 maj_101_U17 ( .A1(maj_101_n26), .A2(maj_101_n27), .ZN(maj_101_n30)
         );
  NAND2_X1 maj_101_U16 ( .A1(maj_101_n30), .A2(maj_101_n29), .ZN(maj_101_n31)
         );
  NAND2_X1 maj_101_U15 ( .A1(v_1_0[5]), .A2(maj_101_n25), .ZN(maj_101_n18) );
  NAND2_X1 maj_101_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_101_n19) );
  NAND2_X1 maj_101_U13 ( .A1(maj_101_n19), .A2(maj_101_n18), .ZN(maj_101_n22)
         );
  NAND2_X1 maj_101_U12 ( .A1(v_1_0[2]), .A2(maj_101_n24), .ZN(maj_101_n20) );
  NAND2_X1 maj_101_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_101_n21) );
  NAND2_X1 maj_101_U10 ( .A1(maj_101_n21), .A2(maj_101_n20), .ZN(maj_101_n23)
         );
  XOR2_X1 maj_101_U9 ( .A(v_1_0[2]), .B(maj_101_n24), .Z(maj_101_n26) );
  XOR2_X1 maj_101_U8 ( .A(v_1_0[5]), .B(maj_101_n25), .Z(maj_101_n27) );
  XOR2_X1 maj_101_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_101_n24) );
  XOR2_X1 maj_101_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_101_n25) );
  OR2_X1 maj_101_U5 ( .A1(maj_101_n23), .A2(maj_101_n22), .ZN(maj_101_n32) );
  NAND2_X1 maj_101_U4 ( .A1(maj_101_n22), .A2(maj_101_n23), .ZN(maj_101_n34)
         );
  NAND2_X1 maj_101_U3 ( .A1(maj_101_n32), .A2(maj_101_n31), .ZN(maj_101_n33)
         );
  NAND2_X1 maj_101_U2 ( .A1(maj_101_n34), .A2(maj_101_n33), .ZN(maj_101_port_o) );
  OR2_X1 maj_102_U19 ( .A1(maj_102_n27), .A2(maj_102_n26), .ZN(maj_102_n28) );
  NAND2_X1 maj_102_U18 ( .A1(u_1_1[6]), .A2(maj_102_n28), .ZN(maj_102_n29) );
  NAND2_X1 maj_102_U17 ( .A1(maj_102_n26), .A2(maj_102_n27), .ZN(maj_102_n30)
         );
  NAND2_X1 maj_102_U16 ( .A1(maj_102_n30), .A2(maj_102_n29), .ZN(maj_102_n31)
         );
  NAND2_X1 maj_102_U15 ( .A1(u_1_1[5]), .A2(maj_102_n25), .ZN(maj_102_n18) );
  NAND2_X1 maj_102_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_102_n19) );
  NAND2_X1 maj_102_U13 ( .A1(maj_102_n19), .A2(maj_102_n18), .ZN(maj_102_n22)
         );
  NAND2_X1 maj_102_U12 ( .A1(u_1_1[2]), .A2(maj_102_n24), .ZN(maj_102_n20) );
  NAND2_X1 maj_102_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_102_n21) );
  NAND2_X1 maj_102_U10 ( .A1(maj_102_n21), .A2(maj_102_n20), .ZN(maj_102_n23)
         );
  XOR2_X1 maj_102_U9 ( .A(u_1_1[2]), .B(maj_102_n24), .Z(maj_102_n26) );
  XOR2_X1 maj_102_U8 ( .A(u_1_1[5]), .B(maj_102_n25), .Z(maj_102_n27) );
  XOR2_X1 maj_102_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_102_n24) );
  XOR2_X1 maj_102_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_102_n25) );
  OR2_X1 maj_102_U5 ( .A1(maj_102_n23), .A2(maj_102_n22), .ZN(maj_102_n32) );
  NAND2_X1 maj_102_U4 ( .A1(maj_102_n22), .A2(maj_102_n23), .ZN(maj_102_n34)
         );
  NAND2_X1 maj_102_U3 ( .A1(maj_102_n32), .A2(maj_102_n31), .ZN(maj_102_n33)
         );
  NAND2_X1 maj_102_U2 ( .A1(maj_102_n34), .A2(maj_102_n33), .ZN(maj_102_port_o) );
  OR2_X1 maj_103_U19 ( .A1(maj_103_n27), .A2(maj_103_n26), .ZN(maj_103_n28) );
  NAND2_X1 maj_103_U18 ( .A1(v_1_1[6]), .A2(maj_103_n28), .ZN(maj_103_n29) );
  NAND2_X1 maj_103_U17 ( .A1(maj_103_n26), .A2(maj_103_n27), .ZN(maj_103_n30)
         );
  NAND2_X1 maj_103_U16 ( .A1(maj_103_n30), .A2(maj_103_n29), .ZN(maj_103_n31)
         );
  NAND2_X1 maj_103_U15 ( .A1(v_1_1[5]), .A2(maj_103_n25), .ZN(maj_103_n18) );
  NAND2_X1 maj_103_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_103_n19) );
  NAND2_X1 maj_103_U13 ( .A1(maj_103_n19), .A2(maj_103_n18), .ZN(maj_103_n22)
         );
  NAND2_X1 maj_103_U12 ( .A1(v_1_1[2]), .A2(maj_103_n24), .ZN(maj_103_n20) );
  NAND2_X1 maj_103_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_103_n21) );
  NAND2_X1 maj_103_U10 ( .A1(maj_103_n21), .A2(maj_103_n20), .ZN(maj_103_n23)
         );
  XOR2_X1 maj_103_U9 ( .A(v_1_1[2]), .B(maj_103_n24), .Z(maj_103_n26) );
  XOR2_X1 maj_103_U8 ( .A(v_1_1[5]), .B(maj_103_n25), .Z(maj_103_n27) );
  XOR2_X1 maj_103_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_103_n24) );
  XOR2_X1 maj_103_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_103_n25) );
  OR2_X1 maj_103_U5 ( .A1(maj_103_n23), .A2(maj_103_n22), .ZN(maj_103_n32) );
  NAND2_X1 maj_103_U4 ( .A1(maj_103_n22), .A2(maj_103_n23), .ZN(maj_103_n34)
         );
  NAND2_X1 maj_103_U3 ( .A1(maj_103_n32), .A2(maj_103_n31), .ZN(maj_103_n33)
         );
  NAND2_X1 maj_103_U2 ( .A1(maj_103_n34), .A2(maj_103_n33), .ZN(maj_103_port_o) );
  OR2_X1 maj_104_U19 ( .A1(maj_104_n27), .A2(maj_104_n26), .ZN(maj_104_n28) );
  NAND2_X1 maj_104_U18 ( .A1(u_2_0[6]), .A2(maj_104_n28), .ZN(maj_104_n29) );
  NAND2_X1 maj_104_U17 ( .A1(maj_104_n26), .A2(maj_104_n27), .ZN(maj_104_n30)
         );
  NAND2_X1 maj_104_U16 ( .A1(maj_104_n30), .A2(maj_104_n29), .ZN(maj_104_n31)
         );
  NAND2_X1 maj_104_U15 ( .A1(u_2_0[5]), .A2(maj_104_n25), .ZN(maj_104_n18) );
  NAND2_X1 maj_104_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_104_n19) );
  NAND2_X1 maj_104_U13 ( .A1(maj_104_n19), .A2(maj_104_n18), .ZN(maj_104_n22)
         );
  NAND2_X1 maj_104_U12 ( .A1(u_2_0[2]), .A2(maj_104_n24), .ZN(maj_104_n20) );
  NAND2_X1 maj_104_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_104_n21) );
  NAND2_X1 maj_104_U10 ( .A1(maj_104_n21), .A2(maj_104_n20), .ZN(maj_104_n23)
         );
  XOR2_X1 maj_104_U9 ( .A(u_2_0[2]), .B(maj_104_n24), .Z(maj_104_n26) );
  XOR2_X1 maj_104_U8 ( .A(u_2_0[5]), .B(maj_104_n25), .Z(maj_104_n27) );
  XOR2_X1 maj_104_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_104_n24) );
  XOR2_X1 maj_104_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_104_n25) );
  OR2_X1 maj_104_U5 ( .A1(maj_104_n23), .A2(maj_104_n22), .ZN(maj_104_n32) );
  NAND2_X1 maj_104_U4 ( .A1(maj_104_n22), .A2(maj_104_n23), .ZN(maj_104_n34)
         );
  NAND2_X1 maj_104_U3 ( .A1(maj_104_n32), .A2(maj_104_n31), .ZN(maj_104_n33)
         );
  NAND2_X1 maj_104_U2 ( .A1(maj_104_n34), .A2(maj_104_n33), .ZN(maj_104_port_o) );
  OR2_X1 maj_105_U19 ( .A1(maj_105_n27), .A2(maj_105_n26), .ZN(maj_105_n28) );
  NAND2_X1 maj_105_U18 ( .A1(v_2_0[6]), .A2(maj_105_n28), .ZN(maj_105_n29) );
  NAND2_X1 maj_105_U17 ( .A1(maj_105_n26), .A2(maj_105_n27), .ZN(maj_105_n30)
         );
  NAND2_X1 maj_105_U16 ( .A1(maj_105_n30), .A2(maj_105_n29), .ZN(maj_105_n31)
         );
  NAND2_X1 maj_105_U15 ( .A1(v_2_0[5]), .A2(maj_105_n25), .ZN(maj_105_n18) );
  NAND2_X1 maj_105_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_105_n19) );
  NAND2_X1 maj_105_U13 ( .A1(maj_105_n19), .A2(maj_105_n18), .ZN(maj_105_n22)
         );
  NAND2_X1 maj_105_U12 ( .A1(v_2_0[2]), .A2(maj_105_n24), .ZN(maj_105_n20) );
  NAND2_X1 maj_105_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_105_n21) );
  NAND2_X1 maj_105_U10 ( .A1(maj_105_n21), .A2(maj_105_n20), .ZN(maj_105_n23)
         );
  XOR2_X1 maj_105_U9 ( .A(v_2_0[2]), .B(maj_105_n24), .Z(maj_105_n26) );
  XOR2_X1 maj_105_U8 ( .A(v_2_0[5]), .B(maj_105_n25), .Z(maj_105_n27) );
  XOR2_X1 maj_105_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_105_n24) );
  XOR2_X1 maj_105_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_105_n25) );
  OR2_X1 maj_105_U5 ( .A1(maj_105_n23), .A2(maj_105_n22), .ZN(maj_105_n32) );
  NAND2_X1 maj_105_U4 ( .A1(maj_105_n22), .A2(maj_105_n23), .ZN(maj_105_n34)
         );
  NAND2_X1 maj_105_U3 ( .A1(maj_105_n32), .A2(maj_105_n31), .ZN(maj_105_n33)
         );
  NAND2_X1 maj_105_U2 ( .A1(maj_105_n34), .A2(maj_105_n33), .ZN(maj_105_port_o) );
  OR2_X1 maj_106_U19 ( .A1(maj_106_n27), .A2(maj_106_n26), .ZN(maj_106_n28) );
  NAND2_X1 maj_106_U18 ( .A1(u_2_1[6]), .A2(maj_106_n28), .ZN(maj_106_n29) );
  NAND2_X1 maj_106_U17 ( .A1(maj_106_n26), .A2(maj_106_n27), .ZN(maj_106_n30)
         );
  NAND2_X1 maj_106_U16 ( .A1(maj_106_n30), .A2(maj_106_n29), .ZN(maj_106_n31)
         );
  NAND2_X1 maj_106_U15 ( .A1(u_2_1[5]), .A2(maj_106_n25), .ZN(maj_106_n18) );
  NAND2_X1 maj_106_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_106_n19) );
  NAND2_X1 maj_106_U13 ( .A1(maj_106_n19), .A2(maj_106_n18), .ZN(maj_106_n22)
         );
  NAND2_X1 maj_106_U12 ( .A1(u_2_1[2]), .A2(maj_106_n24), .ZN(maj_106_n20) );
  NAND2_X1 maj_106_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_106_n21) );
  NAND2_X1 maj_106_U10 ( .A1(maj_106_n21), .A2(maj_106_n20), .ZN(maj_106_n23)
         );
  XOR2_X1 maj_106_U9 ( .A(u_2_1[2]), .B(maj_106_n24), .Z(maj_106_n26) );
  XOR2_X1 maj_106_U8 ( .A(u_2_1[5]), .B(maj_106_n25), .Z(maj_106_n27) );
  XOR2_X1 maj_106_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_106_n24) );
  XOR2_X1 maj_106_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_106_n25) );
  OR2_X1 maj_106_U5 ( .A1(maj_106_n23), .A2(maj_106_n22), .ZN(maj_106_n32) );
  NAND2_X1 maj_106_U4 ( .A1(maj_106_n22), .A2(maj_106_n23), .ZN(maj_106_n34)
         );
  NAND2_X1 maj_106_U3 ( .A1(maj_106_n32), .A2(maj_106_n31), .ZN(maj_106_n33)
         );
  NAND2_X1 maj_106_U2 ( .A1(maj_106_n34), .A2(maj_106_n33), .ZN(maj_106_port_o) );
  OR2_X1 maj_107_U19 ( .A1(maj_107_n27), .A2(maj_107_n26), .ZN(maj_107_n28) );
  NAND2_X1 maj_107_U18 ( .A1(v_2_1[6]), .A2(maj_107_n28), .ZN(maj_107_n29) );
  NAND2_X1 maj_107_U17 ( .A1(maj_107_n26), .A2(maj_107_n27), .ZN(maj_107_n30)
         );
  NAND2_X1 maj_107_U16 ( .A1(maj_107_n30), .A2(maj_107_n29), .ZN(maj_107_n31)
         );
  NAND2_X1 maj_107_U15 ( .A1(v_2_1[5]), .A2(maj_107_n25), .ZN(maj_107_n18) );
  NAND2_X1 maj_107_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_107_n19) );
  NAND2_X1 maj_107_U13 ( .A1(maj_107_n19), .A2(maj_107_n18), .ZN(maj_107_n22)
         );
  NAND2_X1 maj_107_U12 ( .A1(v_2_1[2]), .A2(maj_107_n24), .ZN(maj_107_n20) );
  NAND2_X1 maj_107_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_107_n21) );
  NAND2_X1 maj_107_U10 ( .A1(maj_107_n21), .A2(maj_107_n20), .ZN(maj_107_n23)
         );
  XOR2_X1 maj_107_U9 ( .A(v_2_1[2]), .B(maj_107_n24), .Z(maj_107_n26) );
  XOR2_X1 maj_107_U8 ( .A(v_2_1[5]), .B(maj_107_n25), .Z(maj_107_n27) );
  XOR2_X1 maj_107_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_107_n24) );
  XOR2_X1 maj_107_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_107_n25) );
  OR2_X1 maj_107_U5 ( .A1(maj_107_n23), .A2(maj_107_n22), .ZN(maj_107_n32) );
  NAND2_X1 maj_107_U4 ( .A1(maj_107_n22), .A2(maj_107_n23), .ZN(maj_107_n34)
         );
  NAND2_X1 maj_107_U3 ( .A1(maj_107_n32), .A2(maj_107_n31), .ZN(maj_107_n33)
         );
  NAND2_X1 maj_107_U2 ( .A1(maj_107_n34), .A2(maj_107_n33), .ZN(maj_107_port_o) );
  OR2_X1 maj_108_U19 ( .A1(maj_108_n27), .A2(maj_108_n26), .ZN(maj_108_n28) );
  NAND2_X1 maj_108_U18 ( .A1(u_0_0[6]), .A2(maj_108_n28), .ZN(maj_108_n29) );
  NAND2_X1 maj_108_U17 ( .A1(maj_108_n26), .A2(maj_108_n27), .ZN(maj_108_n30)
         );
  NAND2_X1 maj_108_U16 ( .A1(maj_108_n30), .A2(maj_108_n29), .ZN(maj_108_n31)
         );
  NAND2_X1 maj_108_U15 ( .A1(u_0_0[5]), .A2(maj_108_n25), .ZN(maj_108_n18) );
  NAND2_X1 maj_108_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_108_n19) );
  NAND2_X1 maj_108_U13 ( .A1(maj_108_n19), .A2(maj_108_n18), .ZN(maj_108_n22)
         );
  NAND2_X1 maj_108_U12 ( .A1(u_0_0[2]), .A2(maj_108_n24), .ZN(maj_108_n20) );
  NAND2_X1 maj_108_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_108_n21) );
  NAND2_X1 maj_108_U10 ( .A1(maj_108_n21), .A2(maj_108_n20), .ZN(maj_108_n23)
         );
  XOR2_X1 maj_108_U9 ( .A(u_0_0[2]), .B(maj_108_n24), .Z(maj_108_n26) );
  XOR2_X1 maj_108_U8 ( .A(u_0_0[5]), .B(maj_108_n25), .Z(maj_108_n27) );
  XOR2_X1 maj_108_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_108_n24) );
  XOR2_X1 maj_108_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_108_n25) );
  OR2_X1 maj_108_U5 ( .A1(maj_108_n23), .A2(maj_108_n22), .ZN(maj_108_n32) );
  NAND2_X1 maj_108_U4 ( .A1(maj_108_n22), .A2(maj_108_n23), .ZN(maj_108_n34)
         );
  NAND2_X1 maj_108_U3 ( .A1(maj_108_n32), .A2(maj_108_n31), .ZN(maj_108_n33)
         );
  NAND2_X1 maj_108_U2 ( .A1(maj_108_n34), .A2(maj_108_n33), .ZN(maj_108_port_o) );
  OR2_X1 maj_109_U19 ( .A1(maj_109_n27), .A2(maj_109_n26), .ZN(maj_109_n28) );
  NAND2_X1 maj_109_U18 ( .A1(v_0_0[6]), .A2(maj_109_n28), .ZN(maj_109_n29) );
  NAND2_X1 maj_109_U17 ( .A1(maj_109_n26), .A2(maj_109_n27), .ZN(maj_109_n30)
         );
  NAND2_X1 maj_109_U16 ( .A1(maj_109_n30), .A2(maj_109_n29), .ZN(maj_109_n31)
         );
  NAND2_X1 maj_109_U15 ( .A1(v_0_0[5]), .A2(maj_109_n25), .ZN(maj_109_n18) );
  NAND2_X1 maj_109_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_109_n19) );
  NAND2_X1 maj_109_U13 ( .A1(maj_109_n19), .A2(maj_109_n18), .ZN(maj_109_n22)
         );
  NAND2_X1 maj_109_U12 ( .A1(v_0_0[2]), .A2(maj_109_n24), .ZN(maj_109_n20) );
  NAND2_X1 maj_109_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_109_n21) );
  NAND2_X1 maj_109_U10 ( .A1(maj_109_n21), .A2(maj_109_n20), .ZN(maj_109_n23)
         );
  XOR2_X1 maj_109_U9 ( .A(v_0_0[2]), .B(maj_109_n24), .Z(maj_109_n26) );
  XOR2_X1 maj_109_U8 ( .A(v_0_0[5]), .B(maj_109_n25), .Z(maj_109_n27) );
  XOR2_X1 maj_109_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_109_n24) );
  XOR2_X1 maj_109_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_109_n25) );
  OR2_X1 maj_109_U5 ( .A1(maj_109_n23), .A2(maj_109_n22), .ZN(maj_109_n32) );
  NAND2_X1 maj_109_U4 ( .A1(maj_109_n22), .A2(maj_109_n23), .ZN(maj_109_n34)
         );
  NAND2_X1 maj_109_U3 ( .A1(maj_109_n32), .A2(maj_109_n31), .ZN(maj_109_n33)
         );
  NAND2_X1 maj_109_U2 ( .A1(maj_109_n34), .A2(maj_109_n33), .ZN(maj_109_port_o) );
  OR2_X1 maj_110_U19 ( .A1(maj_110_n27), .A2(maj_110_n26), .ZN(maj_110_n28) );
  NAND2_X1 maj_110_U18 ( .A1(u_0_1[6]), .A2(maj_110_n28), .ZN(maj_110_n29) );
  NAND2_X1 maj_110_U17 ( .A1(maj_110_n26), .A2(maj_110_n27), .ZN(maj_110_n30)
         );
  NAND2_X1 maj_110_U16 ( .A1(maj_110_n30), .A2(maj_110_n29), .ZN(maj_110_n31)
         );
  NAND2_X1 maj_110_U15 ( .A1(u_0_1[5]), .A2(maj_110_n25), .ZN(maj_110_n18) );
  NAND2_X1 maj_110_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_110_n19) );
  NAND2_X1 maj_110_U13 ( .A1(maj_110_n19), .A2(maj_110_n18), .ZN(maj_110_n22)
         );
  NAND2_X1 maj_110_U12 ( .A1(u_0_1[2]), .A2(maj_110_n24), .ZN(maj_110_n20) );
  NAND2_X1 maj_110_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_110_n21) );
  NAND2_X1 maj_110_U10 ( .A1(maj_110_n21), .A2(maj_110_n20), .ZN(maj_110_n23)
         );
  XOR2_X1 maj_110_U9 ( .A(u_0_1[2]), .B(maj_110_n24), .Z(maj_110_n26) );
  XOR2_X1 maj_110_U8 ( .A(u_0_1[5]), .B(maj_110_n25), .Z(maj_110_n27) );
  XOR2_X1 maj_110_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_110_n24) );
  XOR2_X1 maj_110_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_110_n25) );
  OR2_X1 maj_110_U5 ( .A1(maj_110_n23), .A2(maj_110_n22), .ZN(maj_110_n32) );
  NAND2_X1 maj_110_U4 ( .A1(maj_110_n22), .A2(maj_110_n23), .ZN(maj_110_n34)
         );
  NAND2_X1 maj_110_U3 ( .A1(maj_110_n32), .A2(maj_110_n31), .ZN(maj_110_n33)
         );
  NAND2_X1 maj_110_U2 ( .A1(maj_110_n34), .A2(maj_110_n33), .ZN(maj_110_port_o) );
  OR2_X1 maj_111_U19 ( .A1(maj_111_n27), .A2(maj_111_n26), .ZN(maj_111_n28) );
  NAND2_X1 maj_111_U18 ( .A1(v_0_1[6]), .A2(maj_111_n28), .ZN(maj_111_n29) );
  NAND2_X1 maj_111_U17 ( .A1(maj_111_n26), .A2(maj_111_n27), .ZN(maj_111_n30)
         );
  NAND2_X1 maj_111_U16 ( .A1(maj_111_n30), .A2(maj_111_n29), .ZN(maj_111_n31)
         );
  NAND2_X1 maj_111_U15 ( .A1(v_0_1[5]), .A2(maj_111_n25), .ZN(maj_111_n18) );
  NAND2_X1 maj_111_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_111_n19) );
  NAND2_X1 maj_111_U13 ( .A1(maj_111_n19), .A2(maj_111_n18), .ZN(maj_111_n22)
         );
  NAND2_X1 maj_111_U12 ( .A1(v_0_1[2]), .A2(maj_111_n24), .ZN(maj_111_n20) );
  NAND2_X1 maj_111_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_111_n21) );
  NAND2_X1 maj_111_U10 ( .A1(maj_111_n21), .A2(maj_111_n20), .ZN(maj_111_n23)
         );
  XOR2_X1 maj_111_U9 ( .A(v_0_1[2]), .B(maj_111_n24), .Z(maj_111_n26) );
  XOR2_X1 maj_111_U8 ( .A(v_0_1[5]), .B(maj_111_n25), .Z(maj_111_n27) );
  XOR2_X1 maj_111_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_111_n24) );
  XOR2_X1 maj_111_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_111_n25) );
  OR2_X1 maj_111_U5 ( .A1(maj_111_n23), .A2(maj_111_n22), .ZN(maj_111_n32) );
  NAND2_X1 maj_111_U4 ( .A1(maj_111_n22), .A2(maj_111_n23), .ZN(maj_111_n34)
         );
  NAND2_X1 maj_111_U3 ( .A1(maj_111_n32), .A2(maj_111_n31), .ZN(maj_111_n33)
         );
  NAND2_X1 maj_111_U2 ( .A1(maj_111_n34), .A2(maj_111_n33), .ZN(maj_111_port_o) );
  OR2_X1 maj_112_U19 ( .A1(maj_112_n27), .A2(maj_112_n26), .ZN(maj_112_n28) );
  NAND2_X1 maj_112_U18 ( .A1(u_1_0[6]), .A2(maj_112_n28), .ZN(maj_112_n29) );
  NAND2_X1 maj_112_U17 ( .A1(maj_112_n26), .A2(maj_112_n27), .ZN(maj_112_n30)
         );
  NAND2_X1 maj_112_U16 ( .A1(maj_112_n30), .A2(maj_112_n29), .ZN(maj_112_n31)
         );
  NAND2_X1 maj_112_U15 ( .A1(u_1_0[5]), .A2(maj_112_n25), .ZN(maj_112_n18) );
  NAND2_X1 maj_112_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_112_n19) );
  NAND2_X1 maj_112_U13 ( .A1(maj_112_n19), .A2(maj_112_n18), .ZN(maj_112_n22)
         );
  NAND2_X1 maj_112_U12 ( .A1(u_1_0[2]), .A2(maj_112_n24), .ZN(maj_112_n20) );
  NAND2_X1 maj_112_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_112_n21) );
  NAND2_X1 maj_112_U10 ( .A1(maj_112_n21), .A2(maj_112_n20), .ZN(maj_112_n23)
         );
  XOR2_X1 maj_112_U9 ( .A(u_1_0[2]), .B(maj_112_n24), .Z(maj_112_n26) );
  XOR2_X1 maj_112_U8 ( .A(u_1_0[5]), .B(maj_112_n25), .Z(maj_112_n27) );
  XOR2_X1 maj_112_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_112_n24) );
  XOR2_X1 maj_112_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_112_n25) );
  OR2_X1 maj_112_U5 ( .A1(maj_112_n23), .A2(maj_112_n22), .ZN(maj_112_n32) );
  NAND2_X1 maj_112_U4 ( .A1(maj_112_n22), .A2(maj_112_n23), .ZN(maj_112_n34)
         );
  NAND2_X1 maj_112_U3 ( .A1(maj_112_n32), .A2(maj_112_n31), .ZN(maj_112_n33)
         );
  NAND2_X1 maj_112_U2 ( .A1(maj_112_n34), .A2(maj_112_n33), .ZN(maj_112_port_o) );
  OR2_X1 maj_113_U19 ( .A1(maj_113_n27), .A2(maj_113_n26), .ZN(maj_113_n28) );
  NAND2_X1 maj_113_U18 ( .A1(v_1_0[6]), .A2(maj_113_n28), .ZN(maj_113_n29) );
  NAND2_X1 maj_113_U17 ( .A1(maj_113_n26), .A2(maj_113_n27), .ZN(maj_113_n30)
         );
  NAND2_X1 maj_113_U16 ( .A1(maj_113_n30), .A2(maj_113_n29), .ZN(maj_113_n31)
         );
  NAND2_X1 maj_113_U15 ( .A1(v_1_0[5]), .A2(maj_113_n25), .ZN(maj_113_n18) );
  NAND2_X1 maj_113_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_113_n19) );
  NAND2_X1 maj_113_U13 ( .A1(maj_113_n19), .A2(maj_113_n18), .ZN(maj_113_n22)
         );
  NAND2_X1 maj_113_U12 ( .A1(v_1_0[2]), .A2(maj_113_n24), .ZN(maj_113_n20) );
  NAND2_X1 maj_113_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_113_n21) );
  NAND2_X1 maj_113_U10 ( .A1(maj_113_n21), .A2(maj_113_n20), .ZN(maj_113_n23)
         );
  XOR2_X1 maj_113_U9 ( .A(v_1_0[2]), .B(maj_113_n24), .Z(maj_113_n26) );
  XOR2_X1 maj_113_U8 ( .A(v_1_0[5]), .B(maj_113_n25), .Z(maj_113_n27) );
  XOR2_X1 maj_113_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_113_n24) );
  XOR2_X1 maj_113_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_113_n25) );
  OR2_X1 maj_113_U5 ( .A1(maj_113_n23), .A2(maj_113_n22), .ZN(maj_113_n32) );
  NAND2_X1 maj_113_U4 ( .A1(maj_113_n22), .A2(maj_113_n23), .ZN(maj_113_n34)
         );
  NAND2_X1 maj_113_U3 ( .A1(maj_113_n32), .A2(maj_113_n31), .ZN(maj_113_n33)
         );
  NAND2_X1 maj_113_U2 ( .A1(maj_113_n34), .A2(maj_113_n33), .ZN(maj_113_port_o) );
  OR2_X1 maj_114_U19 ( .A1(maj_114_n27), .A2(maj_114_n26), .ZN(maj_114_n28) );
  NAND2_X1 maj_114_U18 ( .A1(u_1_1[6]), .A2(maj_114_n28), .ZN(maj_114_n29) );
  NAND2_X1 maj_114_U17 ( .A1(maj_114_n26), .A2(maj_114_n27), .ZN(maj_114_n30)
         );
  NAND2_X1 maj_114_U16 ( .A1(maj_114_n30), .A2(maj_114_n29), .ZN(maj_114_n31)
         );
  NAND2_X1 maj_114_U15 ( .A1(u_1_1[5]), .A2(maj_114_n25), .ZN(maj_114_n18) );
  NAND2_X1 maj_114_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_114_n19) );
  NAND2_X1 maj_114_U13 ( .A1(maj_114_n19), .A2(maj_114_n18), .ZN(maj_114_n22)
         );
  NAND2_X1 maj_114_U12 ( .A1(u_1_1[2]), .A2(maj_114_n24), .ZN(maj_114_n20) );
  NAND2_X1 maj_114_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_114_n21) );
  NAND2_X1 maj_114_U10 ( .A1(maj_114_n21), .A2(maj_114_n20), .ZN(maj_114_n23)
         );
  XOR2_X1 maj_114_U9 ( .A(u_1_1[2]), .B(maj_114_n24), .Z(maj_114_n26) );
  XOR2_X1 maj_114_U8 ( .A(u_1_1[5]), .B(maj_114_n25), .Z(maj_114_n27) );
  XOR2_X1 maj_114_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_114_n24) );
  XOR2_X1 maj_114_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_114_n25) );
  OR2_X1 maj_114_U5 ( .A1(maj_114_n23), .A2(maj_114_n22), .ZN(maj_114_n32) );
  NAND2_X1 maj_114_U4 ( .A1(maj_114_n22), .A2(maj_114_n23), .ZN(maj_114_n34)
         );
  NAND2_X1 maj_114_U3 ( .A1(maj_114_n32), .A2(maj_114_n31), .ZN(maj_114_n33)
         );
  NAND2_X1 maj_114_U2 ( .A1(maj_114_n34), .A2(maj_114_n33), .ZN(maj_114_port_o) );
  OR2_X1 maj_115_U19 ( .A1(maj_115_n27), .A2(maj_115_n26), .ZN(maj_115_n28) );
  NAND2_X1 maj_115_U18 ( .A1(v_1_1[6]), .A2(maj_115_n28), .ZN(maj_115_n29) );
  NAND2_X1 maj_115_U17 ( .A1(maj_115_n26), .A2(maj_115_n27), .ZN(maj_115_n30)
         );
  NAND2_X1 maj_115_U16 ( .A1(maj_115_n30), .A2(maj_115_n29), .ZN(maj_115_n31)
         );
  NAND2_X1 maj_115_U15 ( .A1(v_1_1[5]), .A2(maj_115_n25), .ZN(maj_115_n18) );
  NAND2_X1 maj_115_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_115_n19) );
  NAND2_X1 maj_115_U13 ( .A1(maj_115_n19), .A2(maj_115_n18), .ZN(maj_115_n22)
         );
  NAND2_X1 maj_115_U12 ( .A1(v_1_1[2]), .A2(maj_115_n24), .ZN(maj_115_n20) );
  NAND2_X1 maj_115_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_115_n21) );
  NAND2_X1 maj_115_U10 ( .A1(maj_115_n21), .A2(maj_115_n20), .ZN(maj_115_n23)
         );
  XOR2_X1 maj_115_U9 ( .A(v_1_1[2]), .B(maj_115_n24), .Z(maj_115_n26) );
  XOR2_X1 maj_115_U8 ( .A(v_1_1[5]), .B(maj_115_n25), .Z(maj_115_n27) );
  XOR2_X1 maj_115_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_115_n24) );
  XOR2_X1 maj_115_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_115_n25) );
  OR2_X1 maj_115_U5 ( .A1(maj_115_n23), .A2(maj_115_n22), .ZN(maj_115_n32) );
  NAND2_X1 maj_115_U4 ( .A1(maj_115_n22), .A2(maj_115_n23), .ZN(maj_115_n34)
         );
  NAND2_X1 maj_115_U3 ( .A1(maj_115_n32), .A2(maj_115_n31), .ZN(maj_115_n33)
         );
  NAND2_X1 maj_115_U2 ( .A1(maj_115_n34), .A2(maj_115_n33), .ZN(maj_115_port_o) );
  OR2_X1 maj_116_U19 ( .A1(maj_116_n27), .A2(maj_116_n26), .ZN(maj_116_n28) );
  NAND2_X1 maj_116_U18 ( .A1(u_2_0[6]), .A2(maj_116_n28), .ZN(maj_116_n29) );
  NAND2_X1 maj_116_U17 ( .A1(maj_116_n26), .A2(maj_116_n27), .ZN(maj_116_n30)
         );
  NAND2_X1 maj_116_U16 ( .A1(maj_116_n30), .A2(maj_116_n29), .ZN(maj_116_n31)
         );
  NAND2_X1 maj_116_U15 ( .A1(u_2_0[5]), .A2(maj_116_n25), .ZN(maj_116_n18) );
  NAND2_X1 maj_116_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_116_n19) );
  NAND2_X1 maj_116_U13 ( .A1(maj_116_n19), .A2(maj_116_n18), .ZN(maj_116_n22)
         );
  NAND2_X1 maj_116_U12 ( .A1(u_2_0[2]), .A2(maj_116_n24), .ZN(maj_116_n20) );
  NAND2_X1 maj_116_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_116_n21) );
  NAND2_X1 maj_116_U10 ( .A1(maj_116_n21), .A2(maj_116_n20), .ZN(maj_116_n23)
         );
  XOR2_X1 maj_116_U9 ( .A(u_2_0[2]), .B(maj_116_n24), .Z(maj_116_n26) );
  XOR2_X1 maj_116_U8 ( .A(u_2_0[5]), .B(maj_116_n25), .Z(maj_116_n27) );
  XOR2_X1 maj_116_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_116_n24) );
  XOR2_X1 maj_116_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_116_n25) );
  OR2_X1 maj_116_U5 ( .A1(maj_116_n23), .A2(maj_116_n22), .ZN(maj_116_n32) );
  NAND2_X1 maj_116_U4 ( .A1(maj_116_n22), .A2(maj_116_n23), .ZN(maj_116_n34)
         );
  NAND2_X1 maj_116_U3 ( .A1(maj_116_n32), .A2(maj_116_n31), .ZN(maj_116_n33)
         );
  NAND2_X1 maj_116_U2 ( .A1(maj_116_n34), .A2(maj_116_n33), .ZN(maj_116_port_o) );
  OR2_X1 maj_117_U19 ( .A1(maj_117_n27), .A2(maj_117_n26), .ZN(maj_117_n28) );
  NAND2_X1 maj_117_U18 ( .A1(v_2_0[6]), .A2(maj_117_n28), .ZN(maj_117_n29) );
  NAND2_X1 maj_117_U17 ( .A1(maj_117_n26), .A2(maj_117_n27), .ZN(maj_117_n30)
         );
  NAND2_X1 maj_117_U16 ( .A1(maj_117_n30), .A2(maj_117_n29), .ZN(maj_117_n31)
         );
  NAND2_X1 maj_117_U15 ( .A1(v_2_0[5]), .A2(maj_117_n25), .ZN(maj_117_n18) );
  NAND2_X1 maj_117_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_117_n19) );
  NAND2_X1 maj_117_U13 ( .A1(maj_117_n19), .A2(maj_117_n18), .ZN(maj_117_n22)
         );
  NAND2_X1 maj_117_U12 ( .A1(v_2_0[2]), .A2(maj_117_n24), .ZN(maj_117_n20) );
  NAND2_X1 maj_117_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_117_n21) );
  NAND2_X1 maj_117_U10 ( .A1(maj_117_n21), .A2(maj_117_n20), .ZN(maj_117_n23)
         );
  XOR2_X1 maj_117_U9 ( .A(v_2_0[2]), .B(maj_117_n24), .Z(maj_117_n26) );
  XOR2_X1 maj_117_U8 ( .A(v_2_0[5]), .B(maj_117_n25), .Z(maj_117_n27) );
  XOR2_X1 maj_117_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_117_n24) );
  XOR2_X1 maj_117_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_117_n25) );
  OR2_X1 maj_117_U5 ( .A1(maj_117_n23), .A2(maj_117_n22), .ZN(maj_117_n32) );
  NAND2_X1 maj_117_U4 ( .A1(maj_117_n22), .A2(maj_117_n23), .ZN(maj_117_n34)
         );
  NAND2_X1 maj_117_U3 ( .A1(maj_117_n32), .A2(maj_117_n31), .ZN(maj_117_n33)
         );
  NAND2_X1 maj_117_U2 ( .A1(maj_117_n34), .A2(maj_117_n33), .ZN(maj_117_port_o) );
  OR2_X1 maj_118_U19 ( .A1(maj_118_n27), .A2(maj_118_n26), .ZN(maj_118_n28) );
  NAND2_X1 maj_118_U18 ( .A1(u_2_1[6]), .A2(maj_118_n28), .ZN(maj_118_n29) );
  NAND2_X1 maj_118_U17 ( .A1(maj_118_n26), .A2(maj_118_n27), .ZN(maj_118_n30)
         );
  NAND2_X1 maj_118_U16 ( .A1(maj_118_n30), .A2(maj_118_n29), .ZN(maj_118_n31)
         );
  NAND2_X1 maj_118_U15 ( .A1(u_2_1[5]), .A2(maj_118_n25), .ZN(maj_118_n18) );
  NAND2_X1 maj_118_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_118_n19) );
  NAND2_X1 maj_118_U13 ( .A1(maj_118_n19), .A2(maj_118_n18), .ZN(maj_118_n22)
         );
  NAND2_X1 maj_118_U12 ( .A1(u_2_1[2]), .A2(maj_118_n24), .ZN(maj_118_n20) );
  NAND2_X1 maj_118_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_118_n21) );
  NAND2_X1 maj_118_U10 ( .A1(maj_118_n21), .A2(maj_118_n20), .ZN(maj_118_n23)
         );
  XOR2_X1 maj_118_U9 ( .A(u_2_1[2]), .B(maj_118_n24), .Z(maj_118_n26) );
  XOR2_X1 maj_118_U8 ( .A(u_2_1[5]), .B(maj_118_n25), .Z(maj_118_n27) );
  XOR2_X1 maj_118_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_118_n24) );
  XOR2_X1 maj_118_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_118_n25) );
  OR2_X1 maj_118_U5 ( .A1(maj_118_n23), .A2(maj_118_n22), .ZN(maj_118_n32) );
  NAND2_X1 maj_118_U4 ( .A1(maj_118_n22), .A2(maj_118_n23), .ZN(maj_118_n34)
         );
  NAND2_X1 maj_118_U3 ( .A1(maj_118_n32), .A2(maj_118_n31), .ZN(maj_118_n33)
         );
  NAND2_X1 maj_118_U2 ( .A1(maj_118_n34), .A2(maj_118_n33), .ZN(maj_118_port_o) );
  OR2_X1 maj_119_U19 ( .A1(maj_119_n27), .A2(maj_119_n26), .ZN(maj_119_n28) );
  NAND2_X1 maj_119_U18 ( .A1(v_2_1[6]), .A2(maj_119_n28), .ZN(maj_119_n29) );
  NAND2_X1 maj_119_U17 ( .A1(maj_119_n26), .A2(maj_119_n27), .ZN(maj_119_n30)
         );
  NAND2_X1 maj_119_U16 ( .A1(maj_119_n30), .A2(maj_119_n29), .ZN(maj_119_n31)
         );
  NAND2_X1 maj_119_U15 ( .A1(v_2_1[5]), .A2(maj_119_n25), .ZN(maj_119_n18) );
  NAND2_X1 maj_119_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_119_n19) );
  NAND2_X1 maj_119_U13 ( .A1(maj_119_n19), .A2(maj_119_n18), .ZN(maj_119_n22)
         );
  NAND2_X1 maj_119_U12 ( .A1(v_2_1[2]), .A2(maj_119_n24), .ZN(maj_119_n20) );
  NAND2_X1 maj_119_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_119_n21) );
  NAND2_X1 maj_119_U10 ( .A1(maj_119_n21), .A2(maj_119_n20), .ZN(maj_119_n23)
         );
  XOR2_X1 maj_119_U9 ( .A(v_2_1[2]), .B(maj_119_n24), .Z(maj_119_n26) );
  XOR2_X1 maj_119_U8 ( .A(v_2_1[5]), .B(maj_119_n25), .Z(maj_119_n27) );
  XOR2_X1 maj_119_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_119_n24) );
  XOR2_X1 maj_119_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_119_n25) );
  OR2_X1 maj_119_U5 ( .A1(maj_119_n23), .A2(maj_119_n22), .ZN(maj_119_n32) );
  NAND2_X1 maj_119_U4 ( .A1(maj_119_n22), .A2(maj_119_n23), .ZN(maj_119_n34)
         );
  NAND2_X1 maj_119_U3 ( .A1(maj_119_n32), .A2(maj_119_n31), .ZN(maj_119_n33)
         );
  NAND2_X1 maj_119_U2 ( .A1(maj_119_n34), .A2(maj_119_n33), .ZN(maj_119_port_o) );
  OR2_X1 maj_120_U19 ( .A1(maj_120_n27), .A2(maj_120_n26), .ZN(maj_120_n28) );
  NAND2_X1 maj_120_U18 ( .A1(u_0_0[6]), .A2(maj_120_n28), .ZN(maj_120_n29) );
  NAND2_X1 maj_120_U17 ( .A1(maj_120_n26), .A2(maj_120_n27), .ZN(maj_120_n30)
         );
  NAND2_X1 maj_120_U16 ( .A1(maj_120_n30), .A2(maj_120_n29), .ZN(maj_120_n31)
         );
  NAND2_X1 maj_120_U15 ( .A1(u_0_0[5]), .A2(maj_120_n25), .ZN(maj_120_n18) );
  NAND2_X1 maj_120_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_120_n19) );
  NAND2_X1 maj_120_U13 ( .A1(maj_120_n19), .A2(maj_120_n18), .ZN(maj_120_n22)
         );
  NAND2_X1 maj_120_U12 ( .A1(u_0_0[2]), .A2(maj_120_n24), .ZN(maj_120_n20) );
  NAND2_X1 maj_120_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_120_n21) );
  NAND2_X1 maj_120_U10 ( .A1(maj_120_n21), .A2(maj_120_n20), .ZN(maj_120_n23)
         );
  XOR2_X1 maj_120_U9 ( .A(u_0_0[2]), .B(maj_120_n24), .Z(maj_120_n26) );
  XOR2_X1 maj_120_U8 ( .A(u_0_0[5]), .B(maj_120_n25), .Z(maj_120_n27) );
  XOR2_X1 maj_120_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_120_n24) );
  XOR2_X1 maj_120_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_120_n25) );
  OR2_X1 maj_120_U5 ( .A1(maj_120_n23), .A2(maj_120_n22), .ZN(maj_120_n32) );
  NAND2_X1 maj_120_U4 ( .A1(maj_120_n22), .A2(maj_120_n23), .ZN(maj_120_n34)
         );
  NAND2_X1 maj_120_U3 ( .A1(maj_120_n32), .A2(maj_120_n31), .ZN(maj_120_n33)
         );
  NAND2_X1 maj_120_U2 ( .A1(maj_120_n34), .A2(maj_120_n33), .ZN(maj_120_port_o) );
  OR2_X1 maj_121_U19 ( .A1(maj_121_n27), .A2(maj_121_n26), .ZN(maj_121_n28) );
  NAND2_X1 maj_121_U18 ( .A1(v_0_0[6]), .A2(maj_121_n28), .ZN(maj_121_n29) );
  NAND2_X1 maj_121_U17 ( .A1(maj_121_n26), .A2(maj_121_n27), .ZN(maj_121_n30)
         );
  NAND2_X1 maj_121_U16 ( .A1(maj_121_n30), .A2(maj_121_n29), .ZN(maj_121_n31)
         );
  NAND2_X1 maj_121_U15 ( .A1(v_0_0[5]), .A2(maj_121_n25), .ZN(maj_121_n18) );
  NAND2_X1 maj_121_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_121_n19) );
  NAND2_X1 maj_121_U13 ( .A1(maj_121_n19), .A2(maj_121_n18), .ZN(maj_121_n22)
         );
  NAND2_X1 maj_121_U12 ( .A1(v_0_0[2]), .A2(maj_121_n24), .ZN(maj_121_n20) );
  NAND2_X1 maj_121_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_121_n21) );
  NAND2_X1 maj_121_U10 ( .A1(maj_121_n21), .A2(maj_121_n20), .ZN(maj_121_n23)
         );
  XOR2_X1 maj_121_U9 ( .A(v_0_0[2]), .B(maj_121_n24), .Z(maj_121_n26) );
  XOR2_X1 maj_121_U8 ( .A(v_0_0[5]), .B(maj_121_n25), .Z(maj_121_n27) );
  XOR2_X1 maj_121_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_121_n24) );
  XOR2_X1 maj_121_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_121_n25) );
  OR2_X1 maj_121_U5 ( .A1(maj_121_n23), .A2(maj_121_n22), .ZN(maj_121_n32) );
  NAND2_X1 maj_121_U4 ( .A1(maj_121_n22), .A2(maj_121_n23), .ZN(maj_121_n34)
         );
  NAND2_X1 maj_121_U3 ( .A1(maj_121_n32), .A2(maj_121_n31), .ZN(maj_121_n33)
         );
  NAND2_X1 maj_121_U2 ( .A1(maj_121_n34), .A2(maj_121_n33), .ZN(maj_121_port_o) );
  OR2_X1 maj_122_U19 ( .A1(maj_122_n27), .A2(maj_122_n26), .ZN(maj_122_n28) );
  NAND2_X1 maj_122_U18 ( .A1(u_0_1[6]), .A2(maj_122_n28), .ZN(maj_122_n29) );
  NAND2_X1 maj_122_U17 ( .A1(maj_122_n26), .A2(maj_122_n27), .ZN(maj_122_n30)
         );
  NAND2_X1 maj_122_U16 ( .A1(maj_122_n30), .A2(maj_122_n29), .ZN(maj_122_n31)
         );
  NAND2_X1 maj_122_U15 ( .A1(u_0_1[5]), .A2(maj_122_n25), .ZN(maj_122_n18) );
  NAND2_X1 maj_122_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_122_n19) );
  NAND2_X1 maj_122_U13 ( .A1(maj_122_n19), .A2(maj_122_n18), .ZN(maj_122_n22)
         );
  NAND2_X1 maj_122_U12 ( .A1(u_0_1[2]), .A2(maj_122_n24), .ZN(maj_122_n20) );
  NAND2_X1 maj_122_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_122_n21) );
  NAND2_X1 maj_122_U10 ( .A1(maj_122_n21), .A2(maj_122_n20), .ZN(maj_122_n23)
         );
  XOR2_X1 maj_122_U9 ( .A(u_0_1[2]), .B(maj_122_n24), .Z(maj_122_n26) );
  XOR2_X1 maj_122_U8 ( .A(u_0_1[5]), .B(maj_122_n25), .Z(maj_122_n27) );
  XOR2_X1 maj_122_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_122_n24) );
  XOR2_X1 maj_122_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_122_n25) );
  OR2_X1 maj_122_U5 ( .A1(maj_122_n23), .A2(maj_122_n22), .ZN(maj_122_n32) );
  NAND2_X1 maj_122_U4 ( .A1(maj_122_n22), .A2(maj_122_n23), .ZN(maj_122_n34)
         );
  NAND2_X1 maj_122_U3 ( .A1(maj_122_n32), .A2(maj_122_n31), .ZN(maj_122_n33)
         );
  NAND2_X1 maj_122_U2 ( .A1(maj_122_n34), .A2(maj_122_n33), .ZN(maj_122_port_o) );
  OR2_X1 maj_123_U19 ( .A1(maj_123_n27), .A2(maj_123_n26), .ZN(maj_123_n28) );
  NAND2_X1 maj_123_U18 ( .A1(v_0_1[6]), .A2(maj_123_n28), .ZN(maj_123_n29) );
  NAND2_X1 maj_123_U17 ( .A1(maj_123_n26), .A2(maj_123_n27), .ZN(maj_123_n30)
         );
  NAND2_X1 maj_123_U16 ( .A1(maj_123_n30), .A2(maj_123_n29), .ZN(maj_123_n31)
         );
  NAND2_X1 maj_123_U15 ( .A1(v_0_1[5]), .A2(maj_123_n25), .ZN(maj_123_n18) );
  NAND2_X1 maj_123_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_123_n19) );
  NAND2_X1 maj_123_U13 ( .A1(maj_123_n19), .A2(maj_123_n18), .ZN(maj_123_n22)
         );
  NAND2_X1 maj_123_U12 ( .A1(v_0_1[2]), .A2(maj_123_n24), .ZN(maj_123_n20) );
  NAND2_X1 maj_123_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_123_n21) );
  NAND2_X1 maj_123_U10 ( .A1(maj_123_n21), .A2(maj_123_n20), .ZN(maj_123_n23)
         );
  XOR2_X1 maj_123_U9 ( .A(v_0_1[2]), .B(maj_123_n24), .Z(maj_123_n26) );
  XOR2_X1 maj_123_U8 ( .A(v_0_1[5]), .B(maj_123_n25), .Z(maj_123_n27) );
  XOR2_X1 maj_123_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_123_n24) );
  XOR2_X1 maj_123_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_123_n25) );
  OR2_X1 maj_123_U5 ( .A1(maj_123_n23), .A2(maj_123_n22), .ZN(maj_123_n32) );
  NAND2_X1 maj_123_U4 ( .A1(maj_123_n22), .A2(maj_123_n23), .ZN(maj_123_n34)
         );
  NAND2_X1 maj_123_U3 ( .A1(maj_123_n32), .A2(maj_123_n31), .ZN(maj_123_n33)
         );
  NAND2_X1 maj_123_U2 ( .A1(maj_123_n34), .A2(maj_123_n33), .ZN(maj_123_port_o) );
  OR2_X1 maj_124_U19 ( .A1(maj_124_n27), .A2(maj_124_n26), .ZN(maj_124_n28) );
  NAND2_X1 maj_124_U18 ( .A1(u_1_0[6]), .A2(maj_124_n28), .ZN(maj_124_n29) );
  NAND2_X1 maj_124_U17 ( .A1(maj_124_n26), .A2(maj_124_n27), .ZN(maj_124_n30)
         );
  NAND2_X1 maj_124_U16 ( .A1(maj_124_n30), .A2(maj_124_n29), .ZN(maj_124_n31)
         );
  NAND2_X1 maj_124_U15 ( .A1(u_1_0[5]), .A2(maj_124_n25), .ZN(maj_124_n18) );
  NAND2_X1 maj_124_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_124_n19) );
  NAND2_X1 maj_124_U13 ( .A1(maj_124_n19), .A2(maj_124_n18), .ZN(maj_124_n22)
         );
  NAND2_X1 maj_124_U12 ( .A1(u_1_0[2]), .A2(maj_124_n24), .ZN(maj_124_n20) );
  NAND2_X1 maj_124_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_124_n21) );
  NAND2_X1 maj_124_U10 ( .A1(maj_124_n21), .A2(maj_124_n20), .ZN(maj_124_n23)
         );
  XOR2_X1 maj_124_U9 ( .A(u_1_0[2]), .B(maj_124_n24), .Z(maj_124_n26) );
  XOR2_X1 maj_124_U8 ( .A(u_1_0[5]), .B(maj_124_n25), .Z(maj_124_n27) );
  XOR2_X1 maj_124_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_124_n24) );
  XOR2_X1 maj_124_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_124_n25) );
  OR2_X1 maj_124_U5 ( .A1(maj_124_n23), .A2(maj_124_n22), .ZN(maj_124_n32) );
  NAND2_X1 maj_124_U4 ( .A1(maj_124_n22), .A2(maj_124_n23), .ZN(maj_124_n34)
         );
  NAND2_X1 maj_124_U3 ( .A1(maj_124_n32), .A2(maj_124_n31), .ZN(maj_124_n33)
         );
  NAND2_X1 maj_124_U2 ( .A1(maj_124_n34), .A2(maj_124_n33), .ZN(maj_124_port_o) );
  OR2_X1 maj_125_U19 ( .A1(maj_125_n27), .A2(maj_125_n26), .ZN(maj_125_n28) );
  NAND2_X1 maj_125_U18 ( .A1(v_1_0[6]), .A2(maj_125_n28), .ZN(maj_125_n29) );
  NAND2_X1 maj_125_U17 ( .A1(maj_125_n26), .A2(maj_125_n27), .ZN(maj_125_n30)
         );
  NAND2_X1 maj_125_U16 ( .A1(maj_125_n30), .A2(maj_125_n29), .ZN(maj_125_n31)
         );
  NAND2_X1 maj_125_U15 ( .A1(v_1_0[5]), .A2(maj_125_n25), .ZN(maj_125_n18) );
  NAND2_X1 maj_125_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_125_n19) );
  NAND2_X1 maj_125_U13 ( .A1(maj_125_n19), .A2(maj_125_n18), .ZN(maj_125_n22)
         );
  NAND2_X1 maj_125_U12 ( .A1(v_1_0[2]), .A2(maj_125_n24), .ZN(maj_125_n20) );
  NAND2_X1 maj_125_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_125_n21) );
  NAND2_X1 maj_125_U10 ( .A1(maj_125_n21), .A2(maj_125_n20), .ZN(maj_125_n23)
         );
  XOR2_X1 maj_125_U9 ( .A(v_1_0[2]), .B(maj_125_n24), .Z(maj_125_n26) );
  XOR2_X1 maj_125_U8 ( .A(v_1_0[5]), .B(maj_125_n25), .Z(maj_125_n27) );
  XOR2_X1 maj_125_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_125_n24) );
  XOR2_X1 maj_125_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_125_n25) );
  OR2_X1 maj_125_U5 ( .A1(maj_125_n23), .A2(maj_125_n22), .ZN(maj_125_n32) );
  NAND2_X1 maj_125_U4 ( .A1(maj_125_n22), .A2(maj_125_n23), .ZN(maj_125_n34)
         );
  NAND2_X1 maj_125_U3 ( .A1(maj_125_n32), .A2(maj_125_n31), .ZN(maj_125_n33)
         );
  NAND2_X1 maj_125_U2 ( .A1(maj_125_n34), .A2(maj_125_n33), .ZN(maj_125_port_o) );
  OR2_X1 maj_126_U19 ( .A1(maj_126_n27), .A2(maj_126_n26), .ZN(maj_126_n28) );
  NAND2_X1 maj_126_U18 ( .A1(u_1_1[6]), .A2(maj_126_n28), .ZN(maj_126_n29) );
  NAND2_X1 maj_126_U17 ( .A1(maj_126_n26), .A2(maj_126_n27), .ZN(maj_126_n30)
         );
  NAND2_X1 maj_126_U16 ( .A1(maj_126_n30), .A2(maj_126_n29), .ZN(maj_126_n31)
         );
  NAND2_X1 maj_126_U15 ( .A1(u_1_1[5]), .A2(maj_126_n25), .ZN(maj_126_n18) );
  NAND2_X1 maj_126_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_126_n19) );
  NAND2_X1 maj_126_U13 ( .A1(maj_126_n19), .A2(maj_126_n18), .ZN(maj_126_n22)
         );
  NAND2_X1 maj_126_U12 ( .A1(u_1_1[2]), .A2(maj_126_n24), .ZN(maj_126_n20) );
  NAND2_X1 maj_126_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_126_n21) );
  NAND2_X1 maj_126_U10 ( .A1(maj_126_n21), .A2(maj_126_n20), .ZN(maj_126_n23)
         );
  XOR2_X1 maj_126_U9 ( .A(u_1_1[2]), .B(maj_126_n24), .Z(maj_126_n26) );
  XOR2_X1 maj_126_U8 ( .A(u_1_1[5]), .B(maj_126_n25), .Z(maj_126_n27) );
  XOR2_X1 maj_126_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_126_n24) );
  XOR2_X1 maj_126_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_126_n25) );
  OR2_X1 maj_126_U5 ( .A1(maj_126_n23), .A2(maj_126_n22), .ZN(maj_126_n32) );
  NAND2_X1 maj_126_U4 ( .A1(maj_126_n22), .A2(maj_126_n23), .ZN(maj_126_n34)
         );
  NAND2_X1 maj_126_U3 ( .A1(maj_126_n32), .A2(maj_126_n31), .ZN(maj_126_n33)
         );
  NAND2_X1 maj_126_U2 ( .A1(maj_126_n34), .A2(maj_126_n33), .ZN(maj_126_port_o) );
  OR2_X1 maj_127_U19 ( .A1(maj_127_n27), .A2(maj_127_n26), .ZN(maj_127_n28) );
  NAND2_X1 maj_127_U18 ( .A1(v_1_1[6]), .A2(maj_127_n28), .ZN(maj_127_n29) );
  NAND2_X1 maj_127_U17 ( .A1(maj_127_n26), .A2(maj_127_n27), .ZN(maj_127_n30)
         );
  NAND2_X1 maj_127_U16 ( .A1(maj_127_n30), .A2(maj_127_n29), .ZN(maj_127_n31)
         );
  NAND2_X1 maj_127_U15 ( .A1(v_1_1[5]), .A2(maj_127_n25), .ZN(maj_127_n18) );
  NAND2_X1 maj_127_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_127_n19) );
  NAND2_X1 maj_127_U13 ( .A1(maj_127_n19), .A2(maj_127_n18), .ZN(maj_127_n22)
         );
  NAND2_X1 maj_127_U12 ( .A1(v_1_1[2]), .A2(maj_127_n24), .ZN(maj_127_n20) );
  NAND2_X1 maj_127_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_127_n21) );
  NAND2_X1 maj_127_U10 ( .A1(maj_127_n21), .A2(maj_127_n20), .ZN(maj_127_n23)
         );
  XOR2_X1 maj_127_U9 ( .A(v_1_1[2]), .B(maj_127_n24), .Z(maj_127_n26) );
  XOR2_X1 maj_127_U8 ( .A(v_1_1[5]), .B(maj_127_n25), .Z(maj_127_n27) );
  XOR2_X1 maj_127_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_127_n24) );
  XOR2_X1 maj_127_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_127_n25) );
  OR2_X1 maj_127_U5 ( .A1(maj_127_n23), .A2(maj_127_n22), .ZN(maj_127_n32) );
  NAND2_X1 maj_127_U4 ( .A1(maj_127_n22), .A2(maj_127_n23), .ZN(maj_127_n34)
         );
  NAND2_X1 maj_127_U3 ( .A1(maj_127_n32), .A2(maj_127_n31), .ZN(maj_127_n33)
         );
  NAND2_X1 maj_127_U2 ( .A1(maj_127_n34), .A2(maj_127_n33), .ZN(maj_127_port_o) );
  OR2_X1 maj_128_U19 ( .A1(maj_128_n27), .A2(maj_128_n26), .ZN(maj_128_n28) );
  NAND2_X1 maj_128_U18 ( .A1(u_2_0[6]), .A2(maj_128_n28), .ZN(maj_128_n29) );
  NAND2_X1 maj_128_U17 ( .A1(maj_128_n26), .A2(maj_128_n27), .ZN(maj_128_n30)
         );
  NAND2_X1 maj_128_U16 ( .A1(maj_128_n30), .A2(maj_128_n29), .ZN(maj_128_n31)
         );
  NAND2_X1 maj_128_U15 ( .A1(u_2_0[5]), .A2(maj_128_n25), .ZN(maj_128_n18) );
  NAND2_X1 maj_128_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_128_n19) );
  NAND2_X1 maj_128_U13 ( .A1(maj_128_n19), .A2(maj_128_n18), .ZN(maj_128_n22)
         );
  NAND2_X1 maj_128_U12 ( .A1(u_2_0[2]), .A2(maj_128_n24), .ZN(maj_128_n20) );
  NAND2_X1 maj_128_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_128_n21) );
  NAND2_X1 maj_128_U10 ( .A1(maj_128_n21), .A2(maj_128_n20), .ZN(maj_128_n23)
         );
  XOR2_X1 maj_128_U9 ( .A(u_2_0[2]), .B(maj_128_n24), .Z(maj_128_n26) );
  XOR2_X1 maj_128_U8 ( .A(u_2_0[5]), .B(maj_128_n25), .Z(maj_128_n27) );
  XOR2_X1 maj_128_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_128_n24) );
  XOR2_X1 maj_128_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_128_n25) );
  OR2_X1 maj_128_U5 ( .A1(maj_128_n23), .A2(maj_128_n22), .ZN(maj_128_n32) );
  NAND2_X1 maj_128_U4 ( .A1(maj_128_n22), .A2(maj_128_n23), .ZN(maj_128_n34)
         );
  NAND2_X1 maj_128_U3 ( .A1(maj_128_n32), .A2(maj_128_n31), .ZN(maj_128_n33)
         );
  NAND2_X1 maj_128_U2 ( .A1(maj_128_n34), .A2(maj_128_n33), .ZN(maj_128_port_o) );
  OR2_X1 maj_129_U19 ( .A1(maj_129_n27), .A2(maj_129_n26), .ZN(maj_129_n28) );
  NAND2_X1 maj_129_U18 ( .A1(v_2_0[6]), .A2(maj_129_n28), .ZN(maj_129_n29) );
  NAND2_X1 maj_129_U17 ( .A1(maj_129_n26), .A2(maj_129_n27), .ZN(maj_129_n30)
         );
  NAND2_X1 maj_129_U16 ( .A1(maj_129_n30), .A2(maj_129_n29), .ZN(maj_129_n31)
         );
  NAND2_X1 maj_129_U15 ( .A1(v_2_0[5]), .A2(maj_129_n25), .ZN(maj_129_n18) );
  NAND2_X1 maj_129_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_129_n19) );
  NAND2_X1 maj_129_U13 ( .A1(maj_129_n19), .A2(maj_129_n18), .ZN(maj_129_n22)
         );
  NAND2_X1 maj_129_U12 ( .A1(v_2_0[2]), .A2(maj_129_n24), .ZN(maj_129_n20) );
  NAND2_X1 maj_129_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_129_n21) );
  NAND2_X1 maj_129_U10 ( .A1(maj_129_n21), .A2(maj_129_n20), .ZN(maj_129_n23)
         );
  XOR2_X1 maj_129_U9 ( .A(v_2_0[2]), .B(maj_129_n24), .Z(maj_129_n26) );
  XOR2_X1 maj_129_U8 ( .A(v_2_0[5]), .B(maj_129_n25), .Z(maj_129_n27) );
  XOR2_X1 maj_129_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_129_n24) );
  XOR2_X1 maj_129_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_129_n25) );
  OR2_X1 maj_129_U5 ( .A1(maj_129_n23), .A2(maj_129_n22), .ZN(maj_129_n32) );
  NAND2_X1 maj_129_U4 ( .A1(maj_129_n22), .A2(maj_129_n23), .ZN(maj_129_n34)
         );
  NAND2_X1 maj_129_U3 ( .A1(maj_129_n32), .A2(maj_129_n31), .ZN(maj_129_n33)
         );
  NAND2_X1 maj_129_U2 ( .A1(maj_129_n34), .A2(maj_129_n33), .ZN(maj_129_port_o) );
  OR2_X1 maj_130_U19 ( .A1(maj_130_n27), .A2(maj_130_n26), .ZN(maj_130_n28) );
  NAND2_X1 maj_130_U18 ( .A1(u_2_1[6]), .A2(maj_130_n28), .ZN(maj_130_n29) );
  NAND2_X1 maj_130_U17 ( .A1(maj_130_n26), .A2(maj_130_n27), .ZN(maj_130_n30)
         );
  NAND2_X1 maj_130_U16 ( .A1(maj_130_n30), .A2(maj_130_n29), .ZN(maj_130_n31)
         );
  NAND2_X1 maj_130_U15 ( .A1(u_2_1[5]), .A2(maj_130_n25), .ZN(maj_130_n18) );
  NAND2_X1 maj_130_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_130_n19) );
  NAND2_X1 maj_130_U13 ( .A1(maj_130_n19), .A2(maj_130_n18), .ZN(maj_130_n22)
         );
  NAND2_X1 maj_130_U12 ( .A1(u_2_1[2]), .A2(maj_130_n24), .ZN(maj_130_n20) );
  NAND2_X1 maj_130_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_130_n21) );
  NAND2_X1 maj_130_U10 ( .A1(maj_130_n21), .A2(maj_130_n20), .ZN(maj_130_n23)
         );
  XOR2_X1 maj_130_U9 ( .A(u_2_1[2]), .B(maj_130_n24), .Z(maj_130_n26) );
  XOR2_X1 maj_130_U8 ( .A(u_2_1[5]), .B(maj_130_n25), .Z(maj_130_n27) );
  XOR2_X1 maj_130_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_130_n24) );
  XOR2_X1 maj_130_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_130_n25) );
  OR2_X1 maj_130_U5 ( .A1(maj_130_n23), .A2(maj_130_n22), .ZN(maj_130_n32) );
  NAND2_X1 maj_130_U4 ( .A1(maj_130_n22), .A2(maj_130_n23), .ZN(maj_130_n34)
         );
  NAND2_X1 maj_130_U3 ( .A1(maj_130_n32), .A2(maj_130_n31), .ZN(maj_130_n33)
         );
  NAND2_X1 maj_130_U2 ( .A1(maj_130_n34), .A2(maj_130_n33), .ZN(maj_130_port_o) );
  OR2_X1 maj_131_U19 ( .A1(maj_131_n27), .A2(maj_131_n26), .ZN(maj_131_n28) );
  NAND2_X1 maj_131_U18 ( .A1(v_2_1[6]), .A2(maj_131_n28), .ZN(maj_131_n29) );
  NAND2_X1 maj_131_U17 ( .A1(maj_131_n26), .A2(maj_131_n27), .ZN(maj_131_n30)
         );
  NAND2_X1 maj_131_U16 ( .A1(maj_131_n30), .A2(maj_131_n29), .ZN(maj_131_n31)
         );
  NAND2_X1 maj_131_U15 ( .A1(v_2_1[5]), .A2(maj_131_n25), .ZN(maj_131_n18) );
  NAND2_X1 maj_131_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_131_n19) );
  NAND2_X1 maj_131_U13 ( .A1(maj_131_n19), .A2(maj_131_n18), .ZN(maj_131_n22)
         );
  NAND2_X1 maj_131_U12 ( .A1(v_2_1[2]), .A2(maj_131_n24), .ZN(maj_131_n20) );
  NAND2_X1 maj_131_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_131_n21) );
  NAND2_X1 maj_131_U10 ( .A1(maj_131_n21), .A2(maj_131_n20), .ZN(maj_131_n23)
         );
  XOR2_X1 maj_131_U9 ( .A(v_2_1[2]), .B(maj_131_n24), .Z(maj_131_n26) );
  XOR2_X1 maj_131_U8 ( .A(v_2_1[5]), .B(maj_131_n25), .Z(maj_131_n27) );
  XOR2_X1 maj_131_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_131_n24) );
  XOR2_X1 maj_131_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_131_n25) );
  OR2_X1 maj_131_U5 ( .A1(maj_131_n23), .A2(maj_131_n22), .ZN(maj_131_n32) );
  NAND2_X1 maj_131_U4 ( .A1(maj_131_n22), .A2(maj_131_n23), .ZN(maj_131_n34)
         );
  NAND2_X1 maj_131_U3 ( .A1(maj_131_n32), .A2(maj_131_n31), .ZN(maj_131_n33)
         );
  NAND2_X1 maj_131_U2 ( .A1(maj_131_n34), .A2(maj_131_n33), .ZN(maj_131_port_o) );
  OR2_X1 maj_132_U19 ( .A1(maj_132_n27), .A2(maj_132_n26), .ZN(maj_132_n28) );
  NAND2_X1 maj_132_U18 ( .A1(u_0_0[6]), .A2(maj_132_n28), .ZN(maj_132_n29) );
  NAND2_X1 maj_132_U17 ( .A1(maj_132_n26), .A2(maj_132_n27), .ZN(maj_132_n30)
         );
  NAND2_X1 maj_132_U16 ( .A1(maj_132_n30), .A2(maj_132_n29), .ZN(maj_132_n31)
         );
  NAND2_X1 maj_132_U15 ( .A1(u_0_0[5]), .A2(maj_132_n25), .ZN(maj_132_n18) );
  NAND2_X1 maj_132_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_132_n19) );
  NAND2_X1 maj_132_U13 ( .A1(maj_132_n19), .A2(maj_132_n18), .ZN(maj_132_n22)
         );
  NAND2_X1 maj_132_U12 ( .A1(u_0_0[2]), .A2(maj_132_n24), .ZN(maj_132_n20) );
  NAND2_X1 maj_132_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_132_n21) );
  NAND2_X1 maj_132_U10 ( .A1(maj_132_n21), .A2(maj_132_n20), .ZN(maj_132_n23)
         );
  XOR2_X1 maj_132_U9 ( .A(u_0_0[2]), .B(maj_132_n24), .Z(maj_132_n26) );
  XOR2_X1 maj_132_U8 ( .A(u_0_0[5]), .B(maj_132_n25), .Z(maj_132_n27) );
  XOR2_X1 maj_132_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_132_n24) );
  XOR2_X1 maj_132_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_132_n25) );
  OR2_X1 maj_132_U5 ( .A1(maj_132_n23), .A2(maj_132_n22), .ZN(maj_132_n32) );
  NAND2_X1 maj_132_U4 ( .A1(maj_132_n22), .A2(maj_132_n23), .ZN(maj_132_n34)
         );
  NAND2_X1 maj_132_U3 ( .A1(maj_132_n32), .A2(maj_132_n31), .ZN(maj_132_n33)
         );
  NAND2_X1 maj_132_U2 ( .A1(maj_132_n34), .A2(maj_132_n33), .ZN(maj_132_port_o) );
  OR2_X1 maj_133_U19 ( .A1(maj_133_n27), .A2(maj_133_n26), .ZN(maj_133_n28) );
  NAND2_X1 maj_133_U18 ( .A1(v_0_0[6]), .A2(maj_133_n28), .ZN(maj_133_n29) );
  NAND2_X1 maj_133_U17 ( .A1(maj_133_n26), .A2(maj_133_n27), .ZN(maj_133_n30)
         );
  NAND2_X1 maj_133_U16 ( .A1(maj_133_n30), .A2(maj_133_n29), .ZN(maj_133_n31)
         );
  NAND2_X1 maj_133_U15 ( .A1(v_0_0[5]), .A2(maj_133_n25), .ZN(maj_133_n18) );
  NAND2_X1 maj_133_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_133_n19) );
  NAND2_X1 maj_133_U13 ( .A1(maj_133_n19), .A2(maj_133_n18), .ZN(maj_133_n22)
         );
  NAND2_X1 maj_133_U12 ( .A1(v_0_0[2]), .A2(maj_133_n24), .ZN(maj_133_n20) );
  NAND2_X1 maj_133_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_133_n21) );
  NAND2_X1 maj_133_U10 ( .A1(maj_133_n21), .A2(maj_133_n20), .ZN(maj_133_n23)
         );
  XOR2_X1 maj_133_U9 ( .A(v_0_0[2]), .B(maj_133_n24), .Z(maj_133_n26) );
  XOR2_X1 maj_133_U8 ( .A(v_0_0[5]), .B(maj_133_n25), .Z(maj_133_n27) );
  XOR2_X1 maj_133_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_133_n24) );
  XOR2_X1 maj_133_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_133_n25) );
  OR2_X1 maj_133_U5 ( .A1(maj_133_n23), .A2(maj_133_n22), .ZN(maj_133_n32) );
  NAND2_X1 maj_133_U4 ( .A1(maj_133_n22), .A2(maj_133_n23), .ZN(maj_133_n34)
         );
  NAND2_X1 maj_133_U3 ( .A1(maj_133_n32), .A2(maj_133_n31), .ZN(maj_133_n33)
         );
  NAND2_X1 maj_133_U2 ( .A1(maj_133_n34), .A2(maj_133_n33), .ZN(maj_133_port_o) );
  OR2_X1 maj_134_U19 ( .A1(maj_134_n27), .A2(maj_134_n26), .ZN(maj_134_n28) );
  NAND2_X1 maj_134_U18 ( .A1(u_0_1[6]), .A2(maj_134_n28), .ZN(maj_134_n29) );
  NAND2_X1 maj_134_U17 ( .A1(maj_134_n26), .A2(maj_134_n27), .ZN(maj_134_n30)
         );
  NAND2_X1 maj_134_U16 ( .A1(maj_134_n30), .A2(maj_134_n29), .ZN(maj_134_n31)
         );
  NAND2_X1 maj_134_U15 ( .A1(u_0_1[5]), .A2(maj_134_n25), .ZN(maj_134_n18) );
  NAND2_X1 maj_134_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_134_n19) );
  NAND2_X1 maj_134_U13 ( .A1(maj_134_n19), .A2(maj_134_n18), .ZN(maj_134_n22)
         );
  NAND2_X1 maj_134_U12 ( .A1(u_0_1[2]), .A2(maj_134_n24), .ZN(maj_134_n20) );
  NAND2_X1 maj_134_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_134_n21) );
  NAND2_X1 maj_134_U10 ( .A1(maj_134_n21), .A2(maj_134_n20), .ZN(maj_134_n23)
         );
  XOR2_X1 maj_134_U9 ( .A(u_0_1[2]), .B(maj_134_n24), .Z(maj_134_n26) );
  XOR2_X1 maj_134_U8 ( .A(u_0_1[5]), .B(maj_134_n25), .Z(maj_134_n27) );
  XOR2_X1 maj_134_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_134_n24) );
  XOR2_X1 maj_134_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_134_n25) );
  OR2_X1 maj_134_U5 ( .A1(maj_134_n23), .A2(maj_134_n22), .ZN(maj_134_n32) );
  NAND2_X1 maj_134_U4 ( .A1(maj_134_n22), .A2(maj_134_n23), .ZN(maj_134_n34)
         );
  NAND2_X1 maj_134_U3 ( .A1(maj_134_n32), .A2(maj_134_n31), .ZN(maj_134_n33)
         );
  NAND2_X1 maj_134_U2 ( .A1(maj_134_n34), .A2(maj_134_n33), .ZN(maj_134_port_o) );
  OR2_X1 maj_135_U19 ( .A1(maj_135_n27), .A2(maj_135_n26), .ZN(maj_135_n28) );
  NAND2_X1 maj_135_U18 ( .A1(v_0_1[6]), .A2(maj_135_n28), .ZN(maj_135_n29) );
  NAND2_X1 maj_135_U17 ( .A1(maj_135_n26), .A2(maj_135_n27), .ZN(maj_135_n30)
         );
  NAND2_X1 maj_135_U16 ( .A1(maj_135_n30), .A2(maj_135_n29), .ZN(maj_135_n31)
         );
  NAND2_X1 maj_135_U15 ( .A1(v_0_1[5]), .A2(maj_135_n25), .ZN(maj_135_n18) );
  NAND2_X1 maj_135_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_135_n19) );
  NAND2_X1 maj_135_U13 ( .A1(maj_135_n19), .A2(maj_135_n18), .ZN(maj_135_n22)
         );
  NAND2_X1 maj_135_U12 ( .A1(v_0_1[2]), .A2(maj_135_n24), .ZN(maj_135_n20) );
  NAND2_X1 maj_135_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_135_n21) );
  NAND2_X1 maj_135_U10 ( .A1(maj_135_n21), .A2(maj_135_n20), .ZN(maj_135_n23)
         );
  XOR2_X1 maj_135_U9 ( .A(v_0_1[2]), .B(maj_135_n24), .Z(maj_135_n26) );
  XOR2_X1 maj_135_U8 ( .A(v_0_1[5]), .B(maj_135_n25), .Z(maj_135_n27) );
  XOR2_X1 maj_135_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_135_n24) );
  XOR2_X1 maj_135_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_135_n25) );
  OR2_X1 maj_135_U5 ( .A1(maj_135_n23), .A2(maj_135_n22), .ZN(maj_135_n32) );
  NAND2_X1 maj_135_U4 ( .A1(maj_135_n22), .A2(maj_135_n23), .ZN(maj_135_n34)
         );
  NAND2_X1 maj_135_U3 ( .A1(maj_135_n32), .A2(maj_135_n31), .ZN(maj_135_n33)
         );
  NAND2_X1 maj_135_U2 ( .A1(maj_135_n34), .A2(maj_135_n33), .ZN(maj_135_port_o) );
  OR2_X1 maj_136_U19 ( .A1(maj_136_n27), .A2(maj_136_n26), .ZN(maj_136_n28) );
  NAND2_X1 maj_136_U18 ( .A1(u_1_0[6]), .A2(maj_136_n28), .ZN(maj_136_n29) );
  NAND2_X1 maj_136_U17 ( .A1(maj_136_n26), .A2(maj_136_n27), .ZN(maj_136_n30)
         );
  NAND2_X1 maj_136_U16 ( .A1(maj_136_n30), .A2(maj_136_n29), .ZN(maj_136_n31)
         );
  NAND2_X1 maj_136_U15 ( .A1(u_1_0[5]), .A2(maj_136_n25), .ZN(maj_136_n18) );
  NAND2_X1 maj_136_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_136_n19) );
  NAND2_X1 maj_136_U13 ( .A1(maj_136_n19), .A2(maj_136_n18), .ZN(maj_136_n22)
         );
  NAND2_X1 maj_136_U12 ( .A1(u_1_0[2]), .A2(maj_136_n24), .ZN(maj_136_n20) );
  NAND2_X1 maj_136_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_136_n21) );
  NAND2_X1 maj_136_U10 ( .A1(maj_136_n21), .A2(maj_136_n20), .ZN(maj_136_n23)
         );
  XOR2_X1 maj_136_U9 ( .A(u_1_0[2]), .B(maj_136_n24), .Z(maj_136_n26) );
  XOR2_X1 maj_136_U8 ( .A(u_1_0[5]), .B(maj_136_n25), .Z(maj_136_n27) );
  XOR2_X1 maj_136_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_136_n24) );
  XOR2_X1 maj_136_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_136_n25) );
  OR2_X1 maj_136_U5 ( .A1(maj_136_n23), .A2(maj_136_n22), .ZN(maj_136_n32) );
  NAND2_X1 maj_136_U4 ( .A1(maj_136_n22), .A2(maj_136_n23), .ZN(maj_136_n34)
         );
  NAND2_X1 maj_136_U3 ( .A1(maj_136_n32), .A2(maj_136_n31), .ZN(maj_136_n33)
         );
  NAND2_X1 maj_136_U2 ( .A1(maj_136_n34), .A2(maj_136_n33), .ZN(maj_136_port_o) );
  OR2_X1 maj_137_U19 ( .A1(maj_137_n27), .A2(maj_137_n26), .ZN(maj_137_n28) );
  NAND2_X1 maj_137_U18 ( .A1(v_1_0[6]), .A2(maj_137_n28), .ZN(maj_137_n29) );
  NAND2_X1 maj_137_U17 ( .A1(maj_137_n26), .A2(maj_137_n27), .ZN(maj_137_n30)
         );
  NAND2_X1 maj_137_U16 ( .A1(maj_137_n30), .A2(maj_137_n29), .ZN(maj_137_n31)
         );
  NAND2_X1 maj_137_U15 ( .A1(v_1_0[5]), .A2(maj_137_n25), .ZN(maj_137_n18) );
  NAND2_X1 maj_137_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_137_n19) );
  NAND2_X1 maj_137_U13 ( .A1(maj_137_n19), .A2(maj_137_n18), .ZN(maj_137_n22)
         );
  NAND2_X1 maj_137_U12 ( .A1(v_1_0[2]), .A2(maj_137_n24), .ZN(maj_137_n20) );
  NAND2_X1 maj_137_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_137_n21) );
  NAND2_X1 maj_137_U10 ( .A1(maj_137_n21), .A2(maj_137_n20), .ZN(maj_137_n23)
         );
  XOR2_X1 maj_137_U9 ( .A(v_1_0[2]), .B(maj_137_n24), .Z(maj_137_n26) );
  XOR2_X1 maj_137_U8 ( .A(v_1_0[5]), .B(maj_137_n25), .Z(maj_137_n27) );
  XOR2_X1 maj_137_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_137_n24) );
  XOR2_X1 maj_137_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_137_n25) );
  OR2_X1 maj_137_U5 ( .A1(maj_137_n23), .A2(maj_137_n22), .ZN(maj_137_n32) );
  NAND2_X1 maj_137_U4 ( .A1(maj_137_n22), .A2(maj_137_n23), .ZN(maj_137_n34)
         );
  NAND2_X1 maj_137_U3 ( .A1(maj_137_n32), .A2(maj_137_n31), .ZN(maj_137_n33)
         );
  NAND2_X1 maj_137_U2 ( .A1(maj_137_n34), .A2(maj_137_n33), .ZN(maj_137_port_o) );
  OR2_X1 maj_138_U19 ( .A1(maj_138_n27), .A2(maj_138_n26), .ZN(maj_138_n28) );
  NAND2_X1 maj_138_U18 ( .A1(u_1_1[6]), .A2(maj_138_n28), .ZN(maj_138_n29) );
  NAND2_X1 maj_138_U17 ( .A1(maj_138_n26), .A2(maj_138_n27), .ZN(maj_138_n30)
         );
  NAND2_X1 maj_138_U16 ( .A1(maj_138_n30), .A2(maj_138_n29), .ZN(maj_138_n31)
         );
  NAND2_X1 maj_138_U15 ( .A1(u_1_1[5]), .A2(maj_138_n25), .ZN(maj_138_n18) );
  NAND2_X1 maj_138_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_138_n19) );
  NAND2_X1 maj_138_U13 ( .A1(maj_138_n19), .A2(maj_138_n18), .ZN(maj_138_n22)
         );
  NAND2_X1 maj_138_U12 ( .A1(u_1_1[2]), .A2(maj_138_n24), .ZN(maj_138_n20) );
  NAND2_X1 maj_138_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_138_n21) );
  NAND2_X1 maj_138_U10 ( .A1(maj_138_n21), .A2(maj_138_n20), .ZN(maj_138_n23)
         );
  XOR2_X1 maj_138_U9 ( .A(u_1_1[2]), .B(maj_138_n24), .Z(maj_138_n26) );
  XOR2_X1 maj_138_U8 ( .A(u_1_1[5]), .B(maj_138_n25), .Z(maj_138_n27) );
  XOR2_X1 maj_138_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_138_n24) );
  XOR2_X1 maj_138_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_138_n25) );
  OR2_X1 maj_138_U5 ( .A1(maj_138_n23), .A2(maj_138_n22), .ZN(maj_138_n32) );
  NAND2_X1 maj_138_U4 ( .A1(maj_138_n22), .A2(maj_138_n23), .ZN(maj_138_n34)
         );
  NAND2_X1 maj_138_U3 ( .A1(maj_138_n32), .A2(maj_138_n31), .ZN(maj_138_n33)
         );
  NAND2_X1 maj_138_U2 ( .A1(maj_138_n34), .A2(maj_138_n33), .ZN(maj_138_port_o) );
  OR2_X1 maj_139_U19 ( .A1(maj_139_n27), .A2(maj_139_n26), .ZN(maj_139_n28) );
  NAND2_X1 maj_139_U18 ( .A1(v_1_1[6]), .A2(maj_139_n28), .ZN(maj_139_n29) );
  NAND2_X1 maj_139_U17 ( .A1(maj_139_n26), .A2(maj_139_n27), .ZN(maj_139_n30)
         );
  NAND2_X1 maj_139_U16 ( .A1(maj_139_n30), .A2(maj_139_n29), .ZN(maj_139_n31)
         );
  NAND2_X1 maj_139_U15 ( .A1(v_1_1[5]), .A2(maj_139_n25), .ZN(maj_139_n18) );
  NAND2_X1 maj_139_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_139_n19) );
  NAND2_X1 maj_139_U13 ( .A1(maj_139_n19), .A2(maj_139_n18), .ZN(maj_139_n22)
         );
  NAND2_X1 maj_139_U12 ( .A1(v_1_1[2]), .A2(maj_139_n24), .ZN(maj_139_n20) );
  NAND2_X1 maj_139_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_139_n21) );
  NAND2_X1 maj_139_U10 ( .A1(maj_139_n21), .A2(maj_139_n20), .ZN(maj_139_n23)
         );
  XOR2_X1 maj_139_U9 ( .A(v_1_1[2]), .B(maj_139_n24), .Z(maj_139_n26) );
  XOR2_X1 maj_139_U8 ( .A(v_1_1[5]), .B(maj_139_n25), .Z(maj_139_n27) );
  XOR2_X1 maj_139_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_139_n24) );
  XOR2_X1 maj_139_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_139_n25) );
  OR2_X1 maj_139_U5 ( .A1(maj_139_n23), .A2(maj_139_n22), .ZN(maj_139_n32) );
  NAND2_X1 maj_139_U4 ( .A1(maj_139_n22), .A2(maj_139_n23), .ZN(maj_139_n34)
         );
  NAND2_X1 maj_139_U3 ( .A1(maj_139_n32), .A2(maj_139_n31), .ZN(maj_139_n33)
         );
  NAND2_X1 maj_139_U2 ( .A1(maj_139_n34), .A2(maj_139_n33), .ZN(maj_139_port_o) );
  OR2_X1 maj_140_U19 ( .A1(maj_140_n27), .A2(maj_140_n26), .ZN(maj_140_n28) );
  NAND2_X1 maj_140_U18 ( .A1(u_2_0[6]), .A2(maj_140_n28), .ZN(maj_140_n29) );
  NAND2_X1 maj_140_U17 ( .A1(maj_140_n26), .A2(maj_140_n27), .ZN(maj_140_n30)
         );
  NAND2_X1 maj_140_U16 ( .A1(maj_140_n30), .A2(maj_140_n29), .ZN(maj_140_n31)
         );
  NAND2_X1 maj_140_U15 ( .A1(u_2_0[5]), .A2(maj_140_n25), .ZN(maj_140_n18) );
  NAND2_X1 maj_140_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_140_n19) );
  NAND2_X1 maj_140_U13 ( .A1(maj_140_n19), .A2(maj_140_n18), .ZN(maj_140_n22)
         );
  NAND2_X1 maj_140_U12 ( .A1(u_2_0[2]), .A2(maj_140_n24), .ZN(maj_140_n20) );
  NAND2_X1 maj_140_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_140_n21) );
  NAND2_X1 maj_140_U10 ( .A1(maj_140_n21), .A2(maj_140_n20), .ZN(maj_140_n23)
         );
  XOR2_X1 maj_140_U9 ( .A(u_2_0[2]), .B(maj_140_n24), .Z(maj_140_n26) );
  XOR2_X1 maj_140_U8 ( .A(u_2_0[5]), .B(maj_140_n25), .Z(maj_140_n27) );
  XOR2_X1 maj_140_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_140_n24) );
  XOR2_X1 maj_140_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_140_n25) );
  OR2_X1 maj_140_U5 ( .A1(maj_140_n23), .A2(maj_140_n22), .ZN(maj_140_n32) );
  NAND2_X1 maj_140_U4 ( .A1(maj_140_n22), .A2(maj_140_n23), .ZN(maj_140_n34)
         );
  NAND2_X1 maj_140_U3 ( .A1(maj_140_n32), .A2(maj_140_n31), .ZN(maj_140_n33)
         );
  NAND2_X1 maj_140_U2 ( .A1(maj_140_n34), .A2(maj_140_n33), .ZN(maj_140_port_o) );
  OR2_X1 maj_141_U19 ( .A1(maj_141_n27), .A2(maj_141_n26), .ZN(maj_141_n28) );
  NAND2_X1 maj_141_U18 ( .A1(v_2_0[6]), .A2(maj_141_n28), .ZN(maj_141_n29) );
  NAND2_X1 maj_141_U17 ( .A1(maj_141_n26), .A2(maj_141_n27), .ZN(maj_141_n30)
         );
  NAND2_X1 maj_141_U16 ( .A1(maj_141_n30), .A2(maj_141_n29), .ZN(maj_141_n31)
         );
  NAND2_X1 maj_141_U15 ( .A1(v_2_0[5]), .A2(maj_141_n25), .ZN(maj_141_n18) );
  NAND2_X1 maj_141_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_141_n19) );
  NAND2_X1 maj_141_U13 ( .A1(maj_141_n19), .A2(maj_141_n18), .ZN(maj_141_n22)
         );
  NAND2_X1 maj_141_U12 ( .A1(v_2_0[2]), .A2(maj_141_n24), .ZN(maj_141_n20) );
  NAND2_X1 maj_141_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_141_n21) );
  NAND2_X1 maj_141_U10 ( .A1(maj_141_n21), .A2(maj_141_n20), .ZN(maj_141_n23)
         );
  XOR2_X1 maj_141_U9 ( .A(v_2_0[2]), .B(maj_141_n24), .Z(maj_141_n26) );
  XOR2_X1 maj_141_U8 ( .A(v_2_0[5]), .B(maj_141_n25), .Z(maj_141_n27) );
  XOR2_X1 maj_141_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_141_n24) );
  XOR2_X1 maj_141_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_141_n25) );
  OR2_X1 maj_141_U5 ( .A1(maj_141_n23), .A2(maj_141_n22), .ZN(maj_141_n32) );
  NAND2_X1 maj_141_U4 ( .A1(maj_141_n22), .A2(maj_141_n23), .ZN(maj_141_n34)
         );
  NAND2_X1 maj_141_U3 ( .A1(maj_141_n32), .A2(maj_141_n31), .ZN(maj_141_n33)
         );
  NAND2_X1 maj_141_U2 ( .A1(maj_141_n34), .A2(maj_141_n33), .ZN(maj_141_port_o) );
  OR2_X1 maj_142_U19 ( .A1(maj_142_n27), .A2(maj_142_n26), .ZN(maj_142_n28) );
  NAND2_X1 maj_142_U18 ( .A1(u_2_1[6]), .A2(maj_142_n28), .ZN(maj_142_n29) );
  NAND2_X1 maj_142_U17 ( .A1(maj_142_n26), .A2(maj_142_n27), .ZN(maj_142_n30)
         );
  NAND2_X1 maj_142_U16 ( .A1(maj_142_n30), .A2(maj_142_n29), .ZN(maj_142_n31)
         );
  NAND2_X1 maj_142_U15 ( .A1(u_2_1[5]), .A2(maj_142_n25), .ZN(maj_142_n18) );
  NAND2_X1 maj_142_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_142_n19) );
  NAND2_X1 maj_142_U13 ( .A1(maj_142_n19), .A2(maj_142_n18), .ZN(maj_142_n22)
         );
  NAND2_X1 maj_142_U12 ( .A1(u_2_1[2]), .A2(maj_142_n24), .ZN(maj_142_n20) );
  NAND2_X1 maj_142_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_142_n21) );
  NAND2_X1 maj_142_U10 ( .A1(maj_142_n21), .A2(maj_142_n20), .ZN(maj_142_n23)
         );
  XOR2_X1 maj_142_U9 ( .A(u_2_1[2]), .B(maj_142_n24), .Z(maj_142_n26) );
  XOR2_X1 maj_142_U8 ( .A(u_2_1[5]), .B(maj_142_n25), .Z(maj_142_n27) );
  XOR2_X1 maj_142_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_142_n24) );
  XOR2_X1 maj_142_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_142_n25) );
  OR2_X1 maj_142_U5 ( .A1(maj_142_n23), .A2(maj_142_n22), .ZN(maj_142_n32) );
  NAND2_X1 maj_142_U4 ( .A1(maj_142_n22), .A2(maj_142_n23), .ZN(maj_142_n34)
         );
  NAND2_X1 maj_142_U3 ( .A1(maj_142_n32), .A2(maj_142_n31), .ZN(maj_142_n33)
         );
  NAND2_X1 maj_142_U2 ( .A1(maj_142_n34), .A2(maj_142_n33), .ZN(maj_142_port_o) );
  OR2_X1 maj_143_U19 ( .A1(maj_143_n27), .A2(maj_143_n26), .ZN(maj_143_n28) );
  NAND2_X1 maj_143_U18 ( .A1(v_2_1[6]), .A2(maj_143_n28), .ZN(maj_143_n29) );
  NAND2_X1 maj_143_U17 ( .A1(maj_143_n26), .A2(maj_143_n27), .ZN(maj_143_n30)
         );
  NAND2_X1 maj_143_U16 ( .A1(maj_143_n30), .A2(maj_143_n29), .ZN(maj_143_n31)
         );
  NAND2_X1 maj_143_U15 ( .A1(v_2_1[5]), .A2(maj_143_n25), .ZN(maj_143_n18) );
  NAND2_X1 maj_143_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_143_n19) );
  NAND2_X1 maj_143_U13 ( .A1(maj_143_n19), .A2(maj_143_n18), .ZN(maj_143_n22)
         );
  NAND2_X1 maj_143_U12 ( .A1(v_2_1[2]), .A2(maj_143_n24), .ZN(maj_143_n20) );
  NAND2_X1 maj_143_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_143_n21) );
  NAND2_X1 maj_143_U10 ( .A1(maj_143_n21), .A2(maj_143_n20), .ZN(maj_143_n23)
         );
  XOR2_X1 maj_143_U9 ( .A(v_2_1[2]), .B(maj_143_n24), .Z(maj_143_n26) );
  XOR2_X1 maj_143_U8 ( .A(v_2_1[5]), .B(maj_143_n25), .Z(maj_143_n27) );
  XOR2_X1 maj_143_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_143_n24) );
  XOR2_X1 maj_143_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_143_n25) );
  OR2_X1 maj_143_U5 ( .A1(maj_143_n23), .A2(maj_143_n22), .ZN(maj_143_n32) );
  NAND2_X1 maj_143_U4 ( .A1(maj_143_n22), .A2(maj_143_n23), .ZN(maj_143_n34)
         );
  NAND2_X1 maj_143_U3 ( .A1(maj_143_n32), .A2(maj_143_n31), .ZN(maj_143_n33)
         );
  NAND2_X1 maj_143_U2 ( .A1(maj_143_n34), .A2(maj_143_n33), .ZN(maj_143_port_o) );
  OR2_X1 maj_144_U19 ( .A1(maj_144_n27), .A2(maj_144_n26), .ZN(maj_144_n28) );
  NAND2_X1 maj_144_U18 ( .A1(u_0_0[6]), .A2(maj_144_n28), .ZN(maj_144_n29) );
  NAND2_X1 maj_144_U17 ( .A1(maj_144_n26), .A2(maj_144_n27), .ZN(maj_144_n30)
         );
  NAND2_X1 maj_144_U16 ( .A1(maj_144_n30), .A2(maj_144_n29), .ZN(maj_144_n31)
         );
  NAND2_X1 maj_144_U15 ( .A1(u_0_0[5]), .A2(maj_144_n25), .ZN(maj_144_n18) );
  NAND2_X1 maj_144_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_144_n19) );
  NAND2_X1 maj_144_U13 ( .A1(maj_144_n19), .A2(maj_144_n18), .ZN(maj_144_n22)
         );
  NAND2_X1 maj_144_U12 ( .A1(u_0_0[2]), .A2(maj_144_n24), .ZN(maj_144_n20) );
  NAND2_X1 maj_144_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_144_n21) );
  NAND2_X1 maj_144_U10 ( .A1(maj_144_n21), .A2(maj_144_n20), .ZN(maj_144_n23)
         );
  XOR2_X1 maj_144_U9 ( .A(u_0_0[2]), .B(maj_144_n24), .Z(maj_144_n26) );
  XOR2_X1 maj_144_U8 ( .A(u_0_0[5]), .B(maj_144_n25), .Z(maj_144_n27) );
  XOR2_X1 maj_144_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_144_n24) );
  XOR2_X1 maj_144_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_144_n25) );
  OR2_X1 maj_144_U5 ( .A1(maj_144_n23), .A2(maj_144_n22), .ZN(maj_144_n32) );
  NAND2_X1 maj_144_U4 ( .A1(maj_144_n22), .A2(maj_144_n23), .ZN(maj_144_n34)
         );
  NAND2_X1 maj_144_U3 ( .A1(maj_144_n32), .A2(maj_144_n31), .ZN(maj_144_n33)
         );
  NAND2_X1 maj_144_U2 ( .A1(maj_144_n34), .A2(maj_144_n33), .ZN(maj_144_port_o) );
  OR2_X1 maj_145_U19 ( .A1(maj_145_n27), .A2(maj_145_n26), .ZN(maj_145_n28) );
  NAND2_X1 maj_145_U18 ( .A1(v_0_0[6]), .A2(maj_145_n28), .ZN(maj_145_n29) );
  NAND2_X1 maj_145_U17 ( .A1(maj_145_n26), .A2(maj_145_n27), .ZN(maj_145_n30)
         );
  NAND2_X1 maj_145_U16 ( .A1(maj_145_n30), .A2(maj_145_n29), .ZN(maj_145_n31)
         );
  NAND2_X1 maj_145_U15 ( .A1(v_0_0[5]), .A2(maj_145_n25), .ZN(maj_145_n18) );
  NAND2_X1 maj_145_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_145_n19) );
  NAND2_X1 maj_145_U13 ( .A1(maj_145_n19), .A2(maj_145_n18), .ZN(maj_145_n22)
         );
  NAND2_X1 maj_145_U12 ( .A1(v_0_0[2]), .A2(maj_145_n24), .ZN(maj_145_n20) );
  NAND2_X1 maj_145_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_145_n21) );
  NAND2_X1 maj_145_U10 ( .A1(maj_145_n21), .A2(maj_145_n20), .ZN(maj_145_n23)
         );
  XOR2_X1 maj_145_U9 ( .A(v_0_0[2]), .B(maj_145_n24), .Z(maj_145_n26) );
  XOR2_X1 maj_145_U8 ( .A(v_0_0[5]), .B(maj_145_n25), .Z(maj_145_n27) );
  XOR2_X1 maj_145_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_145_n24) );
  XOR2_X1 maj_145_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_145_n25) );
  OR2_X1 maj_145_U5 ( .A1(maj_145_n23), .A2(maj_145_n22), .ZN(maj_145_n32) );
  NAND2_X1 maj_145_U4 ( .A1(maj_145_n22), .A2(maj_145_n23), .ZN(maj_145_n34)
         );
  NAND2_X1 maj_145_U3 ( .A1(maj_145_n32), .A2(maj_145_n31), .ZN(maj_145_n33)
         );
  NAND2_X1 maj_145_U2 ( .A1(maj_145_n34), .A2(maj_145_n33), .ZN(maj_145_port_o) );
  OR2_X1 maj_146_U19 ( .A1(maj_146_n27), .A2(maj_146_n26), .ZN(maj_146_n28) );
  NAND2_X1 maj_146_U18 ( .A1(u_0_1[6]), .A2(maj_146_n28), .ZN(maj_146_n29) );
  NAND2_X1 maj_146_U17 ( .A1(maj_146_n26), .A2(maj_146_n27), .ZN(maj_146_n30)
         );
  NAND2_X1 maj_146_U16 ( .A1(maj_146_n30), .A2(maj_146_n29), .ZN(maj_146_n31)
         );
  NAND2_X1 maj_146_U15 ( .A1(u_0_1[5]), .A2(maj_146_n25), .ZN(maj_146_n18) );
  NAND2_X1 maj_146_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_146_n19) );
  NAND2_X1 maj_146_U13 ( .A1(maj_146_n19), .A2(maj_146_n18), .ZN(maj_146_n22)
         );
  NAND2_X1 maj_146_U12 ( .A1(u_0_1[2]), .A2(maj_146_n24), .ZN(maj_146_n20) );
  NAND2_X1 maj_146_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_146_n21) );
  NAND2_X1 maj_146_U10 ( .A1(maj_146_n21), .A2(maj_146_n20), .ZN(maj_146_n23)
         );
  XOR2_X1 maj_146_U9 ( .A(u_0_1[2]), .B(maj_146_n24), .Z(maj_146_n26) );
  XOR2_X1 maj_146_U8 ( .A(u_0_1[5]), .B(maj_146_n25), .Z(maj_146_n27) );
  XOR2_X1 maj_146_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_146_n24) );
  XOR2_X1 maj_146_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_146_n25) );
  OR2_X1 maj_146_U5 ( .A1(maj_146_n23), .A2(maj_146_n22), .ZN(maj_146_n32) );
  NAND2_X1 maj_146_U4 ( .A1(maj_146_n22), .A2(maj_146_n23), .ZN(maj_146_n34)
         );
  NAND2_X1 maj_146_U3 ( .A1(maj_146_n32), .A2(maj_146_n31), .ZN(maj_146_n33)
         );
  NAND2_X1 maj_146_U2 ( .A1(maj_146_n34), .A2(maj_146_n33), .ZN(maj_146_port_o) );
  OR2_X1 maj_147_U19 ( .A1(maj_147_n27), .A2(maj_147_n26), .ZN(maj_147_n28) );
  NAND2_X1 maj_147_U18 ( .A1(v_0_1[6]), .A2(maj_147_n28), .ZN(maj_147_n29) );
  NAND2_X1 maj_147_U17 ( .A1(maj_147_n26), .A2(maj_147_n27), .ZN(maj_147_n30)
         );
  NAND2_X1 maj_147_U16 ( .A1(maj_147_n30), .A2(maj_147_n29), .ZN(maj_147_n31)
         );
  NAND2_X1 maj_147_U15 ( .A1(v_0_1[5]), .A2(maj_147_n25), .ZN(maj_147_n18) );
  NAND2_X1 maj_147_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_147_n19) );
  NAND2_X1 maj_147_U13 ( .A1(maj_147_n19), .A2(maj_147_n18), .ZN(maj_147_n22)
         );
  NAND2_X1 maj_147_U12 ( .A1(v_0_1[2]), .A2(maj_147_n24), .ZN(maj_147_n20) );
  NAND2_X1 maj_147_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_147_n21) );
  NAND2_X1 maj_147_U10 ( .A1(maj_147_n21), .A2(maj_147_n20), .ZN(maj_147_n23)
         );
  XOR2_X1 maj_147_U9 ( .A(v_0_1[2]), .B(maj_147_n24), .Z(maj_147_n26) );
  XOR2_X1 maj_147_U8 ( .A(v_0_1[5]), .B(maj_147_n25), .Z(maj_147_n27) );
  XOR2_X1 maj_147_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_147_n24) );
  XOR2_X1 maj_147_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_147_n25) );
  OR2_X1 maj_147_U5 ( .A1(maj_147_n23), .A2(maj_147_n22), .ZN(maj_147_n32) );
  NAND2_X1 maj_147_U4 ( .A1(maj_147_n22), .A2(maj_147_n23), .ZN(maj_147_n34)
         );
  NAND2_X1 maj_147_U3 ( .A1(maj_147_n32), .A2(maj_147_n31), .ZN(maj_147_n33)
         );
  NAND2_X1 maj_147_U2 ( .A1(maj_147_n34), .A2(maj_147_n33), .ZN(maj_147_port_o) );
  OR2_X1 maj_148_U19 ( .A1(maj_148_n27), .A2(maj_148_n26), .ZN(maj_148_n28) );
  NAND2_X1 maj_148_U18 ( .A1(u_1_0[6]), .A2(maj_148_n28), .ZN(maj_148_n29) );
  NAND2_X1 maj_148_U17 ( .A1(maj_148_n26), .A2(maj_148_n27), .ZN(maj_148_n30)
         );
  NAND2_X1 maj_148_U16 ( .A1(maj_148_n30), .A2(maj_148_n29), .ZN(maj_148_n31)
         );
  NAND2_X1 maj_148_U15 ( .A1(u_1_0[5]), .A2(maj_148_n25), .ZN(maj_148_n18) );
  NAND2_X1 maj_148_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_148_n19) );
  NAND2_X1 maj_148_U13 ( .A1(maj_148_n19), .A2(maj_148_n18), .ZN(maj_148_n22)
         );
  NAND2_X1 maj_148_U12 ( .A1(u_1_0[2]), .A2(maj_148_n24), .ZN(maj_148_n20) );
  NAND2_X1 maj_148_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_148_n21) );
  NAND2_X1 maj_148_U10 ( .A1(maj_148_n21), .A2(maj_148_n20), .ZN(maj_148_n23)
         );
  XOR2_X1 maj_148_U9 ( .A(u_1_0[2]), .B(maj_148_n24), .Z(maj_148_n26) );
  XOR2_X1 maj_148_U8 ( .A(u_1_0[5]), .B(maj_148_n25), .Z(maj_148_n27) );
  XOR2_X1 maj_148_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_148_n24) );
  XOR2_X1 maj_148_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_148_n25) );
  OR2_X1 maj_148_U5 ( .A1(maj_148_n23), .A2(maj_148_n22), .ZN(maj_148_n32) );
  NAND2_X1 maj_148_U4 ( .A1(maj_148_n22), .A2(maj_148_n23), .ZN(maj_148_n34)
         );
  NAND2_X1 maj_148_U3 ( .A1(maj_148_n32), .A2(maj_148_n31), .ZN(maj_148_n33)
         );
  NAND2_X1 maj_148_U2 ( .A1(maj_148_n34), .A2(maj_148_n33), .ZN(maj_148_port_o) );
  OR2_X1 maj_149_U19 ( .A1(maj_149_n27), .A2(maj_149_n26), .ZN(maj_149_n28) );
  NAND2_X1 maj_149_U18 ( .A1(v_1_0[6]), .A2(maj_149_n28), .ZN(maj_149_n29) );
  NAND2_X1 maj_149_U17 ( .A1(maj_149_n26), .A2(maj_149_n27), .ZN(maj_149_n30)
         );
  NAND2_X1 maj_149_U16 ( .A1(maj_149_n30), .A2(maj_149_n29), .ZN(maj_149_n31)
         );
  NAND2_X1 maj_149_U15 ( .A1(v_1_0[5]), .A2(maj_149_n25), .ZN(maj_149_n18) );
  NAND2_X1 maj_149_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_149_n19) );
  NAND2_X1 maj_149_U13 ( .A1(maj_149_n19), .A2(maj_149_n18), .ZN(maj_149_n22)
         );
  NAND2_X1 maj_149_U12 ( .A1(v_1_0[2]), .A2(maj_149_n24), .ZN(maj_149_n20) );
  NAND2_X1 maj_149_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_149_n21) );
  NAND2_X1 maj_149_U10 ( .A1(maj_149_n21), .A2(maj_149_n20), .ZN(maj_149_n23)
         );
  XOR2_X1 maj_149_U9 ( .A(v_1_0[2]), .B(maj_149_n24), .Z(maj_149_n26) );
  XOR2_X1 maj_149_U8 ( .A(v_1_0[5]), .B(maj_149_n25), .Z(maj_149_n27) );
  XOR2_X1 maj_149_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_149_n24) );
  XOR2_X1 maj_149_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_149_n25) );
  OR2_X1 maj_149_U5 ( .A1(maj_149_n23), .A2(maj_149_n22), .ZN(maj_149_n32) );
  NAND2_X1 maj_149_U4 ( .A1(maj_149_n22), .A2(maj_149_n23), .ZN(maj_149_n34)
         );
  NAND2_X1 maj_149_U3 ( .A1(maj_149_n32), .A2(maj_149_n31), .ZN(maj_149_n33)
         );
  NAND2_X1 maj_149_U2 ( .A1(maj_149_n34), .A2(maj_149_n33), .ZN(maj_149_port_o) );
  OR2_X1 maj_150_U19 ( .A1(maj_150_n27), .A2(maj_150_n26), .ZN(maj_150_n28) );
  NAND2_X1 maj_150_U18 ( .A1(u_1_1[6]), .A2(maj_150_n28), .ZN(maj_150_n29) );
  NAND2_X1 maj_150_U17 ( .A1(maj_150_n26), .A2(maj_150_n27), .ZN(maj_150_n30)
         );
  NAND2_X1 maj_150_U16 ( .A1(maj_150_n30), .A2(maj_150_n29), .ZN(maj_150_n31)
         );
  NAND2_X1 maj_150_U15 ( .A1(u_1_1[5]), .A2(maj_150_n25), .ZN(maj_150_n18) );
  NAND2_X1 maj_150_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_150_n19) );
  NAND2_X1 maj_150_U13 ( .A1(maj_150_n19), .A2(maj_150_n18), .ZN(maj_150_n22)
         );
  NAND2_X1 maj_150_U12 ( .A1(u_1_1[2]), .A2(maj_150_n24), .ZN(maj_150_n20) );
  NAND2_X1 maj_150_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_150_n21) );
  NAND2_X1 maj_150_U10 ( .A1(maj_150_n21), .A2(maj_150_n20), .ZN(maj_150_n23)
         );
  XOR2_X1 maj_150_U9 ( .A(u_1_1[2]), .B(maj_150_n24), .Z(maj_150_n26) );
  XOR2_X1 maj_150_U8 ( .A(u_1_1[5]), .B(maj_150_n25), .Z(maj_150_n27) );
  XOR2_X1 maj_150_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_150_n24) );
  XOR2_X1 maj_150_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_150_n25) );
  OR2_X1 maj_150_U5 ( .A1(maj_150_n23), .A2(maj_150_n22), .ZN(maj_150_n32) );
  NAND2_X1 maj_150_U4 ( .A1(maj_150_n22), .A2(maj_150_n23), .ZN(maj_150_n34)
         );
  NAND2_X1 maj_150_U3 ( .A1(maj_150_n32), .A2(maj_150_n31), .ZN(maj_150_n33)
         );
  NAND2_X1 maj_150_U2 ( .A1(maj_150_n34), .A2(maj_150_n33), .ZN(maj_150_port_o) );
  OR2_X1 maj_151_U19 ( .A1(maj_151_n27), .A2(maj_151_n26), .ZN(maj_151_n28) );
  NAND2_X1 maj_151_U18 ( .A1(v_1_1[6]), .A2(maj_151_n28), .ZN(maj_151_n29) );
  NAND2_X1 maj_151_U17 ( .A1(maj_151_n26), .A2(maj_151_n27), .ZN(maj_151_n30)
         );
  NAND2_X1 maj_151_U16 ( .A1(maj_151_n30), .A2(maj_151_n29), .ZN(maj_151_n31)
         );
  NAND2_X1 maj_151_U15 ( .A1(v_1_1[5]), .A2(maj_151_n25), .ZN(maj_151_n18) );
  NAND2_X1 maj_151_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_151_n19) );
  NAND2_X1 maj_151_U13 ( .A1(maj_151_n19), .A2(maj_151_n18), .ZN(maj_151_n22)
         );
  NAND2_X1 maj_151_U12 ( .A1(v_1_1[2]), .A2(maj_151_n24), .ZN(maj_151_n20) );
  NAND2_X1 maj_151_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_151_n21) );
  NAND2_X1 maj_151_U10 ( .A1(maj_151_n21), .A2(maj_151_n20), .ZN(maj_151_n23)
         );
  XOR2_X1 maj_151_U9 ( .A(v_1_1[2]), .B(maj_151_n24), .Z(maj_151_n26) );
  XOR2_X1 maj_151_U8 ( .A(v_1_1[5]), .B(maj_151_n25), .Z(maj_151_n27) );
  XOR2_X1 maj_151_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_151_n24) );
  XOR2_X1 maj_151_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_151_n25) );
  OR2_X1 maj_151_U5 ( .A1(maj_151_n23), .A2(maj_151_n22), .ZN(maj_151_n32) );
  NAND2_X1 maj_151_U4 ( .A1(maj_151_n22), .A2(maj_151_n23), .ZN(maj_151_n34)
         );
  NAND2_X1 maj_151_U3 ( .A1(maj_151_n32), .A2(maj_151_n31), .ZN(maj_151_n33)
         );
  NAND2_X1 maj_151_U2 ( .A1(maj_151_n34), .A2(maj_151_n33), .ZN(maj_151_port_o) );
  OR2_X1 maj_152_U19 ( .A1(maj_152_n27), .A2(maj_152_n26), .ZN(maj_152_n28) );
  NAND2_X1 maj_152_U18 ( .A1(u_2_0[6]), .A2(maj_152_n28), .ZN(maj_152_n29) );
  NAND2_X1 maj_152_U17 ( .A1(maj_152_n26), .A2(maj_152_n27), .ZN(maj_152_n30)
         );
  NAND2_X1 maj_152_U16 ( .A1(maj_152_n30), .A2(maj_152_n29), .ZN(maj_152_n31)
         );
  NAND2_X1 maj_152_U15 ( .A1(u_2_0[5]), .A2(maj_152_n25), .ZN(maj_152_n18) );
  NAND2_X1 maj_152_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_152_n19) );
  NAND2_X1 maj_152_U13 ( .A1(maj_152_n19), .A2(maj_152_n18), .ZN(maj_152_n22)
         );
  NAND2_X1 maj_152_U12 ( .A1(u_2_0[2]), .A2(maj_152_n24), .ZN(maj_152_n20) );
  NAND2_X1 maj_152_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_152_n21) );
  NAND2_X1 maj_152_U10 ( .A1(maj_152_n21), .A2(maj_152_n20), .ZN(maj_152_n23)
         );
  XOR2_X1 maj_152_U9 ( .A(u_2_0[2]), .B(maj_152_n24), .Z(maj_152_n26) );
  XOR2_X1 maj_152_U8 ( .A(u_2_0[5]), .B(maj_152_n25), .Z(maj_152_n27) );
  XOR2_X1 maj_152_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_152_n24) );
  XOR2_X1 maj_152_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_152_n25) );
  OR2_X1 maj_152_U5 ( .A1(maj_152_n23), .A2(maj_152_n22), .ZN(maj_152_n32) );
  NAND2_X1 maj_152_U4 ( .A1(maj_152_n22), .A2(maj_152_n23), .ZN(maj_152_n34)
         );
  NAND2_X1 maj_152_U3 ( .A1(maj_152_n32), .A2(maj_152_n31), .ZN(maj_152_n33)
         );
  NAND2_X1 maj_152_U2 ( .A1(maj_152_n34), .A2(maj_152_n33), .ZN(maj_152_port_o) );
  OR2_X1 maj_153_U19 ( .A1(maj_153_n27), .A2(maj_153_n26), .ZN(maj_153_n28) );
  NAND2_X1 maj_153_U18 ( .A1(v_2_0[6]), .A2(maj_153_n28), .ZN(maj_153_n29) );
  NAND2_X1 maj_153_U17 ( .A1(maj_153_n26), .A2(maj_153_n27), .ZN(maj_153_n30)
         );
  NAND2_X1 maj_153_U16 ( .A1(maj_153_n30), .A2(maj_153_n29), .ZN(maj_153_n31)
         );
  NAND2_X1 maj_153_U15 ( .A1(v_2_0[5]), .A2(maj_153_n25), .ZN(maj_153_n18) );
  NAND2_X1 maj_153_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_153_n19) );
  NAND2_X1 maj_153_U13 ( .A1(maj_153_n19), .A2(maj_153_n18), .ZN(maj_153_n22)
         );
  NAND2_X1 maj_153_U12 ( .A1(v_2_0[2]), .A2(maj_153_n24), .ZN(maj_153_n20) );
  NAND2_X1 maj_153_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_153_n21) );
  NAND2_X1 maj_153_U10 ( .A1(maj_153_n21), .A2(maj_153_n20), .ZN(maj_153_n23)
         );
  XOR2_X1 maj_153_U9 ( .A(v_2_0[2]), .B(maj_153_n24), .Z(maj_153_n26) );
  XOR2_X1 maj_153_U8 ( .A(v_2_0[5]), .B(maj_153_n25), .Z(maj_153_n27) );
  XOR2_X1 maj_153_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_153_n24) );
  XOR2_X1 maj_153_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_153_n25) );
  OR2_X1 maj_153_U5 ( .A1(maj_153_n23), .A2(maj_153_n22), .ZN(maj_153_n32) );
  NAND2_X1 maj_153_U4 ( .A1(maj_153_n22), .A2(maj_153_n23), .ZN(maj_153_n34)
         );
  NAND2_X1 maj_153_U3 ( .A1(maj_153_n32), .A2(maj_153_n31), .ZN(maj_153_n33)
         );
  NAND2_X1 maj_153_U2 ( .A1(maj_153_n34), .A2(maj_153_n33), .ZN(maj_153_port_o) );
  OR2_X1 maj_154_U19 ( .A1(maj_154_n27), .A2(maj_154_n26), .ZN(maj_154_n28) );
  NAND2_X1 maj_154_U18 ( .A1(u_2_1[6]), .A2(maj_154_n28), .ZN(maj_154_n29) );
  NAND2_X1 maj_154_U17 ( .A1(maj_154_n26), .A2(maj_154_n27), .ZN(maj_154_n30)
         );
  NAND2_X1 maj_154_U16 ( .A1(maj_154_n30), .A2(maj_154_n29), .ZN(maj_154_n31)
         );
  NAND2_X1 maj_154_U15 ( .A1(u_2_1[5]), .A2(maj_154_n25), .ZN(maj_154_n18) );
  NAND2_X1 maj_154_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_154_n19) );
  NAND2_X1 maj_154_U13 ( .A1(maj_154_n19), .A2(maj_154_n18), .ZN(maj_154_n22)
         );
  NAND2_X1 maj_154_U12 ( .A1(u_2_1[2]), .A2(maj_154_n24), .ZN(maj_154_n20) );
  NAND2_X1 maj_154_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_154_n21) );
  NAND2_X1 maj_154_U10 ( .A1(maj_154_n21), .A2(maj_154_n20), .ZN(maj_154_n23)
         );
  XOR2_X1 maj_154_U9 ( .A(u_2_1[2]), .B(maj_154_n24), .Z(maj_154_n26) );
  XOR2_X1 maj_154_U8 ( .A(u_2_1[5]), .B(maj_154_n25), .Z(maj_154_n27) );
  XOR2_X1 maj_154_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_154_n24) );
  XOR2_X1 maj_154_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_154_n25) );
  OR2_X1 maj_154_U5 ( .A1(maj_154_n23), .A2(maj_154_n22), .ZN(maj_154_n32) );
  NAND2_X1 maj_154_U4 ( .A1(maj_154_n22), .A2(maj_154_n23), .ZN(maj_154_n34)
         );
  NAND2_X1 maj_154_U3 ( .A1(maj_154_n32), .A2(maj_154_n31), .ZN(maj_154_n33)
         );
  NAND2_X1 maj_154_U2 ( .A1(maj_154_n34), .A2(maj_154_n33), .ZN(maj_154_port_o) );
  OR2_X1 maj_155_U19 ( .A1(maj_155_n27), .A2(maj_155_n26), .ZN(maj_155_n28) );
  NAND2_X1 maj_155_U18 ( .A1(v_2_1[6]), .A2(maj_155_n28), .ZN(maj_155_n29) );
  NAND2_X1 maj_155_U17 ( .A1(maj_155_n26), .A2(maj_155_n27), .ZN(maj_155_n30)
         );
  NAND2_X1 maj_155_U16 ( .A1(maj_155_n30), .A2(maj_155_n29), .ZN(maj_155_n31)
         );
  NAND2_X1 maj_155_U15 ( .A1(v_2_1[5]), .A2(maj_155_n25), .ZN(maj_155_n18) );
  NAND2_X1 maj_155_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_155_n19) );
  NAND2_X1 maj_155_U13 ( .A1(maj_155_n19), .A2(maj_155_n18), .ZN(maj_155_n22)
         );
  NAND2_X1 maj_155_U12 ( .A1(v_2_1[2]), .A2(maj_155_n24), .ZN(maj_155_n20) );
  NAND2_X1 maj_155_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_155_n21) );
  NAND2_X1 maj_155_U10 ( .A1(maj_155_n21), .A2(maj_155_n20), .ZN(maj_155_n23)
         );
  XOR2_X1 maj_155_U9 ( .A(v_2_1[2]), .B(maj_155_n24), .Z(maj_155_n26) );
  XOR2_X1 maj_155_U8 ( .A(v_2_1[5]), .B(maj_155_n25), .Z(maj_155_n27) );
  XOR2_X1 maj_155_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_155_n24) );
  XOR2_X1 maj_155_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_155_n25) );
  OR2_X1 maj_155_U5 ( .A1(maj_155_n23), .A2(maj_155_n22), .ZN(maj_155_n32) );
  NAND2_X1 maj_155_U4 ( .A1(maj_155_n22), .A2(maj_155_n23), .ZN(maj_155_n34)
         );
  NAND2_X1 maj_155_U3 ( .A1(maj_155_n32), .A2(maj_155_n31), .ZN(maj_155_n33)
         );
  NAND2_X1 maj_155_U2 ( .A1(maj_155_n34), .A2(maj_155_n33), .ZN(maj_155_port_o) );
  OR2_X1 maj_156_U19 ( .A1(maj_156_n27), .A2(maj_156_n26), .ZN(maj_156_n28) );
  NAND2_X1 maj_156_U18 ( .A1(u_0_0[6]), .A2(maj_156_n28), .ZN(maj_156_n29) );
  NAND2_X1 maj_156_U17 ( .A1(maj_156_n26), .A2(maj_156_n27), .ZN(maj_156_n30)
         );
  NAND2_X1 maj_156_U16 ( .A1(maj_156_n30), .A2(maj_156_n29), .ZN(maj_156_n31)
         );
  NAND2_X1 maj_156_U15 ( .A1(u_0_0[5]), .A2(maj_156_n25), .ZN(maj_156_n18) );
  NAND2_X1 maj_156_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_156_n19) );
  NAND2_X1 maj_156_U13 ( .A1(maj_156_n19), .A2(maj_156_n18), .ZN(maj_156_n22)
         );
  NAND2_X1 maj_156_U12 ( .A1(u_0_0[2]), .A2(maj_156_n24), .ZN(maj_156_n20) );
  NAND2_X1 maj_156_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_156_n21) );
  NAND2_X1 maj_156_U10 ( .A1(maj_156_n21), .A2(maj_156_n20), .ZN(maj_156_n23)
         );
  XOR2_X1 maj_156_U9 ( .A(u_0_0[2]), .B(maj_156_n24), .Z(maj_156_n26) );
  XOR2_X1 maj_156_U8 ( .A(u_0_0[5]), .B(maj_156_n25), .Z(maj_156_n27) );
  XOR2_X1 maj_156_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_156_n24) );
  XOR2_X1 maj_156_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_156_n25) );
  OR2_X1 maj_156_U5 ( .A1(maj_156_n23), .A2(maj_156_n22), .ZN(maj_156_n32) );
  NAND2_X1 maj_156_U4 ( .A1(maj_156_n22), .A2(maj_156_n23), .ZN(maj_156_n34)
         );
  NAND2_X1 maj_156_U3 ( .A1(maj_156_n32), .A2(maj_156_n31), .ZN(maj_156_n33)
         );
  NAND2_X1 maj_156_U2 ( .A1(maj_156_n34), .A2(maj_156_n33), .ZN(maj_156_port_o) );
  OR2_X1 maj_157_U19 ( .A1(maj_157_n27), .A2(maj_157_n26), .ZN(maj_157_n28) );
  NAND2_X1 maj_157_U18 ( .A1(v_0_0[6]), .A2(maj_157_n28), .ZN(maj_157_n29) );
  NAND2_X1 maj_157_U17 ( .A1(maj_157_n26), .A2(maj_157_n27), .ZN(maj_157_n30)
         );
  NAND2_X1 maj_157_U16 ( .A1(maj_157_n30), .A2(maj_157_n29), .ZN(maj_157_n31)
         );
  NAND2_X1 maj_157_U15 ( .A1(v_0_0[5]), .A2(maj_157_n25), .ZN(maj_157_n18) );
  NAND2_X1 maj_157_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_157_n19) );
  NAND2_X1 maj_157_U13 ( .A1(maj_157_n19), .A2(maj_157_n18), .ZN(maj_157_n22)
         );
  NAND2_X1 maj_157_U12 ( .A1(v_0_0[2]), .A2(maj_157_n24), .ZN(maj_157_n20) );
  NAND2_X1 maj_157_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_157_n21) );
  NAND2_X1 maj_157_U10 ( .A1(maj_157_n21), .A2(maj_157_n20), .ZN(maj_157_n23)
         );
  XOR2_X1 maj_157_U9 ( .A(v_0_0[2]), .B(maj_157_n24), .Z(maj_157_n26) );
  XOR2_X1 maj_157_U8 ( .A(v_0_0[5]), .B(maj_157_n25), .Z(maj_157_n27) );
  XOR2_X1 maj_157_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_157_n24) );
  XOR2_X1 maj_157_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_157_n25) );
  OR2_X1 maj_157_U5 ( .A1(maj_157_n23), .A2(maj_157_n22), .ZN(maj_157_n32) );
  NAND2_X1 maj_157_U4 ( .A1(maj_157_n22), .A2(maj_157_n23), .ZN(maj_157_n34)
         );
  NAND2_X1 maj_157_U3 ( .A1(maj_157_n32), .A2(maj_157_n31), .ZN(maj_157_n33)
         );
  NAND2_X1 maj_157_U2 ( .A1(maj_157_n34), .A2(maj_157_n33), .ZN(maj_157_port_o) );
  OR2_X1 maj_158_U19 ( .A1(maj_158_n27), .A2(maj_158_n26), .ZN(maj_158_n28) );
  NAND2_X1 maj_158_U18 ( .A1(u_0_1[6]), .A2(maj_158_n28), .ZN(maj_158_n29) );
  NAND2_X1 maj_158_U17 ( .A1(maj_158_n26), .A2(maj_158_n27), .ZN(maj_158_n30)
         );
  NAND2_X1 maj_158_U16 ( .A1(maj_158_n30), .A2(maj_158_n29), .ZN(maj_158_n31)
         );
  NAND2_X1 maj_158_U15 ( .A1(u_0_1[5]), .A2(maj_158_n25), .ZN(maj_158_n18) );
  NAND2_X1 maj_158_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_158_n19) );
  NAND2_X1 maj_158_U13 ( .A1(maj_158_n19), .A2(maj_158_n18), .ZN(maj_158_n22)
         );
  NAND2_X1 maj_158_U12 ( .A1(u_0_1[2]), .A2(maj_158_n24), .ZN(maj_158_n20) );
  NAND2_X1 maj_158_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_158_n21) );
  NAND2_X1 maj_158_U10 ( .A1(maj_158_n21), .A2(maj_158_n20), .ZN(maj_158_n23)
         );
  XOR2_X1 maj_158_U9 ( .A(u_0_1[2]), .B(maj_158_n24), .Z(maj_158_n26) );
  XOR2_X1 maj_158_U8 ( .A(u_0_1[5]), .B(maj_158_n25), .Z(maj_158_n27) );
  XOR2_X1 maj_158_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_158_n24) );
  XOR2_X1 maj_158_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_158_n25) );
  OR2_X1 maj_158_U5 ( .A1(maj_158_n23), .A2(maj_158_n22), .ZN(maj_158_n32) );
  NAND2_X1 maj_158_U4 ( .A1(maj_158_n22), .A2(maj_158_n23), .ZN(maj_158_n34)
         );
  NAND2_X1 maj_158_U3 ( .A1(maj_158_n32), .A2(maj_158_n31), .ZN(maj_158_n33)
         );
  NAND2_X1 maj_158_U2 ( .A1(maj_158_n34), .A2(maj_158_n33), .ZN(maj_158_port_o) );
  OR2_X1 maj_159_U19 ( .A1(maj_159_n27), .A2(maj_159_n26), .ZN(maj_159_n28) );
  NAND2_X1 maj_159_U18 ( .A1(v_0_1[6]), .A2(maj_159_n28), .ZN(maj_159_n29) );
  NAND2_X1 maj_159_U17 ( .A1(maj_159_n26), .A2(maj_159_n27), .ZN(maj_159_n30)
         );
  NAND2_X1 maj_159_U16 ( .A1(maj_159_n30), .A2(maj_159_n29), .ZN(maj_159_n31)
         );
  NAND2_X1 maj_159_U15 ( .A1(v_0_1[5]), .A2(maj_159_n25), .ZN(maj_159_n18) );
  NAND2_X1 maj_159_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_159_n19) );
  NAND2_X1 maj_159_U13 ( .A1(maj_159_n19), .A2(maj_159_n18), .ZN(maj_159_n22)
         );
  NAND2_X1 maj_159_U12 ( .A1(v_0_1[2]), .A2(maj_159_n24), .ZN(maj_159_n20) );
  NAND2_X1 maj_159_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_159_n21) );
  NAND2_X1 maj_159_U10 ( .A1(maj_159_n21), .A2(maj_159_n20), .ZN(maj_159_n23)
         );
  XOR2_X1 maj_159_U9 ( .A(v_0_1[2]), .B(maj_159_n24), .Z(maj_159_n26) );
  XOR2_X1 maj_159_U8 ( .A(v_0_1[5]), .B(maj_159_n25), .Z(maj_159_n27) );
  XOR2_X1 maj_159_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_159_n24) );
  XOR2_X1 maj_159_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_159_n25) );
  OR2_X1 maj_159_U5 ( .A1(maj_159_n23), .A2(maj_159_n22), .ZN(maj_159_n32) );
  NAND2_X1 maj_159_U4 ( .A1(maj_159_n22), .A2(maj_159_n23), .ZN(maj_159_n34)
         );
  NAND2_X1 maj_159_U3 ( .A1(maj_159_n32), .A2(maj_159_n31), .ZN(maj_159_n33)
         );
  NAND2_X1 maj_159_U2 ( .A1(maj_159_n34), .A2(maj_159_n33), .ZN(maj_159_port_o) );
  OR2_X1 maj_160_U19 ( .A1(maj_160_n27), .A2(maj_160_n26), .ZN(maj_160_n28) );
  NAND2_X1 maj_160_U18 ( .A1(u_1_0[6]), .A2(maj_160_n28), .ZN(maj_160_n29) );
  NAND2_X1 maj_160_U17 ( .A1(maj_160_n26), .A2(maj_160_n27), .ZN(maj_160_n30)
         );
  NAND2_X1 maj_160_U16 ( .A1(maj_160_n30), .A2(maj_160_n29), .ZN(maj_160_n31)
         );
  NAND2_X1 maj_160_U15 ( .A1(u_1_0[5]), .A2(maj_160_n25), .ZN(maj_160_n18) );
  NAND2_X1 maj_160_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_160_n19) );
  NAND2_X1 maj_160_U13 ( .A1(maj_160_n19), .A2(maj_160_n18), .ZN(maj_160_n22)
         );
  NAND2_X1 maj_160_U12 ( .A1(u_1_0[2]), .A2(maj_160_n24), .ZN(maj_160_n20) );
  NAND2_X1 maj_160_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_160_n21) );
  NAND2_X1 maj_160_U10 ( .A1(maj_160_n21), .A2(maj_160_n20), .ZN(maj_160_n23)
         );
  XOR2_X1 maj_160_U9 ( .A(u_1_0[2]), .B(maj_160_n24), .Z(maj_160_n26) );
  XOR2_X1 maj_160_U8 ( .A(u_1_0[5]), .B(maj_160_n25), .Z(maj_160_n27) );
  XOR2_X1 maj_160_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_160_n24) );
  XOR2_X1 maj_160_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_160_n25) );
  OR2_X1 maj_160_U5 ( .A1(maj_160_n23), .A2(maj_160_n22), .ZN(maj_160_n32) );
  NAND2_X1 maj_160_U4 ( .A1(maj_160_n22), .A2(maj_160_n23), .ZN(maj_160_n34)
         );
  NAND2_X1 maj_160_U3 ( .A1(maj_160_n32), .A2(maj_160_n31), .ZN(maj_160_n33)
         );
  NAND2_X1 maj_160_U2 ( .A1(maj_160_n34), .A2(maj_160_n33), .ZN(maj_160_port_o) );
  OR2_X1 maj_161_U19 ( .A1(maj_161_n27), .A2(maj_161_n26), .ZN(maj_161_n28) );
  NAND2_X1 maj_161_U18 ( .A1(v_1_0[6]), .A2(maj_161_n28), .ZN(maj_161_n29) );
  NAND2_X1 maj_161_U17 ( .A1(maj_161_n26), .A2(maj_161_n27), .ZN(maj_161_n30)
         );
  NAND2_X1 maj_161_U16 ( .A1(maj_161_n30), .A2(maj_161_n29), .ZN(maj_161_n31)
         );
  NAND2_X1 maj_161_U15 ( .A1(v_1_0[5]), .A2(maj_161_n25), .ZN(maj_161_n18) );
  NAND2_X1 maj_161_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_161_n19) );
  NAND2_X1 maj_161_U13 ( .A1(maj_161_n19), .A2(maj_161_n18), .ZN(maj_161_n22)
         );
  NAND2_X1 maj_161_U12 ( .A1(v_1_0[2]), .A2(maj_161_n24), .ZN(maj_161_n20) );
  NAND2_X1 maj_161_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_161_n21) );
  NAND2_X1 maj_161_U10 ( .A1(maj_161_n21), .A2(maj_161_n20), .ZN(maj_161_n23)
         );
  XOR2_X1 maj_161_U9 ( .A(v_1_0[2]), .B(maj_161_n24), .Z(maj_161_n26) );
  XOR2_X1 maj_161_U8 ( .A(v_1_0[5]), .B(maj_161_n25), .Z(maj_161_n27) );
  XOR2_X1 maj_161_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_161_n24) );
  XOR2_X1 maj_161_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_161_n25) );
  OR2_X1 maj_161_U5 ( .A1(maj_161_n23), .A2(maj_161_n22), .ZN(maj_161_n32) );
  NAND2_X1 maj_161_U4 ( .A1(maj_161_n22), .A2(maj_161_n23), .ZN(maj_161_n34)
         );
  NAND2_X1 maj_161_U3 ( .A1(maj_161_n32), .A2(maj_161_n31), .ZN(maj_161_n33)
         );
  NAND2_X1 maj_161_U2 ( .A1(maj_161_n34), .A2(maj_161_n33), .ZN(maj_161_port_o) );
  OR2_X1 maj_162_U19 ( .A1(maj_162_n27), .A2(maj_162_n26), .ZN(maj_162_n28) );
  NAND2_X1 maj_162_U18 ( .A1(u_1_1[6]), .A2(maj_162_n28), .ZN(maj_162_n29) );
  NAND2_X1 maj_162_U17 ( .A1(maj_162_n26), .A2(maj_162_n27), .ZN(maj_162_n30)
         );
  NAND2_X1 maj_162_U16 ( .A1(maj_162_n30), .A2(maj_162_n29), .ZN(maj_162_n31)
         );
  NAND2_X1 maj_162_U15 ( .A1(u_1_1[5]), .A2(maj_162_n25), .ZN(maj_162_n18) );
  NAND2_X1 maj_162_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_162_n19) );
  NAND2_X1 maj_162_U13 ( .A1(maj_162_n19), .A2(maj_162_n18), .ZN(maj_162_n22)
         );
  NAND2_X1 maj_162_U12 ( .A1(u_1_1[2]), .A2(maj_162_n24), .ZN(maj_162_n20) );
  NAND2_X1 maj_162_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_162_n21) );
  NAND2_X1 maj_162_U10 ( .A1(maj_162_n21), .A2(maj_162_n20), .ZN(maj_162_n23)
         );
  XOR2_X1 maj_162_U9 ( .A(u_1_1[2]), .B(maj_162_n24), .Z(maj_162_n26) );
  XOR2_X1 maj_162_U8 ( .A(u_1_1[5]), .B(maj_162_n25), .Z(maj_162_n27) );
  XOR2_X1 maj_162_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_162_n24) );
  XOR2_X1 maj_162_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_162_n25) );
  OR2_X1 maj_162_U5 ( .A1(maj_162_n23), .A2(maj_162_n22), .ZN(maj_162_n32) );
  NAND2_X1 maj_162_U4 ( .A1(maj_162_n22), .A2(maj_162_n23), .ZN(maj_162_n34)
         );
  NAND2_X1 maj_162_U3 ( .A1(maj_162_n32), .A2(maj_162_n31), .ZN(maj_162_n33)
         );
  NAND2_X1 maj_162_U2 ( .A1(maj_162_n34), .A2(maj_162_n33), .ZN(maj_162_port_o) );
  OR2_X1 maj_163_U19 ( .A1(maj_163_n27), .A2(maj_163_n26), .ZN(maj_163_n28) );
  NAND2_X1 maj_163_U18 ( .A1(v_1_1[6]), .A2(maj_163_n28), .ZN(maj_163_n29) );
  NAND2_X1 maj_163_U17 ( .A1(maj_163_n26), .A2(maj_163_n27), .ZN(maj_163_n30)
         );
  NAND2_X1 maj_163_U16 ( .A1(maj_163_n30), .A2(maj_163_n29), .ZN(maj_163_n31)
         );
  NAND2_X1 maj_163_U15 ( .A1(v_1_1[5]), .A2(maj_163_n25), .ZN(maj_163_n18) );
  NAND2_X1 maj_163_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_163_n19) );
  NAND2_X1 maj_163_U13 ( .A1(maj_163_n19), .A2(maj_163_n18), .ZN(maj_163_n22)
         );
  NAND2_X1 maj_163_U12 ( .A1(v_1_1[2]), .A2(maj_163_n24), .ZN(maj_163_n20) );
  NAND2_X1 maj_163_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_163_n21) );
  NAND2_X1 maj_163_U10 ( .A1(maj_163_n21), .A2(maj_163_n20), .ZN(maj_163_n23)
         );
  XOR2_X1 maj_163_U9 ( .A(v_1_1[2]), .B(maj_163_n24), .Z(maj_163_n26) );
  XOR2_X1 maj_163_U8 ( .A(v_1_1[5]), .B(maj_163_n25), .Z(maj_163_n27) );
  XOR2_X1 maj_163_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_163_n24) );
  XOR2_X1 maj_163_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_163_n25) );
  OR2_X1 maj_163_U5 ( .A1(maj_163_n23), .A2(maj_163_n22), .ZN(maj_163_n32) );
  NAND2_X1 maj_163_U4 ( .A1(maj_163_n22), .A2(maj_163_n23), .ZN(maj_163_n34)
         );
  NAND2_X1 maj_163_U3 ( .A1(maj_163_n32), .A2(maj_163_n31), .ZN(maj_163_n33)
         );
  NAND2_X1 maj_163_U2 ( .A1(maj_163_n34), .A2(maj_163_n33), .ZN(maj_163_port_o) );
  OR2_X1 maj_164_U19 ( .A1(maj_164_n27), .A2(maj_164_n26), .ZN(maj_164_n28) );
  NAND2_X1 maj_164_U18 ( .A1(u_2_0[6]), .A2(maj_164_n28), .ZN(maj_164_n29) );
  NAND2_X1 maj_164_U17 ( .A1(maj_164_n26), .A2(maj_164_n27), .ZN(maj_164_n30)
         );
  NAND2_X1 maj_164_U16 ( .A1(maj_164_n30), .A2(maj_164_n29), .ZN(maj_164_n31)
         );
  NAND2_X1 maj_164_U15 ( .A1(u_2_0[5]), .A2(maj_164_n25), .ZN(maj_164_n18) );
  NAND2_X1 maj_164_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_164_n19) );
  NAND2_X1 maj_164_U13 ( .A1(maj_164_n19), .A2(maj_164_n18), .ZN(maj_164_n22)
         );
  NAND2_X1 maj_164_U12 ( .A1(u_2_0[2]), .A2(maj_164_n24), .ZN(maj_164_n20) );
  NAND2_X1 maj_164_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_164_n21) );
  NAND2_X1 maj_164_U10 ( .A1(maj_164_n21), .A2(maj_164_n20), .ZN(maj_164_n23)
         );
  XOR2_X1 maj_164_U9 ( .A(u_2_0[2]), .B(maj_164_n24), .Z(maj_164_n26) );
  XOR2_X1 maj_164_U8 ( .A(u_2_0[5]), .B(maj_164_n25), .Z(maj_164_n27) );
  XOR2_X1 maj_164_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_164_n24) );
  XOR2_X1 maj_164_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_164_n25) );
  OR2_X1 maj_164_U5 ( .A1(maj_164_n23), .A2(maj_164_n22), .ZN(maj_164_n32) );
  NAND2_X1 maj_164_U4 ( .A1(maj_164_n22), .A2(maj_164_n23), .ZN(maj_164_n34)
         );
  NAND2_X1 maj_164_U3 ( .A1(maj_164_n32), .A2(maj_164_n31), .ZN(maj_164_n33)
         );
  NAND2_X1 maj_164_U2 ( .A1(maj_164_n34), .A2(maj_164_n33), .ZN(maj_164_port_o) );
  OR2_X1 maj_165_U19 ( .A1(maj_165_n27), .A2(maj_165_n26), .ZN(maj_165_n28) );
  NAND2_X1 maj_165_U18 ( .A1(v_2_0[6]), .A2(maj_165_n28), .ZN(maj_165_n29) );
  NAND2_X1 maj_165_U17 ( .A1(maj_165_n26), .A2(maj_165_n27), .ZN(maj_165_n30)
         );
  NAND2_X1 maj_165_U16 ( .A1(maj_165_n30), .A2(maj_165_n29), .ZN(maj_165_n31)
         );
  NAND2_X1 maj_165_U15 ( .A1(v_2_0[5]), .A2(maj_165_n25), .ZN(maj_165_n18) );
  NAND2_X1 maj_165_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_165_n19) );
  NAND2_X1 maj_165_U13 ( .A1(maj_165_n19), .A2(maj_165_n18), .ZN(maj_165_n22)
         );
  NAND2_X1 maj_165_U12 ( .A1(v_2_0[2]), .A2(maj_165_n24), .ZN(maj_165_n20) );
  NAND2_X1 maj_165_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_165_n21) );
  NAND2_X1 maj_165_U10 ( .A1(maj_165_n21), .A2(maj_165_n20), .ZN(maj_165_n23)
         );
  XOR2_X1 maj_165_U9 ( .A(v_2_0[2]), .B(maj_165_n24), .Z(maj_165_n26) );
  XOR2_X1 maj_165_U8 ( .A(v_2_0[5]), .B(maj_165_n25), .Z(maj_165_n27) );
  XOR2_X1 maj_165_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_165_n24) );
  XOR2_X1 maj_165_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_165_n25) );
  OR2_X1 maj_165_U5 ( .A1(maj_165_n23), .A2(maj_165_n22), .ZN(maj_165_n32) );
  NAND2_X1 maj_165_U4 ( .A1(maj_165_n22), .A2(maj_165_n23), .ZN(maj_165_n34)
         );
  NAND2_X1 maj_165_U3 ( .A1(maj_165_n32), .A2(maj_165_n31), .ZN(maj_165_n33)
         );
  NAND2_X1 maj_165_U2 ( .A1(maj_165_n34), .A2(maj_165_n33), .ZN(maj_165_port_o) );
  OR2_X1 maj_166_U19 ( .A1(maj_166_n27), .A2(maj_166_n26), .ZN(maj_166_n28) );
  NAND2_X1 maj_166_U18 ( .A1(u_2_1[6]), .A2(maj_166_n28), .ZN(maj_166_n29) );
  NAND2_X1 maj_166_U17 ( .A1(maj_166_n26), .A2(maj_166_n27), .ZN(maj_166_n30)
         );
  NAND2_X1 maj_166_U16 ( .A1(maj_166_n30), .A2(maj_166_n29), .ZN(maj_166_n31)
         );
  NAND2_X1 maj_166_U15 ( .A1(u_2_1[5]), .A2(maj_166_n25), .ZN(maj_166_n18) );
  NAND2_X1 maj_166_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_166_n19) );
  NAND2_X1 maj_166_U13 ( .A1(maj_166_n19), .A2(maj_166_n18), .ZN(maj_166_n22)
         );
  NAND2_X1 maj_166_U12 ( .A1(u_2_1[2]), .A2(maj_166_n24), .ZN(maj_166_n20) );
  NAND2_X1 maj_166_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_166_n21) );
  NAND2_X1 maj_166_U10 ( .A1(maj_166_n21), .A2(maj_166_n20), .ZN(maj_166_n23)
         );
  XOR2_X1 maj_166_U9 ( .A(u_2_1[2]), .B(maj_166_n24), .Z(maj_166_n26) );
  XOR2_X1 maj_166_U8 ( .A(u_2_1[5]), .B(maj_166_n25), .Z(maj_166_n27) );
  XOR2_X1 maj_166_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_166_n24) );
  XOR2_X1 maj_166_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_166_n25) );
  OR2_X1 maj_166_U5 ( .A1(maj_166_n23), .A2(maj_166_n22), .ZN(maj_166_n32) );
  NAND2_X1 maj_166_U4 ( .A1(maj_166_n22), .A2(maj_166_n23), .ZN(maj_166_n34)
         );
  NAND2_X1 maj_166_U3 ( .A1(maj_166_n32), .A2(maj_166_n31), .ZN(maj_166_n33)
         );
  NAND2_X1 maj_166_U2 ( .A1(maj_166_n34), .A2(maj_166_n33), .ZN(maj_166_port_o) );
  OR2_X1 maj_167_U19 ( .A1(maj_167_n27), .A2(maj_167_n26), .ZN(maj_167_n28) );
  NAND2_X1 maj_167_U18 ( .A1(v_2_1[6]), .A2(maj_167_n28), .ZN(maj_167_n29) );
  NAND2_X1 maj_167_U17 ( .A1(maj_167_n26), .A2(maj_167_n27), .ZN(maj_167_n30)
         );
  NAND2_X1 maj_167_U16 ( .A1(maj_167_n30), .A2(maj_167_n29), .ZN(maj_167_n31)
         );
  NAND2_X1 maj_167_U15 ( .A1(v_2_1[5]), .A2(maj_167_n25), .ZN(maj_167_n18) );
  NAND2_X1 maj_167_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_167_n19) );
  NAND2_X1 maj_167_U13 ( .A1(maj_167_n19), .A2(maj_167_n18), .ZN(maj_167_n22)
         );
  NAND2_X1 maj_167_U12 ( .A1(v_2_1[2]), .A2(maj_167_n24), .ZN(maj_167_n20) );
  NAND2_X1 maj_167_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_167_n21) );
  NAND2_X1 maj_167_U10 ( .A1(maj_167_n21), .A2(maj_167_n20), .ZN(maj_167_n23)
         );
  XOR2_X1 maj_167_U9 ( .A(v_2_1[2]), .B(maj_167_n24), .Z(maj_167_n26) );
  XOR2_X1 maj_167_U8 ( .A(v_2_1[5]), .B(maj_167_n25), .Z(maj_167_n27) );
  XOR2_X1 maj_167_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_167_n24) );
  XOR2_X1 maj_167_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_167_n25) );
  OR2_X1 maj_167_U5 ( .A1(maj_167_n23), .A2(maj_167_n22), .ZN(maj_167_n32) );
  NAND2_X1 maj_167_U4 ( .A1(maj_167_n22), .A2(maj_167_n23), .ZN(maj_167_n34)
         );
  NAND2_X1 maj_167_U3 ( .A1(maj_167_n32), .A2(maj_167_n31), .ZN(maj_167_n33)
         );
  NAND2_X1 maj_167_U2 ( .A1(maj_167_n34), .A2(maj_167_n33), .ZN(maj_167_port_o) );
endmodule

