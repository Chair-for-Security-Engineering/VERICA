
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i0_s5, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, 
        io_i1_s5, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, 
        p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, 
        p_rand_12, p_rand_13, p_rand_14, p_rand_15, p_rand_16, p_rand_17, 
        p_rand_18, p_rand_19, p_rand_20, p_rand_21, p_rand_22, p_rand_23, 
        p_rand_24, p_rand_25, p_rand_26, p_rand_27, p_rand_28, p_rand_29, 
        io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i0_s5, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, io_i1_s5,
         p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6,
         p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12,
         p_rand_13, p_rand_14, p_rand_15, p_rand_16, p_rand_17, p_rand_18,
         p_rand_19, p_rand_20, p_rand_21, p_rand_22, p_rand_23, p_rand_24,
         p_rand_25, p_rand_26, p_rand_27, p_rand_28, p_rand_29;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4, io_o0_s5;
  wire   n_hpc2_0_n108, n_hpc2_0_n107, n_hpc2_0_n106, n_hpc2_0_n105,
         n_hpc2_0_n104, n_hpc2_0_n103, n_hpc2_0_n102, n_hpc2_0_n101,
         n_hpc2_0_n100, n_hpc2_0_n99, n_hpc2_0_n98, n_hpc2_0_n97, n_hpc2_0_n96,
         n_hpc2_0_n95, n_hpc2_0_n94, n_hpc2_0_n93, n_hpc2_0_n92, n_hpc2_0_n91,
         n_hpc2_0_n90, n_hpc2_0_n89, n_hpc2_0_n88, n_hpc2_0_n87, n_hpc2_0_n86,
         n_hpc2_0_n85, n_hpc2_0_n84, n_hpc2_0_n83, n_hpc2_0_n82, n_hpc2_0_n81,
         n_hpc2_0_n80, n_hpc2_0_n79, n_hpc2_0_n78, n_hpc2_0_n77, n_hpc2_0_n76,
         n_hpc2_0_n75, n_hpc2_0_n74, n_hpc2_0_n73, n_hpc2_0_n72, n_hpc2_0_n71,
         n_hpc2_0_n70, n_hpc2_0_n69, n_hpc2_0_n68, n_hpc2_0_n67, n_hpc2_0_n66,
         n_hpc2_0_n65, n_hpc2_0_n64, n_hpc2_0_n63, n_hpc2_0_n62, n_hpc2_0_n61,
         n_hpc2_0_n60, n_hpc2_0_n59, n_hpc2_0_n58, n_hpc2_0_n57, n_hpc2_0_n56,
         n_hpc2_0_n55, n_hpc2_0_n54, n_hpc2_0_n53, n_hpc2_0_n52, n_hpc2_0_n51,
         n_hpc2_0_n50, n_hpc2_0_n49, n_hpc2_0_n48, n_hpc2_0_n47, n_hpc2_0_n46,
         n_hpc2_0_n45, n_hpc2_0_n44, n_hpc2_0_n43, n_hpc2_0_n42, n_hpc2_0_n41,
         n_hpc2_0_n40, n_hpc2_0_n39, n_hpc2_0_n38, n_hpc2_0_n37, n_hpc2_0_n36,
         n_hpc2_0_n35, n_hpc2_0_n34, n_hpc2_0_n33, n_hpc2_0_n32, n_hpc2_0_n31,
         n_hpc2_0_n30, n_hpc2_0_n29, n_hpc2_0_n28, n_hpc2_0_n27, n_hpc2_0_n26,
         n_hpc2_0_n25, n_hpc2_0_n24, n_hpc2_0_n23, n_hpc2_0_n22, n_hpc2_0_n21,
         n_hpc2_0_n20, n_hpc2_0_n19, n_hpc2_0_n18, n_hpc2_0_n17, n_hpc2_0_n16,
         n_hpc2_0_n15, n_hpc2_0_n14, n_hpc2_0_n13, n_hpc2_0_n12, n_hpc2_0_n11,
         n_hpc2_0_n10, n_hpc2_0_n9, n_hpc2_0_n8, n_hpc2_0_n7, n_hpc2_0_n6,
         n_hpc2_0_n5, n_hpc2_0_n4, n_hpc2_0_n3, n_hpc2_0_n2, n_hpc2_0_n1,
         n_hpc2_0_N41, n_hpc2_0_N40, n_hpc2_0_N39, n_hpc2_0_N38, n_hpc2_0_N37,
         n_hpc2_0_N36, n_hpc2_0_N35, n_hpc2_0_N34, n_hpc2_0_N33, n_hpc2_0_N32,
         n_hpc2_0_N31, n_hpc2_0_N30, n_hpc2_0_N29, n_hpc2_0_N28, n_hpc2_0_N27,
         n_hpc2_0_N26, n_hpc2_0_N25, n_hpc2_0_N24, n_hpc2_0_N23, n_hpc2_0_N22,
         n_hpc2_0_N21, n_hpc2_0_N20, n_hpc2_0_N19, n_hpc2_0_N18, n_hpc2_0_N17,
         n_hpc2_0_N16, n_hpc2_0_N15, n_hpc2_0_N14, n_hpc2_0_N13, n_hpc2_0_N12,
         n_hpc2_0_N11, n_hpc2_0_N10, n_hpc2_0_N9, n_hpc2_0_N8, n_hpc2_0_N7,
         n_hpc2_0_N6, n_hpc2_0_reg_pipeline_19, n_hpc2_0_reg_pipeline_18,
         n_hpc2_0_reg_pipeline_17, n_hpc2_0_reg_pipeline_16,
         n_hpc2_0_reg_pipeline_15, n_hpc2_0_reg_pipeline_14,
         n_hpc2_0_reg_pipeline_13, n_hpc2_0_reg_pipeline_12,
         n_hpc2_0_reg_pipeline_11, n_hpc2_0_reg_pipeline_10,
         n_hpc2_0_reg_pipeline_9, n_hpc2_0_reg_pipeline_8,
         n_hpc2_0_reg_pipeline_7, n_hpc2_0_reg_pipeline_6,
         n_hpc2_0_reg_pipeline_5, n_hpc2_0_reg_pipeline_4,
         n_hpc2_0_reg_pipeline_3, n_hpc2_0_reg_pipeline_2,
         n_hpc2_0_reg_pipeline_1, n_hpc2_0_reg_pipeline_0,
         n_hpc2_0_reg_pipeline, n_hpc2_0_N5, n_hpc2_0_N4, n_hpc2_0_N3,
         n_hpc2_0_N2, n_hpc2_0_N1, n_hpc2_0_N0, n_hpc2_0__hpc1_z54,
         n_hpc2_0__hpc1_z51, n_hpc2_0__hpc1_z41, n_hpc2_0__hpc1_z44,
         n_hpc2_0__hpc1_z34, n_hpc2_0__hpc1_z31, n_hpc2_0__hpc1_z24,
         n_hpc2_0__hpc1_z21, n_hpc2_0__hpc1_z14, n_hpc2_0__hpc1_z11,
         n_hpc2_0__hpc1_z04, n_hpc2_0__hpc1_z01;

  XOR2_X1 u_hpc2_0_U128 ( .A(io_i1_s0), .B(p_rand_4), .Z(n_hpc2_0_n84) );
  XOR2_X1 u_hpc2_0_U127 ( .A(p_rand_3), .B(n_hpc2_0_n84), .Z(n_hpc2_0_n81) );
  XOR2_X1 u_hpc2_0_U126 ( .A(p_rand_2), .B(p_rand_1), .Z(n_hpc2_0_n83) );
  XOR2_X1 u_hpc2_0_U125 ( .A(p_rand_0), .B(n_hpc2_0_n83), .Z(n_hpc2_0_n82) );
  XOR2_X1 u_hpc2_0_U124 ( .A(n_hpc2_0_n81), .B(n_hpc2_0_n82), .Z(n_hpc2_0_N0)
         );
  XOR2_X1 u_hpc2_0_U123 ( .A(io_i1_s1), .B(p_rand_8), .Z(n_hpc2_0_n80) );
  XOR2_X1 u_hpc2_0_U122 ( .A(p_rand_7), .B(n_hpc2_0_n80), .Z(n_hpc2_0_n77) );
  XOR2_X1 u_hpc2_0_U121 ( .A(p_rand_6), .B(p_rand_5), .Z(n_hpc2_0_n79) );
  XOR2_X1 u_hpc2_0_U120 ( .A(p_rand_0), .B(n_hpc2_0_n79), .Z(n_hpc2_0_n78) );
  XOR2_X1 u_hpc2_0_U119 ( .A(n_hpc2_0_n77), .B(n_hpc2_0_n78), .Z(n_hpc2_0_N1)
         );
  NAND2_X1 u_hpc2_0_U118 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n6), .ZN(
        n_hpc2_0_n76) );
  XNOR2_X1 u_hpc2_0_U117 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n76), .ZN(
        n_hpc2_0_N10) );
  NAND2_X1 u_hpc2_0_U116 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n5), .ZN(
        n_hpc2_0_n75) );
  XNOR2_X1 u_hpc2_0_U115 ( .A(n_hpc2_0_reg_pipeline_4), .B(n_hpc2_0_n75), .ZN(
        n_hpc2_0_N11) );
  NAND2_X1 u_hpc2_0_U114 ( .A1(n_hpc2_0_reg_pipeline_5), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n74) );
  XNOR2_X1 u_hpc2_0_U113 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n74), .ZN(
        n_hpc2_0_N12) );
  AND2_X1 u_hpc2_0_U112 ( .A1(n_hpc2_0_n3), .A2(n_hpc2_0_reg_pipeline_5), .ZN(
        n_hpc2_0_N13) );
  NAND2_X1 u_hpc2_0_U111 ( .A1(n_hpc2_0_reg_pipeline_5), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n73) );
  XNOR2_X1 u_hpc2_0_U110 ( .A(n_hpc2_0_reg_pipeline_6), .B(n_hpc2_0_n73), .ZN(
        n_hpc2_0_N14) );
  NAND2_X1 u_hpc2_0_U109 ( .A1(n_hpc2_0_reg_pipeline_5), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n72) );
  XNOR2_X1 u_hpc2_0_U108 ( .A(n_hpc2_0_reg_pipeline_7), .B(n_hpc2_0_n72), .ZN(
        n_hpc2_0_N15) );
  NAND2_X1 u_hpc2_0_U107 ( .A1(n_hpc2_0_reg_pipeline_5), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n71) );
  XNOR2_X1 u_hpc2_0_U106 ( .A(n_hpc2_0_reg_pipeline_8), .B(n_hpc2_0_n71), .ZN(
        n_hpc2_0_N16) );
  NAND2_X1 u_hpc2_0_U105 ( .A1(n_hpc2_0_reg_pipeline_5), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n70) );
  XNOR2_X1 u_hpc2_0_U104 ( .A(n_hpc2_0_reg_pipeline_9), .B(n_hpc2_0_n70), .ZN(
        n_hpc2_0_N17) );
  NAND2_X1 u_hpc2_0_U103 ( .A1(n_hpc2_0_reg_pipeline_10), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n69) );
  XNOR2_X1 u_hpc2_0_U102 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n69), .ZN(
        n_hpc2_0_N18) );
  NAND2_X1 u_hpc2_0_U101 ( .A1(n_hpc2_0_reg_pipeline_10), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n68) );
  XNOR2_X1 u_hpc2_0_U100 ( .A(n_hpc2_0_reg_pipeline_6), .B(n_hpc2_0_n68), .ZN(
        n_hpc2_0_N19) );
  XOR2_X1 u_hpc2_0_U99 ( .A(io_i1_s2), .B(p_rand_9), .Z(n_hpc2_0_n67) );
  XOR2_X1 u_hpc2_0_U98 ( .A(p_rand_5), .B(n_hpc2_0_n67), .Z(n_hpc2_0_n64) );
  XOR2_X1 u_hpc2_0_U97 ( .A(p_rand_11), .B(p_rand_10), .Z(n_hpc2_0_n66) );
  XOR2_X1 u_hpc2_0_U96 ( .A(p_rand_1), .B(n_hpc2_0_n66), .Z(n_hpc2_0_n65) );
  XOR2_X1 u_hpc2_0_U95 ( .A(n_hpc2_0_n64), .B(n_hpc2_0_n65), .Z(n_hpc2_0_N2)
         );
  AND2_X1 u_hpc2_0_U94 ( .A1(n_hpc2_0_n2), .A2(n_hpc2_0_reg_pipeline_10), .ZN(
        n_hpc2_0_N20) );
  NAND2_X1 u_hpc2_0_U93 ( .A1(n_hpc2_0_reg_pipeline_10), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n63) );
  XNOR2_X1 u_hpc2_0_U92 ( .A(n_hpc2_0_reg_pipeline_11), .B(n_hpc2_0_n63), .ZN(
        n_hpc2_0_N21) );
  NAND2_X1 u_hpc2_0_U91 ( .A1(n_hpc2_0_reg_pipeline_10), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n62) );
  XNOR2_X1 u_hpc2_0_U90 ( .A(n_hpc2_0_reg_pipeline_12), .B(n_hpc2_0_n62), .ZN(
        n_hpc2_0_N22) );
  NAND2_X1 u_hpc2_0_U89 ( .A1(n_hpc2_0_reg_pipeline_10), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n61) );
  XNOR2_X1 u_hpc2_0_U88 ( .A(n_hpc2_0_reg_pipeline_13), .B(n_hpc2_0_n61), .ZN(
        n_hpc2_0_N23) );
  NAND2_X1 u_hpc2_0_U87 ( .A1(n_hpc2_0_reg_pipeline_14), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n60) );
  XNOR2_X1 u_hpc2_0_U86 ( .A(n_hpc2_0_reg_pipeline_2), .B(n_hpc2_0_n60), .ZN(
        n_hpc2_0_N24) );
  NAND2_X1 u_hpc2_0_U85 ( .A1(n_hpc2_0_reg_pipeline_14), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n59) );
  XNOR2_X1 u_hpc2_0_U84 ( .A(n_hpc2_0_reg_pipeline_7), .B(n_hpc2_0_n59), .ZN(
        n_hpc2_0_N25) );
  NAND2_X1 u_hpc2_0_U83 ( .A1(n_hpc2_0_reg_pipeline_14), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n58) );
  XNOR2_X1 u_hpc2_0_U82 ( .A(n_hpc2_0_reg_pipeline_11), .B(n_hpc2_0_n58), .ZN(
        n_hpc2_0_N26) );
  AND2_X1 u_hpc2_0_U81 ( .A1(n_hpc2_0_n1), .A2(n_hpc2_0_reg_pipeline_14), .ZN(
        n_hpc2_0_N27) );
  NAND2_X1 u_hpc2_0_U80 ( .A1(n_hpc2_0_reg_pipeline_14), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n57) );
  XNOR2_X1 u_hpc2_0_U79 ( .A(n_hpc2_0_reg_pipeline_15), .B(n_hpc2_0_n57), .ZN(
        n_hpc2_0_N28) );
  NAND2_X1 u_hpc2_0_U78 ( .A1(n_hpc2_0_reg_pipeline_14), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n56) );
  XNOR2_X1 u_hpc2_0_U77 ( .A(n_hpc2_0_reg_pipeline_16), .B(n_hpc2_0_n56), .ZN(
        n_hpc2_0_N29) );
  XOR2_X1 u_hpc2_0_U76 ( .A(io_i1_s3), .B(p_rand_9), .Z(n_hpc2_0_n55) );
  XOR2_X1 u_hpc2_0_U75 ( .A(p_rand_6), .B(n_hpc2_0_n55), .Z(n_hpc2_0_n52) );
  XOR2_X1 u_hpc2_0_U74 ( .A(p_rand_2), .B(p_rand_13), .Z(n_hpc2_0_n54) );
  XOR2_X1 u_hpc2_0_U73 ( .A(p_rand_12), .B(n_hpc2_0_n54), .Z(n_hpc2_0_n53) );
  XOR2_X1 u_hpc2_0_U72 ( .A(n_hpc2_0_n52), .B(n_hpc2_0_n53), .Z(n_hpc2_0_N3)
         );
  NAND2_X1 u_hpc2_0_U71 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n51) );
  XNOR2_X1 u_hpc2_0_U70 ( .A(n_hpc2_0_reg_pipeline_3), .B(n_hpc2_0_n51), .ZN(
        n_hpc2_0_N30) );
  NAND2_X1 u_hpc2_0_U69 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n50) );
  XNOR2_X1 u_hpc2_0_U68 ( .A(n_hpc2_0_reg_pipeline_8), .B(n_hpc2_0_n50), .ZN(
        n_hpc2_0_N31) );
  NAND2_X1 u_hpc2_0_U67 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n49) );
  XNOR2_X1 u_hpc2_0_U66 ( .A(n_hpc2_0_reg_pipeline_12), .B(n_hpc2_0_n49), .ZN(
        n_hpc2_0_N32) );
  NAND2_X1 u_hpc2_0_U65 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n48) );
  XNOR2_X1 u_hpc2_0_U64 ( .A(n_hpc2_0_reg_pipeline_15), .B(n_hpc2_0_n48), .ZN(
        n_hpc2_0_N33) );
  AND2_X1 u_hpc2_0_U63 ( .A1(n_hpc2_0_n6), .A2(n_hpc2_0_reg_pipeline_17), .ZN(
        n_hpc2_0_N34) );
  NAND2_X1 u_hpc2_0_U62 ( .A1(n_hpc2_0_reg_pipeline_17), .A2(n_hpc2_0_n5), 
        .ZN(n_hpc2_0_n47) );
  XNOR2_X1 u_hpc2_0_U61 ( .A(n_hpc2_0_reg_pipeline_18), .B(n_hpc2_0_n47), .ZN(
        n_hpc2_0_N35) );
  NAND2_X1 u_hpc2_0_U60 ( .A1(n_hpc2_0_reg_pipeline_19), .A2(n_hpc2_0_n4), 
        .ZN(n_hpc2_0_n46) );
  XNOR2_X1 u_hpc2_0_U59 ( .A(n_hpc2_0_reg_pipeline_4), .B(n_hpc2_0_n46), .ZN(
        n_hpc2_0_N36) );
  NAND2_X1 u_hpc2_0_U58 ( .A1(n_hpc2_0_reg_pipeline_19), .A2(n_hpc2_0_n3), 
        .ZN(n_hpc2_0_n45) );
  XNOR2_X1 u_hpc2_0_U57 ( .A(n_hpc2_0_reg_pipeline_9), .B(n_hpc2_0_n45), .ZN(
        n_hpc2_0_N37) );
  NAND2_X1 u_hpc2_0_U56 ( .A1(n_hpc2_0_reg_pipeline_19), .A2(n_hpc2_0_n2), 
        .ZN(n_hpc2_0_n44) );
  XNOR2_X1 u_hpc2_0_U55 ( .A(n_hpc2_0_reg_pipeline_13), .B(n_hpc2_0_n44), .ZN(
        n_hpc2_0_N38) );
  NAND2_X1 u_hpc2_0_U54 ( .A1(n_hpc2_0_reg_pipeline_19), .A2(n_hpc2_0_n1), 
        .ZN(n_hpc2_0_n43) );
  XNOR2_X1 u_hpc2_0_U53 ( .A(n_hpc2_0_reg_pipeline_16), .B(n_hpc2_0_n43), .ZN(
        n_hpc2_0_N39) );
  XOR2_X1 u_hpc2_0_U52 ( .A(io_i1_s4), .B(p_rand_7), .Z(n_hpc2_0_n42) );
  XOR2_X1 u_hpc2_0_U51 ( .A(p_rand_3), .B(n_hpc2_0_n42), .Z(n_hpc2_0_n39) );
  XOR2_X1 u_hpc2_0_U50 ( .A(p_rand_14), .B(p_rand_12), .Z(n_hpc2_0_n41) );
  XOR2_X1 u_hpc2_0_U49 ( .A(p_rand_10), .B(n_hpc2_0_n41), .Z(n_hpc2_0_n40) );
  XOR2_X1 u_hpc2_0_U48 ( .A(n_hpc2_0_n39), .B(n_hpc2_0_n40), .Z(n_hpc2_0_N4)
         );
  NAND2_X1 u_hpc2_0_U47 ( .A1(n_hpc2_0_reg_pipeline_19), .A2(n_hpc2_0_n6), 
        .ZN(n_hpc2_0_n38) );
  XNOR2_X1 u_hpc2_0_U46 ( .A(n_hpc2_0_reg_pipeline_18), .B(n_hpc2_0_n38), .ZN(
        n_hpc2_0_N40) );
  AND2_X1 u_hpc2_0_U45 ( .A1(n_hpc2_0_n5), .A2(n_hpc2_0_reg_pipeline_19), .ZN(
        n_hpc2_0_N41) );
  XOR2_X1 u_hpc2_0_U44 ( .A(io_i1_s5), .B(p_rand_8), .Z(n_hpc2_0_n37) );
  XOR2_X1 u_hpc2_0_U43 ( .A(p_rand_4), .B(n_hpc2_0_n37), .Z(n_hpc2_0_n34) );
  XOR2_X1 u_hpc2_0_U42 ( .A(p_rand_14), .B(p_rand_13), .Z(n_hpc2_0_n36) );
  XOR2_X1 u_hpc2_0_U41 ( .A(p_rand_11), .B(n_hpc2_0_n36), .Z(n_hpc2_0_n35) );
  XOR2_X1 u_hpc2_0_U40 ( .A(n_hpc2_0_n34), .B(n_hpc2_0_n35), .Z(n_hpc2_0_N5)
         );
  AND2_X1 u_hpc2_0_U39 ( .A1(n_hpc2_0_n4), .A2(n_hpc2_0_reg_pipeline), .ZN(
        n_hpc2_0_N6) );
  NAND2_X1 u_hpc2_0_U38 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n3), .ZN(
        n_hpc2_0_n33) );
  XNOR2_X1 u_hpc2_0_U37 ( .A(n_hpc2_0_reg_pipeline_0), .B(n_hpc2_0_n33), .ZN(
        n_hpc2_0_N7) );
  NAND2_X1 u_hpc2_0_U36 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n2), .ZN(
        n_hpc2_0_n32) );
  XNOR2_X1 u_hpc2_0_U35 ( .A(n_hpc2_0_reg_pipeline_1), .B(n_hpc2_0_n32), .ZN(
        n_hpc2_0_N8) );
  NAND2_X1 u_hpc2_0_U34 ( .A1(n_hpc2_0_reg_pipeline), .A2(n_hpc2_0_n1), .ZN(
        n_hpc2_0_n31) );
  XNOR2_X1 u_hpc2_0_U33 ( .A(n_hpc2_0_reg_pipeline_2), .B(n_hpc2_0_n31), .ZN(
        n_hpc2_0_N9) );
  XOR2_X1 u_hpc2_0_U32 ( .A(n_hpc2_0__hpc1_z01), .B(n_hpc2_0_n105), .Z(
        n_hpc2_0_n30) );
  XOR2_X1 u_hpc2_0_U31 ( .A(n_hpc2_0_n30), .B(n_hpc2_0_n106), .Z(n_hpc2_0_n27)
         );
  XOR2_X1 u_hpc2_0_U30 ( .A(n_hpc2_0__hpc1_z04), .B(n_hpc2_0_n107), .Z(
        n_hpc2_0_n29) );
  XOR2_X1 u_hpc2_0_U29 ( .A(n_hpc2_0_n29), .B(n_hpc2_0_n108), .Z(n_hpc2_0_n28)
         );
  XOR2_X1 u_hpc2_0_U28 ( .A(n_hpc2_0_n27), .B(n_hpc2_0_n28), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U27 ( .A(n_hpc2_0__hpc1_z11), .B(n_hpc2_0_n101), .Z(
        n_hpc2_0_n26) );
  XOR2_X1 u_hpc2_0_U26 ( .A(n_hpc2_0_n26), .B(n_hpc2_0_n102), .Z(n_hpc2_0_n23)
         );
  XOR2_X1 u_hpc2_0_U25 ( .A(n_hpc2_0__hpc1_z14), .B(n_hpc2_0_n103), .Z(
        n_hpc2_0_n25) );
  XOR2_X1 u_hpc2_0_U24 ( .A(n_hpc2_0_n25), .B(n_hpc2_0_n104), .Z(n_hpc2_0_n24)
         );
  XOR2_X1 u_hpc2_0_U23 ( .A(n_hpc2_0_n23), .B(n_hpc2_0_n24), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U22 ( .A(n_hpc2_0__hpc1_z21), .B(n_hpc2_0_n97), .Z(
        n_hpc2_0_n22) );
  XOR2_X1 u_hpc2_0_U21 ( .A(n_hpc2_0_n22), .B(n_hpc2_0_n98), .Z(n_hpc2_0_n19)
         );
  XOR2_X1 u_hpc2_0_U20 ( .A(n_hpc2_0__hpc1_z24), .B(n_hpc2_0_n99), .Z(
        n_hpc2_0_n21) );
  XOR2_X1 u_hpc2_0_U19 ( .A(n_hpc2_0_n21), .B(n_hpc2_0_n100), .Z(n_hpc2_0_n20)
         );
  XOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0_n19), .B(n_hpc2_0_n20), .Z(io_o0_s2) );
  XOR2_X1 u_hpc2_0_U17 ( .A(n_hpc2_0__hpc1_z31), .B(n_hpc2_0_n93), .Z(
        n_hpc2_0_n18) );
  XOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_n18), .B(n_hpc2_0_n94), .Z(n_hpc2_0_n15)
         );
  XOR2_X1 u_hpc2_0_U15 ( .A(n_hpc2_0__hpc1_z34), .B(n_hpc2_0_n95), .Z(
        n_hpc2_0_n17) );
  XOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0_n17), .B(n_hpc2_0_n96), .Z(n_hpc2_0_n16)
         );
  XOR2_X1 u_hpc2_0_U13 ( .A(n_hpc2_0_n15), .B(n_hpc2_0_n16), .Z(io_o0_s3) );
  XOR2_X1 u_hpc2_0_U12 ( .A(n_hpc2_0__hpc1_z41), .B(n_hpc2_0_n89), .Z(
        n_hpc2_0_n14) );
  XOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_n14), .B(n_hpc2_0_n90), .Z(n_hpc2_0_n11)
         );
  XOR2_X1 u_hpc2_0_U10 ( .A(n_hpc2_0__hpc1_z44), .B(n_hpc2_0_n91), .Z(
        n_hpc2_0_n13) );
  XOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_n13), .B(n_hpc2_0_n92), .Z(n_hpc2_0_n12)
         );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0_n11), .B(n_hpc2_0_n12), .Z(io_o0_s4) );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0__hpc1_z51), .B(n_hpc2_0_n85), .Z(
        n_hpc2_0_n10) );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0_n10), .B(n_hpc2_0_n86), .Z(n_hpc2_0_n7) );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0__hpc1_z54), .B(n_hpc2_0_n87), .Z(
        n_hpc2_0_n9) );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0_n9), .B(n_hpc2_0_n88), .Z(n_hpc2_0_n8) );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n7), .B(n_hpc2_0_n8), .Z(io_o0_s5) );
  DFF_X1 u_hpc2_0__hpc1_z45_reg ( .D(n_hpc2_0_N35), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n92) );
  DFF_X1 u_hpc2_0__hpc1_z44_reg ( .D(n_hpc2_0_N34), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z44), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z43_reg ( .D(n_hpc2_0_N33), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n91) );
  DFF_X1 u_hpc2_0__hpc1_z42_reg ( .D(n_hpc2_0_N32), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n90) );
  DFF_X1 u_hpc2_0__hpc1_z41_reg ( .D(n_hpc2_0_N31), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z41), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z40_reg ( .D(n_hpc2_0_N30), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n89) );
  DFF_X1 u_hpc2_0__hpc1_z35_reg ( .D(n_hpc2_0_N29), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n96) );
  DFF_X1 u_hpc2_0__hpc1_z34_reg ( .D(n_hpc2_0_N28), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z34), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z33_reg ( .D(n_hpc2_0_N27), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n95) );
  DFF_X1 u_hpc2_0__hpc1_z32_reg ( .D(n_hpc2_0_N26), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n94) );
  DFF_X1 u_hpc2_0__hpc1_z31_reg ( .D(n_hpc2_0_N25), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z31), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z30_reg ( .D(n_hpc2_0_N24), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n93) );
  DFF_X1 u_hpc2_0__hpc1_z25_reg ( .D(n_hpc2_0_N23), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n100) );
  DFF_X1 u_hpc2_0__hpc1_z24_reg ( .D(n_hpc2_0_N22), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z24), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z23_reg ( .D(n_hpc2_0_N21), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n99) );
  DFF_X1 u_hpc2_0__hpc1_z22_reg ( .D(n_hpc2_0_N20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n98) );
  DFF_X1 u_hpc2_0__hpc1_z21_reg ( .D(n_hpc2_0_N19), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z21), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z20_reg ( .D(n_hpc2_0_N18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n97) );
  DFF_X1 u_hpc2_0__hpc1_z15_reg ( .D(n_hpc2_0_N17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n104) );
  DFF_X1 u_hpc2_0__hpc1_z14_reg ( .D(n_hpc2_0_N16), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z14), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z13_reg ( .D(n_hpc2_0_N15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n103) );
  DFF_X1 u_hpc2_0__hpc1_z12_reg ( .D(n_hpc2_0_N14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n102) );
  DFF_X1 u_hpc2_0__hpc1_z11_reg ( .D(n_hpc2_0_N13), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z11), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z10_reg ( .D(n_hpc2_0_N12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n101) );
  DFF_X1 u_hpc2_0__hpc1_z05_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n108) );
  DFF_X1 u_hpc2_0__hpc1_z04_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z04), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z03_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n107) );
  DFF_X1 u_hpc2_0__hpc1_z02_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n106) );
  DFF_X1 u_hpc2_0__hpc1_z01_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z01), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z00_reg ( .D(n_hpc2_0_N6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n105) );
  DFF_X1 u_hpc2_0__hpc1_z54_reg ( .D(n_hpc2_0_N40), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z54), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_18_reg ( .D(p_rand_29), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_18), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(io_i0_s0), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_5_reg ( .D(io_i0_s1), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_5), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(p_rand_16), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_1), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z51_reg ( .D(n_hpc2_0_N37), .CK(clock_0), .Q(
        n_hpc2_0__hpc1_z51), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_9_reg ( .D(p_rand_23), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_9), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_11_reg ( .D(p_rand_24), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_11), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z53_reg ( .D(n_hpc2_0_N39), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n87) );
  DFF_X1 u_hpc2_0__hpc1_ref_v3_reg ( .D(n_hpc2_0_N3), .CK(clock_0), .Q(
        n_hpc2_0_n1), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z52_reg ( .D(n_hpc2_0_N38), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n86) );
  DFF_X1 u_hpc2_0_reg_pipeline_13_reg ( .D(p_rand_26), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_13), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v1_reg ( .D(n_hpc2_0_N1), .CK(clock_0), .Q(
        n_hpc2_0_n3), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_15_reg ( .D(p_rand_27), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_15), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_17_reg ( .D(io_i0_s4), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_17), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z50_reg ( .D(n_hpc2_0_N36), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n85) );
  DFF_X1 u_hpc2_0__hpc1_ref_v0_reg ( .D(n_hpc2_0_N0), .CK(clock_0), .Q(
        n_hpc2_0_n4), .QN() );
  DFF_X1 u_hpc2_0__hpc1_z55_reg ( .D(n_hpc2_0_N41), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n88) );
  DFF_X1 u_hpc2_0_reg_pipeline_16_reg ( .D(p_rand_28), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_16), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(p_rand_19), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_4), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_14_reg ( .D(io_i0_s3), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_14), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_8_reg ( .D(p_rand_22), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_8), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(p_rand_18), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_3), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_12_reg ( .D(p_rand_25), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_12), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v4_reg ( .D(n_hpc2_0_N4), .CK(clock_0), .Q(
        n_hpc2_0_n6), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_7_reg ( .D(p_rand_21), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_7), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(p_rand_17), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_2), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_10_reg ( .D(io_i0_s2), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_10), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v2_reg ( .D(n_hpc2_0_N2), .CK(clock_0), .Q(
        n_hpc2_0_n2), .QN() );
  DFF_X1 u_hpc2_0__hpc1_ref_v5_reg ( .D(n_hpc2_0_N5), .CK(clock_0), .Q(
        n_hpc2_0_n5), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_6_reg ( .D(p_rand_20), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_6), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_19_reg ( .D(io_i0_s5), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_19), .QN() );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(p_rand_15), .CK(clock_0), .Q(
        n_hpc2_0_reg_pipeline_0), .QN() );
endmodule

