
module keccak_b25_r10_i1_o1 ( clock, reset, io_block_i0, io_block_o0 );
  input [9:0] io_block_i0;
  output [9:0] io_block_o0;
  input clock, reset;
  wire   n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320;

  XOR2_X1 U1166 ( .A(n1156), .B(n1157), .Z(io_block_o0[9]) );
  NAND2_X1 U1167 ( .A1(n1158), .A2(n1159), .ZN(n1156) );
  XOR2_X1 U1168 ( .A(n1160), .B(n1161), .Z(io_block_o0[8]) );
  NAND2_X1 U1169 ( .A1(n1158), .A2(n1157), .ZN(n1160) );
  XOR2_X1 U1170 ( .A(n1162), .B(n1163), .Z(io_block_o0[7]) );
  NAND2_X1 U1171 ( .A1(n1161), .A2(n1157), .ZN(n1162) );
  XNOR2_X1 U1172 ( .A(n1164), .B(n1165), .ZN(n1157) );
  XOR2_X1 U1173 ( .A(n1166), .B(n1159), .Z(io_block_o0[6]) );
  NAND2_X1 U1174 ( .A1(n1163), .A2(n1161), .ZN(n1166) );
  XOR2_X1 U1175 ( .A(n1167), .B(n1168), .Z(n1161) );
  XOR2_X1 U1176 ( .A(n1169), .B(n1158), .Z(io_block_o0[5]) );
  XNOR2_X1 U1177 ( .A(n1170), .B(n1171), .ZN(n1158) );
  NAND2_X1 U1178 ( .A1(n1163), .A2(n1159), .ZN(n1169) );
  XOR2_X1 U1179 ( .A(n1172), .B(n1173), .Z(n1159) );
  XNOR2_X1 U1180 ( .A(n1174), .B(n1175), .ZN(n1163) );
  XOR2_X1 U1181 ( .A(n1176), .B(n1177), .Z(io_block_o0[4]) );
  NAND2_X1 U1182 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
  XOR2_X1 U1183 ( .A(n1180), .B(n1181), .Z(io_block_o0[3]) );
  NAND2_X1 U1184 ( .A1(n1177), .A2(n1179), .ZN(n1180) );
  XOR2_X1 U1185 ( .A(n1182), .B(n1183), .Z(io_block_o0[2]) );
  NAND2_X1 U1186 ( .A1(n1181), .A2(n1177), .ZN(n1182) );
  XNOR2_X1 U1187 ( .A(n1172), .B(n1184), .ZN(n1177) );
  XNOR2_X1 U1188 ( .A(n1185), .B(n1186), .ZN(n1172) );
  XOR2_X1 U1189 ( .A(n1187), .B(n1178), .Z(io_block_o0[1]) );
  NAND2_X1 U1190 ( .A1(n1183), .A2(n1181), .ZN(n1187) );
  XNOR2_X1 U1191 ( .A(n1170), .B(n1188), .ZN(n1181) );
  XOR2_X1 U1192 ( .A(n1189), .B(n1190), .Z(n1170) );
  XOR2_X1 U1193 ( .A(n1191), .B(n1179), .Z(io_block_o0[0]) );
  XOR2_X1 U1194 ( .A(n1174), .B(n1192), .Z(n1179) );
  XOR2_X1 U1195 ( .A(n1193), .B(n1190), .Z(n1174) );
  XNOR2_X1 U1196 ( .A(n1194), .B(n1195), .ZN(n1190) );
  XOR2_X1 U1197 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR2_X1 U1198 ( .A(n1198), .B(n1199), .Z(n1197) );
  NAND2_X1 U1199 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
  XOR2_X1 U1200 ( .A(n1202), .B(n1203), .Z(n1196) );
  XOR2_X1 U1201 ( .A(n1204), .B(n1205), .Z(n1194) );
  XOR2_X1 U1202 ( .A(n1206), .B(n1207), .Z(n1205) );
  XNOR2_X1 U1203 ( .A(n1184), .B(n1173), .ZN(n1204) );
  XNOR2_X1 U1204 ( .A(n1208), .B(n1209), .ZN(n1173) );
  NAND2_X1 U1205 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
  INV_X1 U1206 ( .A(n1212), .ZN(n1210) );
  XNOR2_X1 U1207 ( .A(n1213), .B(n1214), .ZN(n1184) );
  OR2_X1 U1208 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
  NAND2_X1 U1209 ( .A1(n1183), .A2(n1178), .ZN(n1191) );
  XNOR2_X1 U1210 ( .A(n1167), .B(n1217), .ZN(n1178) );
  XOR2_X1 U1211 ( .A(n1189), .B(n1185), .Z(n1167) );
  XNOR2_X1 U1212 ( .A(n1218), .B(n1219), .ZN(n1185) );
  XOR2_X1 U1213 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR2_X1 U1214 ( .A(n1215), .B(n1201), .Z(n1221) );
  XNOR2_X1 U1215 ( .A(n1222), .B(n1211), .ZN(n1220) );
  NAND2_X1 U1216 ( .A1(n1200), .A2(n1223), .ZN(n1222) );
  XOR2_X1 U1217 ( .A(n1224), .B(n1225), .Z(n1218) );
  XNOR2_X1 U1218 ( .A(n1226), .B(n1192), .ZN(n1225) );
  NAND2_X1 U1219 ( .A1(n1227), .A2(n1228), .ZN(n1192) );
  NAND2_X1 U1220 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
  NAND2_X1 U1221 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
  INV_X1 U1222 ( .A(n1233), .ZN(n1231) );
  NAND2_X1 U1223 ( .A1(n1202), .A2(n1232), .ZN(n1227) );
  NOR2_X1 U1224 ( .A1(n1233), .A2(n1229), .ZN(n1202) );
  XOR2_X1 U1225 ( .A(n1175), .B(n1234), .Z(n1224) );
  NOR2_X1 U1226 ( .A1(n1216), .A2(n1235), .ZN(n1234) );
  NAND2_X1 U1227 ( .A1(n1236), .A2(n1237), .ZN(n1175) );
  NAND2_X1 U1228 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
  OR2_X1 U1229 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
  NAND2_X1 U1230 ( .A1(n1203), .A2(n1242), .ZN(n1236) );
  NOR2_X1 U1231 ( .A1(n1238), .A2(n1240), .ZN(n1203) );
  XOR2_X1 U1232 ( .A(n1243), .B(n1244), .Z(n1189) );
  XOR2_X1 U1233 ( .A(n1245), .B(n1246), .Z(n1244) );
  XNOR2_X1 U1234 ( .A(n1247), .B(n1248), .ZN(n1246) );
  AND2_X1 U1235 ( .A1(n1207), .A2(n1249), .ZN(n1248) );
  XNOR2_X1 U1236 ( .A(n1250), .B(n1251), .ZN(n1245) );
  AND2_X1 U1237 ( .A1(n1209), .A2(n1252), .ZN(n1251) );
  XOR2_X1 U1238 ( .A(n1253), .B(n1254), .Z(n1243) );
  XNOR2_X1 U1239 ( .A(n1255), .B(n1223), .ZN(n1254) );
  XNOR2_X1 U1240 ( .A(n1165), .B(n1232), .ZN(n1253) );
  XOR2_X1 U1241 ( .A(n1256), .B(n1235), .Z(n1165) );
  OR2_X1 U1242 ( .A1(n1257), .A2(n1214), .ZN(n1256) );
  XNOR2_X1 U1243 ( .A(n1164), .B(n1247), .ZN(n1183) );
  AND2_X1 U1244 ( .A1(n1258), .A2(n1259), .ZN(n1247) );
  NAND2_X1 U1245 ( .A1(n1241), .A2(n1260), .ZN(n1259) );
  NAND2_X1 U1246 ( .A1(n1261), .A2(n1206), .ZN(n1260) );
  INV_X1 U1247 ( .A(n1242), .ZN(n1241) );
  NAND2_X1 U1248 ( .A1(n1262), .A2(n1206), .ZN(n1258) );
  XOR2_X1 U1249 ( .A(n1193), .B(n1186), .Z(n1164) );
  XNOR2_X1 U1250 ( .A(n1263), .B(n1264), .ZN(n1186) );
  XOR2_X1 U1251 ( .A(n1265), .B(n1266), .Z(n1264) );
  XNOR2_X1 U1252 ( .A(n1252), .B(n1261), .ZN(n1266) );
  XNOR2_X1 U1253 ( .A(n1188), .B(n1257), .ZN(n1265) );
  XOR2_X1 U1254 ( .A(n1267), .B(n1249), .Z(n1188) );
  NAND2_X1 U1255 ( .A1(n1207), .A2(n1201), .ZN(n1267) );
  XNOR2_X1 U1256 ( .A(n1268), .B(n1269), .ZN(n1201) );
  XOR2_X1 U1257 ( .A(n1270), .B(n1271), .Z(n1207) );
  XOR2_X1 U1258 ( .A(n1272), .B(n1273), .Z(n1263) );
  XOR2_X1 U1259 ( .A(n1171), .B(n1274), .Z(n1273) );
  NAND2_X1 U1260 ( .A1(n1209), .A2(n1211), .ZN(n1274) );
  XNOR2_X1 U1261 ( .A(n1270), .B(n1275), .ZN(n1211) );
  XNOR2_X1 U1262 ( .A(n1276), .B(n1277), .ZN(n1209) );
  NAND2_X1 U1263 ( .A1(n1278), .A2(n1279), .ZN(n1171) );
  NAND2_X1 U1264 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
  OR2_X1 U1265 ( .A1(n1229), .A2(n1199), .ZN(n1281) );
  INV_X1 U1266 ( .A(n1282), .ZN(n1229) );
  NAND2_X1 U1267 ( .A1(n1250), .A2(n1282), .ZN(n1278) );
  XNOR2_X1 U1268 ( .A(n1283), .B(n1284), .ZN(n1282) );
  NOR2_X1 U1269 ( .A1(n1280), .A2(n1199), .ZN(n1250) );
  XOR2_X1 U1270 ( .A(n1268), .B(n1285), .Z(n1199) );
  INV_X1 U1271 ( .A(n1286), .ZN(n1280) );
  XOR2_X1 U1272 ( .A(n1287), .B(n1288), .Z(n1272) );
  NOR2_X1 U1273 ( .A1(n1215), .A2(n1214), .ZN(n1288) );
  XNOR2_X1 U1274 ( .A(n1289), .B(n1290), .ZN(n1214) );
  XNOR2_X1 U1275 ( .A(n1276), .B(n1291), .ZN(n1215) );
  NAND2_X1 U1276 ( .A1(n1206), .A2(n1292), .ZN(n1287) );
  INV_X1 U1277 ( .A(n1238), .ZN(n1292) );
  XNOR2_X1 U1278 ( .A(n1289), .B(n1293), .ZN(n1238) );
  XOR2_X1 U1279 ( .A(n1283), .B(n1294), .Z(n1206) );
  XOR2_X1 U1280 ( .A(n1295), .B(n1296), .Z(n1193) );
  XOR2_X1 U1281 ( .A(n1297), .B(n1298), .Z(n1296) );
  XNOR2_X1 U1282 ( .A(n1262), .B(n1299), .ZN(n1298) );
  NOR2_X1 U1283 ( .A1(n1235), .A2(n1257), .ZN(n1299) );
  XOR2_X1 U1284 ( .A(n1283), .B(n1300), .Z(n1257) );
  INV_X1 U1285 ( .A(n1301), .ZN(n1300) );
  XOR2_X1 U1286 ( .A(n1268), .B(n1302), .Z(n1235) );
  AND2_X1 U1287 ( .A1(n1261), .A2(n1242), .ZN(n1262) );
  XNOR2_X1 U1288 ( .A(n1270), .B(n1303), .ZN(n1242) );
  XOR2_X1 U1289 ( .A(n1268), .B(n1304), .Z(n1261) );
  XOR2_X1 U1290 ( .A(n1305), .B(n1217), .Z(n1297) );
  AND2_X1 U1291 ( .A1(n1306), .A2(n1307), .ZN(n1217) );
  NAND2_X1 U1292 ( .A1(n1212), .A2(n1308), .ZN(n1307) );
  NAND2_X1 U1293 ( .A1(n1255), .A2(n1252), .ZN(n1308) );
  INV_X1 U1294 ( .A(n1309), .ZN(n1255) );
  NAND2_X1 U1295 ( .A1(n1226), .A2(n1252), .ZN(n1306) );
  XOR2_X1 U1296 ( .A(n1289), .B(n1310), .Z(n1252) );
  NOR2_X1 U1297 ( .A1(n1309), .A2(n1212), .ZN(n1226) );
  XNOR2_X1 U1298 ( .A(n1268), .B(n1311), .ZN(n1212) );
  XOR2_X1 U1299 ( .A(n1312), .B(n1313), .Z(n1268) );
  XNOR2_X1 U1300 ( .A(n1283), .B(n1314), .ZN(n1309) );
  NAND2_X1 U1301 ( .A1(n1232), .A2(n1286), .ZN(n1305) );
  XNOR2_X1 U1302 ( .A(n1270), .B(n1315), .ZN(n1286) );
  XNOR2_X1 U1303 ( .A(n1276), .B(n1316), .ZN(n1232) );
  XOR2_X1 U1304 ( .A(n1317), .B(n1318), .Z(n1295) );
  XNOR2_X1 U1305 ( .A(n1216), .B(n1233), .ZN(n1318) );
  XNOR2_X1 U1306 ( .A(n1289), .B(n1319), .ZN(n1233) );
  XOR2_X1 U1307 ( .A(n1270), .B(n1320), .Z(n1216) );
  XNOR2_X1 U1308 ( .A(n1321), .B(n1322), .ZN(n1270) );
  XNOR2_X1 U1309 ( .A(n1168), .B(n1240), .ZN(n1317) );
  XNOR2_X1 U1310 ( .A(n1276), .B(n1323), .ZN(n1240) );
  XOR2_X1 U1311 ( .A(n1324), .B(n1200), .Z(n1168) );
  XOR2_X1 U1312 ( .A(n1283), .B(n1325), .Z(n1200) );
  XNOR2_X1 U1313 ( .A(n1326), .B(n1321), .ZN(n1283) );
  XNOR2_X1 U1314 ( .A(n1327), .B(n1328), .ZN(n1321) );
  XOR2_X1 U1315 ( .A(n1311), .B(n1304), .Z(n1328) );
  XOR2_X1 U1316 ( .A(n1329), .B(n1330), .Z(n1304) );
  NAND2_X1 U1317 ( .A1(n1331), .A2(n1332), .ZN(n1329) );
  XOR2_X1 U1318 ( .A(n1333), .B(n1334), .Z(n1311) );
  NAND2_X1 U1319 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
  XOR2_X1 U1320 ( .A(n1337), .B(n1285), .Z(n1327) );
  XNOR2_X1 U1321 ( .A(n1338), .B(n1339), .ZN(n1285) );
  NAND2_X1 U1322 ( .A1(n1340), .A2(n1341), .ZN(n1338) );
  XNOR2_X1 U1323 ( .A(n1302), .B(n1269), .ZN(n1337) );
  XNOR2_X1 U1324 ( .A(n1342), .B(n1343), .ZN(n1269) );
  NAND2_X1 U1325 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
  XNOR2_X1 U1326 ( .A(n1346), .B(n1347), .ZN(n1302) );
  NAND2_X1 U1327 ( .A1(n1348), .A2(n1349), .ZN(n1346) );
  NAND2_X1 U1328 ( .A1(n1249), .A2(n1223), .ZN(n1324) );
  XNOR2_X1 U1329 ( .A(n1289), .B(n1350), .ZN(n1223) );
  XNOR2_X1 U1330 ( .A(n1322), .B(n1313), .ZN(n1289) );
  XNOR2_X1 U1331 ( .A(n1351), .B(n1352), .ZN(n1313) );
  XOR2_X1 U1332 ( .A(n1314), .B(n1284), .Z(n1352) );
  XOR2_X1 U1333 ( .A(n1353), .B(n1345), .Z(n1284) );
  NAND2_X1 U1334 ( .A1(n1344), .A2(n1354), .ZN(n1353) );
  XNOR2_X1 U1335 ( .A(n1355), .B(n1349), .ZN(n1314) );
  NAND2_X1 U1336 ( .A1(n1356), .A2(n1348), .ZN(n1355) );
  XOR2_X1 U1337 ( .A(n1357), .B(n1325), .Z(n1351) );
  XNOR2_X1 U1338 ( .A(n1358), .B(n1336), .ZN(n1325) );
  NAND2_X1 U1339 ( .A1(n1335), .A2(n1359), .ZN(n1358) );
  XNOR2_X1 U1340 ( .A(n1301), .B(n1294), .ZN(n1357) );
  XNOR2_X1 U1341 ( .A(n1360), .B(n1341), .ZN(n1294) );
  NAND2_X1 U1342 ( .A1(n1340), .A2(n1361), .ZN(n1360) );
  XNOR2_X1 U1343 ( .A(n1362), .B(n1332), .ZN(n1301) );
  NAND2_X1 U1344 ( .A1(n1331), .A2(n1363), .ZN(n1362) );
  XNOR2_X1 U1345 ( .A(n1364), .B(n1365), .ZN(n1322) );
  XOR2_X1 U1346 ( .A(n1323), .B(n1316), .Z(n1365) );
  XOR2_X1 U1347 ( .A(n1366), .B(n1356), .Z(n1316) );
  NAND2_X1 U1348 ( .A1(n1367), .A2(n1347), .ZN(n1366) );
  XNOR2_X1 U1349 ( .A(n1368), .B(n1359), .ZN(n1323) );
  NAND2_X1 U1350 ( .A1(n1369), .A2(n1334), .ZN(n1368) );
  XOR2_X1 U1351 ( .A(n1370), .B(n1291), .Z(n1364) );
  XNOR2_X1 U1352 ( .A(n1371), .B(n1354), .ZN(n1291) );
  NAND2_X1 U1353 ( .A1(n1372), .A2(n1343), .ZN(n1371) );
  XNOR2_X1 U1354 ( .A(n1277), .B(n1373), .ZN(n1370) );
  XOR2_X1 U1355 ( .A(n1374), .B(n1361), .Z(n1277) );
  NAND2_X1 U1356 ( .A1(n1375), .A2(n1339), .ZN(n1374) );
  XOR2_X1 U1357 ( .A(n1276), .B(n1373), .Z(n1249) );
  XNOR2_X1 U1358 ( .A(n1376), .B(n1363), .ZN(n1373) );
  NAND2_X1 U1359 ( .A1(n1377), .A2(n1330), .ZN(n1376) );
  XOR2_X1 U1360 ( .A(n1312), .B(n1326), .Z(n1276) );
  XNOR2_X1 U1361 ( .A(n1378), .B(n1379), .ZN(n1326) );
  XOR2_X1 U1362 ( .A(n1319), .B(n1350), .Z(n1379) );
  XNOR2_X1 U1363 ( .A(n1380), .B(n1348), .ZN(n1350) );
  XNOR2_X1 U1364 ( .A(n1381), .B(n1382), .ZN(n1348) );
  NAND2_X1 U1365 ( .A1(n1356), .A2(n1367), .ZN(n1380) );
  XOR2_X1 U1366 ( .A(n1383), .B(n1384), .Z(n1356) );
  XOR2_X1 U1367 ( .A(n1385), .B(n1335), .Z(n1319) );
  XOR2_X1 U1368 ( .A(n1386), .B(n1387), .Z(n1335) );
  NAND2_X1 U1369 ( .A1(n1369), .A2(n1359), .ZN(n1385) );
  XNOR2_X1 U1370 ( .A(n1388), .B(n1389), .ZN(n1359) );
  XOR2_X1 U1371 ( .A(n1390), .B(n1310), .Z(n1378) );
  XOR2_X1 U1372 ( .A(n1391), .B(n1331), .Z(n1310) );
  XOR2_X1 U1373 ( .A(n1388), .B(n1392), .Z(n1331) );
  NAND2_X1 U1374 ( .A1(n1377), .A2(n1363), .ZN(n1391) );
  XNOR2_X1 U1375 ( .A(n1393), .B(n1394), .ZN(n1363) );
  XNOR2_X1 U1376 ( .A(n1293), .B(n1290), .ZN(n1390) );
  XOR2_X1 U1377 ( .A(n1395), .B(n1340), .Z(n1290) );
  XOR2_X1 U1378 ( .A(n1383), .B(n1396), .Z(n1340) );
  NAND2_X1 U1379 ( .A1(n1361), .A2(n1375), .ZN(n1395) );
  XOR2_X1 U1380 ( .A(n1386), .B(n1397), .Z(n1361) );
  XOR2_X1 U1381 ( .A(n1398), .B(n1344), .Z(n1293) );
  XOR2_X1 U1382 ( .A(n1393), .B(n1399), .Z(n1344) );
  NAND2_X1 U1383 ( .A1(n1372), .A2(n1354), .ZN(n1398) );
  XNOR2_X1 U1384 ( .A(n1381), .B(n1400), .ZN(n1354) );
  XOR2_X1 U1385 ( .A(n1401), .B(n1402), .Z(n1312) );
  XOR2_X1 U1386 ( .A(n1303), .B(n1320), .Z(n1402) );
  XOR2_X1 U1387 ( .A(n1403), .B(n1369), .Z(n1320) );
  XOR2_X1 U1388 ( .A(n1393), .B(n1404), .Z(n1369) );
  NAND2_X1 U1389 ( .A1(n1334), .A2(n1336), .ZN(n1403) );
  XNOR2_X1 U1390 ( .A(n1383), .B(n1405), .ZN(n1336) );
  XOR2_X1 U1391 ( .A(n1381), .B(n1406), .Z(n1334) );
  XOR2_X1 U1392 ( .A(n1407), .B(n1367), .Z(n1303) );
  XOR2_X1 U1393 ( .A(n1386), .B(n1408), .Z(n1367) );
  NAND2_X1 U1394 ( .A1(n1347), .A2(n1349), .ZN(n1407) );
  XNOR2_X1 U1395 ( .A(n1393), .B(n1409), .ZN(n1349) );
  XNOR2_X1 U1396 ( .A(n1388), .B(n1410), .ZN(n1347) );
  XOR2_X1 U1397 ( .A(n1411), .B(n1271), .Z(n1401) );
  XNOR2_X1 U1398 ( .A(n1412), .B(n1375), .ZN(n1271) );
  XNOR2_X1 U1399 ( .A(n1388), .B(n1413), .ZN(n1375) );
  NAND2_X1 U1400 ( .A1(n1341), .A2(n1339), .ZN(n1412) );
  XNOR2_X1 U1401 ( .A(n1393), .B(n1414), .ZN(n1339) );
  XNOR2_X1 U1402 ( .A(n1415), .B(n1416), .ZN(n1393) );
  XNOR2_X1 U1403 ( .A(n1381), .B(n1417), .ZN(n1341) );
  XNOR2_X1 U1404 ( .A(n1275), .B(n1315), .ZN(n1411) );
  XOR2_X1 U1405 ( .A(n1418), .B(n1377), .Z(n1315) );
  XOR2_X1 U1406 ( .A(n1381), .B(n1419), .Z(n1377) );
  XOR2_X1 U1407 ( .A(n1420), .B(n1421), .Z(n1381) );
  NAND2_X1 U1408 ( .A1(n1330), .A2(n1332), .ZN(n1418) );
  XNOR2_X1 U1409 ( .A(n1386), .B(n1422), .ZN(n1332) );
  XOR2_X1 U1410 ( .A(n1383), .B(n1423), .Z(n1330) );
  XOR2_X1 U1411 ( .A(n1424), .B(n1372), .Z(n1275) );
  XNOR2_X1 U1412 ( .A(n1383), .B(n1425), .ZN(n1372) );
  XNOR2_X1 U1413 ( .A(n1426), .B(n1427), .ZN(n1383) );
  INV_X1 U1414 ( .A(n1415), .ZN(n1427) );
  XNOR2_X1 U1415 ( .A(n1428), .B(n1429), .ZN(n1415) );
  XOR2_X1 U1416 ( .A(n1400), .B(n1382), .Z(n1429) );
  XNOR2_X1 U1417 ( .A(n1430), .B(n1431), .ZN(n1382) );
  NAND2_X1 U1418 ( .A1(n1432), .A2(n1433), .ZN(n1430) );
  XNOR2_X1 U1419 ( .A(n1434), .B(n1435), .ZN(n1400) );
  NAND2_X1 U1420 ( .A1(n1436), .A2(n1437), .ZN(n1434) );
  XOR2_X1 U1421 ( .A(n1438), .B(n1406), .Z(n1428) );
  XOR2_X1 U1422 ( .A(n1439), .B(n1440), .Z(n1406) );
  NAND2_X1 U1423 ( .A1(n1441), .A2(n1442), .ZN(n1439) );
  XNOR2_X1 U1424 ( .A(n1419), .B(n1417), .ZN(n1438) );
  XNOR2_X1 U1425 ( .A(n1443), .B(n1444), .ZN(n1417) );
  NAND2_X1 U1426 ( .A1(n1445), .A2(n1446), .ZN(n1443) );
  XOR2_X1 U1427 ( .A(n1447), .B(n1448), .Z(n1419) );
  NAND2_X1 U1428 ( .A1(n1449), .A2(n1450), .ZN(n1447) );
  NAND2_X1 U1429 ( .A1(n1345), .A2(n1343), .ZN(n1424) );
  XNOR2_X1 U1430 ( .A(n1386), .B(n1451), .ZN(n1343) );
  XOR2_X1 U1431 ( .A(n1420), .B(n1416), .Z(n1386) );
  XNOR2_X1 U1432 ( .A(n1452), .B(n1453), .ZN(n1416) );
  XOR2_X1 U1433 ( .A(n1389), .B(n1454), .Z(n1453) );
  XOR2_X1 U1434 ( .A(n1455), .B(n1456), .Z(n1389) );
  NAND2_X1 U1435 ( .A1(n1457), .A2(n1435), .ZN(n1455) );
  XOR2_X1 U1436 ( .A(n1458), .B(n1392), .Z(n1452) );
  XNOR2_X1 U1437 ( .A(n1459), .B(n1460), .ZN(n1392) );
  NAND2_X1 U1438 ( .A1(n1461), .A2(n1431), .ZN(n1459) );
  XNOR2_X1 U1439 ( .A(n1413), .B(n1410), .ZN(n1458) );
  XOR2_X1 U1440 ( .A(n1462), .B(n1463), .Z(n1410) );
  NAND2_X1 U1441 ( .A1(n1440), .A2(n1464), .ZN(n1462) );
  XOR2_X1 U1442 ( .A(n1465), .B(n1466), .Z(n1413) );
  NAND2_X1 U1443 ( .A1(n1467), .A2(n1448), .ZN(n1465) );
  XOR2_X1 U1444 ( .A(n1468), .B(n1469), .Z(n1420) );
  XOR2_X1 U1445 ( .A(n1396), .B(n1384), .Z(n1469) );
  XNOR2_X1 U1446 ( .A(n1470), .B(n1436), .ZN(n1384) );
  NAND2_X1 U1447 ( .A1(n1456), .A2(n1437), .ZN(n1470) );
  XNOR2_X1 U1448 ( .A(n1471), .B(n1432), .ZN(n1396) );
  NAND2_X1 U1449 ( .A1(n1460), .A2(n1433), .ZN(n1471) );
  XOR2_X1 U1450 ( .A(n1472), .B(n1423), .Z(n1468) );
  XNOR2_X1 U1451 ( .A(n1473), .B(n1442), .ZN(n1423) );
  NAND2_X1 U1452 ( .A1(n1441), .A2(n1463), .ZN(n1473) );
  XOR2_X1 U1453 ( .A(n1425), .B(n1405), .Z(n1472) );
  XOR2_X1 U1454 ( .A(n1474), .B(n1445), .Z(n1405) );
  NAND2_X1 U1455 ( .A1(n1446), .A2(n1475), .ZN(n1474) );
  XOR2_X1 U1456 ( .A(n1476), .B(n1449), .Z(n1425) );
  NAND2_X1 U1457 ( .A1(n1466), .A2(n1450), .ZN(n1476) );
  XOR2_X1 U1458 ( .A(n1388), .B(n1454), .Z(n1345) );
  XNOR2_X1 U1459 ( .A(n1477), .B(n1475), .ZN(n1454) );
  NAND2_X1 U1460 ( .A1(n1444), .A2(n1478), .ZN(n1477) );
  XOR2_X1 U1461 ( .A(n1426), .B(n1421), .Z(n1388) );
  XNOR2_X1 U1462 ( .A(n1479), .B(n1480), .ZN(n1421) );
  XOR2_X1 U1463 ( .A(n1394), .B(n1399), .Z(n1480) );
  XOR2_X1 U1464 ( .A(n1481), .B(n1461), .Z(n1399) );
  NAND2_X1 U1465 ( .A1(n1431), .A2(n1432), .ZN(n1481) );
  XNOR2_X1 U1466 ( .A(n1482), .B(n1483), .ZN(n1432) );
  XNOR2_X1 U1467 ( .A(n1484), .B(n1485), .ZN(n1431) );
  XNOR2_X1 U1468 ( .A(n1486), .B(n1457), .ZN(n1394) );
  NAND2_X1 U1469 ( .A1(n1435), .A2(n1436), .ZN(n1486) );
  XNOR2_X1 U1470 ( .A(n1487), .B(n1488), .ZN(n1436) );
  XNOR2_X1 U1471 ( .A(n1489), .B(n1490), .ZN(n1435) );
  XOR2_X1 U1472 ( .A(n1491), .B(n1414), .Z(n1479) );
  XNOR2_X1 U1473 ( .A(n1492), .B(n1464), .ZN(n1414) );
  NAND2_X1 U1474 ( .A1(n1440), .A2(n1442), .ZN(n1492) );
  XNOR2_X1 U1475 ( .A(n1484), .B(n1493), .ZN(n1442) );
  XOR2_X1 U1476 ( .A(n1487), .B(n1494), .Z(n1440) );
  XNOR2_X1 U1477 ( .A(n1404), .B(n1409), .ZN(n1491) );
  XNOR2_X1 U1478 ( .A(n1495), .B(n1478), .ZN(n1409) );
  NAND2_X1 U1479 ( .A1(n1445), .A2(n1444), .ZN(n1495) );
  XNOR2_X1 U1480 ( .A(n1496), .B(n1497), .ZN(n1444) );
  XOR2_X1 U1481 ( .A(n1489), .B(n1498), .Z(n1445) );
  XOR2_X1 U1482 ( .A(n1499), .B(n1467), .Z(n1404) );
  NAND2_X1 U1483 ( .A1(n1448), .A2(n1449), .ZN(n1499) );
  XNOR2_X1 U1484 ( .A(n1496), .B(n1500), .ZN(n1449) );
  XOR2_X1 U1485 ( .A(n1482), .B(n1501), .Z(n1448) );
  XOR2_X1 U1486 ( .A(n1502), .B(n1503), .Z(n1426) );
  XOR2_X1 U1487 ( .A(n1387), .B(n1397), .Z(n1503) );
  XNOR2_X1 U1488 ( .A(n1504), .B(n1437), .ZN(n1397) );
  XNOR2_X1 U1489 ( .A(n1484), .B(n1505), .ZN(n1437) );
  NAND2_X1 U1490 ( .A1(n1456), .A2(n1457), .ZN(n1504) );
  XNOR2_X1 U1491 ( .A(n1496), .B(n1506), .ZN(n1457) );
  XOR2_X1 U1492 ( .A(n1482), .B(n1507), .Z(n1456) );
  XNOR2_X1 U1493 ( .A(n1508), .B(n1433), .ZN(n1387) );
  XNOR2_X1 U1494 ( .A(n1496), .B(n1509), .ZN(n1433) );
  NAND2_X1 U1495 ( .A1(n1461), .A2(n1460), .ZN(n1508) );
  XNOR2_X1 U1496 ( .A(n1489), .B(n1510), .ZN(n1460) );
  XOR2_X1 U1497 ( .A(n1487), .B(n1511), .Z(n1461) );
  XOR2_X1 U1498 ( .A(n1512), .B(n1451), .Z(n1502) );
  XOR2_X1 U1499 ( .A(n1513), .B(n1441), .Z(n1451) );
  XOR2_X1 U1500 ( .A(n1482), .B(n1514), .Z(n1441) );
  NAND2_X1 U1501 ( .A1(n1463), .A2(n1464), .ZN(n1513) );
  XNOR2_X1 U1502 ( .A(n1489), .B(n1515), .ZN(n1464) );
  XOR2_X1 U1503 ( .A(n1496), .B(n1516), .Z(n1463) );
  XOR2_X1 U1504 ( .A(n1517), .B(n1518), .Z(n1496) );
  XNOR2_X1 U1505 ( .A(n1408), .B(n1422), .ZN(n1512) );
  XOR2_X1 U1506 ( .A(n1519), .B(n1446), .Z(n1422) );
  XOR2_X1 U1507 ( .A(n1487), .B(n1520), .Z(n1446) );
  NAND2_X1 U1508 ( .A1(n1478), .A2(n1475), .ZN(n1519) );
  XNOR2_X1 U1509 ( .A(n1484), .B(n1521), .ZN(n1475) );
  XNOR2_X1 U1510 ( .A(n1482), .B(n1522), .ZN(n1478) );
  XNOR2_X1 U1511 ( .A(n1523), .B(n1524), .ZN(n1482) );
  XNOR2_X1 U1512 ( .A(n1525), .B(n1450), .ZN(n1408) );
  XNOR2_X1 U1513 ( .A(n1489), .B(n1526), .ZN(n1450) );
  XNOR2_X1 U1514 ( .A(n1527), .B(n1523), .ZN(n1489) );
  XNOR2_X1 U1515 ( .A(n1528), .B(n1529), .ZN(n1523) );
  XOR2_X1 U1516 ( .A(n1516), .B(n1506), .Z(n1529) );
  XNOR2_X1 U1517 ( .A(n1530), .B(n1531), .ZN(n1506) );
  NAND2_X1 U1518 ( .A1(n1532), .A2(n1533), .ZN(n1530) );
  XOR2_X1 U1519 ( .A(n1534), .B(n1535), .Z(n1516) );
  NAND2_X1 U1520 ( .A1(n1536), .A2(n1537), .ZN(n1534) );
  XOR2_X1 U1521 ( .A(n1538), .B(n1500), .Z(n1528) );
  XNOR2_X1 U1522 ( .A(n1539), .B(n1540), .ZN(n1500) );
  NAND2_X1 U1523 ( .A1(n1541), .A2(n1542), .ZN(n1539) );
  XNOR2_X1 U1524 ( .A(n1509), .B(n1497), .ZN(n1538) );
  XNOR2_X1 U1525 ( .A(n1543), .B(n1544), .ZN(n1497) );
  NAND2_X1 U1526 ( .A1(n1545), .A2(n1546), .ZN(n1543) );
  XNOR2_X1 U1527 ( .A(n1547), .B(n1548), .ZN(n1509) );
  NAND2_X1 U1528 ( .A1(n1549), .A2(n1550), .ZN(n1547) );
  NAND2_X1 U1529 ( .A1(n1467), .A2(n1466), .ZN(n1525) );
  XOR2_X1 U1530 ( .A(n1487), .B(n1551), .Z(n1466) );
  XOR2_X1 U1531 ( .A(n1517), .B(n1524), .Z(n1487) );
  XNOR2_X1 U1532 ( .A(n1552), .B(n1553), .ZN(n1524) );
  XOR2_X1 U1533 ( .A(n1521), .B(n1554), .Z(n1553) );
  XNOR2_X1 U1534 ( .A(n1555), .B(n1556), .ZN(n1521) );
  NAND2_X1 U1535 ( .A1(n1557), .A2(n1535), .ZN(n1555) );
  XOR2_X1 U1536 ( .A(n1558), .B(n1505), .Z(n1552) );
  XOR2_X1 U1537 ( .A(n1559), .B(n1560), .Z(n1505) );
  NAND2_X1 U1538 ( .A1(n1561), .A2(n1548), .ZN(n1559) );
  XNOR2_X1 U1539 ( .A(n1493), .B(n1485), .ZN(n1558) );
  XOR2_X1 U1540 ( .A(n1562), .B(n1563), .Z(n1485) );
  NAND2_X1 U1541 ( .A1(n1564), .A2(n1544), .ZN(n1562) );
  XOR2_X1 U1542 ( .A(n1565), .B(n1566), .Z(n1493) );
  NAND2_X1 U1543 ( .A1(n1567), .A2(n1540), .ZN(n1565) );
  XOR2_X1 U1544 ( .A(n1568), .B(n1569), .Z(n1517) );
  XOR2_X1 U1545 ( .A(n1510), .B(n1515), .Z(n1569) );
  XOR2_X1 U1546 ( .A(n1570), .B(n1532), .Z(n1515) );
  NAND2_X1 U1547 ( .A1(n1533), .A2(n1571), .ZN(n1570) );
  XOR2_X1 U1548 ( .A(n1572), .B(n1536), .Z(n1510) );
  NAND2_X1 U1549 ( .A1(n1537), .A2(n1556), .ZN(n1572) );
  XOR2_X1 U1550 ( .A(n1573), .B(n1498), .Z(n1568) );
  XNOR2_X1 U1551 ( .A(n1574), .B(n1542), .ZN(n1498) );
  NAND2_X1 U1552 ( .A1(n1541), .A2(n1566), .ZN(n1574) );
  XNOR2_X1 U1553 ( .A(n1490), .B(n1526), .ZN(n1573) );
  XOR2_X1 U1554 ( .A(n1575), .B(n1549), .Z(n1526) );
  NAND2_X1 U1555 ( .A1(n1560), .A2(n1550), .ZN(n1575) );
  XOR2_X1 U1556 ( .A(n1576), .B(n1545), .Z(n1490) );
  NAND2_X1 U1557 ( .A1(n1563), .A2(n1546), .ZN(n1576) );
  XOR2_X1 U1558 ( .A(n1484), .B(n1554), .Z(n1467) );
  XNOR2_X1 U1559 ( .A(n1577), .B(n1571), .ZN(n1554) );
  NAND2_X1 U1560 ( .A1(n1578), .A2(n1531), .ZN(n1577) );
  XNOR2_X1 U1561 ( .A(n1518), .B(n1527), .ZN(n1484) );
  XNOR2_X1 U1562 ( .A(n1579), .B(n1580), .ZN(n1527) );
  XOR2_X1 U1563 ( .A(n1494), .B(n1511), .Z(n1580) );
  XNOR2_X1 U1564 ( .A(n1581), .B(n1533), .ZN(n1511) );
  XNOR2_X1 U1565 ( .A(n1582), .B(n1583), .ZN(n1533) );
  NAND2_X1 U1566 ( .A1(n1571), .A2(n1578), .ZN(n1581) );
  XNOR2_X1 U1567 ( .A(n1584), .B(n1585), .ZN(n1571) );
  XNOR2_X1 U1568 ( .A(n1586), .B(n1546), .ZN(n1494) );
  XNOR2_X1 U1569 ( .A(n1587), .B(n1588), .ZN(n1546) );
  NAND2_X1 U1570 ( .A1(n1563), .A2(n1564), .ZN(n1586) );
  XOR2_X1 U1571 ( .A(n1589), .B(n1590), .Z(n1563) );
  XOR2_X1 U1572 ( .A(n1591), .B(n1551), .Z(n1579) );
  XNOR2_X1 U1573 ( .A(n1592), .B(n1537), .ZN(n1551) );
  XNOR2_X1 U1574 ( .A(n1593), .B(n1594), .ZN(n1537) );
  NAND2_X1 U1575 ( .A1(n1557), .A2(n1556), .ZN(n1592) );
  XNOR2_X1 U1576 ( .A(n1587), .B(n1595), .ZN(n1556) );
  XNOR2_X1 U1577 ( .A(n1520), .B(n1488), .ZN(n1591) );
  XOR2_X1 U1578 ( .A(n1596), .B(n1541), .Z(n1488) );
  XOR2_X1 U1579 ( .A(n1584), .B(n1597), .Z(n1541) );
  NAND2_X1 U1580 ( .A1(n1566), .A2(n1567), .ZN(n1596) );
  XOR2_X1 U1581 ( .A(n1593), .B(n1598), .Z(n1566) );
  XNOR2_X1 U1582 ( .A(n1599), .B(n1550), .ZN(n1520) );
  XNOR2_X1 U1583 ( .A(n1589), .B(n1600), .ZN(n1550) );
  NAND2_X1 U1584 ( .A1(n1560), .A2(n1561), .ZN(n1599) );
  XOR2_X1 U1585 ( .A(n1582), .B(n1601), .Z(n1560) );
  XNOR2_X1 U1586 ( .A(n1602), .B(n1603), .ZN(n1518) );
  XOR2_X1 U1587 ( .A(n1514), .B(n1522), .Z(n1603) );
  XNOR2_X1 U1588 ( .A(n1604), .B(n1578), .ZN(n1522) );
  XNOR2_X1 U1589 ( .A(n1593), .B(n1605), .ZN(n1578) );
  NAND2_X1 U1590 ( .A1(n1532), .A2(n1531), .ZN(n1604) );
  XNOR2_X1 U1591 ( .A(n1587), .B(n1606), .ZN(n1531) );
  XOR2_X1 U1592 ( .A(n1589), .B(n1607), .Z(n1532) );
  XOR2_X1 U1593 ( .A(n1608), .B(n1561), .Z(n1514) );
  XOR2_X1 U1594 ( .A(n1584), .B(n1609), .Z(n1561) );
  NAND2_X1 U1595 ( .A1(n1549), .A2(n1548), .ZN(n1608) );
  XNOR2_X1 U1596 ( .A(n1593), .B(n1610), .ZN(n1548) );
  XOR2_X1 U1597 ( .A(n1587), .B(n1611), .Z(n1549) );
  XOR2_X1 U1598 ( .A(n1612), .B(n1507), .Z(n1602) );
  XOR2_X1 U1599 ( .A(n1613), .B(n1557), .Z(n1507) );
  XOR2_X1 U1600 ( .A(n1589), .B(n1614), .Z(n1557) );
  NAND2_X1 U1601 ( .A1(n1536), .A2(n1535), .ZN(n1613) );
  XOR2_X1 U1602 ( .A(n1582), .B(n1615), .Z(n1535) );
  XOR2_X1 U1603 ( .A(n1584), .B(n1616), .Z(n1536) );
  XNOR2_X1 U1604 ( .A(n1483), .B(n1501), .ZN(n1612) );
  XOR2_X1 U1605 ( .A(n1617), .B(n1564), .Z(n1501) );
  XOR2_X1 U1606 ( .A(n1582), .B(n1618), .Z(n1564) );
  NAND2_X1 U1607 ( .A1(n1545), .A2(n1544), .ZN(n1617) );
  XNOR2_X1 U1608 ( .A(n1584), .B(n1619), .ZN(n1544) );
  XNOR2_X1 U1609 ( .A(n1620), .B(n1621), .ZN(n1584) );
  XOR2_X1 U1610 ( .A(n1593), .B(n1622), .Z(n1545) );
  XOR2_X1 U1611 ( .A(n1623), .B(n1624), .Z(n1593) );
  XNOR2_X1 U1612 ( .A(n1625), .B(n1567), .ZN(n1483) );
  XNOR2_X1 U1613 ( .A(n1587), .B(n1626), .ZN(n1567) );
  XOR2_X1 U1614 ( .A(n1627), .B(n1621), .Z(n1587) );
  XNOR2_X1 U1615 ( .A(n1628), .B(n1629), .ZN(n1621) );
  XOR2_X1 U1616 ( .A(n1605), .B(n1610), .Z(n1629) );
  XOR2_X1 U1617 ( .A(n1630), .B(n1631), .Z(n1610) );
  NAND2_X1 U1618 ( .A1(n1632), .A2(n1633), .ZN(n1630) );
  XOR2_X1 U1619 ( .A(n1634), .B(n1635), .Z(n1605) );
  NAND2_X1 U1620 ( .A1(n1636), .A2(n1637), .ZN(n1634) );
  XOR2_X1 U1621 ( .A(n1638), .B(n1622), .Z(n1628) );
  XNOR2_X1 U1622 ( .A(n1639), .B(n1640), .ZN(n1622) );
  NAND2_X1 U1623 ( .A1(n1641), .A2(n1642), .ZN(n1639) );
  XNOR2_X1 U1624 ( .A(n1598), .B(n1594), .ZN(n1638) );
  XOR2_X1 U1625 ( .A(n1643), .B(n1644), .Z(n1594) );
  NAND2_X1 U1626 ( .A1(n1645), .A2(n1646), .ZN(n1643) );
  XNOR2_X1 U1627 ( .A(n1647), .B(n1648), .ZN(n1598) );
  NAND2_X1 U1628 ( .A1(n1649), .A2(n1650), .ZN(n1647) );
  NAND2_X1 U1629 ( .A1(n1542), .A2(n1540), .ZN(n1625) );
  XNOR2_X1 U1630 ( .A(n1589), .B(n1651), .ZN(n1540) );
  XNOR2_X1 U1631 ( .A(n1623), .B(n1652), .ZN(n1589) );
  INV_X1 U1632 ( .A(n1620), .ZN(n1652) );
  XNOR2_X1 U1633 ( .A(n1653), .B(n1654), .ZN(n1620) );
  XOR2_X1 U1634 ( .A(n1655), .B(n1583), .Z(n1654) );
  XNOR2_X1 U1635 ( .A(n1656), .B(n1657), .ZN(n1583) );
  NAND2_X1 U1636 ( .A1(n1644), .A2(n1658), .ZN(n1656) );
  XOR2_X1 U1637 ( .A(n1659), .B(n1601), .Z(n1653) );
  XOR2_X1 U1638 ( .A(n1660), .B(n1661), .Z(n1601) );
  NAND2_X1 U1639 ( .A1(n1662), .A2(n1648), .ZN(n1660) );
  XNOR2_X1 U1640 ( .A(n1618), .B(n1615), .ZN(n1659) );
  XOR2_X1 U1641 ( .A(n1663), .B(n1664), .Z(n1615) );
  NAND2_X1 U1642 ( .A1(n1665), .A2(n1631), .ZN(n1663) );
  XOR2_X1 U1643 ( .A(n1666), .B(n1667), .Z(n1618) );
  NAND2_X1 U1644 ( .A1(n1635), .A2(n1668), .ZN(n1666) );
  XOR2_X1 U1645 ( .A(n1669), .B(n1670), .Z(n1623) );
  XOR2_X1 U1646 ( .A(n1626), .B(n1595), .Z(n1670) );
  XNOR2_X1 U1647 ( .A(n1671), .B(n1650), .ZN(n1595) );
  NAND2_X1 U1648 ( .A1(n1649), .A2(n1661), .ZN(n1671) );
  XOR2_X1 U1649 ( .A(n1672), .B(n1636), .Z(n1626) );
  NAND2_X1 U1650 ( .A1(n1637), .A2(n1667), .ZN(n1672) );
  XOR2_X1 U1651 ( .A(n1673), .B(n1588), .Z(n1669) );
  XOR2_X1 U1652 ( .A(n1674), .B(n1645), .Z(n1588) );
  NAND2_X1 U1653 ( .A1(n1657), .A2(n1646), .ZN(n1674) );
  XNOR2_X1 U1654 ( .A(n1611), .B(n1606), .ZN(n1673) );
  XOR2_X1 U1655 ( .A(n1675), .B(n1632), .Z(n1606) );
  NAND2_X1 U1656 ( .A1(n1664), .A2(n1633), .ZN(n1675) );
  XNOR2_X1 U1657 ( .A(n1676), .B(n1642), .ZN(n1611) );
  NAND2_X1 U1658 ( .A1(n1641), .A2(n1677), .ZN(n1676) );
  XNOR2_X1 U1659 ( .A(n1582), .B(n1655), .ZN(n1542) );
  XNOR2_X1 U1660 ( .A(n1678), .B(n1677), .ZN(n1655) );
  NAND2_X1 U1661 ( .A1(n1640), .A2(n1679), .ZN(n1678) );
  XOR2_X1 U1662 ( .A(n1627), .B(n1624), .Z(n1582) );
  XNOR2_X1 U1663 ( .A(n1680), .B(n1681), .ZN(n1624) );
  XOR2_X1 U1664 ( .A(n1619), .B(n1609), .Z(n1681) );
  XNOR2_X1 U1665 ( .A(n1682), .B(n1668), .ZN(n1609) );
  NAND2_X1 U1666 ( .A1(n1635), .A2(n1636), .ZN(n1682) );
  XOR2_X1 U1667 ( .A(n1683), .B(n1684), .Z(n1636) );
  XOR2_X1 U1668 ( .A(n1685), .B(n1686), .Z(n1635) );
  XOR2_X1 U1669 ( .A(n1687), .B(n1665), .Z(n1619) );
  NAND2_X1 U1670 ( .A1(n1631), .A2(n1632), .ZN(n1687) );
  XOR2_X1 U1671 ( .A(n1688), .B(n1689), .Z(n1632) );
  XOR2_X1 U1672 ( .A(n1690), .B(n1691), .Z(n1631) );
  XOR2_X1 U1673 ( .A(n1692), .B(n1616), .Z(n1680) );
  XNOR2_X1 U1674 ( .A(n1693), .B(n1679), .ZN(n1616) );
  NAND2_X1 U1675 ( .A1(n1640), .A2(n1642), .ZN(n1693) );
  XNOR2_X1 U1676 ( .A(n1694), .B(n1695), .ZN(n1642) );
  XNOR2_X1 U1677 ( .A(n1683), .B(n1696), .ZN(n1640) );
  XNOR2_X1 U1678 ( .A(n1585), .B(n1597), .ZN(n1692) );
  XNOR2_X1 U1679 ( .A(n1697), .B(n1658), .ZN(n1597) );
  NAND2_X1 U1680 ( .A1(n1644), .A2(n1645), .ZN(n1697) );
  XOR2_X1 U1681 ( .A(n1685), .B(n1698), .Z(n1645) );
  XOR2_X1 U1682 ( .A(n1688), .B(n1699), .Z(n1644) );
  XOR2_X1 U1683 ( .A(n1700), .B(n1662), .Z(n1585) );
  NAND2_X1 U1684 ( .A1(n1648), .A2(n1650), .ZN(n1700) );
  XNOR2_X1 U1685 ( .A(n1690), .B(n1701), .ZN(n1650) );
  XNOR2_X1 U1686 ( .A(n1694), .B(n1702), .ZN(n1648) );
  XOR2_X1 U1687 ( .A(n1703), .B(n1704), .Z(n1627) );
  XOR2_X1 U1688 ( .A(n1590), .B(n1651), .Z(n1704) );
  XNOR2_X1 U1689 ( .A(n1705), .B(n1633), .ZN(n1651) );
  XNOR2_X1 U1690 ( .A(n1685), .B(n1706), .ZN(n1633) );
  NAND2_X1 U1691 ( .A1(n1665), .A2(n1664), .ZN(n1705) );
  XOR2_X1 U1692 ( .A(n1683), .B(n1707), .Z(n1664) );
  XOR2_X1 U1693 ( .A(n1694), .B(n1708), .Z(n1665) );
  XOR2_X1 U1694 ( .A(n1709), .B(n1649), .Z(n1590) );
  XOR2_X1 U1695 ( .A(n1688), .B(n1710), .Z(n1649) );
  NAND2_X1 U1696 ( .A1(n1662), .A2(n1661), .ZN(n1709) );
  XOR2_X1 U1697 ( .A(n1685), .B(n1711), .Z(n1661) );
  XOR2_X1 U1698 ( .A(n1683), .B(n1712), .Z(n1662) );
  XOR2_X1 U1699 ( .A(n1713), .B(n1607), .Z(n1703) );
  XOR2_X1 U1700 ( .A(n1714), .B(n1641), .Z(n1607) );
  XOR2_X1 U1701 ( .A(n1690), .B(n1715), .Z(n1641) );
  NAND2_X1 U1702 ( .A1(n1679), .A2(n1677), .ZN(n1714) );
  XNOR2_X1 U1703 ( .A(n1688), .B(n1716), .ZN(n1677) );
  XNOR2_X1 U1704 ( .A(n1685), .B(n1717), .ZN(n1679) );
  XOR2_X1 U1705 ( .A(n1718), .B(n1719), .Z(n1685) );
  XNOR2_X1 U1706 ( .A(n1614), .B(n1600), .ZN(n1713) );
  XNOR2_X1 U1707 ( .A(n1720), .B(n1646), .ZN(n1600) );
  XNOR2_X1 U1708 ( .A(n1683), .B(n1721), .ZN(n1646) );
  XNOR2_X1 U1709 ( .A(n1722), .B(n1723), .ZN(n1683) );
  NAND2_X1 U1710 ( .A1(n1658), .A2(n1657), .ZN(n1720) );
  XNOR2_X1 U1711 ( .A(n1694), .B(n1724), .ZN(n1657) );
  XNOR2_X1 U1712 ( .A(n1690), .B(n1725), .ZN(n1658) );
  XOR2_X1 U1713 ( .A(n1726), .B(n1637), .Z(n1614) );
  XOR2_X1 U1714 ( .A(n1694), .B(n1727), .Z(n1637) );
  XOR2_X1 U1715 ( .A(n1728), .B(n1719), .Z(n1694) );
  XNOR2_X1 U1716 ( .A(n1729), .B(n1730), .ZN(n1719) );
  XOR2_X1 U1717 ( .A(n1721), .B(n1696), .Z(n1730) );
  XOR2_X1 U1718 ( .A(n1731), .B(n1732), .Z(n1696) );
  NAND2_X1 U1719 ( .A1(n1733), .A2(n1734), .ZN(n1731) );
  XOR2_X1 U1720 ( .A(n1735), .B(n1736), .Z(n1721) );
  NAND2_X1 U1721 ( .A1(n1737), .A2(n1738), .ZN(n1735) );
  XOR2_X1 U1722 ( .A(n1739), .B(n1712), .Z(n1729) );
  XNOR2_X1 U1723 ( .A(n1740), .B(n1741), .ZN(n1712) );
  NAND2_X1 U1724 ( .A1(n1742), .A2(n1743), .ZN(n1740) );
  XNOR2_X1 U1725 ( .A(n1684), .B(n1707), .ZN(n1739) );
  XNOR2_X1 U1726 ( .A(n1744), .B(n1745), .ZN(n1707) );
  NAND2_X1 U1727 ( .A1(n1746), .A2(n1747), .ZN(n1744) );
  XNOR2_X1 U1728 ( .A(n1748), .B(n1749), .ZN(n1684) );
  NAND2_X1 U1729 ( .A1(n1750), .A2(n1751), .ZN(n1748) );
  NAND2_X1 U1730 ( .A1(n1667), .A2(n1668), .ZN(n1726) );
  XNOR2_X1 U1731 ( .A(n1688), .B(n1752), .ZN(n1668) );
  XNOR2_X1 U1732 ( .A(n1728), .B(n1753), .ZN(n1688) );
  INV_X1 U1733 ( .A(n1722), .ZN(n1753) );
  XNOR2_X1 U1734 ( .A(n1754), .B(n1755), .ZN(n1722) );
  XOR2_X1 U1735 ( .A(n1706), .B(n1711), .Z(n1755) );
  XOR2_X1 U1736 ( .A(n1756), .B(n1757), .Z(n1711) );
  NAND2_X1 U1737 ( .A1(n1746), .A2(n1745), .ZN(n1756) );
  XNOR2_X1 U1738 ( .A(n1758), .B(n1759), .ZN(n1706) );
  NAND2_X1 U1739 ( .A1(n1736), .A2(n1738), .ZN(n1758) );
  XOR2_X1 U1740 ( .A(n1760), .B(n1686), .Z(n1754) );
  XOR2_X1 U1741 ( .A(n1761), .B(n1762), .Z(n1686) );
  NAND2_X1 U1742 ( .A1(n1732), .A2(n1733), .ZN(n1761) );
  XNOR2_X1 U1743 ( .A(n1717), .B(n1698), .ZN(n1760) );
  XOR2_X1 U1744 ( .A(n1763), .B(n1764), .Z(n1698) );
  NAND2_X1 U1745 ( .A1(n1750), .A2(n1749), .ZN(n1763) );
  XNOR2_X1 U1746 ( .A(n1765), .B(n1766), .ZN(n1717) );
  NAND2_X1 U1747 ( .A1(n1741), .A2(n1743), .ZN(n1765) );
  XOR2_X1 U1748 ( .A(n1767), .B(n1768), .Z(n1728) );
  XOR2_X1 U1749 ( .A(n1701), .B(n1691), .Z(n1768) );
  XNOR2_X1 U1750 ( .A(n1769), .B(n1734), .ZN(n1691) );
  NAND2_X1 U1751 ( .A1(n1770), .A2(n1762), .ZN(n1769) );
  XNOR2_X1 U1752 ( .A(n1771), .B(n1751), .ZN(n1701) );
  NAND2_X1 U1753 ( .A1(n1772), .A2(n1764), .ZN(n1771) );
  XOR2_X1 U1754 ( .A(n1773), .B(n1715), .Z(n1767) );
  XNOR2_X1 U1755 ( .A(n1774), .B(n1737), .ZN(n1715) );
  NAND2_X1 U1756 ( .A1(n1775), .A2(n1759), .ZN(n1774) );
  XNOR2_X1 U1757 ( .A(n1725), .B(n1776), .ZN(n1773) );
  XOR2_X1 U1758 ( .A(n1777), .B(n1742), .Z(n1725) );
  NAND2_X1 U1759 ( .A1(n1778), .A2(n1766), .ZN(n1777) );
  XOR2_X1 U1760 ( .A(n1690), .B(n1776), .Z(n1667) );
  XNOR2_X1 U1761 ( .A(n1779), .B(n1747), .ZN(n1776) );
  NAND2_X1 U1762 ( .A1(n1757), .A2(n1780), .ZN(n1779) );
  XOR2_X1 U1763 ( .A(n1718), .B(n1723), .Z(n1690) );
  XNOR2_X1 U1764 ( .A(n1781), .B(n1782), .ZN(n1723) );
  XOR2_X1 U1765 ( .A(n1724), .B(n1727), .Z(n1782) );
  XNOR2_X1 U1766 ( .A(n1783), .B(n1738), .ZN(n1727) );
  XNOR2_X1 U1767 ( .A(n1784), .B(n1785), .ZN(n1738) );
  NAND2_X1 U1768 ( .A1(n1775), .A2(n1737), .ZN(n1783) );
  XNOR2_X1 U1769 ( .A(n1786), .B(n1787), .ZN(n1737) );
  XOR2_X1 U1770 ( .A(n1788), .B(n1746), .Z(n1724) );
  XOR2_X1 U1771 ( .A(n1789), .B(n1790), .Z(n1746) );
  NAND2_X1 U1772 ( .A1(n1780), .A2(n1747), .ZN(n1788) );
  XNOR2_X1 U1773 ( .A(n1791), .B(n1792), .ZN(n1747) );
  XOR2_X1 U1774 ( .A(n1793), .B(n1702), .Z(n1781) );
  XOR2_X1 U1775 ( .A(n1794), .B(n1733), .Z(n1702) );
  XOR2_X1 U1776 ( .A(n1791), .B(n1795), .Z(n1733) );
  NAND2_X1 U1777 ( .A1(n1770), .A2(n1734), .ZN(n1794) );
  XNOR2_X1 U1778 ( .A(n1784), .B(n1796), .ZN(n1734) );
  XNOR2_X1 U1779 ( .A(n1708), .B(n1695), .ZN(n1793) );
  XOR2_X1 U1780 ( .A(n1797), .B(n1750), .Z(n1695) );
  XOR2_X1 U1781 ( .A(n1798), .B(n1799), .Z(n1750) );
  NAND2_X1 U1782 ( .A1(n1772), .A2(n1751), .ZN(n1797) );
  XNOR2_X1 U1783 ( .A(n1789), .B(n1800), .ZN(n1751) );
  XNOR2_X1 U1784 ( .A(n1801), .B(n1743), .ZN(n1708) );
  XNOR2_X1 U1785 ( .A(n1786), .B(n1802), .ZN(n1743) );
  NAND2_X1 U1786 ( .A1(n1742), .A2(n1778), .ZN(n1801) );
  XOR2_X1 U1787 ( .A(n1798), .B(n1803), .Z(n1742) );
  XOR2_X1 U1788 ( .A(n1804), .B(n1805), .Z(n1718) );
  XOR2_X1 U1789 ( .A(n1710), .B(n1689), .Z(n1805) );
  XOR2_X1 U1790 ( .A(n1806), .B(n1772), .Z(n1689) );
  XOR2_X1 U1791 ( .A(n1791), .B(n1807), .Z(n1772) );
  NAND2_X1 U1792 ( .A1(n1764), .A2(n1749), .ZN(n1806) );
  XNOR2_X1 U1793 ( .A(n1786), .B(n1808), .ZN(n1749) );
  XOR2_X1 U1794 ( .A(n1784), .B(n1809), .Z(n1764) );
  XOR2_X1 U1795 ( .A(n1810), .B(n1775), .Z(n1710) );
  XOR2_X1 U1796 ( .A(n1798), .B(n1811), .Z(n1775) );
  NAND2_X1 U1797 ( .A1(n1736), .A2(n1759), .ZN(n1810) );
  XNOR2_X1 U1798 ( .A(n1789), .B(n1812), .ZN(n1759) );
  XOR2_X1 U1799 ( .A(n1791), .B(n1813), .Z(n1736) );
  XOR2_X1 U1800 ( .A(n1814), .B(n1716), .Z(n1804) );
  XNOR2_X1 U1801 ( .A(n1815), .B(n1780), .ZN(n1716) );
  XNOR2_X1 U1802 ( .A(n1784), .B(n1816), .ZN(n1780) );
  NAND2_X1 U1803 ( .A1(n1757), .A2(n1745), .ZN(n1815) );
  XNOR2_X1 U1804 ( .A(n1798), .B(n1817), .ZN(n1745) );
  XOR2_X1 U1805 ( .A(n1786), .B(n1818), .Z(n1757) );
  XNOR2_X1 U1806 ( .A(n1699), .B(n1752), .ZN(n1814) );
  XNOR2_X1 U1807 ( .A(n1819), .B(n1778), .ZN(n1752) );
  XNOR2_X1 U1808 ( .A(n1789), .B(n1820), .ZN(n1778) );
  NAND2_X1 U1809 ( .A1(n1766), .A2(n1741), .ZN(n1819) );
  XNOR2_X1 U1810 ( .A(n1784), .B(n1821), .ZN(n1741) );
  XOR2_X1 U1811 ( .A(n1822), .B(n1823), .Z(n1784) );
  XNOR2_X1 U1812 ( .A(n1791), .B(n1824), .ZN(n1766) );
  XNOR2_X1 U1813 ( .A(n1825), .B(n1826), .ZN(n1791) );
  XOR2_X1 U1814 ( .A(n1827), .B(n1770), .Z(n1699) );
  XOR2_X1 U1815 ( .A(n1786), .B(n1828), .Z(n1770) );
  XNOR2_X1 U1816 ( .A(n1826), .B(n1829), .ZN(n1786) );
  XNOR2_X1 U1817 ( .A(n1830), .B(n1831), .ZN(n1826) );
  XOR2_X1 U1818 ( .A(n1816), .B(n1821), .Z(n1831) );
  XOR2_X1 U1819 ( .A(n1832), .B(n1833), .Z(n1821) );
  NAND2_X1 U1820 ( .A1(n1834), .A2(n1835), .ZN(n1832) );
  XOR2_X1 U1821 ( .A(n1836), .B(n1837), .Z(n1816) );
  NAND2_X1 U1822 ( .A1(n1838), .A2(n1839), .ZN(n1836) );
  XOR2_X1 U1823 ( .A(n1840), .B(n1809), .Z(n1830) );
  XNOR2_X1 U1824 ( .A(n1841), .B(n1842), .ZN(n1809) );
  NAND2_X1 U1825 ( .A1(n1843), .A2(n1844), .ZN(n1841) );
  XNOR2_X1 U1826 ( .A(n1796), .B(n1785), .ZN(n1840) );
  XOR2_X1 U1827 ( .A(n1845), .B(n1846), .Z(n1785) );
  NAND2_X1 U1828 ( .A1(n1847), .A2(n1848), .ZN(n1845) );
  XOR2_X1 U1829 ( .A(n1849), .B(n1850), .Z(n1796) );
  NAND2_X1 U1830 ( .A1(n1851), .A2(n1852), .ZN(n1849) );
  NAND2_X1 U1831 ( .A1(n1762), .A2(n1732), .ZN(n1827) );
  XOR2_X1 U1832 ( .A(n1789), .B(n1853), .Z(n1732) );
  XNOR2_X1 U1833 ( .A(n1823), .B(n1829), .ZN(n1789) );
  XNOR2_X1 U1834 ( .A(n1854), .B(n1855), .ZN(n1829) );
  XNOR2_X1 U1835 ( .A(n1856), .B(n1811), .ZN(n1855) );
  XNOR2_X1 U1836 ( .A(n1857), .B(n1839), .ZN(n1811) );
  NAND2_X1 U1837 ( .A1(n1858), .A2(n1859), .ZN(n1857) );
  XOR2_X1 U1838 ( .A(n1860), .B(n1803), .Z(n1854) );
  XNOR2_X1 U1839 ( .A(n1861), .B(n1851), .ZN(n1803) );
  NAND2_X1 U1840 ( .A1(n1862), .A2(n1863), .ZN(n1861) );
  XNOR2_X1 U1841 ( .A(n1799), .B(n1817), .ZN(n1860) );
  XOR2_X1 U1842 ( .A(n1864), .B(n1834), .Z(n1817) );
  NAND2_X1 U1843 ( .A1(n1865), .A2(n1866), .ZN(n1864) );
  XNOR2_X1 U1844 ( .A(n1867), .B(n1847), .ZN(n1799) );
  NAND2_X1 U1845 ( .A1(n1868), .A2(n1869), .ZN(n1867) );
  XNOR2_X1 U1846 ( .A(n1870), .B(n1871), .ZN(n1823) );
  XOR2_X1 U1847 ( .A(n1807), .B(n1824), .Z(n1871) );
  XOR2_X1 U1848 ( .A(n1872), .B(n1873), .Z(n1824) );
  NAND2_X1 U1849 ( .A1(n1843), .A2(n1842), .ZN(n1872) );
  XNOR2_X1 U1850 ( .A(n1874), .B(n1859), .ZN(n1807) );
  NAND2_X1 U1851 ( .A1(n1838), .A2(n1837), .ZN(n1874) );
  XOR2_X1 U1852 ( .A(n1875), .B(n1795), .Z(n1870) );
  XNOR2_X1 U1853 ( .A(n1876), .B(n1869), .ZN(n1795) );
  NAND2_X1 U1854 ( .A1(n1846), .A2(n1848), .ZN(n1876) );
  XNOR2_X1 U1855 ( .A(n1813), .B(n1792), .ZN(n1875) );
  XOR2_X1 U1856 ( .A(n1877), .B(n1863), .Z(n1792) );
  NAND2_X1 U1857 ( .A1(n1850), .A2(n1852), .ZN(n1877) );
  XNOR2_X1 U1858 ( .A(n1878), .B(n1866), .ZN(n1813) );
  NAND2_X1 U1859 ( .A1(n1833), .A2(n1835), .ZN(n1878) );
  XNOR2_X1 U1860 ( .A(n1798), .B(n1856), .ZN(n1762) );
  XOR2_X1 U1861 ( .A(n1879), .B(n1844), .Z(n1856) );
  NAND2_X1 U1862 ( .A1(n1873), .A2(n1880), .ZN(n1879) );
  XNOR2_X1 U1863 ( .A(n1822), .B(n1881), .ZN(n1798) );
  INV_X1 U1864 ( .A(n1825), .ZN(n1881) );
  XNOR2_X1 U1865 ( .A(n1882), .B(n1883), .ZN(n1825) );
  XOR2_X1 U1866 ( .A(n1853), .B(n1790), .Z(n1883) );
  XOR2_X1 U1867 ( .A(n1884), .B(n1868), .Z(n1790) );
  NAND2_X1 U1868 ( .A1(n1846), .A2(n1869), .ZN(n1884) );
  XNOR2_X1 U1869 ( .A(n1885), .B(n1886), .ZN(n1869) );
  XOR2_X1 U1870 ( .A(n1887), .B(n1888), .Z(n1846) );
  XOR2_X1 U1871 ( .A(n1889), .B(n1865), .Z(n1853) );
  NAND2_X1 U1872 ( .A1(n1833), .A2(n1866), .ZN(n1889) );
  XNOR2_X1 U1873 ( .A(n1890), .B(n1891), .ZN(n1866) );
  XOR2_X1 U1874 ( .A(n1892), .B(n1893), .Z(n1833) );
  XOR2_X1 U1875 ( .A(n1894), .B(n1800), .Z(n1882) );
  XOR2_X1 U1876 ( .A(n1895), .B(n1862), .Z(n1800) );
  NAND2_X1 U1877 ( .A1(n1850), .A2(n1863), .ZN(n1895) );
  XOR2_X1 U1878 ( .A(n1892), .B(n1896), .Z(n1863) );
  XOR2_X1 U1879 ( .A(n1897), .B(n1898), .Z(n1850) );
  XNOR2_X1 U1880 ( .A(n1820), .B(n1812), .ZN(n1894) );
  XNOR2_X1 U1881 ( .A(n1899), .B(n1880), .ZN(n1812) );
  NAND2_X1 U1882 ( .A1(n1873), .A2(n1842), .ZN(n1899) );
  XNOR2_X1 U1883 ( .A(n1885), .B(n1900), .ZN(n1842) );
  XOR2_X1 U1884 ( .A(n1897), .B(n1901), .Z(n1873) );
  XNOR2_X1 U1885 ( .A(n1902), .B(n1858), .ZN(n1820) );
  NAND2_X1 U1886 ( .A1(n1837), .A2(n1859), .ZN(n1902) );
  XNOR2_X1 U1887 ( .A(n1887), .B(n1903), .ZN(n1859) );
  XOR2_X1 U1888 ( .A(n1890), .B(n1904), .Z(n1837) );
  XOR2_X1 U1889 ( .A(n1905), .B(n1906), .Z(n1822) );
  XOR2_X1 U1890 ( .A(n1818), .B(n1828), .Z(n1906) );
  XOR2_X1 U1891 ( .A(n1907), .B(n1838), .Z(n1828) );
  XOR2_X1 U1892 ( .A(n1892), .B(n1908), .Z(n1838) );
  NAND2_X1 U1893 ( .A1(n1839), .A2(n1858), .ZN(n1907) );
  XNOR2_X1 U1894 ( .A(n1885), .B(n1909), .ZN(n1858) );
  XNOR2_X1 U1895 ( .A(n1897), .B(n1910), .ZN(n1839) );
  XOR2_X1 U1896 ( .A(n1911), .B(n1843), .Z(n1818) );
  XOR2_X1 U1897 ( .A(n1887), .B(n1912), .Z(n1843) );
  NAND2_X1 U1898 ( .A1(n1844), .A2(n1880), .ZN(n1911) );
  XNOR2_X1 U1899 ( .A(n1892), .B(n1913), .ZN(n1880) );
  XNOR2_X1 U1900 ( .A(n1890), .B(n1914), .ZN(n1844) );
  XOR2_X1 U1901 ( .A(n1915), .B(n1802), .Z(n1905) );
  XNOR2_X1 U1902 ( .A(n1916), .B(n1848), .ZN(n1802) );
  XNOR2_X1 U1903 ( .A(n1890), .B(n1917), .ZN(n1848) );
  NAND2_X1 U1904 ( .A1(n1868), .A2(n1847), .ZN(n1916) );
  XNOR2_X1 U1905 ( .A(n1892), .B(n1918), .ZN(n1847) );
  XNOR2_X1 U1906 ( .A(n1919), .B(n1920), .ZN(n1892) );
  XOR2_X1 U1907 ( .A(n1897), .B(n1921), .Z(n1868) );
  XNOR2_X1 U1908 ( .A(n1787), .B(n1808), .ZN(n1915) );
  XNOR2_X1 U1909 ( .A(n1922), .B(n1835), .ZN(n1808) );
  XNOR2_X1 U1910 ( .A(n1897), .B(n1923), .ZN(n1835) );
  XOR2_X1 U1911 ( .A(n1924), .B(n1925), .Z(n1897) );
  NAND2_X1 U1912 ( .A1(n1834), .A2(n1865), .ZN(n1922) );
  XOR2_X1 U1913 ( .A(n1887), .B(n1926), .Z(n1865) );
  XOR2_X1 U1914 ( .A(n1885), .B(n1927), .Z(n1834) );
  XNOR2_X1 U1915 ( .A(n1928), .B(n1852), .ZN(n1787) );
  XNOR2_X1 U1916 ( .A(n1885), .B(n1929), .ZN(n1852) );
  XNOR2_X1 U1917 ( .A(n1930), .B(n1919), .ZN(n1885) );
  XNOR2_X1 U1918 ( .A(n1931), .B(n1932), .ZN(n1919) );
  XOR2_X1 U1919 ( .A(n1901), .B(n1923), .Z(n1932) );
  XNOR2_X1 U1920 ( .A(n1933), .B(n1934), .ZN(n1923) );
  NAND2_X1 U1921 ( .A1(n1935), .A2(n1936), .ZN(n1933) );
  XOR2_X1 U1922 ( .A(n1937), .B(n1938), .Z(n1901) );
  NAND2_X1 U1923 ( .A1(n1939), .A2(n1940), .ZN(n1937) );
  XOR2_X1 U1924 ( .A(n1941), .B(n1898), .Z(n1931) );
  XOR2_X1 U1925 ( .A(n1942), .B(n1943), .Z(n1898) );
  NAND2_X1 U1926 ( .A1(n1944), .A2(n1945), .ZN(n1942) );
  XNOR2_X1 U1927 ( .A(n1921), .B(n1910), .ZN(n1941) );
  XNOR2_X1 U1928 ( .A(n1946), .B(n1947), .ZN(n1910) );
  NAND2_X1 U1929 ( .A1(n1948), .A2(n1949), .ZN(n1946) );
  XOR2_X1 U1930 ( .A(n1950), .B(n1951), .Z(n1921) );
  NAND2_X1 U1931 ( .A1(n1952), .A2(n1953), .ZN(n1950) );
  NAND2_X1 U1932 ( .A1(n1862), .A2(n1851), .ZN(n1928) );
  XNOR2_X1 U1933 ( .A(n1887), .B(n1954), .ZN(n1851) );
  XNOR2_X1 U1934 ( .A(n1925), .B(n1920), .ZN(n1887) );
  XNOR2_X1 U1935 ( .A(n1955), .B(n1956), .ZN(n1920) );
  XOR2_X1 U1936 ( .A(n1904), .B(n1891), .Z(n1956) );
  XOR2_X1 U1937 ( .A(n1957), .B(n1958), .Z(n1891) );
  NAND2_X1 U1938 ( .A1(n1938), .A2(n1959), .ZN(n1957) );
  XNOR2_X1 U1939 ( .A(n1960), .B(n1961), .ZN(n1904) );
  NAND2_X1 U1940 ( .A1(n1943), .A2(n1962), .ZN(n1960) );
  XOR2_X1 U1941 ( .A(n1963), .B(n1964), .Z(n1955) );
  XNOR2_X1 U1942 ( .A(n1917), .B(n1914), .ZN(n1963) );
  XOR2_X1 U1943 ( .A(n1965), .B(n1966), .Z(n1914) );
  NAND2_X1 U1944 ( .A1(n1967), .A2(n1947), .ZN(n1965) );
  XOR2_X1 U1945 ( .A(n1968), .B(n1969), .Z(n1917) );
  NAND2_X1 U1946 ( .A1(n1934), .A2(n1970), .ZN(n1968) );
  XNOR2_X1 U1947 ( .A(n1971), .B(n1972), .ZN(n1925) );
  XOR2_X1 U1948 ( .A(n1927), .B(n1886), .Z(n1972) );
  XNOR2_X1 U1949 ( .A(n1973), .B(n1940), .ZN(n1886) );
  NAND2_X1 U1950 ( .A1(n1939), .A2(n1958), .ZN(n1973) );
  XOR2_X1 U1951 ( .A(n1974), .B(n1948), .Z(n1927) );
  NAND2_X1 U1952 ( .A1(n1949), .A2(n1966), .ZN(n1974) );
  XOR2_X1 U1953 ( .A(n1975), .B(n1909), .Z(n1971) );
  XNOR2_X1 U1954 ( .A(n1976), .B(n1953), .ZN(n1909) );
  NAND2_X1 U1955 ( .A1(n1952), .A2(n1977), .ZN(n1976) );
  XNOR2_X1 U1956 ( .A(n1900), .B(n1929), .ZN(n1975) );
  XNOR2_X1 U1957 ( .A(n1978), .B(n1935), .ZN(n1929) );
  NAND2_X1 U1958 ( .A1(n1969), .A2(n1936), .ZN(n1978) );
  XNOR2_X1 U1959 ( .A(n1979), .B(n1945), .ZN(n1900) );
  NAND2_X1 U1960 ( .A1(n1944), .A2(n1961), .ZN(n1979) );
  XOR2_X1 U1961 ( .A(n1890), .B(n1964), .Z(n1862) );
  XNOR2_X1 U1962 ( .A(n1980), .B(n1977), .ZN(n1964) );
  NAND2_X1 U1963 ( .A1(n1981), .A2(n1951), .ZN(n1980) );
  XNOR2_X1 U1964 ( .A(n1924), .B(n1982), .ZN(n1890) );
  INV_X1 U1965 ( .A(n1930), .ZN(n1982) );
  XNOR2_X1 U1966 ( .A(n1983), .B(n1984), .ZN(n1930) );
  XOR2_X1 U1967 ( .A(n1903), .B(n1888), .Z(n1984) );
  XNOR2_X1 U1968 ( .A(n1985), .B(n1944), .ZN(n1888) );
  XNOR2_X1 U1969 ( .A(n1986), .B(n1987), .ZN(n1944) );
  NAND2_X1 U1970 ( .A1(n1961), .A2(n1962), .ZN(n1985) );
  XNOR2_X1 U1971 ( .A(n1988), .B(n1989), .ZN(n1961) );
  XOR2_X1 U1972 ( .A(n1990), .B(n1939), .Z(n1903) );
  XOR2_X1 U1973 ( .A(n1991), .B(n1992), .Z(n1939) );
  NAND2_X1 U1974 ( .A1(n1958), .A2(n1959), .ZN(n1990) );
  XOR2_X1 U1975 ( .A(n1993), .B(n1994), .Z(n1958) );
  XOR2_X1 U1976 ( .A(n1995), .B(n1926), .Z(n1983) );
  XNOR2_X1 U1977 ( .A(n1996), .B(n1952), .ZN(n1926) );
  XNOR2_X1 U1978 ( .A(n1997), .B(n1998), .ZN(n1952) );
  NAND2_X1 U1979 ( .A1(n1981), .A2(n1977), .ZN(n1996) );
  XNOR2_X1 U1980 ( .A(n1986), .B(n1999), .ZN(n1977) );
  XNOR2_X1 U1981 ( .A(n1912), .B(n1954), .ZN(n1995) );
  XOR2_X1 U1982 ( .A(n2000), .B(n1949), .Z(n1954) );
  XOR2_X1 U1983 ( .A(n1988), .B(n2001), .Z(n1949) );
  NAND2_X1 U1984 ( .A1(n1966), .A2(n1967), .ZN(n2000) );
  XOR2_X1 U1985 ( .A(n1991), .B(n2002), .Z(n1966) );
  XNOR2_X1 U1986 ( .A(n2003), .B(n1936), .ZN(n1912) );
  XNOR2_X1 U1987 ( .A(n1993), .B(n2004), .ZN(n1936) );
  NAND2_X1 U1988 ( .A1(n1969), .A2(n1970), .ZN(n2003) );
  XOR2_X1 U1989 ( .A(n1997), .B(n2005), .Z(n1969) );
  XOR2_X1 U1990 ( .A(n2006), .B(n2007), .Z(n1924) );
  XOR2_X1 U1991 ( .A(n1918), .B(n1893), .Z(n2007) );
  XNOR2_X1 U1992 ( .A(n2008), .B(n1962), .ZN(n1893) );
  XNOR2_X1 U1993 ( .A(n1991), .B(n2009), .ZN(n1962) );
  NAND2_X1 U1994 ( .A1(n1943), .A2(n1945), .ZN(n2008) );
  XNOR2_X1 U1995 ( .A(n1997), .B(n2010), .ZN(n1945) );
  XOR2_X1 U1996 ( .A(n1993), .B(n2011), .Z(n1943) );
  XOR2_X1 U1997 ( .A(n2012), .B(n1967), .Z(n1918) );
  XOR2_X1 U1998 ( .A(n1993), .B(n2013), .Z(n1967) );
  NAND2_X1 U1999 ( .A1(n1948), .A2(n1947), .ZN(n2012) );
  XNOR2_X1 U2000 ( .A(n1997), .B(n2014), .ZN(n1947) );
  XOR2_X1 U2001 ( .A(n1986), .B(n2015), .Z(n1948) );
  XOR2_X1 U2002 ( .A(n2016), .B(n1913), .Z(n2006) );
  XOR2_X1 U2003 ( .A(n2017), .B(n1981), .Z(n1913) );
  XOR2_X1 U2004 ( .A(n1988), .B(n2018), .Z(n1981) );
  NAND2_X1 U2005 ( .A1(n1951), .A2(n1953), .ZN(n2017) );
  XNOR2_X1 U2006 ( .A(n1993), .B(n2019), .ZN(n1953) );
  XOR2_X1 U2007 ( .A(n2020), .B(n2021), .Z(n1993) );
  XOR2_X1 U2008 ( .A(n1991), .B(n2022), .Z(n1951) );
  XNOR2_X1 U2009 ( .A(n1908), .B(n1896), .ZN(n2016) );
  XNOR2_X1 U2010 ( .A(n2023), .B(n1959), .ZN(n1896) );
  XNOR2_X1 U2011 ( .A(n1997), .B(n2024), .ZN(n1959) );
  XNOR2_X1 U2012 ( .A(n2025), .B(n2026), .ZN(n1997) );
  NAND2_X1 U2013 ( .A1(n1938), .A2(n1940), .ZN(n2023) );
  XNOR2_X1 U2014 ( .A(n1988), .B(n2027), .ZN(n1940) );
  XOR2_X1 U2015 ( .A(n1986), .B(n2028), .Z(n1938) );
  XNOR2_X1 U2016 ( .A(n2029), .B(n1970), .ZN(n1908) );
  XNOR2_X1 U2017 ( .A(n1986), .B(n2030), .ZN(n1970) );
  XNOR2_X1 U2018 ( .A(n2021), .B(n2031), .ZN(n1986) );
  XNOR2_X1 U2019 ( .A(n2032), .B(n2033), .ZN(n2021) );
  XOR2_X1 U2020 ( .A(n1998), .B(n2024), .Z(n2033) );
  XNOR2_X1 U2021 ( .A(n2034), .B(n2035), .ZN(n2024) );
  NAND2_X1 U2022 ( .A1(n2036), .A2(n2037), .ZN(n2034) );
  XNOR2_X1 U2023 ( .A(n2038), .B(n2039), .ZN(n1998) );
  NAND2_X1 U2024 ( .A1(n2040), .A2(n2041), .ZN(n2038) );
  XOR2_X1 U2025 ( .A(n2042), .B(n2005), .Z(n2032) );
  XOR2_X1 U2026 ( .A(n2043), .B(n2044), .Z(n2005) );
  NAND2_X1 U2027 ( .A1(n2045), .A2(n2046), .ZN(n2043) );
  XNOR2_X1 U2028 ( .A(n2010), .B(n2014), .ZN(n2042) );
  XNOR2_X1 U2029 ( .A(n2047), .B(n2048), .ZN(n2014) );
  NAND2_X1 U2030 ( .A1(n2049), .A2(n2050), .ZN(n2047) );
  XNOR2_X1 U2031 ( .A(n2051), .B(n2052), .ZN(n2010) );
  NAND2_X1 U2032 ( .A1(n2053), .A2(n2054), .ZN(n2051) );
  NAND2_X1 U2033 ( .A1(n1935), .A2(n1934), .ZN(n2029) );
  XNOR2_X1 U2034 ( .A(n1988), .B(n2055), .ZN(n1934) );
  XNOR2_X1 U2035 ( .A(n2020), .B(n2056), .ZN(n1988) );
  INV_X1 U2036 ( .A(n2025), .ZN(n2056) );
  XNOR2_X1 U2037 ( .A(n2057), .B(n2058), .ZN(n2025) );
  XOR2_X1 U2038 ( .A(n2028), .B(n1999), .Z(n2058) );
  XOR2_X1 U2039 ( .A(n2059), .B(n2046), .Z(n1999) );
  NAND2_X1 U2040 ( .A1(n2060), .A2(n2045), .ZN(n2059) );
  XNOR2_X1 U2041 ( .A(n2061), .B(n2050), .ZN(n2028) );
  NAND2_X1 U2042 ( .A1(n2062), .A2(n2049), .ZN(n2061) );
  XOR2_X1 U2043 ( .A(n2063), .B(n2030), .Z(n2057) );
  XOR2_X1 U2044 ( .A(n2064), .B(n2036), .Z(n2030) );
  NAND2_X1 U2045 ( .A1(n2065), .A2(n2037), .ZN(n2064) );
  XNOR2_X1 U2046 ( .A(n1987), .B(n2015), .ZN(n2063) );
  XNOR2_X1 U2047 ( .A(n2066), .B(n2054), .ZN(n2015) );
  NAND2_X1 U2048 ( .A1(n2053), .A2(n2067), .ZN(n2066) );
  XOR2_X1 U2049 ( .A(n2068), .B(n2040), .Z(n1987) );
  NAND2_X1 U2050 ( .A1(n2069), .A2(n2041), .ZN(n2068) );
  XOR2_X1 U2051 ( .A(n2070), .B(n2071), .Z(n2020) );
  XOR2_X1 U2052 ( .A(n2009), .B(n2022), .Z(n2071) );
  XOR2_X1 U2053 ( .A(n2072), .B(n2062), .Z(n2022) );
  NAND2_X1 U2054 ( .A1(n2073), .A2(n2048), .ZN(n2072) );
  XNOR2_X1 U2055 ( .A(n2074), .B(n2065), .ZN(n2009) );
  NAND2_X1 U2056 ( .A1(n2075), .A2(n2035), .ZN(n2074) );
  XOR2_X1 U2057 ( .A(n2076), .B(n1992), .Z(n2070) );
  XOR2_X1 U2058 ( .A(n2077), .B(n2069), .Z(n1992) );
  NAND2_X1 U2059 ( .A1(n2078), .A2(n2039), .ZN(n2077) );
  XNOR2_X1 U2060 ( .A(n2079), .B(n2002), .ZN(n2076) );
  XOR2_X1 U2061 ( .A(n2080), .B(n2060), .Z(n2002) );
  NAND2_X1 U2062 ( .A1(n2044), .A2(n2081), .ZN(n2080) );
  XNOR2_X1 U2063 ( .A(n1991), .B(n2079), .ZN(n1935) );
  XNOR2_X1 U2064 ( .A(n2082), .B(n2067), .ZN(n2079) );
  NAND2_X1 U2065 ( .A1(n2083), .A2(n2052), .ZN(n2082) );
  XNOR2_X1 U2066 ( .A(n2026), .B(n2031), .ZN(n1991) );
  XNOR2_X1 U2067 ( .A(n2084), .B(n2085), .ZN(n2031) );
  XOR2_X1 U2068 ( .A(n2027), .B(n2018), .Z(n2085) );
  XNOR2_X1 U2069 ( .A(n2086), .B(n2037), .ZN(n2018) );
  XNOR2_X1 U2070 ( .A(n2087), .B(n2088), .ZN(n2037) );
  NAND2_X1 U2071 ( .A1(n2065), .A2(n2075), .ZN(n2086) );
  XNOR2_X1 U2072 ( .A(n2089), .B(n2090), .ZN(n2065) );
  XOR2_X1 U2073 ( .A(n2091), .B(n2053), .Z(n2027) );
  XOR2_X1 U2074 ( .A(n2089), .B(n2092), .Z(n2053) );
  NAND2_X1 U2075 ( .A1(n2083), .A2(n2067), .ZN(n2091) );
  XNOR2_X1 U2076 ( .A(n2093), .B(n2094), .ZN(n2067) );
  XOR2_X1 U2077 ( .A(n2095), .B(n1989), .Z(n2084) );
  XOR2_X1 U2078 ( .A(n2096), .B(n2045), .Z(n1989) );
  XOR2_X1 U2079 ( .A(n2093), .B(n2097), .Z(n2045) );
  NAND2_X1 U2080 ( .A1(n2060), .A2(n2081), .ZN(n2096) );
  XOR2_X1 U2081 ( .A(n2098), .B(n2099), .Z(n2060) );
  XNOR2_X1 U2082 ( .A(n2055), .B(n2001), .ZN(n2095) );
  XNOR2_X1 U2083 ( .A(n2100), .B(n2041), .ZN(n2001) );
  XNOR2_X1 U2084 ( .A(n2101), .B(n2102), .ZN(n2041) );
  NAND2_X1 U2085 ( .A1(n2069), .A2(n2078), .ZN(n2100) );
  XOR2_X1 U2086 ( .A(n2087), .B(n2103), .Z(n2069) );
  XOR2_X1 U2087 ( .A(n2104), .B(n2049), .Z(n2055) );
  XOR2_X1 U2088 ( .A(n2098), .B(n2105), .Z(n2049) );
  NAND2_X1 U2089 ( .A1(n2062), .A2(n2073), .ZN(n2104) );
  XOR2_X1 U2090 ( .A(n2101), .B(n2106), .Z(n2062) );
  XNOR2_X1 U2091 ( .A(n2107), .B(n2108), .ZN(n2026) );
  XOR2_X1 U2092 ( .A(n2013), .B(n2011), .Z(n2108) );
  XNOR2_X1 U2093 ( .A(n2109), .B(n2073), .ZN(n2011) );
  XNOR2_X1 U2094 ( .A(n2087), .B(n2110), .ZN(n2073) );
  NAND2_X1 U2095 ( .A1(n2048), .A2(n2050), .ZN(n2109) );
  XNOR2_X1 U2096 ( .A(n2093), .B(n2111), .ZN(n2050) );
  XNOR2_X1 U2097 ( .A(n2089), .B(n2112), .ZN(n2048) );
  XNOR2_X1 U2098 ( .A(n2113), .B(n2075), .ZN(n2013) );
  XNOR2_X1 U2099 ( .A(n2093), .B(n2114), .ZN(n2075) );
  NAND2_X1 U2100 ( .A1(n2036), .A2(n2035), .ZN(n2113) );
  XNOR2_X1 U2101 ( .A(n2098), .B(n2115), .ZN(n2035) );
  XOR2_X1 U2102 ( .A(n2101), .B(n2116), .Z(n2036) );
  XOR2_X1 U2103 ( .A(n2117), .B(n2004), .Z(n2107) );
  XOR2_X1 U2104 ( .A(n2118), .B(n2078), .Z(n2004) );
  XOR2_X1 U2105 ( .A(n2089), .B(n2119), .Z(n2078) );
  NAND2_X1 U2106 ( .A1(n2040), .A2(n2039), .ZN(n2118) );
  XNOR2_X1 U2107 ( .A(n2093), .B(n2120), .ZN(n2039) );
  XOR2_X1 U2108 ( .A(n2121), .B(n2122), .Z(n2093) );
  XOR2_X1 U2109 ( .A(n2098), .B(n2123), .Z(n2040) );
  XNOR2_X1 U2110 ( .A(n2019), .B(n1994), .ZN(n2117) );
  XNOR2_X1 U2111 ( .A(n2124), .B(n2081), .ZN(n1994) );
  XNOR2_X1 U2112 ( .A(n2101), .B(n2125), .ZN(n2081) );
  NAND2_X1 U2113 ( .A1(n2044), .A2(n2046), .ZN(n2124) );
  XOR2_X1 U2114 ( .A(n2089), .B(n2126), .Z(n2046) );
  XOR2_X1 U2115 ( .A(n2127), .B(n2128), .Z(n2089) );
  XOR2_X1 U2116 ( .A(n2087), .B(n2129), .Z(n2044) );
  XOR2_X1 U2117 ( .A(n2130), .B(n2083), .Z(n2019) );
  XOR2_X1 U2118 ( .A(n2098), .B(n2131), .Z(n2083) );
  XNOR2_X1 U2119 ( .A(n2132), .B(n2128), .ZN(n2098) );
  XNOR2_X1 U2120 ( .A(n2133), .B(n2134), .ZN(n2128) );
  XOR2_X1 U2121 ( .A(n2097), .B(n2094), .Z(n2134) );
  XOR2_X1 U2122 ( .A(n2135), .B(n2136), .Z(n2094) );
  NAND2_X1 U2123 ( .A1(n2137), .A2(n2138), .ZN(n2135) );
  XNOR2_X1 U2124 ( .A(n2139), .B(n2140), .ZN(n2097) );
  NAND2_X1 U2125 ( .A1(n2141), .A2(n2142), .ZN(n2139) );
  XOR2_X1 U2126 ( .A(n2143), .B(n2111), .Z(n2133) );
  XOR2_X1 U2127 ( .A(n2144), .B(n2145), .Z(n2111) );
  NAND2_X1 U2128 ( .A1(n2146), .A2(n2147), .ZN(n2144) );
  XNOR2_X1 U2129 ( .A(n2120), .B(n2114), .ZN(n2143) );
  XOR2_X1 U2130 ( .A(n2148), .B(n2149), .Z(n2114) );
  NAND2_X1 U2131 ( .A1(n2150), .A2(n2151), .ZN(n2148) );
  XOR2_X1 U2132 ( .A(n2152), .B(n2153), .Z(n2120) );
  NAND2_X1 U2133 ( .A1(n2154), .A2(n2155), .ZN(n2152) );
  NAND2_X1 U2134 ( .A1(n2052), .A2(n2054), .ZN(n2130) );
  XNOR2_X1 U2135 ( .A(n2087), .B(n2156), .ZN(n2054) );
  XNOR2_X1 U2136 ( .A(n2121), .B(n2157), .ZN(n2087) );
  INV_X1 U2137 ( .A(n2132), .ZN(n2157) );
  XNOR2_X1 U2138 ( .A(n2158), .B(n2159), .ZN(n2132) );
  XOR2_X1 U2139 ( .A(n2106), .B(n2102), .Z(n2159) );
  XOR2_X1 U2140 ( .A(n2160), .B(n2142), .Z(n2102) );
  NAND2_X1 U2141 ( .A1(n2161), .A2(n2162), .ZN(n2160) );
  XNOR2_X1 U2142 ( .A(n2163), .B(n2138), .ZN(n2106) );
  NAND2_X1 U2143 ( .A1(n2164), .A2(n2165), .ZN(n2163) );
  XOR2_X1 U2144 ( .A(n2166), .B(n2116), .Z(n2158) );
  XNOR2_X1 U2145 ( .A(n2167), .B(n2147), .ZN(n2116) );
  NAND2_X1 U2146 ( .A1(n2168), .A2(n2169), .ZN(n2167) );
  XNOR2_X1 U2147 ( .A(n2125), .B(n2170), .ZN(n2166) );
  XOR2_X1 U2148 ( .A(n2171), .B(n2151), .Z(n2125) );
  NAND2_X1 U2149 ( .A1(n2172), .A2(n2173), .ZN(n2171) );
  XOR2_X1 U2150 ( .A(n2174), .B(n2175), .Z(n2121) );
  XOR2_X1 U2151 ( .A(n2092), .B(n2090), .Z(n2175) );
  XOR2_X1 U2152 ( .A(n2176), .B(n2165), .Z(n2090) );
  NAND2_X1 U2153 ( .A1(n2137), .A2(n2136), .ZN(n2176) );
  XNOR2_X1 U2154 ( .A(n2177), .B(n2162), .ZN(n2092) );
  NAND2_X1 U2155 ( .A1(n2141), .A2(n2140), .ZN(n2177) );
  XOR2_X1 U2156 ( .A(n2178), .B(n2112), .Z(n2174) );
  XOR2_X1 U2157 ( .A(n2179), .B(n2180), .Z(n2112) );
  NAND2_X1 U2158 ( .A1(n2153), .A2(n2155), .ZN(n2179) );
  XNOR2_X1 U2159 ( .A(n2119), .B(n2126), .ZN(n2178) );
  XNOR2_X1 U2160 ( .A(n2181), .B(n2169), .ZN(n2126) );
  NAND2_X1 U2161 ( .A1(n2146), .A2(n2145), .ZN(n2181) );
  XNOR2_X1 U2162 ( .A(n2182), .B(n2173), .ZN(n2119) );
  NAND2_X1 U2163 ( .A1(n2150), .A2(n2149), .ZN(n2182) );
  XNOR2_X1 U2164 ( .A(n2101), .B(n2170), .ZN(n2052) );
  XOR2_X1 U2165 ( .A(n2183), .B(n2154), .Z(n2170) );
  NAND2_X1 U2166 ( .A1(n2184), .A2(n2180), .ZN(n2183) );
  XOR2_X1 U2167 ( .A(n2127), .B(n2122), .Z(n2101) );
  XNOR2_X1 U2168 ( .A(n2185), .B(n2186), .ZN(n2122) );
  XOR2_X1 U2169 ( .A(n2123), .B(n2105), .Z(n2186) );
  XOR2_X1 U2170 ( .A(n2187), .B(n2141), .Z(n2105) );
  XOR2_X1 U2171 ( .A(n2188), .B(n2189), .Z(n2141) );
  NAND2_X1 U2172 ( .A1(n2142), .A2(n2161), .ZN(n2187) );
  XOR2_X1 U2173 ( .A(n2190), .B(n2191), .Z(n2142) );
  XOR2_X1 U2174 ( .A(n2192), .B(n2146), .Z(n2123) );
  XOR2_X1 U2175 ( .A(n2193), .B(n2194), .Z(n2146) );
  NAND2_X1 U2176 ( .A1(n2147), .A2(n2168), .ZN(n2192) );
  XNOR2_X1 U2177 ( .A(n2195), .B(n2196), .ZN(n2147) );
  XOR2_X1 U2178 ( .A(n2197), .B(n2131), .Z(n2185) );
  XOR2_X1 U2179 ( .A(n2198), .B(n2150), .Z(n2131) );
  XOR2_X1 U2180 ( .A(n2190), .B(n2199), .Z(n2150) );
  NAND2_X1 U2181 ( .A1(n2151), .A2(n2172), .ZN(n2198) );
  XOR2_X1 U2182 ( .A(n2193), .B(n2200), .Z(n2151) );
  XNOR2_X1 U2183 ( .A(n2115), .B(n2099), .ZN(n2197) );
  XOR2_X1 U2184 ( .A(n2201), .B(n2137), .Z(n2099) );
  XOR2_X1 U2185 ( .A(n2195), .B(n2202), .Z(n2137) );
  NAND2_X1 U2186 ( .A1(n2164), .A2(n2138), .ZN(n2201) );
  XNOR2_X1 U2187 ( .A(n2203), .B(n2204), .ZN(n2138) );
  XNOR2_X1 U2188 ( .A(n2205), .B(n2155), .ZN(n2115) );
  XNOR2_X1 U2189 ( .A(n2203), .B(n2206), .ZN(n2155) );
  NAND2_X1 U2190 ( .A1(n2154), .A2(n2184), .ZN(n2205) );
  XOR2_X1 U2191 ( .A(n2188), .B(n2207), .Z(n2154) );
  XOR2_X1 U2192 ( .A(n2208), .B(n2209), .Z(n2127) );
  XOR2_X1 U2193 ( .A(n2088), .B(n2103), .Z(n2209) );
  XOR2_X1 U2194 ( .A(n2210), .B(n2164), .Z(n2103) );
  XOR2_X1 U2195 ( .A(n2188), .B(n2211), .Z(n2164) );
  NAND2_X1 U2196 ( .A1(n2165), .A2(n2136), .ZN(n2210) );
  XOR2_X1 U2197 ( .A(n2193), .B(n2212), .Z(n2136) );
  XOR2_X1 U2198 ( .A(n2190), .B(n2213), .Z(n2165) );
  XNOR2_X1 U2199 ( .A(n2214), .B(n2161), .ZN(n2088) );
  XNOR2_X1 U2200 ( .A(n2193), .B(n2215), .ZN(n2161) );
  NAND2_X1 U2201 ( .A1(n2162), .A2(n2140), .ZN(n2214) );
  XNOR2_X1 U2202 ( .A(n2203), .B(n2216), .ZN(n2140) );
  XNOR2_X1 U2203 ( .A(n2195), .B(n2217), .ZN(n2162) );
  XOR2_X1 U2204 ( .A(n2218), .B(n2110), .Z(n2208) );
  XNOR2_X1 U2205 ( .A(n2219), .B(n2172), .ZN(n2110) );
  XNOR2_X1 U2206 ( .A(n2195), .B(n2220), .ZN(n2172) );
  NAND2_X1 U2207 ( .A1(n2149), .A2(n2173), .ZN(n2219) );
  XNOR2_X1 U2208 ( .A(n2203), .B(n2221), .ZN(n2173) );
  XOR2_X1 U2209 ( .A(n2188), .B(n2222), .Z(n2149) );
  XNOR2_X1 U2210 ( .A(n2156), .B(n2129), .ZN(n2218) );
  XOR2_X1 U2211 ( .A(n2223), .B(n2184), .Z(n2129) );
  XOR2_X1 U2212 ( .A(n2190), .B(n2224), .Z(n2184) );
  NAND2_X1 U2213 ( .A1(n2180), .A2(n2153), .ZN(n2223) );
  XOR2_X1 U2214 ( .A(n2195), .B(n2225), .Z(n2153) );
  XOR2_X1 U2215 ( .A(n2226), .B(n2227), .Z(n2195) );
  XOR2_X1 U2216 ( .A(n2193), .B(n2228), .Z(n2180) );
  XNOR2_X1 U2217 ( .A(n2229), .B(n2230), .ZN(n2193) );
  XNOR2_X1 U2218 ( .A(n2231), .B(n2168), .ZN(n2156) );
  XNOR2_X1 U2219 ( .A(n2203), .B(n2232), .ZN(n2168) );
  XNOR2_X1 U2220 ( .A(n2233), .B(n2234), .ZN(n2203) );
  INV_X1 U2221 ( .A(n2229), .ZN(n2234) );
  XNOR2_X1 U2222 ( .A(n2235), .B(n2236), .ZN(n2229) );
  XOR2_X1 U2223 ( .A(n2202), .B(n2225), .Z(n2236) );
  AND2_X1 U2224 ( .A1(n2237), .A2(n2238), .ZN(n2225) );
  NAND2_X1 U2225 ( .A1(n2239), .A2(n2240), .ZN(n2238) );
  NOR2_X1 U2226 ( .A1(n2241), .A2(n2242), .ZN(n2239) );
  NAND2_X1 U2227 ( .A1(n2243), .A2(n2244), .ZN(n2237) );
  NAND2_X1 U2228 ( .A1(n2241), .A2(n2240), .ZN(n2244) );
  AND2_X1 U2229 ( .A1(n2245), .A2(n2246), .ZN(n2202) );
  NAND2_X1 U2230 ( .A1(n2247), .A2(n2248), .ZN(n2246) );
  NOR2_X1 U2231 ( .A1(n2249), .A2(n2250), .ZN(n2247) );
  NAND2_X1 U2232 ( .A1(n2251), .A2(n2252), .ZN(n2245) );
  NAND2_X1 U2233 ( .A1(n2249), .A2(n2248), .ZN(n2252) );
  INV_X1 U2234 ( .A(n2253), .ZN(n2248) );
  XNOR2_X1 U2235 ( .A(n2217), .B(n2254), .ZN(n2235) );
  XOR2_X1 U2236 ( .A(n2196), .B(n2220), .Z(n2254) );
  AND2_X1 U2237 ( .A1(n2255), .A2(n2256), .ZN(n2220) );
  NAND2_X1 U2238 ( .A1(n2250), .A2(n2257), .ZN(n2256) );
  NAND2_X1 U2239 ( .A1(n2258), .A2(n2243), .ZN(n2257) );
  NAND2_X1 U2240 ( .A1(n2259), .A2(n2258), .ZN(n2255) );
  INV_X1 U2241 ( .A(n2260), .ZN(n2258) );
  AND2_X1 U2242 ( .A1(n2261), .A2(n2262), .ZN(n2196) );
  NAND2_X1 U2243 ( .A1(n2242), .A2(n2263), .ZN(n2262) );
  NAND2_X1 U2244 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  NAND2_X1 U2245 ( .A1(n2266), .A2(n2265), .ZN(n2261) );
  INV_X1 U2246 ( .A(n2267), .ZN(n2265) );
  AND2_X1 U2247 ( .A1(n2268), .A2(n2269), .ZN(n2217) );
  NAND2_X1 U2248 ( .A1(n2270), .A2(n2271), .ZN(n2269) );
  NAND2_X1 U2249 ( .A1(n2251), .A2(n2272), .ZN(n2271) );
  NAND2_X1 U2250 ( .A1(n2273), .A2(n2272), .ZN(n2268) );
  INV_X1 U2251 ( .A(n2274), .ZN(n2272) );
  NAND2_X1 U2252 ( .A1(n2145), .A2(n2169), .ZN(n2231) );
  XNOR2_X1 U2253 ( .A(n2188), .B(n2275), .ZN(n2169) );
  XOR2_X1 U2254 ( .A(n2226), .B(n2230), .Z(n2188) );
  XNOR2_X1 U2255 ( .A(n2276), .B(n2277), .ZN(n2230) );
  XNOR2_X1 U2256 ( .A(n2224), .B(n2278), .ZN(n2277) );
  XNOR2_X1 U2257 ( .A(n2213), .B(n2199), .ZN(n2278) );
  XNOR2_X1 U2258 ( .A(n2279), .B(n2273), .ZN(n2199) );
  XNOR2_X1 U2259 ( .A(n2280), .B(n2266), .ZN(n2213) );
  XOR2_X1 U2260 ( .A(n2281), .B(n2282), .Z(n2224) );
  XNOR2_X1 U2261 ( .A(n2283), .B(n2191), .ZN(n2276) );
  XNOR2_X1 U2262 ( .A(n2284), .B(n2241), .ZN(n2191) );
  XOR2_X1 U2263 ( .A(n2285), .B(n2286), .Z(n2226) );
  XOR2_X1 U2264 ( .A(n2216), .B(n2232), .Z(n2286) );
  XNOR2_X1 U2265 ( .A(n2287), .B(n2288), .ZN(n2232) );
  NOR2_X1 U2266 ( .A1(n2260), .A2(n2281), .ZN(n2288) );
  XNOR2_X1 U2267 ( .A(n2242), .B(n2289), .ZN(n2216) );
  NOR2_X1 U2268 ( .A1(n2290), .A2(n2291), .ZN(n2289) );
  XOR2_X1 U2269 ( .A(n2292), .B(n2206), .Z(n2285) );
  XNOR2_X1 U2270 ( .A(n2250), .B(n2293), .ZN(n2206) );
  NOR2_X1 U2271 ( .A1(n2253), .A2(n2279), .ZN(n2293) );
  XNOR2_X1 U2272 ( .A(n2204), .B(n2221), .ZN(n2292) );
  XNOR2_X1 U2273 ( .A(n2294), .B(n2295), .ZN(n2221) );
  NOR2_X1 U2274 ( .A1(n2280), .A2(n2274), .ZN(n2295) );
  XOR2_X1 U2275 ( .A(n2264), .B(n2296), .Z(n2204) );
  NOR2_X1 U2276 ( .A1(n2267), .A2(n2284), .ZN(n2296) );
  XNOR2_X1 U2277 ( .A(n2190), .B(n2297), .ZN(n2145) );
  INV_X1 U2278 ( .A(n2283), .ZN(n2297) );
  XNOR2_X1 U2279 ( .A(n2291), .B(n2259), .ZN(n2283) );
  XOR2_X1 U2280 ( .A(n2233), .B(n2227), .Z(n2190) );
  XNOR2_X1 U2281 ( .A(n2298), .B(n2299), .ZN(n2227) );
  XOR2_X1 U2282 ( .A(n2212), .B(n2194), .Z(n2299) );
  XNOR2_X1 U2283 ( .A(n2282), .B(n2264), .ZN(n2194) );
  XOR2_X1 U2284 ( .A(n2241), .B(n2300), .Z(n2212) );
  XOR2_X1 U2285 ( .A(n2301), .B(n2228), .Z(n2298) );
  XOR2_X1 U2286 ( .A(n2273), .B(n2302), .Z(n2228) );
  NOR2_X1 U2287 ( .A1(n2270), .A2(n2294), .ZN(n2273) );
  XNOR2_X1 U2288 ( .A(n2215), .B(n2200), .ZN(n2301) );
  AND2_X1 U2289 ( .A1(n2303), .A2(n2304), .ZN(n2200) );
  OR2_X1 U2290 ( .A1(n2243), .A2(n2266), .ZN(n2304) );
  NOR2_X1 U2291 ( .A1(n2270), .A2(n2242), .ZN(n2266) );
  NAND2_X1 U2292 ( .A1(n2241), .A2(n2264), .ZN(n2303) );
  NOR2_X1 U2293 ( .A1(n2242), .A2(n2287), .ZN(n2241) );
  AND2_X1 U2294 ( .A1(n2305), .A2(n2306), .ZN(n2215) );
  NAND2_X1 U2295 ( .A1(n2251), .A2(n2307), .ZN(n2306) );
  NAND2_X1 U2296 ( .A1(n2249), .A2(n2243), .ZN(n2307) );
  NAND2_X1 U2297 ( .A1(n2259), .A2(n2282), .ZN(n2305) );
  INV_X1 U2298 ( .A(n2249), .ZN(n2282) );
  NOR2_X1 U2299 ( .A1(n2294), .A2(n2250), .ZN(n2249) );
  NOR2_X1 U2300 ( .A1(n2250), .A2(n2287), .ZN(n2259) );
  XOR2_X1 U2301 ( .A(n2308), .B(n2309), .Z(n2233) );
  XOR2_X1 U2302 ( .A(n2207), .B(n2211), .Z(n2309) );
  XNOR2_X1 U2303 ( .A(n2260), .B(n2310), .ZN(n2211) );
  NOR2_X1 U2304 ( .A1(n2294), .A2(n2281), .ZN(n2310) );
  XNOR2_X1 U2305 ( .A(io_block_i0[8]), .B(n2264), .ZN(n2281) );
  XOR2_X1 U2306 ( .A(io_block_i0[2]), .B(n2242), .Z(n2260) );
  XNOR2_X1 U2307 ( .A(n2267), .B(n2311), .ZN(n2207) );
  NOR2_X1 U2308 ( .A1(n2287), .A2(n2284), .ZN(n2311) );
  XNOR2_X1 U2309 ( .A(io_block_i0[5]), .B(n2300), .ZN(n2284) );
  XOR2_X1 U2310 ( .A(io_block_i0[4]), .B(n2294), .Z(n2267) );
  INV_X1 U2311 ( .A(n2251), .ZN(n2294) );
  XOR2_X1 U2312 ( .A(n2312), .B(n2189), .Z(n2308) );
  XNOR2_X1 U2313 ( .A(n2253), .B(n2313), .ZN(n2189) );
  NOR2_X1 U2314 ( .A1(n2270), .A2(n2279), .ZN(n2313) );
  XNOR2_X1 U2315 ( .A(io_block_i0[7]), .B(n2302), .ZN(n2279) );
  XOR2_X1 U2316 ( .A(io_block_i0[1]), .B(n2287), .Z(n2253) );
  INV_X1 U2317 ( .A(n2243), .ZN(n2287) );
  XNOR2_X1 U2318 ( .A(n2222), .B(n2275), .ZN(n2312) );
  XNOR2_X1 U2319 ( .A(n2274), .B(n2314), .ZN(n2275) );
  NOR2_X1 U2320 ( .A1(n2280), .A2(n2242), .ZN(n2314) );
  INV_X1 U2321 ( .A(n2302), .ZN(n2242) );
  XOR2_X1 U2322 ( .A(n2315), .B(n2316), .Z(n2302) );
  XNOR2_X1 U2323 ( .A(io_block_i0[6]), .B(n2243), .ZN(n2280) );
  XNOR2_X1 U2324 ( .A(n2317), .B(n2318), .ZN(n2243) );
  XOR2_X1 U2325 ( .A(io_block_i0[0]), .B(n2250), .Z(n2274) );
  XOR2_X1 U2326 ( .A(n2240), .B(n2319), .Z(n2222) );
  NOR2_X1 U2327 ( .A1(n2250), .A2(n2291), .ZN(n2319) );
  XNOR2_X1 U2328 ( .A(io_block_i0[9]), .B(n2251), .ZN(n2291) );
  XNOR2_X1 U2329 ( .A(n2317), .B(n2315), .ZN(n2251) );
  XOR2_X1 U2330 ( .A(io_block_i0[3]), .B(io_block_i0[8]), .Z(n2315) );
  XNOR2_X1 U2331 ( .A(io_block_i0[0]), .B(io_block_i0[5]), .ZN(n2317) );
  INV_X1 U2332 ( .A(n2300), .ZN(n2250) );
  XOR2_X1 U2333 ( .A(n2316), .B(n2320), .Z(n2300) );
  XOR2_X1 U2334 ( .A(io_block_i0[1]), .B(io_block_i0[6]), .Z(n2316) );
  INV_X1 U2335 ( .A(n2290), .ZN(n2240) );
  XOR2_X1 U2336 ( .A(io_block_i0[3]), .B(n2270), .Z(n2290) );
  INV_X1 U2337 ( .A(n2264), .ZN(n2270) );
  XOR2_X1 U2338 ( .A(n2318), .B(n2320), .Z(n2264) );
  XOR2_X1 U2339 ( .A(io_block_i0[4]), .B(io_block_i0[9]), .Z(n2320) );
  XOR2_X1 U2340 ( .A(io_block_i0[2]), .B(io_block_i0[7]), .Z(n2318) );
endmodule

