
module PresentSbox_keyAdd_parallel ( clock, reset, io_state, io_key, io_out );
  input [15:0] io_state;
  input [15:0] io_key;
  output [15:0] io_out;
  input clock, reset;
  wire   PresentSbox_keyAdd_sbox_io_o3, PresentSbox_keyAdd_sbox_io_o2,
         PresentSbox_keyAdd_sbox_io_o1, PresentSbox_keyAdd_sbox_io_o0,
         PresentSbox_keyAdd_sbox_n18, PresentSbox_keyAdd_sbox_n17,
         PresentSbox_keyAdd_sbox_n16, PresentSbox_keyAdd_sbox_n15,
         PresentSbox_keyAdd_sbox_n14, PresentSbox_keyAdd_sbox_n13,
         PresentSbox_keyAdd_sbox_n12, PresentSbox_keyAdd_sbox_n11,
         PresentSbox_keyAdd_sbox_n10, PresentSbox_keyAdd_sbox_n9,
         PresentSbox_keyAdd_sbox_n8, PresentSbox_keyAdd_sbox_n7,
         PresentSbox_keyAdd_sbox_n6, PresentSbox_keyAdd_sbox_n5,
         PresentSbox_keyAdd_sbox_n4, PresentSbox_keyAdd_sbox_n3,
         PresentSbox_keyAdd_sbox_n2, PresentSbox_keyAdd_sbox_n1,
         PresentSbox_keyAdd_1_sbox_io_o3, PresentSbox_keyAdd_1_sbox_io_o2,
         PresentSbox_keyAdd_1_sbox_io_o1, PresentSbox_keyAdd_1_sbox_io_o0,
         PresentSbox_keyAdd_1_sbox_n18, PresentSbox_keyAdd_1_sbox_n17,
         PresentSbox_keyAdd_1_sbox_n16, PresentSbox_keyAdd_1_sbox_n15,
         PresentSbox_keyAdd_1_sbox_n14, PresentSbox_keyAdd_1_sbox_n13,
         PresentSbox_keyAdd_1_sbox_n12, PresentSbox_keyAdd_1_sbox_n11,
         PresentSbox_keyAdd_1_sbox_n10, PresentSbox_keyAdd_1_sbox_n9,
         PresentSbox_keyAdd_1_sbox_n8, PresentSbox_keyAdd_1_sbox_n7,
         PresentSbox_keyAdd_1_sbox_n6, PresentSbox_keyAdd_1_sbox_n5,
         PresentSbox_keyAdd_1_sbox_n4, PresentSbox_keyAdd_1_sbox_n3,
         PresentSbox_keyAdd_1_sbox_n2, PresentSbox_keyAdd_1_sbox_n1,
         PresentSbox_keyAdd_2_sbox_io_o3, PresentSbox_keyAdd_2_sbox_io_o2,
         PresentSbox_keyAdd_2_sbox_io_o1, PresentSbox_keyAdd_2_sbox_io_o0,
         PresentSbox_keyAdd_2_sbox_n18, PresentSbox_keyAdd_2_sbox_n17,
         PresentSbox_keyAdd_2_sbox_n16, PresentSbox_keyAdd_2_sbox_n15,
         PresentSbox_keyAdd_2_sbox_n14, PresentSbox_keyAdd_2_sbox_n13,
         PresentSbox_keyAdd_2_sbox_n12, PresentSbox_keyAdd_2_sbox_n11,
         PresentSbox_keyAdd_2_sbox_n10, PresentSbox_keyAdd_2_sbox_n9,
         PresentSbox_keyAdd_2_sbox_n8, PresentSbox_keyAdd_2_sbox_n7,
         PresentSbox_keyAdd_2_sbox_n6, PresentSbox_keyAdd_2_sbox_n5,
         PresentSbox_keyAdd_2_sbox_n4, PresentSbox_keyAdd_2_sbox_n3,
         PresentSbox_keyAdd_2_sbox_n2, PresentSbox_keyAdd_2_sbox_n1,
         PresentSbox_keyAdd_3_sbox_io_o3, PresentSbox_keyAdd_3_sbox_io_o2,
         PresentSbox_keyAdd_3_sbox_io_o1, PresentSbox_keyAdd_3_sbox_io_o0,
         PresentSbox_keyAdd_3_sbox_n18, PresentSbox_keyAdd_3_sbox_n17,
         PresentSbox_keyAdd_3_sbox_n16, PresentSbox_keyAdd_3_sbox_n15,
         PresentSbox_keyAdd_3_sbox_n14, PresentSbox_keyAdd_3_sbox_n13,
         PresentSbox_keyAdd_3_sbox_n12, PresentSbox_keyAdd_3_sbox_n11,
         PresentSbox_keyAdd_3_sbox_n10, PresentSbox_keyAdd_3_sbox_n9,
         PresentSbox_keyAdd_3_sbox_n8, PresentSbox_keyAdd_3_sbox_n7,
         PresentSbox_keyAdd_3_sbox_n6, PresentSbox_keyAdd_3_sbox_n5,
         PresentSbox_keyAdd_3_sbox_n4, PresentSbox_keyAdd_3_sbox_n3,
         PresentSbox_keyAdd_3_sbox_n2, PresentSbox_keyAdd_3_sbox_n1;

  XOR2_X1 PresentSbox_keyAdd_U4 ( .A(PresentSbox_keyAdd_sbox_io_o0), .B(
        io_key[0]), .Z(io_out[0]) );
  XOR2_X1 PresentSbox_keyAdd_U3 ( .A(PresentSbox_keyAdd_sbox_io_o1), .B(
        io_key[1]), .Z(io_out[1]) );
  XOR2_X1 PresentSbox_keyAdd_U2 ( .A(PresentSbox_keyAdd_sbox_io_o2), .B(
        io_key[2]), .Z(io_out[2]) );
  XOR2_X1 PresentSbox_keyAdd_U1 ( .A(PresentSbox_keyAdd_sbox_io_o3), .B(
        io_key[3]), .Z(io_out[3]) );
  INV_X1 PresentSbox_keyAdd_sbox_U22 ( .A(io_state[1]), .ZN(
        PresentSbox_keyAdd_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U21 ( .A1(PresentSbox_keyAdd_sbox_n18), .A2(
        io_state[2]), .ZN(PresentSbox_keyAdd_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_sbox_U20 ( .A1(io_state[2]), .A2(
        PresentSbox_keyAdd_sbox_n18), .ZN(PresentSbox_keyAdd_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_sbox_U19 ( .A1(PresentSbox_keyAdd_sbox_n1), .A2(
        PresentSbox_keyAdd_sbox_n17), .ZN(PresentSbox_keyAdd_sbox_n13) );
  INV_X1 PresentSbox_keyAdd_sbox_U18 ( .A(io_state[3]), .ZN(
        PresentSbox_keyAdd_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U17 ( .A(PresentSbox_keyAdd_sbox_n13), .B(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n15) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U16 ( .A1(PresentSbox_keyAdd_sbox_n13), .A2(
        io_state[0]), .ZN(PresentSbox_keyAdd_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_sbox_U15 ( .A1(PresentSbox_keyAdd_sbox_n11), .A2(
        PresentSbox_keyAdd_sbox_n1), .ZN(PresentSbox_keyAdd_sbox_n14) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U14 ( .A(io_state[0]), .B(io_state[2]), 
        .ZN(PresentSbox_keyAdd_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U13 ( .A(PresentSbox_keyAdd_sbox_n14), .B(
        PresentSbox_keyAdd_sbox_n4), .Z(PresentSbox_keyAdd_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_sbox_U12 ( .A1(PresentSbox_keyAdd_sbox_n15), 
        .A2(PresentSbox_keyAdd_sbox_n16), .ZN(PresentSbox_keyAdd_sbox_n3) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U11 ( .A(PresentSbox_keyAdd_sbox_n14), .B(
        io_state[3]), .ZN(PresentSbox_keyAdd_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U10 ( .A(PresentSbox_keyAdd_sbox_n3), .B(
        PresentSbox_keyAdd_sbox_n6), .Z(PresentSbox_keyAdd_sbox_io_o0) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U9 ( .A(io_state[0]), .B(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U8 ( .A(PresentSbox_keyAdd_sbox_n13), .B(
        PresentSbox_keyAdd_sbox_n2), .Z(PresentSbox_keyAdd_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U7 ( .A1(PresentSbox_keyAdd_sbox_n11), .A2(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n10) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U6 ( .A(PresentSbox_keyAdd_sbox_n4), .B(
        PresentSbox_keyAdd_sbox_n10), .Z(PresentSbox_keyAdd_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_sbox_U5 ( .A1(PresentSbox_keyAdd_sbox_n8), .A2(
        PresentSbox_keyAdd_sbox_n9), .ZN(PresentSbox_keyAdd_sbox_n7) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U4 ( .A(PresentSbox_keyAdd_sbox_n7), .B(
        io_state[2]), .Z(PresentSbox_keyAdd_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U3 ( .A(PresentSbox_keyAdd_sbox_n5), .B(
        PresentSbox_keyAdd_sbox_n6), .Z(PresentSbox_keyAdd_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U2 ( .A(PresentSbox_keyAdd_sbox_n3), .B(
        PresentSbox_keyAdd_sbox_n4), .Z(PresentSbox_keyAdd_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U1 ( .A(PresentSbox_keyAdd_sbox_n1), .B(
        PresentSbox_keyAdd_sbox_n2), .Z(PresentSbox_keyAdd_sbox_io_o3) );
  XOR2_X1 PresentSbox_keyAdd_1_U4 ( .A(PresentSbox_keyAdd_1_sbox_io_o0), .B(
        io_key[4]), .Z(io_out[4]) );
  XOR2_X1 PresentSbox_keyAdd_1_U3 ( .A(PresentSbox_keyAdd_1_sbox_io_o1), .B(
        io_key[5]), .Z(io_out[5]) );
  XOR2_X1 PresentSbox_keyAdd_1_U2 ( .A(PresentSbox_keyAdd_1_sbox_io_o2), .B(
        io_key[6]), .Z(io_out[6]) );
  XOR2_X1 PresentSbox_keyAdd_1_U1 ( .A(PresentSbox_keyAdd_1_sbox_io_o3), .B(
        io_key[7]), .Z(io_out[7]) );
  INV_X1 PresentSbox_keyAdd_1_sbox_U22 ( .A(io_state[5]), .ZN(
        PresentSbox_keyAdd_1_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U21 ( .A1(PresentSbox_keyAdd_1_sbox_n18), 
        .A2(io_state[6]), .ZN(PresentSbox_keyAdd_1_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_1_sbox_U20 ( .A1(io_state[6]), .A2(
        PresentSbox_keyAdd_1_sbox_n18), .ZN(PresentSbox_keyAdd_1_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U19 ( .A1(PresentSbox_keyAdd_1_sbox_n1), 
        .A2(PresentSbox_keyAdd_1_sbox_n17), .ZN(PresentSbox_keyAdd_1_sbox_n13)
         );
  INV_X1 PresentSbox_keyAdd_1_sbox_U18 ( .A(io_state[7]), .ZN(
        PresentSbox_keyAdd_1_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U17 ( .A(PresentSbox_keyAdd_1_sbox_n13), 
        .B(PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n15)
         );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U16 ( .A1(PresentSbox_keyAdd_1_sbox_n13), 
        .A2(io_state[4]), .ZN(PresentSbox_keyAdd_1_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U15 ( .A1(PresentSbox_keyAdd_1_sbox_n11), 
        .A2(PresentSbox_keyAdd_1_sbox_n1), .ZN(PresentSbox_keyAdd_1_sbox_n14)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U14 ( .A(io_state[4]), .B(io_state[6]), 
        .ZN(PresentSbox_keyAdd_1_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U13 ( .A(PresentSbox_keyAdd_1_sbox_n14), 
        .B(PresentSbox_keyAdd_1_sbox_n4), .Z(PresentSbox_keyAdd_1_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U12 ( .A1(PresentSbox_keyAdd_1_sbox_n15), 
        .A2(PresentSbox_keyAdd_1_sbox_n16), .ZN(PresentSbox_keyAdd_1_sbox_n3)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U11 ( .A(PresentSbox_keyAdd_1_sbox_n14), 
        .B(io_state[7]), .ZN(PresentSbox_keyAdd_1_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U10 ( .A(PresentSbox_keyAdd_1_sbox_n3), 
        .B(PresentSbox_keyAdd_1_sbox_n6), .Z(PresentSbox_keyAdd_1_sbox_io_o0)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U9 ( .A(io_state[4]), .B(
        PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U8 ( .A(PresentSbox_keyAdd_1_sbox_n13), 
        .B(PresentSbox_keyAdd_1_sbox_n2), .Z(PresentSbox_keyAdd_1_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U7 ( .A1(PresentSbox_keyAdd_1_sbox_n11), 
        .A2(PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n10)
         );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U6 ( .A(PresentSbox_keyAdd_1_sbox_n4), .B(
        PresentSbox_keyAdd_1_sbox_n10), .Z(PresentSbox_keyAdd_1_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U5 ( .A1(PresentSbox_keyAdd_1_sbox_n8), 
        .A2(PresentSbox_keyAdd_1_sbox_n9), .ZN(PresentSbox_keyAdd_1_sbox_n7)
         );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U4 ( .A(PresentSbox_keyAdd_1_sbox_n7), .B(
        io_state[6]), .Z(PresentSbox_keyAdd_1_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U3 ( .A(PresentSbox_keyAdd_1_sbox_n5), .B(
        PresentSbox_keyAdd_1_sbox_n6), .Z(PresentSbox_keyAdd_1_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U2 ( .A(PresentSbox_keyAdd_1_sbox_n3), .B(
        PresentSbox_keyAdd_1_sbox_n4), .Z(PresentSbox_keyAdd_1_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U1 ( .A(PresentSbox_keyAdd_1_sbox_n1), .B(
        PresentSbox_keyAdd_1_sbox_n2), .Z(PresentSbox_keyAdd_1_sbox_io_o3) );
  XOR2_X1 PresentSbox_keyAdd_2_U4 ( .A(PresentSbox_keyAdd_2_sbox_io_o0), .B(
        io_key[8]), .Z(io_out[8]) );
  XOR2_X1 PresentSbox_keyAdd_2_U3 ( .A(PresentSbox_keyAdd_2_sbox_io_o1), .B(
        io_key[9]), .Z(io_out[9]) );
  XOR2_X1 PresentSbox_keyAdd_2_U2 ( .A(PresentSbox_keyAdd_2_sbox_io_o2), .B(
        io_key[10]), .Z(io_out[10]) );
  XOR2_X1 PresentSbox_keyAdd_2_U1 ( .A(PresentSbox_keyAdd_2_sbox_io_o3), .B(
        io_key[11]), .Z(io_out[11]) );
  INV_X1 PresentSbox_keyAdd_2_sbox_U22 ( .A(io_state[9]), .ZN(
        PresentSbox_keyAdd_2_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_2_sbox_U21 ( .A1(PresentSbox_keyAdd_2_sbox_n18), 
        .A2(io_state[10]), .ZN(PresentSbox_keyAdd_2_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_2_sbox_U20 ( .A1(io_state[10]), .A2(
        PresentSbox_keyAdd_2_sbox_n18), .ZN(PresentSbox_keyAdd_2_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_2_sbox_U19 ( .A1(PresentSbox_keyAdd_2_sbox_n1), 
        .A2(PresentSbox_keyAdd_2_sbox_n17), .ZN(PresentSbox_keyAdd_2_sbox_n13)
         );
  INV_X1 PresentSbox_keyAdd_2_sbox_U18 ( .A(io_state[11]), .ZN(
        PresentSbox_keyAdd_2_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_2_sbox_U17 ( .A(PresentSbox_keyAdd_2_sbox_n13), 
        .B(PresentSbox_keyAdd_2_sbox_n12), .ZN(PresentSbox_keyAdd_2_sbox_n15)
         );
  NOR2_X1 PresentSbox_keyAdd_2_sbox_U16 ( .A1(PresentSbox_keyAdd_2_sbox_n13), 
        .A2(io_state[8]), .ZN(PresentSbox_keyAdd_2_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_2_sbox_U15 ( .A1(PresentSbox_keyAdd_2_sbox_n11), 
        .A2(PresentSbox_keyAdd_2_sbox_n1), .ZN(PresentSbox_keyAdd_2_sbox_n14)
         );
  XNOR2_X1 PresentSbox_keyAdd_2_sbox_U14 ( .A(io_state[8]), .B(io_state[10]), 
        .ZN(PresentSbox_keyAdd_2_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U13 ( .A(PresentSbox_keyAdd_2_sbox_n14), 
        .B(PresentSbox_keyAdd_2_sbox_n4), .Z(PresentSbox_keyAdd_2_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_2_sbox_U12 ( .A1(PresentSbox_keyAdd_2_sbox_n15), 
        .A2(PresentSbox_keyAdd_2_sbox_n16), .ZN(PresentSbox_keyAdd_2_sbox_n3)
         );
  XNOR2_X1 PresentSbox_keyAdd_2_sbox_U11 ( .A(PresentSbox_keyAdd_2_sbox_n14), 
        .B(io_state[11]), .ZN(PresentSbox_keyAdd_2_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U10 ( .A(PresentSbox_keyAdd_2_sbox_n3), 
        .B(PresentSbox_keyAdd_2_sbox_n6), .Z(PresentSbox_keyAdd_2_sbox_io_o0)
         );
  XNOR2_X1 PresentSbox_keyAdd_2_sbox_U9 ( .A(io_state[8]), .B(
        PresentSbox_keyAdd_2_sbox_n12), .ZN(PresentSbox_keyAdd_2_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U8 ( .A(PresentSbox_keyAdd_2_sbox_n13), 
        .B(PresentSbox_keyAdd_2_sbox_n2), .Z(PresentSbox_keyAdd_2_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_2_sbox_U7 ( .A1(PresentSbox_keyAdd_2_sbox_n11), 
        .A2(PresentSbox_keyAdd_2_sbox_n12), .ZN(PresentSbox_keyAdd_2_sbox_n10)
         );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U6 ( .A(PresentSbox_keyAdd_2_sbox_n4), .B(
        PresentSbox_keyAdd_2_sbox_n10), .Z(PresentSbox_keyAdd_2_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_2_sbox_U5 ( .A1(PresentSbox_keyAdd_2_sbox_n8), 
        .A2(PresentSbox_keyAdd_2_sbox_n9), .ZN(PresentSbox_keyAdd_2_sbox_n7)
         );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U4 ( .A(PresentSbox_keyAdd_2_sbox_n7), .B(
        io_state[10]), .Z(PresentSbox_keyAdd_2_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U3 ( .A(PresentSbox_keyAdd_2_sbox_n5), .B(
        PresentSbox_keyAdd_2_sbox_n6), .Z(PresentSbox_keyAdd_2_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U2 ( .A(PresentSbox_keyAdd_2_sbox_n3), .B(
        PresentSbox_keyAdd_2_sbox_n4), .Z(PresentSbox_keyAdd_2_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_2_sbox_U1 ( .A(PresentSbox_keyAdd_2_sbox_n1), .B(
        PresentSbox_keyAdd_2_sbox_n2), .Z(PresentSbox_keyAdd_2_sbox_io_o3) );
  XOR2_X1 PresentSbox_keyAdd_3_U4 ( .A(PresentSbox_keyAdd_3_sbox_io_o0), .B(
        io_key[12]), .Z(io_out[12]) );
  XOR2_X1 PresentSbox_keyAdd_3_U3 ( .A(PresentSbox_keyAdd_3_sbox_io_o1), .B(
        io_key[13]), .Z(io_out[13]) );
  XOR2_X1 PresentSbox_keyAdd_3_U2 ( .A(PresentSbox_keyAdd_3_sbox_io_o2), .B(
        io_key[14]), .Z(io_out[14]) );
  XOR2_X1 PresentSbox_keyAdd_3_U1 ( .A(PresentSbox_keyAdd_3_sbox_io_o3), .B(
        io_key[15]), .Z(io_out[15]) );
  INV_X1 PresentSbox_keyAdd_3_sbox_U22 ( .A(io_state[13]), .ZN(
        PresentSbox_keyAdd_3_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_3_sbox_U21 ( .A1(PresentSbox_keyAdd_3_sbox_n18), 
        .A2(io_state[14]), .ZN(PresentSbox_keyAdd_3_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_3_sbox_U20 ( .A1(io_state[14]), .A2(
        PresentSbox_keyAdd_3_sbox_n18), .ZN(PresentSbox_keyAdd_3_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_3_sbox_U19 ( .A1(PresentSbox_keyAdd_3_sbox_n1), 
        .A2(PresentSbox_keyAdd_3_sbox_n17), .ZN(PresentSbox_keyAdd_3_sbox_n13)
         );
  INV_X1 PresentSbox_keyAdd_3_sbox_U18 ( .A(io_state[15]), .ZN(
        PresentSbox_keyAdd_3_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_3_sbox_U17 ( .A(PresentSbox_keyAdd_3_sbox_n13), 
        .B(PresentSbox_keyAdd_3_sbox_n12), .ZN(PresentSbox_keyAdd_3_sbox_n15)
         );
  NOR2_X1 PresentSbox_keyAdd_3_sbox_U16 ( .A1(PresentSbox_keyAdd_3_sbox_n13), 
        .A2(io_state[12]), .ZN(PresentSbox_keyAdd_3_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_3_sbox_U15 ( .A1(PresentSbox_keyAdd_3_sbox_n11), 
        .A2(PresentSbox_keyAdd_3_sbox_n1), .ZN(PresentSbox_keyAdd_3_sbox_n14)
         );
  XNOR2_X1 PresentSbox_keyAdd_3_sbox_U14 ( .A(io_state[12]), .B(io_state[14]), 
        .ZN(PresentSbox_keyAdd_3_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U13 ( .A(PresentSbox_keyAdd_3_sbox_n14), 
        .B(PresentSbox_keyAdd_3_sbox_n4), .Z(PresentSbox_keyAdd_3_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_3_sbox_U12 ( .A1(PresentSbox_keyAdd_3_sbox_n15), 
        .A2(PresentSbox_keyAdd_3_sbox_n16), .ZN(PresentSbox_keyAdd_3_sbox_n3)
         );
  XNOR2_X1 PresentSbox_keyAdd_3_sbox_U11 ( .A(PresentSbox_keyAdd_3_sbox_n14), 
        .B(io_state[15]), .ZN(PresentSbox_keyAdd_3_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U10 ( .A(PresentSbox_keyAdd_3_sbox_n3), 
        .B(PresentSbox_keyAdd_3_sbox_n6), .Z(PresentSbox_keyAdd_3_sbox_io_o0)
         );
  XNOR2_X1 PresentSbox_keyAdd_3_sbox_U9 ( .A(io_state[12]), .B(
        PresentSbox_keyAdd_3_sbox_n12), .ZN(PresentSbox_keyAdd_3_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U8 ( .A(PresentSbox_keyAdd_3_sbox_n13), 
        .B(PresentSbox_keyAdd_3_sbox_n2), .Z(PresentSbox_keyAdd_3_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_3_sbox_U7 ( .A1(PresentSbox_keyAdd_3_sbox_n11), 
        .A2(PresentSbox_keyAdd_3_sbox_n12), .ZN(PresentSbox_keyAdd_3_sbox_n10)
         );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U6 ( .A(PresentSbox_keyAdd_3_sbox_n4), .B(
        PresentSbox_keyAdd_3_sbox_n10), .Z(PresentSbox_keyAdd_3_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_3_sbox_U5 ( .A1(PresentSbox_keyAdd_3_sbox_n8), 
        .A2(PresentSbox_keyAdd_3_sbox_n9), .ZN(PresentSbox_keyAdd_3_sbox_n7)
         );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U4 ( .A(PresentSbox_keyAdd_3_sbox_n7), .B(
        io_state[14]), .Z(PresentSbox_keyAdd_3_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U3 ( .A(PresentSbox_keyAdd_3_sbox_n5), .B(
        PresentSbox_keyAdd_3_sbox_n6), .Z(PresentSbox_keyAdd_3_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U2 ( .A(PresentSbox_keyAdd_3_sbox_n3), .B(
        PresentSbox_keyAdd_3_sbox_n4), .Z(PresentSbox_keyAdd_3_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_3_sbox_U1 ( .A(PresentSbox_keyAdd_3_sbox_n1), .B(
        PresentSbox_keyAdd_3_sbox_n2), .Z(PresentSbox_keyAdd_3_sbox_io_o3) );
endmodule

