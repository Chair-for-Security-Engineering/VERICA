
module CINI_HPC3 ( port_a_0, port_a_1, port_a_2, port_a_3, port_b_0, port_b_1, 
        port_b_2, port_b_3, port_c_0, port_c_1, port_c_2, port_c_3, 
        port_rand_ref, port_rand_mul, clk, reset );
  input [4:0] port_a_0;
  input [4:0] port_a_1;
  input [4:0] port_a_2;
  input [4:0] port_a_3;
  input [4:0] port_b_0;
  input [4:0] port_b_1;
  input [4:0] port_b_2;
  input [4:0] port_b_3;
  output [4:0] port_c_0;
  output [4:0] port_c_1;
  output [4:0] port_c_2;
  output [4:0] port_c_3;
  input [5:0] port_rand_ref;
  input [5:0] port_rand_mul;
  input clk, reset;
  wire   simpleAnd_60_port_z, simpleAnd_61_port_z, simpleAnd_62_port_z,
         simpleAnd_63_port_z, simpleAnd_64_port_z, simpleAnd_65_port_z,
         simpleAnd_66_port_z, simpleAnd_67_port_z, simpleAnd_68_port_z,
         simpleAnd_69_port_z, simpleAnd_70_port_z, simpleAnd_71_port_z,
         simpleAnd_72_port_z, simpleAnd_73_port_z, simpleAnd_74_port_z,
         simpleAnd_75_port_z, simpleAnd_76_port_z, simpleAnd_77_port_z,
         simpleAnd_78_port_z, simpleAnd_79_port_z, simpleAnd_80_port_z,
         simpleAnd_81_port_z, simpleAnd_82_port_z, simpleAnd_83_port_z,
         simpleAnd_84_port_z, simpleAnd_85_port_z, simpleAnd_86_port_z,
         simpleAnd_87_port_z, simpleAnd_88_port_z, simpleAnd_89_port_z,
         simpleAnd_90_port_z, simpleAnd_91_port_z, simpleAnd_92_port_z,
         simpleAnd_93_port_z, simpleAnd_94_port_z, simpleAnd_95_port_z,
         simpleAnd_96_port_z, simpleAnd_97_port_z, simpleAnd_98_port_z,
         simpleAnd_99_port_z, simpleAnd_100_port_z, simpleAnd_101_port_z,
         simpleAnd_102_port_z, simpleAnd_103_port_z, simpleAnd_104_port_z,
         simpleAnd_105_port_z, simpleAnd_106_port_z, simpleAnd_107_port_z,
         simpleAnd_108_port_z, simpleAnd_109_port_z, simpleAnd_110_port_z,
         simpleAnd_111_port_z, simpleAnd_112_port_z, simpleAnd_113_port_z,
         simpleAnd_114_port_z, simpleAnd_115_port_z, simpleAnd_116_port_z,
         simpleAnd_117_port_z, simpleAnd_118_port_z, simpleAnd_119_port_z,
         maj_120_port_o, maj_121_port_o, maj_122_port_o, maj_123_port_o,
         maj_124_port_o, maj_125_port_o, maj_126_port_o, maj_127_port_o,
         maj_128_port_o, maj_129_port_o, maj_130_port_o, maj_131_port_o,
         maj_132_port_o, maj_133_port_o, maj_134_port_o, maj_135_port_o,
         maj_136_port_o, maj_137_port_o, maj_138_port_o, maj_139_port_o,
         maj_140_port_o, maj_141_port_o, maj_142_port_o, maj_143_port_o,
         maj_144_port_o, maj_145_port_o, maj_146_port_o, maj_147_port_o,
         maj_148_port_o, maj_149_port_o, maj_150_port_o, maj_151_port_o,
         maj_152_port_o, maj_153_port_o, maj_154_port_o, maj_155_port_o,
         maj_156_port_o, maj_157_port_o, maj_158_port_o, maj_159_port_o,
         maj_160_port_o, maj_161_port_o, maj_162_port_o, maj_163_port_o,
         maj_164_port_o, maj_165_port_o, maj_166_port_o, maj_167_port_o,
         maj_168_port_o, maj_169_port_o, maj_170_port_o, maj_171_port_o,
         maj_172_port_o, maj_173_port_o, maj_174_port_o, maj_175_port_o,
         maj_176_port_o, maj_177_port_o, maj_178_port_o, maj_179_port_o,
         maj_180_port_o, maj_181_port_o, maj_182_port_o, maj_183_port_o,
         maj_184_port_o, maj_185_port_o, maj_186_port_o, maj_187_port_o,
         maj_188_port_o, maj_189_port_o, maj_190_port_o, maj_191_port_o,
         maj_192_port_o, maj_193_port_o, maj_194_port_o, maj_195_port_o,
         maj_196_port_o, maj_197_port_o, maj_198_port_o, maj_199_port_o,
         maj_200_port_o, maj_201_port_o, maj_202_port_o, maj_203_port_o,
         maj_204_port_o, maj_205_port_o, maj_206_port_o, maj_207_port_o,
         maj_208_port_o, maj_209_port_o, maj_210_port_o, maj_211_port_o,
         maj_212_port_o, maj_213_port_o, maj_214_port_o, maj_215_port_o,
         maj_216_port_o, maj_217_port_o, maj_218_port_o, maj_219_port_o,
         maj_220_port_o, maj_221_port_o, maj_222_port_o, maj_223_port_o,
         maj_224_port_o, maj_225_port_o, maj_226_port_o, maj_227_port_o,
         maj_228_port_o, maj_229_port_o, maj_230_port_o, maj_231_port_o,
         maj_232_port_o, maj_233_port_o, maj_234_port_o, maj_235_port_o,
         maj_236_port_o, maj_237_port_o, maj_238_port_o, maj_239_port_o, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, maj_120_n13, maj_120_n12, maj_120_n11,
         maj_120_n10, maj_120_n9, maj_120_n8, maj_120_n7, maj_120_n6,
         maj_120_n5, maj_120_n4, maj_120_n3, maj_120_n2, maj_120_n1,
         maj_121_n26, maj_121_n25, maj_121_n24, maj_121_n23, maj_121_n22,
         maj_121_n21, maj_121_n20, maj_121_n19, maj_121_n18, maj_121_n17,
         maj_121_n16, maj_121_n15, maj_121_n14, maj_122_n26, maj_122_n25,
         maj_122_n24, maj_122_n23, maj_122_n22, maj_122_n21, maj_122_n20,
         maj_122_n19, maj_122_n18, maj_122_n17, maj_122_n16, maj_122_n15,
         maj_122_n14, maj_123_n26, maj_123_n25, maj_123_n24, maj_123_n23,
         maj_123_n22, maj_123_n21, maj_123_n20, maj_123_n19, maj_123_n18,
         maj_123_n17, maj_123_n16, maj_123_n15, maj_123_n14, maj_124_n26,
         maj_124_n25, maj_124_n24, maj_124_n23, maj_124_n22, maj_124_n21,
         maj_124_n20, maj_124_n19, maj_124_n18, maj_124_n17, maj_124_n16,
         maj_124_n15, maj_124_n14, maj_125_n26, maj_125_n25, maj_125_n24,
         maj_125_n23, maj_125_n22, maj_125_n21, maj_125_n20, maj_125_n19,
         maj_125_n18, maj_125_n17, maj_125_n16, maj_125_n15, maj_125_n14,
         maj_126_n26, maj_126_n25, maj_126_n24, maj_126_n23, maj_126_n22,
         maj_126_n21, maj_126_n20, maj_126_n19, maj_126_n18, maj_126_n17,
         maj_126_n16, maj_126_n15, maj_126_n14, maj_127_n26, maj_127_n25,
         maj_127_n24, maj_127_n23, maj_127_n22, maj_127_n21, maj_127_n20,
         maj_127_n19, maj_127_n18, maj_127_n17, maj_127_n16, maj_127_n15,
         maj_127_n14, maj_128_n26, maj_128_n25, maj_128_n24, maj_128_n23,
         maj_128_n22, maj_128_n21, maj_128_n20, maj_128_n19, maj_128_n18,
         maj_128_n17, maj_128_n16, maj_128_n15, maj_128_n14, maj_129_n26,
         maj_129_n25, maj_129_n24, maj_129_n23, maj_129_n22, maj_129_n21,
         maj_129_n20, maj_129_n19, maj_129_n18, maj_129_n17, maj_129_n16,
         maj_129_n15, maj_129_n14, maj_130_n26, maj_130_n25, maj_130_n24,
         maj_130_n23, maj_130_n22, maj_130_n21, maj_130_n20, maj_130_n19,
         maj_130_n18, maj_130_n17, maj_130_n16, maj_130_n15, maj_130_n14,
         maj_131_n26, maj_131_n25, maj_131_n24, maj_131_n23, maj_131_n22,
         maj_131_n21, maj_131_n20, maj_131_n19, maj_131_n18, maj_131_n17,
         maj_131_n16, maj_131_n15, maj_131_n14, maj_132_n26, maj_132_n25,
         maj_132_n24, maj_132_n23, maj_132_n22, maj_132_n21, maj_132_n20,
         maj_132_n19, maj_132_n18, maj_132_n17, maj_132_n16, maj_132_n15,
         maj_132_n14, maj_133_n26, maj_133_n25, maj_133_n24, maj_133_n23,
         maj_133_n22, maj_133_n21, maj_133_n20, maj_133_n19, maj_133_n18,
         maj_133_n17, maj_133_n16, maj_133_n15, maj_133_n14, maj_134_n26,
         maj_134_n25, maj_134_n24, maj_134_n23, maj_134_n22, maj_134_n21,
         maj_134_n20, maj_134_n19, maj_134_n18, maj_134_n17, maj_134_n16,
         maj_134_n15, maj_134_n14, maj_135_n26, maj_135_n25, maj_135_n24,
         maj_135_n23, maj_135_n22, maj_135_n21, maj_135_n20, maj_135_n19,
         maj_135_n18, maj_135_n17, maj_135_n16, maj_135_n15, maj_135_n14,
         maj_136_n26, maj_136_n25, maj_136_n24, maj_136_n23, maj_136_n22,
         maj_136_n21, maj_136_n20, maj_136_n19, maj_136_n18, maj_136_n17,
         maj_136_n16, maj_136_n15, maj_136_n14, maj_137_n26, maj_137_n25,
         maj_137_n24, maj_137_n23, maj_137_n22, maj_137_n21, maj_137_n20,
         maj_137_n19, maj_137_n18, maj_137_n17, maj_137_n16, maj_137_n15,
         maj_137_n14, maj_138_n26, maj_138_n25, maj_138_n24, maj_138_n23,
         maj_138_n22, maj_138_n21, maj_138_n20, maj_138_n19, maj_138_n18,
         maj_138_n17, maj_138_n16, maj_138_n15, maj_138_n14, maj_139_n26,
         maj_139_n25, maj_139_n24, maj_139_n23, maj_139_n22, maj_139_n21,
         maj_139_n20, maj_139_n19, maj_139_n18, maj_139_n17, maj_139_n16,
         maj_139_n15, maj_139_n14, maj_140_n26, maj_140_n25, maj_140_n24,
         maj_140_n23, maj_140_n22, maj_140_n21, maj_140_n20, maj_140_n19,
         maj_140_n18, maj_140_n17, maj_140_n16, maj_140_n15, maj_140_n14,
         maj_141_n26, maj_141_n25, maj_141_n24, maj_141_n23, maj_141_n22,
         maj_141_n21, maj_141_n20, maj_141_n19, maj_141_n18, maj_141_n17,
         maj_141_n16, maj_141_n15, maj_141_n14, maj_142_n26, maj_142_n25,
         maj_142_n24, maj_142_n23, maj_142_n22, maj_142_n21, maj_142_n20,
         maj_142_n19, maj_142_n18, maj_142_n17, maj_142_n16, maj_142_n15,
         maj_142_n14, maj_143_n26, maj_143_n25, maj_143_n24, maj_143_n23,
         maj_143_n22, maj_143_n21, maj_143_n20, maj_143_n19, maj_143_n18,
         maj_143_n17, maj_143_n16, maj_143_n15, maj_143_n14, maj_144_n26,
         maj_144_n25, maj_144_n24, maj_144_n23, maj_144_n22, maj_144_n21,
         maj_144_n20, maj_144_n19, maj_144_n18, maj_144_n17, maj_144_n16,
         maj_144_n15, maj_144_n14, maj_145_n26, maj_145_n25, maj_145_n24,
         maj_145_n23, maj_145_n22, maj_145_n21, maj_145_n20, maj_145_n19,
         maj_145_n18, maj_145_n17, maj_145_n16, maj_145_n15, maj_145_n14,
         maj_146_n26, maj_146_n25, maj_146_n24, maj_146_n23, maj_146_n22,
         maj_146_n21, maj_146_n20, maj_146_n19, maj_146_n18, maj_146_n17,
         maj_146_n16, maj_146_n15, maj_146_n14, maj_147_n26, maj_147_n25,
         maj_147_n24, maj_147_n23, maj_147_n22, maj_147_n21, maj_147_n20,
         maj_147_n19, maj_147_n18, maj_147_n17, maj_147_n16, maj_147_n15,
         maj_147_n14, maj_148_n26, maj_148_n25, maj_148_n24, maj_148_n23,
         maj_148_n22, maj_148_n21, maj_148_n20, maj_148_n19, maj_148_n18,
         maj_148_n17, maj_148_n16, maj_148_n15, maj_148_n14, maj_149_n26,
         maj_149_n25, maj_149_n24, maj_149_n23, maj_149_n22, maj_149_n21,
         maj_149_n20, maj_149_n19, maj_149_n18, maj_149_n17, maj_149_n16,
         maj_149_n15, maj_149_n14, maj_150_n26, maj_150_n25, maj_150_n24,
         maj_150_n23, maj_150_n22, maj_150_n21, maj_150_n20, maj_150_n19,
         maj_150_n18, maj_150_n17, maj_150_n16, maj_150_n15, maj_150_n14,
         maj_151_n26, maj_151_n25, maj_151_n24, maj_151_n23, maj_151_n22,
         maj_151_n21, maj_151_n20, maj_151_n19, maj_151_n18, maj_151_n17,
         maj_151_n16, maj_151_n15, maj_151_n14, maj_152_n26, maj_152_n25,
         maj_152_n24, maj_152_n23, maj_152_n22, maj_152_n21, maj_152_n20,
         maj_152_n19, maj_152_n18, maj_152_n17, maj_152_n16, maj_152_n15,
         maj_152_n14, maj_153_n26, maj_153_n25, maj_153_n24, maj_153_n23,
         maj_153_n22, maj_153_n21, maj_153_n20, maj_153_n19, maj_153_n18,
         maj_153_n17, maj_153_n16, maj_153_n15, maj_153_n14, maj_154_n26,
         maj_154_n25, maj_154_n24, maj_154_n23, maj_154_n22, maj_154_n21,
         maj_154_n20, maj_154_n19, maj_154_n18, maj_154_n17, maj_154_n16,
         maj_154_n15, maj_154_n14, maj_155_n26, maj_155_n25, maj_155_n24,
         maj_155_n23, maj_155_n22, maj_155_n21, maj_155_n20, maj_155_n19,
         maj_155_n18, maj_155_n17, maj_155_n16, maj_155_n15, maj_155_n14,
         maj_156_n26, maj_156_n25, maj_156_n24, maj_156_n23, maj_156_n22,
         maj_156_n21, maj_156_n20, maj_156_n19, maj_156_n18, maj_156_n17,
         maj_156_n16, maj_156_n15, maj_156_n14, maj_157_n26, maj_157_n25,
         maj_157_n24, maj_157_n23, maj_157_n22, maj_157_n21, maj_157_n20,
         maj_157_n19, maj_157_n18, maj_157_n17, maj_157_n16, maj_157_n15,
         maj_157_n14, maj_158_n26, maj_158_n25, maj_158_n24, maj_158_n23,
         maj_158_n22, maj_158_n21, maj_158_n20, maj_158_n19, maj_158_n18,
         maj_158_n17, maj_158_n16, maj_158_n15, maj_158_n14, maj_159_n26,
         maj_159_n25, maj_159_n24, maj_159_n23, maj_159_n22, maj_159_n21,
         maj_159_n20, maj_159_n19, maj_159_n18, maj_159_n17, maj_159_n16,
         maj_159_n15, maj_159_n14, maj_160_n26, maj_160_n25, maj_160_n24,
         maj_160_n23, maj_160_n22, maj_160_n21, maj_160_n20, maj_160_n19,
         maj_160_n18, maj_160_n17, maj_160_n16, maj_160_n15, maj_160_n14,
         maj_161_n26, maj_161_n25, maj_161_n24, maj_161_n23, maj_161_n22,
         maj_161_n21, maj_161_n20, maj_161_n19, maj_161_n18, maj_161_n17,
         maj_161_n16, maj_161_n15, maj_161_n14, maj_162_n26, maj_162_n25,
         maj_162_n24, maj_162_n23, maj_162_n22, maj_162_n21, maj_162_n20,
         maj_162_n19, maj_162_n18, maj_162_n17, maj_162_n16, maj_162_n15,
         maj_162_n14, maj_163_n26, maj_163_n25, maj_163_n24, maj_163_n23,
         maj_163_n22, maj_163_n21, maj_163_n20, maj_163_n19, maj_163_n18,
         maj_163_n17, maj_163_n16, maj_163_n15, maj_163_n14, maj_164_n26,
         maj_164_n25, maj_164_n24, maj_164_n23, maj_164_n22, maj_164_n21,
         maj_164_n20, maj_164_n19, maj_164_n18, maj_164_n17, maj_164_n16,
         maj_164_n15, maj_164_n14, maj_165_n26, maj_165_n25, maj_165_n24,
         maj_165_n23, maj_165_n22, maj_165_n21, maj_165_n20, maj_165_n19,
         maj_165_n18, maj_165_n17, maj_165_n16, maj_165_n15, maj_165_n14,
         maj_166_n26, maj_166_n25, maj_166_n24, maj_166_n23, maj_166_n22,
         maj_166_n21, maj_166_n20, maj_166_n19, maj_166_n18, maj_166_n17,
         maj_166_n16, maj_166_n15, maj_166_n14, maj_167_n26, maj_167_n25,
         maj_167_n24, maj_167_n23, maj_167_n22, maj_167_n21, maj_167_n20,
         maj_167_n19, maj_167_n18, maj_167_n17, maj_167_n16, maj_167_n15,
         maj_167_n14, maj_168_n26, maj_168_n25, maj_168_n24, maj_168_n23,
         maj_168_n22, maj_168_n21, maj_168_n20, maj_168_n19, maj_168_n18,
         maj_168_n17, maj_168_n16, maj_168_n15, maj_168_n14, maj_169_n26,
         maj_169_n25, maj_169_n24, maj_169_n23, maj_169_n22, maj_169_n21,
         maj_169_n20, maj_169_n19, maj_169_n18, maj_169_n17, maj_169_n16,
         maj_169_n15, maj_169_n14, maj_170_n26, maj_170_n25, maj_170_n24,
         maj_170_n23, maj_170_n22, maj_170_n21, maj_170_n20, maj_170_n19,
         maj_170_n18, maj_170_n17, maj_170_n16, maj_170_n15, maj_170_n14,
         maj_171_n26, maj_171_n25, maj_171_n24, maj_171_n23, maj_171_n22,
         maj_171_n21, maj_171_n20, maj_171_n19, maj_171_n18, maj_171_n17,
         maj_171_n16, maj_171_n15, maj_171_n14, maj_172_n26, maj_172_n25,
         maj_172_n24, maj_172_n23, maj_172_n22, maj_172_n21, maj_172_n20,
         maj_172_n19, maj_172_n18, maj_172_n17, maj_172_n16, maj_172_n15,
         maj_172_n14, maj_173_n26, maj_173_n25, maj_173_n24, maj_173_n23,
         maj_173_n22, maj_173_n21, maj_173_n20, maj_173_n19, maj_173_n18,
         maj_173_n17, maj_173_n16, maj_173_n15, maj_173_n14, maj_174_n26,
         maj_174_n25, maj_174_n24, maj_174_n23, maj_174_n22, maj_174_n21,
         maj_174_n20, maj_174_n19, maj_174_n18, maj_174_n17, maj_174_n16,
         maj_174_n15, maj_174_n14, maj_175_n26, maj_175_n25, maj_175_n24,
         maj_175_n23, maj_175_n22, maj_175_n21, maj_175_n20, maj_175_n19,
         maj_175_n18, maj_175_n17, maj_175_n16, maj_175_n15, maj_175_n14,
         maj_176_n26, maj_176_n25, maj_176_n24, maj_176_n23, maj_176_n22,
         maj_176_n21, maj_176_n20, maj_176_n19, maj_176_n18, maj_176_n17,
         maj_176_n16, maj_176_n15, maj_176_n14, maj_177_n26, maj_177_n25,
         maj_177_n24, maj_177_n23, maj_177_n22, maj_177_n21, maj_177_n20,
         maj_177_n19, maj_177_n18, maj_177_n17, maj_177_n16, maj_177_n15,
         maj_177_n14, maj_178_n26, maj_178_n25, maj_178_n24, maj_178_n23,
         maj_178_n22, maj_178_n21, maj_178_n20, maj_178_n19, maj_178_n18,
         maj_178_n17, maj_178_n16, maj_178_n15, maj_178_n14, maj_179_n26,
         maj_179_n25, maj_179_n24, maj_179_n23, maj_179_n22, maj_179_n21,
         maj_179_n20, maj_179_n19, maj_179_n18, maj_179_n17, maj_179_n16,
         maj_179_n15, maj_179_n14, maj_180_n26, maj_180_n25, maj_180_n24,
         maj_180_n23, maj_180_n22, maj_180_n21, maj_180_n20, maj_180_n19,
         maj_180_n18, maj_180_n17, maj_180_n16, maj_180_n15, maj_180_n14,
         maj_181_n26, maj_181_n25, maj_181_n24, maj_181_n23, maj_181_n22,
         maj_181_n21, maj_181_n20, maj_181_n19, maj_181_n18, maj_181_n17,
         maj_181_n16, maj_181_n15, maj_181_n14, maj_182_n26, maj_182_n25,
         maj_182_n24, maj_182_n23, maj_182_n22, maj_182_n21, maj_182_n20,
         maj_182_n19, maj_182_n18, maj_182_n17, maj_182_n16, maj_182_n15,
         maj_182_n14, maj_183_n26, maj_183_n25, maj_183_n24, maj_183_n23,
         maj_183_n22, maj_183_n21, maj_183_n20, maj_183_n19, maj_183_n18,
         maj_183_n17, maj_183_n16, maj_183_n15, maj_183_n14, maj_184_n26,
         maj_184_n25, maj_184_n24, maj_184_n23, maj_184_n22, maj_184_n21,
         maj_184_n20, maj_184_n19, maj_184_n18, maj_184_n17, maj_184_n16,
         maj_184_n15, maj_184_n14, maj_185_n26, maj_185_n25, maj_185_n24,
         maj_185_n23, maj_185_n22, maj_185_n21, maj_185_n20, maj_185_n19,
         maj_185_n18, maj_185_n17, maj_185_n16, maj_185_n15, maj_185_n14,
         maj_186_n26, maj_186_n25, maj_186_n24, maj_186_n23, maj_186_n22,
         maj_186_n21, maj_186_n20, maj_186_n19, maj_186_n18, maj_186_n17,
         maj_186_n16, maj_186_n15, maj_186_n14, maj_187_n26, maj_187_n25,
         maj_187_n24, maj_187_n23, maj_187_n22, maj_187_n21, maj_187_n20,
         maj_187_n19, maj_187_n18, maj_187_n17, maj_187_n16, maj_187_n15,
         maj_187_n14, maj_188_n26, maj_188_n25, maj_188_n24, maj_188_n23,
         maj_188_n22, maj_188_n21, maj_188_n20, maj_188_n19, maj_188_n18,
         maj_188_n17, maj_188_n16, maj_188_n15, maj_188_n14, maj_189_n26,
         maj_189_n25, maj_189_n24, maj_189_n23, maj_189_n22, maj_189_n21,
         maj_189_n20, maj_189_n19, maj_189_n18, maj_189_n17, maj_189_n16,
         maj_189_n15, maj_189_n14, maj_190_n26, maj_190_n25, maj_190_n24,
         maj_190_n23, maj_190_n22, maj_190_n21, maj_190_n20, maj_190_n19,
         maj_190_n18, maj_190_n17, maj_190_n16, maj_190_n15, maj_190_n14,
         maj_191_n26, maj_191_n25, maj_191_n24, maj_191_n23, maj_191_n22,
         maj_191_n21, maj_191_n20, maj_191_n19, maj_191_n18, maj_191_n17,
         maj_191_n16, maj_191_n15, maj_191_n14, maj_192_n26, maj_192_n25,
         maj_192_n24, maj_192_n23, maj_192_n22, maj_192_n21, maj_192_n20,
         maj_192_n19, maj_192_n18, maj_192_n17, maj_192_n16, maj_192_n15,
         maj_192_n14, maj_193_n26, maj_193_n25, maj_193_n24, maj_193_n23,
         maj_193_n22, maj_193_n21, maj_193_n20, maj_193_n19, maj_193_n18,
         maj_193_n17, maj_193_n16, maj_193_n15, maj_193_n14, maj_194_n26,
         maj_194_n25, maj_194_n24, maj_194_n23, maj_194_n22, maj_194_n21,
         maj_194_n20, maj_194_n19, maj_194_n18, maj_194_n17, maj_194_n16,
         maj_194_n15, maj_194_n14, maj_195_n26, maj_195_n25, maj_195_n24,
         maj_195_n23, maj_195_n22, maj_195_n21, maj_195_n20, maj_195_n19,
         maj_195_n18, maj_195_n17, maj_195_n16, maj_195_n15, maj_195_n14,
         maj_196_n26, maj_196_n25, maj_196_n24, maj_196_n23, maj_196_n22,
         maj_196_n21, maj_196_n20, maj_196_n19, maj_196_n18, maj_196_n17,
         maj_196_n16, maj_196_n15, maj_196_n14, maj_197_n26, maj_197_n25,
         maj_197_n24, maj_197_n23, maj_197_n22, maj_197_n21, maj_197_n20,
         maj_197_n19, maj_197_n18, maj_197_n17, maj_197_n16, maj_197_n15,
         maj_197_n14, maj_198_n26, maj_198_n25, maj_198_n24, maj_198_n23,
         maj_198_n22, maj_198_n21, maj_198_n20, maj_198_n19, maj_198_n18,
         maj_198_n17, maj_198_n16, maj_198_n15, maj_198_n14, maj_199_n26,
         maj_199_n25, maj_199_n24, maj_199_n23, maj_199_n22, maj_199_n21,
         maj_199_n20, maj_199_n19, maj_199_n18, maj_199_n17, maj_199_n16,
         maj_199_n15, maj_199_n14, maj_200_n26, maj_200_n25, maj_200_n24,
         maj_200_n23, maj_200_n22, maj_200_n21, maj_200_n20, maj_200_n19,
         maj_200_n18, maj_200_n17, maj_200_n16, maj_200_n15, maj_200_n14,
         maj_201_n26, maj_201_n25, maj_201_n24, maj_201_n23, maj_201_n22,
         maj_201_n21, maj_201_n20, maj_201_n19, maj_201_n18, maj_201_n17,
         maj_201_n16, maj_201_n15, maj_201_n14, maj_202_n26, maj_202_n25,
         maj_202_n24, maj_202_n23, maj_202_n22, maj_202_n21, maj_202_n20,
         maj_202_n19, maj_202_n18, maj_202_n17, maj_202_n16, maj_202_n15,
         maj_202_n14, maj_203_n26, maj_203_n25, maj_203_n24, maj_203_n23,
         maj_203_n22, maj_203_n21, maj_203_n20, maj_203_n19, maj_203_n18,
         maj_203_n17, maj_203_n16, maj_203_n15, maj_203_n14, maj_204_n26,
         maj_204_n25, maj_204_n24, maj_204_n23, maj_204_n22, maj_204_n21,
         maj_204_n20, maj_204_n19, maj_204_n18, maj_204_n17, maj_204_n16,
         maj_204_n15, maj_204_n14, maj_205_n26, maj_205_n25, maj_205_n24,
         maj_205_n23, maj_205_n22, maj_205_n21, maj_205_n20, maj_205_n19,
         maj_205_n18, maj_205_n17, maj_205_n16, maj_205_n15, maj_205_n14,
         maj_206_n26, maj_206_n25, maj_206_n24, maj_206_n23, maj_206_n22,
         maj_206_n21, maj_206_n20, maj_206_n19, maj_206_n18, maj_206_n17,
         maj_206_n16, maj_206_n15, maj_206_n14, maj_207_n26, maj_207_n25,
         maj_207_n24, maj_207_n23, maj_207_n22, maj_207_n21, maj_207_n20,
         maj_207_n19, maj_207_n18, maj_207_n17, maj_207_n16, maj_207_n15,
         maj_207_n14, maj_208_n26, maj_208_n25, maj_208_n24, maj_208_n23,
         maj_208_n22, maj_208_n21, maj_208_n20, maj_208_n19, maj_208_n18,
         maj_208_n17, maj_208_n16, maj_208_n15, maj_208_n14, maj_209_n26,
         maj_209_n25, maj_209_n24, maj_209_n23, maj_209_n22, maj_209_n21,
         maj_209_n20, maj_209_n19, maj_209_n18, maj_209_n17, maj_209_n16,
         maj_209_n15, maj_209_n14, maj_210_n26, maj_210_n25, maj_210_n24,
         maj_210_n23, maj_210_n22, maj_210_n21, maj_210_n20, maj_210_n19,
         maj_210_n18, maj_210_n17, maj_210_n16, maj_210_n15, maj_210_n14,
         maj_211_n26, maj_211_n25, maj_211_n24, maj_211_n23, maj_211_n22,
         maj_211_n21, maj_211_n20, maj_211_n19, maj_211_n18, maj_211_n17,
         maj_211_n16, maj_211_n15, maj_211_n14, maj_212_n26, maj_212_n25,
         maj_212_n24, maj_212_n23, maj_212_n22, maj_212_n21, maj_212_n20,
         maj_212_n19, maj_212_n18, maj_212_n17, maj_212_n16, maj_212_n15,
         maj_212_n14, maj_213_n26, maj_213_n25, maj_213_n24, maj_213_n23,
         maj_213_n22, maj_213_n21, maj_213_n20, maj_213_n19, maj_213_n18,
         maj_213_n17, maj_213_n16, maj_213_n15, maj_213_n14, maj_214_n26,
         maj_214_n25, maj_214_n24, maj_214_n23, maj_214_n22, maj_214_n21,
         maj_214_n20, maj_214_n19, maj_214_n18, maj_214_n17, maj_214_n16,
         maj_214_n15, maj_214_n14, maj_215_n26, maj_215_n25, maj_215_n24,
         maj_215_n23, maj_215_n22, maj_215_n21, maj_215_n20, maj_215_n19,
         maj_215_n18, maj_215_n17, maj_215_n16, maj_215_n15, maj_215_n14,
         maj_216_n26, maj_216_n25, maj_216_n24, maj_216_n23, maj_216_n22,
         maj_216_n21, maj_216_n20, maj_216_n19, maj_216_n18, maj_216_n17,
         maj_216_n16, maj_216_n15, maj_216_n14, maj_217_n26, maj_217_n25,
         maj_217_n24, maj_217_n23, maj_217_n22, maj_217_n21, maj_217_n20,
         maj_217_n19, maj_217_n18, maj_217_n17, maj_217_n16, maj_217_n15,
         maj_217_n14, maj_218_n26, maj_218_n25, maj_218_n24, maj_218_n23,
         maj_218_n22, maj_218_n21, maj_218_n20, maj_218_n19, maj_218_n18,
         maj_218_n17, maj_218_n16, maj_218_n15, maj_218_n14, maj_219_n26,
         maj_219_n25, maj_219_n24, maj_219_n23, maj_219_n22, maj_219_n21,
         maj_219_n20, maj_219_n19, maj_219_n18, maj_219_n17, maj_219_n16,
         maj_219_n15, maj_219_n14, maj_220_n26, maj_220_n25, maj_220_n24,
         maj_220_n23, maj_220_n22, maj_220_n21, maj_220_n20, maj_220_n19,
         maj_220_n18, maj_220_n17, maj_220_n16, maj_220_n15, maj_220_n14,
         maj_221_n26, maj_221_n25, maj_221_n24, maj_221_n23, maj_221_n22,
         maj_221_n21, maj_221_n20, maj_221_n19, maj_221_n18, maj_221_n17,
         maj_221_n16, maj_221_n15, maj_221_n14, maj_222_n26, maj_222_n25,
         maj_222_n24, maj_222_n23, maj_222_n22, maj_222_n21, maj_222_n20,
         maj_222_n19, maj_222_n18, maj_222_n17, maj_222_n16, maj_222_n15,
         maj_222_n14, maj_223_n26, maj_223_n25, maj_223_n24, maj_223_n23,
         maj_223_n22, maj_223_n21, maj_223_n20, maj_223_n19, maj_223_n18,
         maj_223_n17, maj_223_n16, maj_223_n15, maj_223_n14, maj_224_n26,
         maj_224_n25, maj_224_n24, maj_224_n23, maj_224_n22, maj_224_n21,
         maj_224_n20, maj_224_n19, maj_224_n18, maj_224_n17, maj_224_n16,
         maj_224_n15, maj_224_n14, maj_225_n26, maj_225_n25, maj_225_n24,
         maj_225_n23, maj_225_n22, maj_225_n21, maj_225_n20, maj_225_n19,
         maj_225_n18, maj_225_n17, maj_225_n16, maj_225_n15, maj_225_n14,
         maj_226_n26, maj_226_n25, maj_226_n24, maj_226_n23, maj_226_n22,
         maj_226_n21, maj_226_n20, maj_226_n19, maj_226_n18, maj_226_n17,
         maj_226_n16, maj_226_n15, maj_226_n14, maj_227_n26, maj_227_n25,
         maj_227_n24, maj_227_n23, maj_227_n22, maj_227_n21, maj_227_n20,
         maj_227_n19, maj_227_n18, maj_227_n17, maj_227_n16, maj_227_n15,
         maj_227_n14, maj_228_n26, maj_228_n25, maj_228_n24, maj_228_n23,
         maj_228_n22, maj_228_n21, maj_228_n20, maj_228_n19, maj_228_n18,
         maj_228_n17, maj_228_n16, maj_228_n15, maj_228_n14, maj_229_n26,
         maj_229_n25, maj_229_n24, maj_229_n23, maj_229_n22, maj_229_n21,
         maj_229_n20, maj_229_n19, maj_229_n18, maj_229_n17, maj_229_n16,
         maj_229_n15, maj_229_n14, maj_230_n26, maj_230_n25, maj_230_n24,
         maj_230_n23, maj_230_n22, maj_230_n21, maj_230_n20, maj_230_n19,
         maj_230_n18, maj_230_n17, maj_230_n16, maj_230_n15, maj_230_n14,
         maj_231_n26, maj_231_n25, maj_231_n24, maj_231_n23, maj_231_n22,
         maj_231_n21, maj_231_n20, maj_231_n19, maj_231_n18, maj_231_n17,
         maj_231_n16, maj_231_n15, maj_231_n14, maj_232_n26, maj_232_n25,
         maj_232_n24, maj_232_n23, maj_232_n22, maj_232_n21, maj_232_n20,
         maj_232_n19, maj_232_n18, maj_232_n17, maj_232_n16, maj_232_n15,
         maj_232_n14, maj_233_n26, maj_233_n25, maj_233_n24, maj_233_n23,
         maj_233_n22, maj_233_n21, maj_233_n20, maj_233_n19, maj_233_n18,
         maj_233_n17, maj_233_n16, maj_233_n15, maj_233_n14, maj_234_n26,
         maj_234_n25, maj_234_n24, maj_234_n23, maj_234_n22, maj_234_n21,
         maj_234_n20, maj_234_n19, maj_234_n18, maj_234_n17, maj_234_n16,
         maj_234_n15, maj_234_n14, maj_235_n26, maj_235_n25, maj_235_n24,
         maj_235_n23, maj_235_n22, maj_235_n21, maj_235_n20, maj_235_n19,
         maj_235_n18, maj_235_n17, maj_235_n16, maj_235_n15, maj_235_n14,
         maj_236_n26, maj_236_n25, maj_236_n24, maj_236_n23, maj_236_n22,
         maj_236_n21, maj_236_n20, maj_236_n19, maj_236_n18, maj_236_n17,
         maj_236_n16, maj_236_n15, maj_236_n14, maj_237_n26, maj_237_n25,
         maj_237_n24, maj_237_n23, maj_237_n22, maj_237_n21, maj_237_n20,
         maj_237_n19, maj_237_n18, maj_237_n17, maj_237_n16, maj_237_n15,
         maj_237_n14, maj_238_n26, maj_238_n25, maj_238_n24, maj_238_n23,
         maj_238_n22, maj_238_n21, maj_238_n20, maj_238_n19, maj_238_n18,
         maj_238_n17, maj_238_n16, maj_238_n15, maj_238_n14, maj_239_n26,
         maj_239_n25, maj_239_n24, maj_239_n23, maj_239_n22, maj_239_n21,
         maj_239_n20, maj_239_n19, maj_239_n18, maj_239_n17, maj_239_n16,
         maj_239_n15, maj_239_n14;
  wire   [4:0] u_0_0;
  wire   [4:0] v_0_0;
  wire   [4:0] u_0_1;
  wire   [4:0] v_0_1;
  wire   [4:0] u_0_2;
  wire   [4:0] v_0_2;
  wire   [4:0] u_1_0;
  wire   [4:0] v_1_0;
  wire   [4:0] u_1_1;
  wire   [4:0] v_1_1;
  wire   [4:0] u_1_2;
  wire   [4:0] v_1_2;
  wire   [4:0] u_2_0;
  wire   [4:0] v_2_0;
  wire   [4:0] u_2_1;
  wire   [4:0] v_2_1;
  wire   [4:0] u_2_2;
  wire   [4:0] v_2_2;
  wire   [4:0] u_3_0;
  wire   [4:0] v_3_0;
  wire   [4:0] u_3_1;
  wire   [4:0] v_3_1;
  wire   [4:0] u_3_2;
  wire   [4:0] v_3_2;
  wire   [4:0] temp_0_0;
  wire   [4:0] a_reg_0;
  wire   [4:0] v_reg_0_0;
  wire   [4:0] u_reg_0_0;
  wire   [4:0] v_reg_0_1;
  wire   [4:0] u_reg_0_1;
  wire   [4:0] v_reg_0_2;
  wire   [4:0] u_reg_0_2;
  wire   [4:0] temp_0_1;
  wire   [4:0] a_reg_1;
  wire   [4:0] v_reg_1_0;
  wire   [4:0] u_reg_1_0;
  wire   [4:0] v_reg_1_1;
  wire   [4:0] u_reg_1_1;
  wire   [4:0] v_reg_1_2;
  wire   [4:0] u_reg_1_2;
  wire   [4:0] temp_0_2;
  wire   [4:0] a_reg_2;
  wire   [4:0] v_reg_2_0;
  wire   [4:0] u_reg_2_0;
  wire   [4:0] v_reg_2_1;
  wire   [4:0] u_reg_2_1;
  wire   [4:0] v_reg_2_2;
  wire   [4:0] u_reg_2_2;
  wire   [4:0] temp_0_3;
  wire   [4:0] a_reg_3;
  wire   [4:0] v_reg_3_0;
  wire   [4:0] u_reg_3_0;
  wire   [4:0] v_reg_3_1;
  wire   [4:0] u_reg_3_1;
  wire   [4:0] v_reg_3_2;
  wire   [4:0] u_reg_3_2;

  DFF_X1 u_reg_1_1_reg_4_ ( .D(maj_224_port_o), .CK(clk), .Q(u_reg_1_1[4]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_3_ ( .D(maj_200_port_o), .CK(clk), .Q(u_reg_1_1[3]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_2_ ( .D(maj_176_port_o), .CK(clk), .Q(u_reg_1_1[2]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_1_ ( .D(maj_152_port_o), .CK(clk), .Q(u_reg_1_1[1]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_0_ ( .D(maj_128_port_o), .CK(clk), .Q(u_reg_1_1[0]), 
        .QN() );
  DFF_X1 a_reg_3_reg_4_ ( .D(port_a_3[4]), .CK(clk), .Q(a_reg_3[4]), .QN() );
  DFF_X1 a_reg_3_reg_3_ ( .D(port_a_3[3]), .CK(clk), .Q(a_reg_3[3]), .QN() );
  DFF_X1 a_reg_3_reg_2_ ( .D(port_a_3[2]), .CK(clk), .Q(a_reg_3[2]), .QN() );
  DFF_X1 a_reg_3_reg_1_ ( .D(port_a_3[1]), .CK(clk), .Q(a_reg_3[1]), .QN() );
  DFF_X1 a_reg_3_reg_0_ ( .D(port_a_3[0]), .CK(clk), .Q(a_reg_3[0]), .QN() );
  DFF_X1 v_reg_2_1_reg_4_ ( .D(maj_231_port_o), .CK(clk), .Q(v_reg_2_1[4]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_3_ ( .D(maj_207_port_o), .CK(clk), .Q(v_reg_2_1[3]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_2_ ( .D(maj_183_port_o), .CK(clk), .Q(v_reg_2_1[2]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_1_ ( .D(maj_159_port_o), .CK(clk), .Q(v_reg_2_1[1]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_0_ ( .D(maj_135_port_o), .CK(clk), .Q(v_reg_2_1[0]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_4_ ( .D(maj_226_port_o), .CK(clk), .Q(u_reg_1_2[4]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_3_ ( .D(maj_202_port_o), .CK(clk), .Q(u_reg_1_2[3]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_2_ ( .D(maj_178_port_o), .CK(clk), .Q(u_reg_1_2[2]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_1_ ( .D(maj_154_port_o), .CK(clk), .Q(u_reg_1_2[1]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_0_ ( .D(maj_130_port_o), .CK(clk), .Q(u_reg_1_2[0]), 
        .QN() );
  DFF_X1 ab_reg_3_reg_4_ ( .D(N19), .CK(clk), .Q(temp_0_3[4]), .QN() );
  DFF_X1 ab_reg_3_reg_3_ ( .D(N15), .CK(clk), .Q(temp_0_3[3]), .QN() );
  DFF_X1 ab_reg_3_reg_2_ ( .D(N11), .CK(clk), .Q(temp_0_3[2]), .QN() );
  DFF_X1 ab_reg_3_reg_1_ ( .D(N7), .CK(clk), .Q(temp_0_3[1]), .QN() );
  DFF_X1 ab_reg_3_reg_0_ ( .D(N3), .CK(clk), .Q(temp_0_3[0]), .QN() );
  DFF_X1 v_reg_2_0_reg_4_ ( .D(maj_229_port_o), .CK(clk), .Q(v_reg_2_0[4]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_3_ ( .D(maj_205_port_o), .CK(clk), .Q(v_reg_2_0[3]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_2_ ( .D(maj_181_port_o), .CK(clk), .Q(v_reg_2_0[2]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_1_ ( .D(maj_157_port_o), .CK(clk), .Q(v_reg_2_0[1]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_0_ ( .D(maj_133_port_o), .CK(clk), .Q(v_reg_2_0[0]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_4_ ( .D(maj_228_port_o), .CK(clk), .Q(u_reg_2_0[4]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_3_ ( .D(maj_204_port_o), .CK(clk), .Q(u_reg_2_0[3]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_2_ ( .D(maj_180_port_o), .CK(clk), .Q(u_reg_2_0[2]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_1_ ( .D(maj_156_port_o), .CK(clk), .Q(u_reg_2_0[1]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_0_ ( .D(maj_132_port_o), .CK(clk), .Q(u_reg_2_0[0]), 
        .QN() );
  DFF_X1 a_reg_2_reg_4_ ( .D(port_a_2[4]), .CK(clk), .Q(a_reg_2[4]), .QN() );
  DFF_X1 a_reg_2_reg_3_ ( .D(port_a_2[3]), .CK(clk), .Q(a_reg_2[3]), .QN() );
  DFF_X1 a_reg_2_reg_2_ ( .D(port_a_2[2]), .CK(clk), .Q(a_reg_2[2]), .QN() );
  DFF_X1 a_reg_2_reg_1_ ( .D(port_a_2[1]), .CK(clk), .Q(a_reg_2[1]), .QN() );
  DFF_X1 a_reg_2_reg_0_ ( .D(port_a_2[0]), .CK(clk), .Q(a_reg_2[0]), .QN() );
  DFF_X1 v_reg_1_2_reg_4_ ( .D(maj_227_port_o), .CK(clk), .Q(v_reg_1_2[4]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_3_ ( .D(maj_203_port_o), .CK(clk), .Q(v_reg_1_2[3]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_2_ ( .D(maj_179_port_o), .CK(clk), .Q(v_reg_1_2[2]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_1_ ( .D(maj_155_port_o), .CK(clk), .Q(v_reg_1_2[1]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_0_ ( .D(maj_131_port_o), .CK(clk), .Q(v_reg_1_2[0]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_4_ ( .D(maj_230_port_o), .CK(clk), .Q(u_reg_2_1[4]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_3_ ( .D(maj_206_port_o), .CK(clk), .Q(u_reg_2_1[3]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_2_ ( .D(maj_182_port_o), .CK(clk), .Q(u_reg_2_1[2]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_1_ ( .D(maj_158_port_o), .CK(clk), .Q(u_reg_2_1[1]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_0_ ( .D(maj_134_port_o), .CK(clk), .Q(u_reg_2_1[0]), 
        .QN() );
  DFF_X1 ab_reg_2_reg_4_ ( .D(N18), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 ab_reg_2_reg_3_ ( .D(N14), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 ab_reg_2_reg_2_ ( .D(N10), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 ab_reg_2_reg_1_ ( .D(N6), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 ab_reg_2_reg_0_ ( .D(N2), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 v_reg_1_1_reg_4_ ( .D(maj_225_port_o), .CK(clk), .Q(v_reg_1_1[4]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_3_ ( .D(maj_201_port_o), .CK(clk), .Q(v_reg_1_1[3]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_2_ ( .D(maj_177_port_o), .CK(clk), .Q(v_reg_1_1[2]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_1_ ( .D(maj_153_port_o), .CK(clk), .Q(v_reg_1_1[1]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_0_ ( .D(maj_129_port_o), .CK(clk), .Q(v_reg_1_1[0]), 
        .QN() );
  DFF_X1 a_reg_1_reg_4_ ( .D(port_a_1[4]), .CK(clk), .Q(a_reg_1[4]), .QN() );
  DFF_X1 a_reg_1_reg_3_ ( .D(port_a_1[3]), .CK(clk), .Q(a_reg_1[3]), .QN() );
  DFF_X1 a_reg_1_reg_2_ ( .D(port_a_1[2]), .CK(clk), .Q(a_reg_1[2]), .QN() );
  DFF_X1 a_reg_1_reg_1_ ( .D(port_a_1[1]), .CK(clk), .Q(a_reg_1[1]), .QN() );
  DFF_X1 a_reg_1_reg_0_ ( .D(port_a_1[0]), .CK(clk), .Q(a_reg_1[0]), .QN() );
  DFF_X1 ab_reg_1_reg_4_ ( .D(N17), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 ab_reg_1_reg_3_ ( .D(N13), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 ab_reg_1_reg_2_ ( .D(N9), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 ab_reg_1_reg_1_ ( .D(N5), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 ab_reg_1_reg_0_ ( .D(N1), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 a_reg_0_reg_4_ ( .D(port_a_0[4]), .CK(clk), .Q(a_reg_0[4]), .QN() );
  DFF_X1 a_reg_0_reg_3_ ( .D(port_a_0[3]), .CK(clk), .Q(a_reg_0[3]), .QN() );
  DFF_X1 a_reg_0_reg_2_ ( .D(port_a_0[2]), .CK(clk), .Q(a_reg_0[2]), .QN() );
  DFF_X1 a_reg_0_reg_1_ ( .D(port_a_0[1]), .CK(clk), .Q(a_reg_0[1]), .QN() );
  DFF_X1 a_reg_0_reg_0_ ( .D(port_a_0[0]), .CK(clk), .Q(a_reg_0[0]), .QN() );
  DFF_X1 ab_reg_0_reg_4_ ( .D(N16), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 ab_reg_0_reg_3_ ( .D(N12), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 ab_reg_0_reg_2_ ( .D(N8), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 ab_reg_0_reg_1_ ( .D(N4), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 ab_reg_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 v_reg_3_2_reg_4_ ( .D(maj_239_port_o), .CK(clk), .Q(v_reg_3_2[4]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_3_ ( .D(maj_215_port_o), .CK(clk), .Q(v_reg_3_2[3]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_2_ ( .D(maj_191_port_o), .CK(clk), .Q(v_reg_3_2[2]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_1_ ( .D(maj_167_port_o), .CK(clk), .Q(v_reg_3_2[1]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_0_ ( .D(maj_143_port_o), .CK(clk), .Q(v_reg_3_2[0]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_4_ ( .D(maj_238_port_o), .CK(clk), .Q(u_reg_3_2[4]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_3_ ( .D(maj_214_port_o), .CK(clk), .Q(u_reg_3_2[3]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_2_ ( .D(maj_190_port_o), .CK(clk), .Q(u_reg_3_2[2]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_1_ ( .D(maj_166_port_o), .CK(clk), .Q(u_reg_3_2[1]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_0_ ( .D(maj_142_port_o), .CK(clk), .Q(u_reg_3_2[0]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_4_ ( .D(maj_237_port_o), .CK(clk), .Q(v_reg_3_1[4]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_3_ ( .D(maj_213_port_o), .CK(clk), .Q(v_reg_3_1[3]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_2_ ( .D(maj_189_port_o), .CK(clk), .Q(v_reg_3_1[2]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_1_ ( .D(maj_165_port_o), .CK(clk), .Q(v_reg_3_1[1]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_0_ ( .D(maj_141_port_o), .CK(clk), .Q(v_reg_3_1[0]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_4_ ( .D(maj_236_port_o), .CK(clk), .Q(u_reg_3_1[4]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_3_ ( .D(maj_212_port_o), .CK(clk), .Q(u_reg_3_1[3]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_2_ ( .D(maj_188_port_o), .CK(clk), .Q(u_reg_3_1[2]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_1_ ( .D(maj_164_port_o), .CK(clk), .Q(u_reg_3_1[1]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_0_ ( .D(maj_140_port_o), .CK(clk), .Q(u_reg_3_1[0]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_4_ ( .D(maj_235_port_o), .CK(clk), .Q(v_reg_3_0[4]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_3_ ( .D(maj_211_port_o), .CK(clk), .Q(v_reg_3_0[3]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_2_ ( .D(maj_187_port_o), .CK(clk), .Q(v_reg_3_0[2]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_1_ ( .D(maj_163_port_o), .CK(clk), .Q(v_reg_3_0[1]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_0_ ( .D(maj_139_port_o), .CK(clk), .Q(v_reg_3_0[0]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_4_ ( .D(maj_234_port_o), .CK(clk), .Q(u_reg_3_0[4]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_3_ ( .D(maj_210_port_o), .CK(clk), .Q(u_reg_3_0[3]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_2_ ( .D(maj_186_port_o), .CK(clk), .Q(u_reg_3_0[2]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_1_ ( .D(maj_162_port_o), .CK(clk), .Q(u_reg_3_0[1]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_0_ ( .D(maj_138_port_o), .CK(clk), .Q(u_reg_3_0[0]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_4_ ( .D(maj_233_port_o), .CK(clk), .Q(v_reg_2_2[4]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_3_ ( .D(maj_209_port_o), .CK(clk), .Q(v_reg_2_2[3]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_2_ ( .D(maj_185_port_o), .CK(clk), .Q(v_reg_2_2[2]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_1_ ( .D(maj_161_port_o), .CK(clk), .Q(v_reg_2_2[1]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_0_ ( .D(maj_137_port_o), .CK(clk), .Q(v_reg_2_2[0]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_4_ ( .D(maj_232_port_o), .CK(clk), .Q(u_reg_2_2[4]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_3_ ( .D(maj_208_port_o), .CK(clk), .Q(u_reg_2_2[3]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_2_ ( .D(maj_184_port_o), .CK(clk), .Q(u_reg_2_2[2]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_1_ ( .D(maj_160_port_o), .CK(clk), .Q(u_reg_2_2[1]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_0_ ( .D(maj_136_port_o), .CK(clk), .Q(u_reg_2_2[0]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_4_ ( .D(maj_216_port_o), .CK(clk), .Q(u_reg_0_0[4]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_3_ ( .D(maj_192_port_o), .CK(clk), .Q(u_reg_0_0[3]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_2_ ( .D(maj_168_port_o), .CK(clk), .Q(u_reg_0_0[2]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_1_ ( .D(maj_144_port_o), .CK(clk), .Q(u_reg_0_0[1]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_0_ ( .D(maj_120_port_o), .CK(clk), .Q(u_reg_0_0[0]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_4_ ( .D(maj_217_port_o), .CK(clk), .Q(v_reg_0_0[4]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_3_ ( .D(maj_193_port_o), .CK(clk), .Q(v_reg_0_0[3]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_2_ ( .D(maj_169_port_o), .CK(clk), .Q(v_reg_0_0[2]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_1_ ( .D(maj_145_port_o), .CK(clk), .Q(v_reg_0_0[1]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_0_ ( .D(maj_121_port_o), .CK(clk), .Q(v_reg_0_0[0]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_4_ ( .D(maj_218_port_o), .CK(clk), .Q(u_reg_0_1[4]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_3_ ( .D(maj_194_port_o), .CK(clk), .Q(u_reg_0_1[3]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_2_ ( .D(maj_170_port_o), .CK(clk), .Q(u_reg_0_1[2]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_1_ ( .D(maj_146_port_o), .CK(clk), .Q(u_reg_0_1[1]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_0_ ( .D(maj_122_port_o), .CK(clk), .Q(u_reg_0_1[0]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_4_ ( .D(maj_219_port_o), .CK(clk), .Q(v_reg_0_1[4]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_3_ ( .D(maj_195_port_o), .CK(clk), .Q(v_reg_0_1[3]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_2_ ( .D(maj_171_port_o), .CK(clk), .Q(v_reg_0_1[2]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_1_ ( .D(maj_147_port_o), .CK(clk), .Q(v_reg_0_1[1]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_0_ ( .D(maj_123_port_o), .CK(clk), .Q(v_reg_0_1[0]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_4_ ( .D(maj_220_port_o), .CK(clk), .Q(u_reg_0_2[4]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_3_ ( .D(maj_196_port_o), .CK(clk), .Q(u_reg_0_2[3]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_2_ ( .D(maj_172_port_o), .CK(clk), .Q(u_reg_0_2[2]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_1_ ( .D(maj_148_port_o), .CK(clk), .Q(u_reg_0_2[1]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_0_ ( .D(maj_124_port_o), .CK(clk), .Q(u_reg_0_2[0]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_4_ ( .D(maj_221_port_o), .CK(clk), .Q(v_reg_0_2[4]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_3_ ( .D(maj_197_port_o), .CK(clk), .Q(v_reg_0_2[3]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_2_ ( .D(maj_173_port_o), .CK(clk), .Q(v_reg_0_2[2]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_1_ ( .D(maj_149_port_o), .CK(clk), .Q(v_reg_0_2[1]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_0_ ( .D(maj_125_port_o), .CK(clk), .Q(v_reg_0_2[0]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_4_ ( .D(maj_222_port_o), .CK(clk), .Q(u_reg_1_0[4]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_3_ ( .D(maj_198_port_o), .CK(clk), .Q(u_reg_1_0[3]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_2_ ( .D(maj_174_port_o), .CK(clk), .Q(u_reg_1_0[2]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_1_ ( .D(maj_150_port_o), .CK(clk), .Q(u_reg_1_0[1]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_0_ ( .D(maj_126_port_o), .CK(clk), .Q(u_reg_1_0[0]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_4_ ( .D(maj_223_port_o), .CK(clk), .Q(v_reg_1_0[4]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_3_ ( .D(maj_199_port_o), .CK(clk), .Q(v_reg_1_0[3]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_2_ ( .D(maj_175_port_o), .CK(clk), .Q(v_reg_1_0[2]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_1_ ( .D(maj_151_port_o), .CK(clk), .Q(v_reg_1_0[1]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_0_ ( .D(maj_127_port_o), .CK(clk), .Q(v_reg_1_0[0]), 
        .QN() );
  XNOR2_X1 U223 ( .A(n57), .B(n58), .ZN(n56) );
  NAND2_X1 U224 ( .A1(v_reg_3_1[0]), .A2(a_reg_3[0]), .ZN(n57) );
  NAND2_X1 U225 ( .A1(v_reg_3_0[0]), .A2(a_reg_3[0]), .ZN(n58) );
  XNOR2_X1 U226 ( .A(n49), .B(n50), .ZN(n48) );
  NAND2_X1 U227 ( .A1(v_reg_3_1[1]), .A2(a_reg_3[1]), .ZN(n49) );
  NAND2_X1 U228 ( .A1(v_reg_3_0[1]), .A2(a_reg_3[1]), .ZN(n50) );
  XNOR2_X1 U229 ( .A(n41), .B(n42), .ZN(n40) );
  NAND2_X1 U230 ( .A1(v_reg_3_1[2]), .A2(a_reg_3[2]), .ZN(n41) );
  NAND2_X1 U231 ( .A1(v_reg_3_0[2]), .A2(a_reg_3[2]), .ZN(n42) );
  XNOR2_X1 U232 ( .A(n33), .B(n34), .ZN(n32) );
  NAND2_X1 U233 ( .A1(v_reg_3_1[3]), .A2(a_reg_3[3]), .ZN(n33) );
  NAND2_X1 U234 ( .A1(v_reg_3_0[3]), .A2(a_reg_3[3]), .ZN(n34) );
  XNOR2_X1 U235 ( .A(n25), .B(n26), .ZN(n24) );
  NAND2_X1 U236 ( .A1(v_reg_3_1[4]), .A2(a_reg_3[4]), .ZN(n25) );
  NAND2_X1 U237 ( .A1(v_reg_3_0[4]), .A2(a_reg_3[4]), .ZN(n26) );
  XNOR2_X1 U238 ( .A(n97), .B(n98), .ZN(n96) );
  NAND2_X1 U239 ( .A1(v_reg_2_1[0]), .A2(a_reg_2[0]), .ZN(n97) );
  NAND2_X1 U240 ( .A1(v_reg_2_0[0]), .A2(a_reg_2[0]), .ZN(n98) );
  XNOR2_X1 U241 ( .A(n89), .B(n90), .ZN(n88) );
  NAND2_X1 U242 ( .A1(v_reg_2_1[1]), .A2(a_reg_2[1]), .ZN(n89) );
  NAND2_X1 U243 ( .A1(v_reg_2_0[1]), .A2(a_reg_2[1]), .ZN(n90) );
  XNOR2_X1 U244 ( .A(n81), .B(n82), .ZN(n80) );
  NAND2_X1 U245 ( .A1(v_reg_2_1[2]), .A2(a_reg_2[2]), .ZN(n81) );
  NAND2_X1 U246 ( .A1(v_reg_2_0[2]), .A2(a_reg_2[2]), .ZN(n82) );
  XNOR2_X1 U247 ( .A(n73), .B(n74), .ZN(n72) );
  NAND2_X1 U248 ( .A1(v_reg_2_1[3]), .A2(a_reg_2[3]), .ZN(n73) );
  NAND2_X1 U249 ( .A1(v_reg_2_0[3]), .A2(a_reg_2[3]), .ZN(n74) );
  XNOR2_X1 U250 ( .A(n65), .B(n66), .ZN(n64) );
  NAND2_X1 U251 ( .A1(v_reg_2_1[4]), .A2(a_reg_2[4]), .ZN(n65) );
  NAND2_X1 U252 ( .A1(v_reg_2_0[4]), .A2(a_reg_2[4]), .ZN(n66) );
  XNOR2_X1 U253 ( .A(n137), .B(n138), .ZN(n136) );
  NAND2_X1 U254 ( .A1(v_reg_1_1[0]), .A2(a_reg_1[0]), .ZN(n137) );
  NAND2_X1 U255 ( .A1(v_reg_1_0[0]), .A2(a_reg_1[0]), .ZN(n138) );
  XNOR2_X1 U256 ( .A(n129), .B(n130), .ZN(n128) );
  NAND2_X1 U257 ( .A1(v_reg_1_1[1]), .A2(a_reg_1[1]), .ZN(n129) );
  NAND2_X1 U258 ( .A1(v_reg_1_0[1]), .A2(a_reg_1[1]), .ZN(n130) );
  XNOR2_X1 U259 ( .A(n121), .B(n122), .ZN(n120) );
  NAND2_X1 U260 ( .A1(v_reg_1_1[2]), .A2(a_reg_1[2]), .ZN(n121) );
  NAND2_X1 U261 ( .A1(v_reg_1_0[2]), .A2(a_reg_1[2]), .ZN(n122) );
  XNOR2_X1 U262 ( .A(n113), .B(n114), .ZN(n112) );
  NAND2_X1 U263 ( .A1(v_reg_1_1[3]), .A2(a_reg_1[3]), .ZN(n113) );
  NAND2_X1 U264 ( .A1(v_reg_1_0[3]), .A2(a_reg_1[3]), .ZN(n114) );
  XNOR2_X1 U265 ( .A(n105), .B(n106), .ZN(n104) );
  NAND2_X1 U266 ( .A1(v_reg_1_1[4]), .A2(a_reg_1[4]), .ZN(n105) );
  NAND2_X1 U267 ( .A1(v_reg_1_0[4]), .A2(a_reg_1[4]), .ZN(n106) );
  XNOR2_X1 U268 ( .A(n177), .B(n178), .ZN(n176) );
  NAND2_X1 U269 ( .A1(v_reg_0_1[0]), .A2(a_reg_0[0]), .ZN(n177) );
  NAND2_X1 U270 ( .A1(v_reg_0_0[0]), .A2(a_reg_0[0]), .ZN(n178) );
  XNOR2_X1 U271 ( .A(n169), .B(n170), .ZN(n168) );
  NAND2_X1 U272 ( .A1(v_reg_0_1[1]), .A2(a_reg_0[1]), .ZN(n169) );
  NAND2_X1 U273 ( .A1(v_reg_0_0[1]), .A2(a_reg_0[1]), .ZN(n170) );
  XNOR2_X1 U274 ( .A(n161), .B(n162), .ZN(n160) );
  NAND2_X1 U275 ( .A1(v_reg_0_1[2]), .A2(a_reg_0[2]), .ZN(n161) );
  NAND2_X1 U276 ( .A1(v_reg_0_0[2]), .A2(a_reg_0[2]), .ZN(n162) );
  XNOR2_X1 U277 ( .A(n153), .B(n154), .ZN(n152) );
  NAND2_X1 U278 ( .A1(v_reg_0_1[3]), .A2(a_reg_0[3]), .ZN(n153) );
  NAND2_X1 U279 ( .A1(v_reg_0_0[3]), .A2(a_reg_0[3]), .ZN(n154) );
  XNOR2_X1 U280 ( .A(n145), .B(n146), .ZN(n144) );
  NAND2_X1 U281 ( .A1(v_reg_0_1[4]), .A2(a_reg_0[4]), .ZN(n145) );
  NAND2_X1 U282 ( .A1(v_reg_0_0[4]), .A2(a_reg_0[4]), .ZN(n146) );
  XNOR2_X1 U283 ( .A(u_reg_3_0[0]), .B(temp_0_3[0]), .ZN(n60) );
  XNOR2_X1 U284 ( .A(u_reg_3_0[1]), .B(temp_0_3[1]), .ZN(n52) );
  XNOR2_X1 U285 ( .A(u_reg_3_0[2]), .B(temp_0_3[2]), .ZN(n44) );
  XNOR2_X1 U286 ( .A(u_reg_3_0[3]), .B(temp_0_3[3]), .ZN(n36) );
  XNOR2_X1 U287 ( .A(u_reg_3_0[4]), .B(temp_0_3[4]), .ZN(n28) );
  XNOR2_X1 U288 ( .A(u_reg_2_0[0]), .B(temp_0_2[0]), .ZN(n100) );
  XNOR2_X1 U289 ( .A(u_reg_2_0[1]), .B(temp_0_2[1]), .ZN(n92) );
  XNOR2_X1 U290 ( .A(u_reg_2_0[2]), .B(temp_0_2[2]), .ZN(n84) );
  XNOR2_X1 U291 ( .A(u_reg_2_0[3]), .B(temp_0_2[3]), .ZN(n76) );
  XNOR2_X1 U292 ( .A(u_reg_2_0[4]), .B(temp_0_2[4]), .ZN(n68) );
  XNOR2_X1 U293 ( .A(u_reg_1_0[0]), .B(temp_0_1[0]), .ZN(n140) );
  XNOR2_X1 U294 ( .A(u_reg_1_0[1]), .B(temp_0_1[1]), .ZN(n132) );
  XNOR2_X1 U295 ( .A(u_reg_1_0[2]), .B(temp_0_1[2]), .ZN(n124) );
  XNOR2_X1 U296 ( .A(u_reg_1_0[3]), .B(temp_0_1[3]), .ZN(n116) );
  XNOR2_X1 U297 ( .A(u_reg_1_0[4]), .B(temp_0_1[4]), .ZN(n108) );
  XNOR2_X1 U298 ( .A(u_reg_0_0[0]), .B(temp_0_0[0]), .ZN(n180) );
  XNOR2_X1 U299 ( .A(u_reg_0_0[1]), .B(temp_0_0[1]), .ZN(n172) );
  XNOR2_X1 U300 ( .A(u_reg_0_0[2]), .B(temp_0_0[2]), .ZN(n164) );
  XNOR2_X1 U301 ( .A(u_reg_0_0[3]), .B(temp_0_0[3]), .ZN(n156) );
  XNOR2_X1 U302 ( .A(u_reg_0_0[4]), .B(temp_0_0[4]), .ZN(n148) );
  INV_X1 U303 ( .A(port_a_0[2]), .ZN(n3) );
  INV_X1 U304 ( .A(port_a_0[1]), .ZN(n4) );
  INV_X1 U305 ( .A(port_a_0[0]), .ZN(n5) );
  INV_X1 U306 ( .A(port_a_0[4]), .ZN(n1) );
  INV_X1 U307 ( .A(port_a_0[3]), .ZN(n2) );
  INV_X1 U308 ( .A(port_a_3[2]), .ZN(n18) );
  INV_X1 U309 ( .A(port_a_3[1]), .ZN(n19) );
  INV_X1 U310 ( .A(port_a_3[0]), .ZN(n20) );
  INV_X1 U311 ( .A(port_a_3[4]), .ZN(n16) );
  INV_X1 U312 ( .A(port_a_3[3]), .ZN(n17) );
  INV_X1 U313 ( .A(port_a_2[2]), .ZN(n13) );
  INV_X1 U314 ( .A(port_a_2[1]), .ZN(n14) );
  INV_X1 U315 ( .A(port_a_2[0]), .ZN(n15) );
  INV_X1 U316 ( .A(port_a_2[4]), .ZN(n11) );
  INV_X1 U317 ( .A(port_a_2[3]), .ZN(n12) );
  INV_X1 U318 ( .A(port_a_1[2]), .ZN(n8) );
  INV_X1 U319 ( .A(port_a_1[1]), .ZN(n9) );
  INV_X1 U320 ( .A(port_a_1[0]), .ZN(n10) );
  INV_X1 U321 ( .A(port_a_1[4]), .ZN(n6) );
  INV_X1 U322 ( .A(port_a_1[3]), .ZN(n7) );
  XOR2_X1 U323 ( .A(n53), .B(n54), .Z(port_c_3[0]) );
  XOR2_X1 U324 ( .A(n59), .B(n60), .Z(n53) );
  XOR2_X1 U325 ( .A(n55), .B(n56), .Z(n54) );
  XNOR2_X1 U326 ( .A(u_reg_3_2[0]), .B(u_reg_3_1[0]), .ZN(n59) );
  XOR2_X1 U327 ( .A(n45), .B(n46), .Z(port_c_3[1]) );
  XOR2_X1 U328 ( .A(n51), .B(n52), .Z(n45) );
  XOR2_X1 U329 ( .A(n47), .B(n48), .Z(n46) );
  XNOR2_X1 U330 ( .A(u_reg_3_2[1]), .B(u_reg_3_1[1]), .ZN(n51) );
  XOR2_X1 U331 ( .A(n37), .B(n38), .Z(port_c_3[2]) );
  XOR2_X1 U332 ( .A(n43), .B(n44), .Z(n37) );
  XOR2_X1 U333 ( .A(n39), .B(n40), .Z(n38) );
  XNOR2_X1 U334 ( .A(u_reg_3_2[2]), .B(u_reg_3_1[2]), .ZN(n43) );
  XOR2_X1 U335 ( .A(n29), .B(n30), .Z(port_c_3[3]) );
  XOR2_X1 U336 ( .A(n35), .B(n36), .Z(n29) );
  XOR2_X1 U337 ( .A(n31), .B(n32), .Z(n30) );
  XNOR2_X1 U338 ( .A(u_reg_3_2[3]), .B(u_reg_3_1[3]), .ZN(n35) );
  XOR2_X1 U339 ( .A(n21), .B(n22), .Z(port_c_3[4]) );
  XOR2_X1 U340 ( .A(n27), .B(n28), .Z(n21) );
  XOR2_X1 U341 ( .A(n23), .B(n24), .Z(n22) );
  XNOR2_X1 U342 ( .A(u_reg_3_2[4]), .B(u_reg_3_1[4]), .ZN(n27) );
  XOR2_X1 U343 ( .A(n93), .B(n94), .Z(port_c_2[0]) );
  XOR2_X1 U344 ( .A(n99), .B(n100), .Z(n93) );
  XOR2_X1 U345 ( .A(n95), .B(n96), .Z(n94) );
  XNOR2_X1 U346 ( .A(u_reg_2_2[0]), .B(u_reg_2_1[0]), .ZN(n99) );
  XOR2_X1 U347 ( .A(n85), .B(n86), .Z(port_c_2[1]) );
  XOR2_X1 U348 ( .A(n91), .B(n92), .Z(n85) );
  XOR2_X1 U349 ( .A(n87), .B(n88), .Z(n86) );
  XNOR2_X1 U350 ( .A(u_reg_2_2[1]), .B(u_reg_2_1[1]), .ZN(n91) );
  XOR2_X1 U351 ( .A(n77), .B(n78), .Z(port_c_2[2]) );
  XOR2_X1 U352 ( .A(n83), .B(n84), .Z(n77) );
  XOR2_X1 U353 ( .A(n79), .B(n80), .Z(n78) );
  XNOR2_X1 U354 ( .A(u_reg_2_2[2]), .B(u_reg_2_1[2]), .ZN(n83) );
  XOR2_X1 U355 ( .A(n69), .B(n70), .Z(port_c_2[3]) );
  XOR2_X1 U356 ( .A(n75), .B(n76), .Z(n69) );
  XOR2_X1 U357 ( .A(n71), .B(n72), .Z(n70) );
  XNOR2_X1 U358 ( .A(u_reg_2_2[3]), .B(u_reg_2_1[3]), .ZN(n75) );
  XOR2_X1 U359 ( .A(n61), .B(n62), .Z(port_c_2[4]) );
  XOR2_X1 U360 ( .A(n67), .B(n68), .Z(n61) );
  XOR2_X1 U361 ( .A(n63), .B(n64), .Z(n62) );
  XNOR2_X1 U362 ( .A(u_reg_2_2[4]), .B(u_reg_2_1[4]), .ZN(n67) );
  XOR2_X1 U363 ( .A(n133), .B(n134), .Z(port_c_1[0]) );
  XOR2_X1 U364 ( .A(n139), .B(n140), .Z(n133) );
  XOR2_X1 U365 ( .A(n135), .B(n136), .Z(n134) );
  XNOR2_X1 U366 ( .A(u_reg_1_2[0]), .B(u_reg_1_1[0]), .ZN(n139) );
  XOR2_X1 U367 ( .A(n125), .B(n126), .Z(port_c_1[1]) );
  XOR2_X1 U368 ( .A(n131), .B(n132), .Z(n125) );
  XOR2_X1 U369 ( .A(n127), .B(n128), .Z(n126) );
  XNOR2_X1 U370 ( .A(u_reg_1_2[1]), .B(u_reg_1_1[1]), .ZN(n131) );
  XOR2_X1 U371 ( .A(n117), .B(n118), .Z(port_c_1[2]) );
  XOR2_X1 U372 ( .A(n123), .B(n124), .Z(n117) );
  XOR2_X1 U373 ( .A(n119), .B(n120), .Z(n118) );
  XNOR2_X1 U374 ( .A(u_reg_1_2[2]), .B(u_reg_1_1[2]), .ZN(n123) );
  XOR2_X1 U375 ( .A(n109), .B(n110), .Z(port_c_1[3]) );
  XOR2_X1 U376 ( .A(n115), .B(n116), .Z(n109) );
  XOR2_X1 U377 ( .A(n111), .B(n112), .Z(n110) );
  XNOR2_X1 U378 ( .A(u_reg_1_2[3]), .B(u_reg_1_1[3]), .ZN(n115) );
  XOR2_X1 U379 ( .A(n101), .B(n102), .Z(port_c_1[4]) );
  XOR2_X1 U380 ( .A(n107), .B(n108), .Z(n101) );
  XOR2_X1 U381 ( .A(n103), .B(n104), .Z(n102) );
  XNOR2_X1 U382 ( .A(u_reg_1_2[4]), .B(u_reg_1_1[4]), .ZN(n107) );
  XOR2_X1 U383 ( .A(n173), .B(n174), .Z(port_c_0[0]) );
  XOR2_X1 U384 ( .A(n179), .B(n180), .Z(n173) );
  XOR2_X1 U385 ( .A(n175), .B(n176), .Z(n174) );
  XNOR2_X1 U386 ( .A(u_reg_0_2[0]), .B(u_reg_0_1[0]), .ZN(n179) );
  XOR2_X1 U387 ( .A(n165), .B(n166), .Z(port_c_0[1]) );
  XOR2_X1 U388 ( .A(n171), .B(n172), .Z(n165) );
  XOR2_X1 U389 ( .A(n167), .B(n168), .Z(n166) );
  XNOR2_X1 U390 ( .A(u_reg_0_2[1]), .B(u_reg_0_1[1]), .ZN(n171) );
  XOR2_X1 U391 ( .A(n157), .B(n158), .Z(port_c_0[2]) );
  XOR2_X1 U392 ( .A(n163), .B(n164), .Z(n157) );
  XOR2_X1 U393 ( .A(n159), .B(n160), .Z(n158) );
  XNOR2_X1 U394 ( .A(u_reg_0_2[2]), .B(u_reg_0_1[2]), .ZN(n163) );
  XOR2_X1 U395 ( .A(n149), .B(n150), .Z(port_c_0[3]) );
  XOR2_X1 U396 ( .A(n155), .B(n156), .Z(n149) );
  XOR2_X1 U397 ( .A(n151), .B(n152), .Z(n150) );
  XNOR2_X1 U398 ( .A(u_reg_0_2[3]), .B(u_reg_0_1[3]), .ZN(n155) );
  XOR2_X1 U399 ( .A(n141), .B(n142), .Z(port_c_0[4]) );
  XOR2_X1 U400 ( .A(n147), .B(n148), .Z(n141) );
  XOR2_X1 U401 ( .A(n143), .B(n144), .Z(n142) );
  XNOR2_X1 U402 ( .A(u_reg_0_2[4]), .B(u_reg_0_1[4]), .ZN(n147) );
  NAND2_X1 U403 ( .A1(v_reg_3_2[0]), .A2(a_reg_3[0]), .ZN(n55) );
  NAND2_X1 U404 ( .A1(v_reg_3_2[1]), .A2(a_reg_3[1]), .ZN(n47) );
  NAND2_X1 U405 ( .A1(v_reg_3_2[2]), .A2(a_reg_3[2]), .ZN(n39) );
  NAND2_X1 U406 ( .A1(v_reg_3_2[3]), .A2(a_reg_3[3]), .ZN(n31) );
  NAND2_X1 U407 ( .A1(v_reg_3_2[4]), .A2(a_reg_3[4]), .ZN(n23) );
  NAND2_X1 U408 ( .A1(v_reg_2_2[0]), .A2(a_reg_2[0]), .ZN(n95) );
  NAND2_X1 U409 ( .A1(v_reg_2_2[1]), .A2(a_reg_2[1]), .ZN(n87) );
  NAND2_X1 U410 ( .A1(v_reg_2_2[2]), .A2(a_reg_2[2]), .ZN(n79) );
  NAND2_X1 U411 ( .A1(v_reg_2_2[3]), .A2(a_reg_2[3]), .ZN(n71) );
  NAND2_X1 U412 ( .A1(v_reg_2_2[4]), .A2(a_reg_2[4]), .ZN(n63) );
  NAND2_X1 U413 ( .A1(v_reg_1_2[0]), .A2(a_reg_1[0]), .ZN(n135) );
  NAND2_X1 U414 ( .A1(v_reg_1_2[1]), .A2(a_reg_1[1]), .ZN(n127) );
  NAND2_X1 U415 ( .A1(v_reg_1_2[2]), .A2(a_reg_1[2]), .ZN(n119) );
  NAND2_X1 U416 ( .A1(v_reg_1_2[3]), .A2(a_reg_1[3]), .ZN(n111) );
  NAND2_X1 U417 ( .A1(v_reg_1_2[4]), .A2(a_reg_1[4]), .ZN(n103) );
  NAND2_X1 U418 ( .A1(v_reg_0_2[0]), .A2(a_reg_0[0]), .ZN(n175) );
  NAND2_X1 U419 ( .A1(v_reg_0_2[1]), .A2(a_reg_0[1]), .ZN(n167) );
  NAND2_X1 U420 ( .A1(v_reg_0_2[2]), .A2(a_reg_0[2]), .ZN(n159) );
  NAND2_X1 U421 ( .A1(v_reg_0_2[3]), .A2(a_reg_0[3]), .ZN(n151) );
  NAND2_X1 U422 ( .A1(v_reg_0_2[4]), .A2(a_reg_0[4]), .ZN(n143) );
  AND2_X1 U423 ( .A1(port_b_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U424 ( .A1(port_b_0[1]), .A2(port_a_0[1]), .ZN(N4) );
  AND2_X1 U425 ( .A1(port_b_0[2]), .A2(port_a_0[2]), .ZN(N8) );
  AND2_X1 U426 ( .A1(port_b_0[3]), .A2(port_a_0[3]), .ZN(N12) );
  AND2_X1 U427 ( .A1(port_b_0[4]), .A2(port_a_0[4]), .ZN(N16) );
  AND2_X1 U428 ( .A1(port_b_1[0]), .A2(port_a_1[0]), .ZN(N1) );
  AND2_X1 U429 ( .A1(port_b_1[1]), .A2(port_a_1[1]), .ZN(N5) );
  AND2_X1 U430 ( .A1(port_b_1[2]), .A2(port_a_1[2]), .ZN(N9) );
  AND2_X1 U431 ( .A1(port_b_1[3]), .A2(port_a_1[3]), .ZN(N13) );
  AND2_X1 U432 ( .A1(port_b_1[4]), .A2(port_a_1[4]), .ZN(N17) );
  AND2_X1 U433 ( .A1(port_b_2[0]), .A2(port_a_2[0]), .ZN(N2) );
  AND2_X1 U434 ( .A1(port_b_2[1]), .A2(port_a_2[1]), .ZN(N6) );
  AND2_X1 U435 ( .A1(port_b_2[2]), .A2(port_a_2[2]), .ZN(N10) );
  AND2_X1 U436 ( .A1(port_b_2[3]), .A2(port_a_2[3]), .ZN(N14) );
  AND2_X1 U437 ( .A1(port_b_2[4]), .A2(port_a_2[4]), .ZN(N18) );
  AND2_X1 U438 ( .A1(port_b_3[0]), .A2(port_a_3[0]), .ZN(N3) );
  AND2_X1 U439 ( .A1(port_b_3[1]), .A2(port_a_3[1]), .ZN(N7) );
  AND2_X1 U440 ( .A1(port_b_3[2]), .A2(port_a_3[2]), .ZN(N11) );
  AND2_X1 U441 ( .A1(port_b_3[3]), .A2(port_a_3[3]), .ZN(N15) );
  AND2_X1 U442 ( .A1(port_b_3[4]), .A2(port_a_3[4]), .ZN(N19) );
  AND2_X1 simpleAnd_60_U1 ( .A1(port_rand_mul[0]), .A2(n5), .ZN(
        simpleAnd_60_port_z) );
  XOR2_X2 simpleXor_120_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_60_port_z), 
        .Z(u_0_0[0]) );
  XOR2_X2 simpleXor_121_U1 ( .A(port_rand_mul[0]), .B(port_b_1[0]), .Z(
        v_0_0[0]) );
  AND2_X1 simpleAnd_61_U1 ( .A1(port_rand_mul[1]), .A2(n5), .ZN(
        simpleAnd_61_port_z) );
  XOR2_X2 simpleXor_122_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_61_port_z), 
        .Z(u_0_1[0]) );
  XOR2_X2 simpleXor_123_U1 ( .A(port_rand_mul[1]), .B(port_b_2[0]), .Z(
        v_0_1[0]) );
  AND2_X1 simpleAnd_62_U1 ( .A1(port_rand_mul[2]), .A2(n5), .ZN(
        simpleAnd_62_port_z) );
  XOR2_X2 simpleXor_124_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_62_port_z), 
        .Z(u_0_2[0]) );
  XOR2_X2 simpleXor_125_U1 ( .A(port_rand_mul[2]), .B(port_b_3[0]), .Z(
        v_0_2[0]) );
  AND2_X1 simpleAnd_63_U1 ( .A1(port_rand_mul[0]), .A2(n10), .ZN(
        simpleAnd_63_port_z) );
  XOR2_X2 simpleXor_126_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_63_port_z), 
        .Z(u_1_0[0]) );
  XOR2_X2 simpleXor_127_U1 ( .A(port_rand_mul[0]), .B(port_b_0[0]), .Z(
        v_1_0[0]) );
  AND2_X1 simpleAnd_64_U1 ( .A1(port_rand_mul[3]), .A2(n10), .ZN(
        simpleAnd_64_port_z) );
  XOR2_X2 simpleXor_128_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_64_port_z), 
        .Z(u_1_1[0]) );
  XOR2_X2 simpleXor_129_U1 ( .A(port_rand_mul[3]), .B(port_b_2[0]), .Z(
        v_1_1[0]) );
  AND2_X1 simpleAnd_65_U1 ( .A1(port_rand_mul[4]), .A2(n10), .ZN(
        simpleAnd_65_port_z) );
  XOR2_X2 simpleXor_130_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_65_port_z), 
        .Z(u_1_2[0]) );
  XOR2_X2 simpleXor_131_U1 ( .A(port_rand_mul[4]), .B(port_b_3[0]), .Z(
        v_1_2[0]) );
  AND2_X1 simpleAnd_66_U1 ( .A1(port_rand_mul[1]), .A2(n15), .ZN(
        simpleAnd_66_port_z) );
  XOR2_X2 simpleXor_132_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_66_port_z), 
        .Z(u_2_0[0]) );
  XOR2_X2 simpleXor_133_U1 ( .A(port_rand_mul[1]), .B(port_b_0[0]), .Z(
        v_2_0[0]) );
  AND2_X1 simpleAnd_67_U1 ( .A1(port_rand_mul[3]), .A2(n15), .ZN(
        simpleAnd_67_port_z) );
  XOR2_X2 simpleXor_134_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_67_port_z), 
        .Z(u_2_1[0]) );
  XOR2_X2 simpleXor_135_U1 ( .A(port_rand_mul[3]), .B(port_b_1[0]), .Z(
        v_2_1[0]) );
  AND2_X1 simpleAnd_68_U1 ( .A1(port_rand_mul[5]), .A2(n15), .ZN(
        simpleAnd_68_port_z) );
  XOR2_X2 simpleXor_136_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_68_port_z), 
        .Z(u_2_2[0]) );
  XOR2_X2 simpleXor_137_U1 ( .A(port_rand_mul[5]), .B(port_b_3[0]), .Z(
        v_2_2[0]) );
  AND2_X1 simpleAnd_69_U1 ( .A1(port_rand_mul[2]), .A2(n20), .ZN(
        simpleAnd_69_port_z) );
  XOR2_X2 simpleXor_138_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_69_port_z), 
        .Z(u_3_0[0]) );
  XOR2_X2 simpleXor_139_U1 ( .A(port_rand_mul[2]), .B(port_b_0[0]), .Z(
        v_3_0[0]) );
  AND2_X1 simpleAnd_70_U1 ( .A1(port_rand_mul[4]), .A2(n20), .ZN(
        simpleAnd_70_port_z) );
  XOR2_X2 simpleXor_140_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_70_port_z), 
        .Z(u_3_1[0]) );
  XOR2_X2 simpleXor_141_U1 ( .A(port_rand_mul[4]), .B(port_b_1[0]), .Z(
        v_3_1[0]) );
  AND2_X1 simpleAnd_71_U1 ( .A1(port_rand_mul[5]), .A2(n20), .ZN(
        simpleAnd_71_port_z) );
  XOR2_X2 simpleXor_142_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_71_port_z), 
        .Z(u_3_2[0]) );
  XOR2_X2 simpleXor_143_U1 ( .A(port_rand_mul[5]), .B(port_b_2[0]), .Z(
        v_3_2[0]) );
  AND2_X1 simpleAnd_72_U1 ( .A1(port_rand_mul[0]), .A2(n4), .ZN(
        simpleAnd_72_port_z) );
  XOR2_X2 simpleXor_144_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_72_port_z), 
        .Z(u_0_0[1]) );
  XOR2_X2 simpleXor_145_U1 ( .A(port_rand_mul[0]), .B(port_b_1[1]), .Z(
        v_0_0[1]) );
  AND2_X1 simpleAnd_73_U1 ( .A1(port_rand_mul[1]), .A2(n4), .ZN(
        simpleAnd_73_port_z) );
  XOR2_X2 simpleXor_146_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_73_port_z), 
        .Z(u_0_1[1]) );
  XOR2_X2 simpleXor_147_U1 ( .A(port_rand_mul[1]), .B(port_b_2[1]), .Z(
        v_0_1[1]) );
  AND2_X1 simpleAnd_74_U1 ( .A1(port_rand_mul[2]), .A2(n4), .ZN(
        simpleAnd_74_port_z) );
  XOR2_X2 simpleXor_148_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_74_port_z), 
        .Z(u_0_2[1]) );
  XOR2_X2 simpleXor_149_U1 ( .A(port_rand_mul[2]), .B(port_b_3[1]), .Z(
        v_0_2[1]) );
  AND2_X1 simpleAnd_75_U1 ( .A1(port_rand_mul[0]), .A2(n9), .ZN(
        simpleAnd_75_port_z) );
  XOR2_X2 simpleXor_150_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_75_port_z), 
        .Z(u_1_0[1]) );
  XOR2_X2 simpleXor_151_U1 ( .A(port_rand_mul[0]), .B(port_b_0[1]), .Z(
        v_1_0[1]) );
  AND2_X1 simpleAnd_76_U1 ( .A1(port_rand_mul[3]), .A2(n9), .ZN(
        simpleAnd_76_port_z) );
  XOR2_X2 simpleXor_152_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_76_port_z), 
        .Z(u_1_1[1]) );
  XOR2_X2 simpleXor_153_U1 ( .A(port_rand_mul[3]), .B(port_b_2[1]), .Z(
        v_1_1[1]) );
  AND2_X1 simpleAnd_77_U1 ( .A1(port_rand_mul[4]), .A2(n9), .ZN(
        simpleAnd_77_port_z) );
  XOR2_X2 simpleXor_154_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_77_port_z), 
        .Z(u_1_2[1]) );
  XOR2_X2 simpleXor_155_U1 ( .A(port_rand_mul[4]), .B(port_b_3[1]), .Z(
        v_1_2[1]) );
  AND2_X1 simpleAnd_78_U1 ( .A1(port_rand_mul[1]), .A2(n14), .ZN(
        simpleAnd_78_port_z) );
  XOR2_X2 simpleXor_156_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_78_port_z), 
        .Z(u_2_0[1]) );
  XOR2_X2 simpleXor_157_U1 ( .A(port_rand_mul[1]), .B(port_b_0[1]), .Z(
        v_2_0[1]) );
  AND2_X1 simpleAnd_79_U1 ( .A1(port_rand_mul[3]), .A2(n14), .ZN(
        simpleAnd_79_port_z) );
  XOR2_X2 simpleXor_158_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_79_port_z), 
        .Z(u_2_1[1]) );
  XOR2_X2 simpleXor_159_U1 ( .A(port_rand_mul[3]), .B(port_b_1[1]), .Z(
        v_2_1[1]) );
  AND2_X1 simpleAnd_80_U1 ( .A1(port_rand_mul[5]), .A2(n14), .ZN(
        simpleAnd_80_port_z) );
  XOR2_X2 simpleXor_160_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_80_port_z), 
        .Z(u_2_2[1]) );
  XOR2_X2 simpleXor_161_U1 ( .A(port_rand_mul[5]), .B(port_b_3[1]), .Z(
        v_2_2[1]) );
  AND2_X1 simpleAnd_81_U1 ( .A1(port_rand_mul[2]), .A2(n19), .ZN(
        simpleAnd_81_port_z) );
  XOR2_X2 simpleXor_162_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_81_port_z), 
        .Z(u_3_0[1]) );
  XOR2_X2 simpleXor_163_U1 ( .A(port_rand_mul[2]), .B(port_b_0[1]), .Z(
        v_3_0[1]) );
  AND2_X1 simpleAnd_82_U1 ( .A1(port_rand_mul[4]), .A2(n19), .ZN(
        simpleAnd_82_port_z) );
  XOR2_X2 simpleXor_164_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_82_port_z), 
        .Z(u_3_1[1]) );
  XOR2_X2 simpleXor_165_U1 ( .A(port_rand_mul[4]), .B(port_b_1[1]), .Z(
        v_3_1[1]) );
  AND2_X1 simpleAnd_83_U1 ( .A1(port_rand_mul[5]), .A2(n19), .ZN(
        simpleAnd_83_port_z) );
  XOR2_X2 simpleXor_166_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_83_port_z), 
        .Z(u_3_2[1]) );
  XOR2_X2 simpleXor_167_U1 ( .A(port_rand_mul[5]), .B(port_b_2[1]), .Z(
        v_3_2[1]) );
  AND2_X1 simpleAnd_84_U1 ( .A1(port_rand_mul[0]), .A2(n3), .ZN(
        simpleAnd_84_port_z) );
  XOR2_X2 simpleXor_168_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_84_port_z), 
        .Z(u_0_0[2]) );
  XOR2_X2 simpleXor_169_U1 ( .A(port_rand_mul[0]), .B(port_b_1[2]), .Z(
        v_0_0[2]) );
  AND2_X1 simpleAnd_85_U1 ( .A1(port_rand_mul[1]), .A2(n3), .ZN(
        simpleAnd_85_port_z) );
  XOR2_X2 simpleXor_170_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_85_port_z), 
        .Z(u_0_1[2]) );
  XOR2_X2 simpleXor_171_U1 ( .A(port_rand_mul[1]), .B(port_b_2[2]), .Z(
        v_0_1[2]) );
  AND2_X1 simpleAnd_86_U1 ( .A1(port_rand_mul[2]), .A2(n3), .ZN(
        simpleAnd_86_port_z) );
  XOR2_X2 simpleXor_172_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_86_port_z), 
        .Z(u_0_2[2]) );
  XOR2_X2 simpleXor_173_U1 ( .A(port_rand_mul[2]), .B(port_b_3[2]), .Z(
        v_0_2[2]) );
  AND2_X1 simpleAnd_87_U1 ( .A1(port_rand_mul[0]), .A2(n8), .ZN(
        simpleAnd_87_port_z) );
  XOR2_X2 simpleXor_174_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_87_port_z), 
        .Z(u_1_0[2]) );
  XOR2_X2 simpleXor_175_U1 ( .A(port_rand_mul[0]), .B(port_b_0[2]), .Z(
        v_1_0[2]) );
  AND2_X1 simpleAnd_88_U1 ( .A1(port_rand_mul[3]), .A2(n8), .ZN(
        simpleAnd_88_port_z) );
  XOR2_X2 simpleXor_176_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_88_port_z), 
        .Z(u_1_1[2]) );
  XOR2_X2 simpleXor_177_U1 ( .A(port_rand_mul[3]), .B(port_b_2[2]), .Z(
        v_1_1[2]) );
  AND2_X1 simpleAnd_89_U1 ( .A1(port_rand_mul[4]), .A2(n8), .ZN(
        simpleAnd_89_port_z) );
  XOR2_X2 simpleXor_178_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_89_port_z), 
        .Z(u_1_2[2]) );
  XOR2_X2 simpleXor_179_U1 ( .A(port_rand_mul[4]), .B(port_b_3[2]), .Z(
        v_1_2[2]) );
  AND2_X1 simpleAnd_90_U1 ( .A1(port_rand_mul[1]), .A2(n13), .ZN(
        simpleAnd_90_port_z) );
  XOR2_X2 simpleXor_180_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_90_port_z), 
        .Z(u_2_0[2]) );
  XOR2_X2 simpleXor_181_U1 ( .A(port_rand_mul[1]), .B(port_b_0[2]), .Z(
        v_2_0[2]) );
  AND2_X1 simpleAnd_91_U1 ( .A1(port_rand_mul[3]), .A2(n13), .ZN(
        simpleAnd_91_port_z) );
  XOR2_X2 simpleXor_182_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_91_port_z), 
        .Z(u_2_1[2]) );
  XOR2_X2 simpleXor_183_U1 ( .A(port_rand_mul[3]), .B(port_b_1[2]), .Z(
        v_2_1[2]) );
  AND2_X1 simpleAnd_92_U1 ( .A1(port_rand_mul[5]), .A2(n13), .ZN(
        simpleAnd_92_port_z) );
  XOR2_X2 simpleXor_184_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_92_port_z), 
        .Z(u_2_2[2]) );
  XOR2_X2 simpleXor_185_U1 ( .A(port_rand_mul[5]), .B(port_b_3[2]), .Z(
        v_2_2[2]) );
  AND2_X1 simpleAnd_93_U1 ( .A1(port_rand_mul[2]), .A2(n18), .ZN(
        simpleAnd_93_port_z) );
  XOR2_X2 simpleXor_186_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_93_port_z), 
        .Z(u_3_0[2]) );
  XOR2_X2 simpleXor_187_U1 ( .A(port_rand_mul[2]), .B(port_b_0[2]), .Z(
        v_3_0[2]) );
  AND2_X1 simpleAnd_94_U1 ( .A1(port_rand_mul[4]), .A2(n18), .ZN(
        simpleAnd_94_port_z) );
  XOR2_X2 simpleXor_188_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_94_port_z), 
        .Z(u_3_1[2]) );
  XOR2_X2 simpleXor_189_U1 ( .A(port_rand_mul[4]), .B(port_b_1[2]), .Z(
        v_3_1[2]) );
  AND2_X1 simpleAnd_95_U1 ( .A1(port_rand_mul[5]), .A2(n18), .ZN(
        simpleAnd_95_port_z) );
  XOR2_X2 simpleXor_190_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_95_port_z), 
        .Z(u_3_2[2]) );
  XOR2_X2 simpleXor_191_U1 ( .A(port_rand_mul[5]), .B(port_b_2[2]), .Z(
        v_3_2[2]) );
  AND2_X1 simpleAnd_96_U1 ( .A1(port_rand_mul[0]), .A2(n2), .ZN(
        simpleAnd_96_port_z) );
  XOR2_X2 simpleXor_192_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_96_port_z), 
        .Z(u_0_0[3]) );
  XOR2_X2 simpleXor_193_U1 ( .A(port_rand_mul[0]), .B(port_b_1[3]), .Z(
        v_0_0[3]) );
  AND2_X1 simpleAnd_97_U1 ( .A1(port_rand_mul[1]), .A2(n2), .ZN(
        simpleAnd_97_port_z) );
  XOR2_X2 simpleXor_194_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_97_port_z), 
        .Z(u_0_1[3]) );
  XOR2_X2 simpleXor_195_U1 ( .A(port_rand_mul[1]), .B(port_b_2[3]), .Z(
        v_0_1[3]) );
  AND2_X1 simpleAnd_98_U1 ( .A1(port_rand_mul[2]), .A2(n2), .ZN(
        simpleAnd_98_port_z) );
  XOR2_X2 simpleXor_196_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_98_port_z), 
        .Z(u_0_2[3]) );
  XOR2_X2 simpleXor_197_U1 ( .A(port_rand_mul[2]), .B(port_b_3[3]), .Z(
        v_0_2[3]) );
  AND2_X1 simpleAnd_99_U1 ( .A1(port_rand_mul[0]), .A2(n7), .ZN(
        simpleAnd_99_port_z) );
  XOR2_X2 simpleXor_198_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_99_port_z), 
        .Z(u_1_0[3]) );
  XOR2_X2 simpleXor_199_U1 ( .A(port_rand_mul[0]), .B(port_b_0[3]), .Z(
        v_1_0[3]) );
  AND2_X1 simpleAnd_100_U1 ( .A1(port_rand_mul[3]), .A2(n7), .ZN(
        simpleAnd_100_port_z) );
  XOR2_X2 simpleXor_200_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_100_port_z), 
        .Z(u_1_1[3]) );
  XOR2_X2 simpleXor_201_U1 ( .A(port_rand_mul[3]), .B(port_b_2[3]), .Z(
        v_1_1[3]) );
  AND2_X1 simpleAnd_101_U1 ( .A1(port_rand_mul[4]), .A2(n7), .ZN(
        simpleAnd_101_port_z) );
  XOR2_X2 simpleXor_202_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_101_port_z), 
        .Z(u_1_2[3]) );
  XOR2_X2 simpleXor_203_U1 ( .A(port_rand_mul[4]), .B(port_b_3[3]), .Z(
        v_1_2[3]) );
  AND2_X1 simpleAnd_102_U1 ( .A1(port_rand_mul[1]), .A2(n12), .ZN(
        simpleAnd_102_port_z) );
  XOR2_X2 simpleXor_204_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_102_port_z), 
        .Z(u_2_0[3]) );
  XOR2_X2 simpleXor_205_U1 ( .A(port_rand_mul[1]), .B(port_b_0[3]), .Z(
        v_2_0[3]) );
  AND2_X1 simpleAnd_103_U1 ( .A1(port_rand_mul[3]), .A2(n12), .ZN(
        simpleAnd_103_port_z) );
  XOR2_X2 simpleXor_206_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_103_port_z), 
        .Z(u_2_1[3]) );
  XOR2_X2 simpleXor_207_U1 ( .A(port_rand_mul[3]), .B(port_b_1[3]), .Z(
        v_2_1[3]) );
  AND2_X1 simpleAnd_104_U1 ( .A1(port_rand_mul[5]), .A2(n12), .ZN(
        simpleAnd_104_port_z) );
  XOR2_X2 simpleXor_208_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_104_port_z), 
        .Z(u_2_2[3]) );
  XOR2_X2 simpleXor_209_U1 ( .A(port_rand_mul[5]), .B(port_b_3[3]), .Z(
        v_2_2[3]) );
  AND2_X1 simpleAnd_105_U1 ( .A1(port_rand_mul[2]), .A2(n17), .ZN(
        simpleAnd_105_port_z) );
  XOR2_X2 simpleXor_210_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_105_port_z), 
        .Z(u_3_0[3]) );
  XOR2_X2 simpleXor_211_U1 ( .A(port_rand_mul[2]), .B(port_b_0[3]), .Z(
        v_3_0[3]) );
  AND2_X1 simpleAnd_106_U1 ( .A1(port_rand_mul[4]), .A2(n17), .ZN(
        simpleAnd_106_port_z) );
  XOR2_X2 simpleXor_212_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_106_port_z), 
        .Z(u_3_1[3]) );
  XOR2_X2 simpleXor_213_U1 ( .A(port_rand_mul[4]), .B(port_b_1[3]), .Z(
        v_3_1[3]) );
  AND2_X1 simpleAnd_107_U1 ( .A1(port_rand_mul[5]), .A2(n17), .ZN(
        simpleAnd_107_port_z) );
  XOR2_X2 simpleXor_214_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_107_port_z), 
        .Z(u_3_2[3]) );
  XOR2_X2 simpleXor_215_U1 ( .A(port_rand_mul[5]), .B(port_b_2[3]), .Z(
        v_3_2[3]) );
  AND2_X1 simpleAnd_108_U1 ( .A1(port_rand_mul[0]), .A2(n1), .ZN(
        simpleAnd_108_port_z) );
  XOR2_X2 simpleXor_216_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_108_port_z), 
        .Z(u_0_0[4]) );
  XOR2_X2 simpleXor_217_U1 ( .A(port_rand_mul[0]), .B(port_b_1[4]), .Z(
        v_0_0[4]) );
  AND2_X1 simpleAnd_109_U1 ( .A1(port_rand_mul[1]), .A2(n1), .ZN(
        simpleAnd_109_port_z) );
  XOR2_X2 simpleXor_218_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_109_port_z), 
        .Z(u_0_1[4]) );
  XOR2_X2 simpleXor_219_U1 ( .A(port_rand_mul[1]), .B(port_b_2[4]), .Z(
        v_0_1[4]) );
  AND2_X1 simpleAnd_110_U1 ( .A1(port_rand_mul[2]), .A2(n1), .ZN(
        simpleAnd_110_port_z) );
  XOR2_X2 simpleXor_220_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_110_port_z), 
        .Z(u_0_2[4]) );
  XOR2_X2 simpleXor_221_U1 ( .A(port_rand_mul[2]), .B(port_b_3[4]), .Z(
        v_0_2[4]) );
  AND2_X1 simpleAnd_111_U1 ( .A1(port_rand_mul[0]), .A2(n6), .ZN(
        simpleAnd_111_port_z) );
  XOR2_X2 simpleXor_222_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_111_port_z), 
        .Z(u_1_0[4]) );
  XOR2_X2 simpleXor_223_U1 ( .A(port_rand_mul[0]), .B(port_b_0[4]), .Z(
        v_1_0[4]) );
  AND2_X1 simpleAnd_112_U1 ( .A1(port_rand_mul[3]), .A2(n6), .ZN(
        simpleAnd_112_port_z) );
  XOR2_X2 simpleXor_224_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_112_port_z), 
        .Z(u_1_1[4]) );
  XOR2_X2 simpleXor_225_U1 ( .A(port_rand_mul[3]), .B(port_b_2[4]), .Z(
        v_1_1[4]) );
  AND2_X1 simpleAnd_113_U1 ( .A1(port_rand_mul[4]), .A2(n6), .ZN(
        simpleAnd_113_port_z) );
  XOR2_X2 simpleXor_226_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_113_port_z), 
        .Z(u_1_2[4]) );
  XOR2_X2 simpleXor_227_U1 ( .A(port_rand_mul[4]), .B(port_b_3[4]), .Z(
        v_1_2[4]) );
  AND2_X1 simpleAnd_114_U1 ( .A1(port_rand_mul[1]), .A2(n11), .ZN(
        simpleAnd_114_port_z) );
  XOR2_X2 simpleXor_228_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_114_port_z), 
        .Z(u_2_0[4]) );
  XOR2_X2 simpleXor_229_U1 ( .A(port_rand_mul[1]), .B(port_b_0[4]), .Z(
        v_2_0[4]) );
  AND2_X1 simpleAnd_115_U1 ( .A1(port_rand_mul[3]), .A2(n11), .ZN(
        simpleAnd_115_port_z) );
  XOR2_X2 simpleXor_230_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_115_port_z), 
        .Z(u_2_1[4]) );
  XOR2_X2 simpleXor_231_U1 ( .A(port_rand_mul[3]), .B(port_b_1[4]), .Z(
        v_2_1[4]) );
  AND2_X1 simpleAnd_116_U1 ( .A1(port_rand_mul[5]), .A2(n11), .ZN(
        simpleAnd_116_port_z) );
  XOR2_X2 simpleXor_232_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_116_port_z), 
        .Z(u_2_2[4]) );
  XOR2_X2 simpleXor_233_U1 ( .A(port_rand_mul[5]), .B(port_b_3[4]), .Z(
        v_2_2[4]) );
  AND2_X1 simpleAnd_117_U1 ( .A1(port_rand_mul[2]), .A2(n16), .ZN(
        simpleAnd_117_port_z) );
  XOR2_X2 simpleXor_234_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_117_port_z), 
        .Z(u_3_0[4]) );
  XOR2_X2 simpleXor_235_U1 ( .A(port_rand_mul[2]), .B(port_b_0[4]), .Z(
        v_3_0[4]) );
  AND2_X1 simpleAnd_118_U1 ( .A1(port_rand_mul[4]), .A2(n16), .ZN(
        simpleAnd_118_port_z) );
  XOR2_X2 simpleXor_236_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_118_port_z), 
        .Z(u_3_1[4]) );
  XOR2_X2 simpleXor_237_U1 ( .A(port_rand_mul[4]), .B(port_b_1[4]), .Z(
        v_3_1[4]) );
  AND2_X1 simpleAnd_119_U1 ( .A1(port_rand_mul[5]), .A2(n16), .ZN(
        simpleAnd_119_port_z) );
  XOR2_X2 simpleXor_238_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_119_port_z), 
        .Z(u_3_2[4]) );
  XOR2_X2 simpleXor_239_U1 ( .A(port_rand_mul[5]), .B(port_b_2[4]), .Z(
        v_3_2[4]) );
  NAND2_X1 maj_120_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_120_n9) );
  NAND2_X1 maj_120_U14 ( .A1(maj_120_n6), .A2(maj_120_n5), .ZN(maj_120_n10) );
  NAND2_X1 maj_120_U13 ( .A1(maj_120_n9), .A2(maj_120_n10), .ZN(maj_120_n8) );
  NAND2_X1 maj_120_U12 ( .A1(u_0_0[2]), .A2(maj_120_n11), .ZN(maj_120_n13) );
  NAND2_X1 maj_120_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_120_n12) );
  NAND2_X1 maj_120_U10 ( .A1(maj_120_n12), .A2(maj_120_n13), .ZN(maj_120_n7)
         );
  XOR2_X1 maj_120_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_120_n5) );
  XOR2_X1 maj_120_U8 ( .A(u_0_0[2]), .B(maj_120_n11), .Z(maj_120_n6) );
  XOR2_X1 maj_120_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_120_n11) );
  OR2_X1 maj_120_U6 ( .A1(maj_120_n7), .A2(maj_120_n8), .ZN(maj_120_n3) );
  NAND2_X1 maj_120_U5 ( .A1(maj_120_n3), .A2(maj_120_n4), .ZN(maj_120_n2) );
  NAND2_X1 maj_120_U4 ( .A1(maj_120_n7), .A2(maj_120_n8), .ZN(maj_120_n1) );
  NAND2_X1 maj_120_U3 ( .A1(maj_120_n1), .A2(maj_120_n2), .ZN(maj_120_port_o)
         );
  XOR2_X1 maj_120_U2 ( .A(maj_120_n5), .B(maj_120_n6), .Z(maj_120_n4) );
  NAND2_X1 maj_121_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_121_n18) );
  NAND2_X1 maj_121_U14 ( .A1(maj_121_n21), .A2(maj_121_n22), .ZN(maj_121_n17)
         );
  NAND2_X1 maj_121_U13 ( .A1(maj_121_n18), .A2(maj_121_n17), .ZN(maj_121_n19)
         );
  NAND2_X1 maj_121_U12 ( .A1(v_0_0[2]), .A2(maj_121_n16), .ZN(maj_121_n14) );
  NAND2_X1 maj_121_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_121_n15) );
  NAND2_X1 maj_121_U10 ( .A1(maj_121_n15), .A2(maj_121_n14), .ZN(maj_121_n20)
         );
  XOR2_X1 maj_121_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_121_n22) );
  XOR2_X1 maj_121_U8 ( .A(v_0_0[2]), .B(maj_121_n16), .Z(maj_121_n21) );
  XOR2_X1 maj_121_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_121_n16) );
  OR2_X1 maj_121_U6 ( .A1(maj_121_n20), .A2(maj_121_n19), .ZN(maj_121_n24) );
  NAND2_X1 maj_121_U5 ( .A1(maj_121_n24), .A2(maj_121_n23), .ZN(maj_121_n25)
         );
  NAND2_X1 maj_121_U4 ( .A1(maj_121_n20), .A2(maj_121_n19), .ZN(maj_121_n26)
         );
  NAND2_X1 maj_121_U3 ( .A1(maj_121_n26), .A2(maj_121_n25), .ZN(maj_121_port_o) );
  XOR2_X1 maj_121_U2 ( .A(maj_121_n22), .B(maj_121_n21), .Z(maj_121_n23) );
  NAND2_X1 maj_122_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_122_n18) );
  NAND2_X1 maj_122_U14 ( .A1(maj_122_n21), .A2(maj_122_n22), .ZN(maj_122_n17)
         );
  NAND2_X1 maj_122_U13 ( .A1(maj_122_n18), .A2(maj_122_n17), .ZN(maj_122_n19)
         );
  NAND2_X1 maj_122_U12 ( .A1(u_0_1[2]), .A2(maj_122_n16), .ZN(maj_122_n14) );
  NAND2_X1 maj_122_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_122_n15) );
  NAND2_X1 maj_122_U10 ( .A1(maj_122_n15), .A2(maj_122_n14), .ZN(maj_122_n20)
         );
  XOR2_X1 maj_122_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_122_n22) );
  XOR2_X1 maj_122_U8 ( .A(u_0_1[2]), .B(maj_122_n16), .Z(maj_122_n21) );
  XOR2_X1 maj_122_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_122_n16) );
  OR2_X1 maj_122_U6 ( .A1(maj_122_n20), .A2(maj_122_n19), .ZN(maj_122_n24) );
  NAND2_X1 maj_122_U5 ( .A1(maj_122_n24), .A2(maj_122_n23), .ZN(maj_122_n25)
         );
  NAND2_X1 maj_122_U4 ( .A1(maj_122_n20), .A2(maj_122_n19), .ZN(maj_122_n26)
         );
  NAND2_X1 maj_122_U3 ( .A1(maj_122_n26), .A2(maj_122_n25), .ZN(maj_122_port_o) );
  XOR2_X1 maj_122_U2 ( .A(maj_122_n22), .B(maj_122_n21), .Z(maj_122_n23) );
  NAND2_X1 maj_123_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_123_n18) );
  NAND2_X1 maj_123_U14 ( .A1(maj_123_n21), .A2(maj_123_n22), .ZN(maj_123_n17)
         );
  NAND2_X1 maj_123_U13 ( .A1(maj_123_n18), .A2(maj_123_n17), .ZN(maj_123_n19)
         );
  NAND2_X1 maj_123_U12 ( .A1(v_0_1[2]), .A2(maj_123_n16), .ZN(maj_123_n14) );
  NAND2_X1 maj_123_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_123_n15) );
  NAND2_X1 maj_123_U10 ( .A1(maj_123_n15), .A2(maj_123_n14), .ZN(maj_123_n20)
         );
  XOR2_X1 maj_123_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_123_n22) );
  XOR2_X1 maj_123_U8 ( .A(v_0_1[2]), .B(maj_123_n16), .Z(maj_123_n21) );
  XOR2_X1 maj_123_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_123_n16) );
  OR2_X1 maj_123_U6 ( .A1(maj_123_n20), .A2(maj_123_n19), .ZN(maj_123_n24) );
  NAND2_X1 maj_123_U5 ( .A1(maj_123_n24), .A2(maj_123_n23), .ZN(maj_123_n25)
         );
  NAND2_X1 maj_123_U4 ( .A1(maj_123_n20), .A2(maj_123_n19), .ZN(maj_123_n26)
         );
  NAND2_X1 maj_123_U3 ( .A1(maj_123_n26), .A2(maj_123_n25), .ZN(maj_123_port_o) );
  XOR2_X1 maj_123_U2 ( .A(maj_123_n22), .B(maj_123_n21), .Z(maj_123_n23) );
  NAND2_X1 maj_124_U15 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_124_n18) );
  NAND2_X1 maj_124_U14 ( .A1(maj_124_n21), .A2(maj_124_n22), .ZN(maj_124_n17)
         );
  NAND2_X1 maj_124_U13 ( .A1(maj_124_n18), .A2(maj_124_n17), .ZN(maj_124_n19)
         );
  NAND2_X1 maj_124_U12 ( .A1(u_0_2[2]), .A2(maj_124_n16), .ZN(maj_124_n14) );
  NAND2_X1 maj_124_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_124_n15) );
  NAND2_X1 maj_124_U10 ( .A1(maj_124_n15), .A2(maj_124_n14), .ZN(maj_124_n20)
         );
  XOR2_X1 maj_124_U9 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_124_n22) );
  XOR2_X1 maj_124_U8 ( .A(u_0_2[2]), .B(maj_124_n16), .Z(maj_124_n21) );
  XOR2_X1 maj_124_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_124_n16) );
  OR2_X1 maj_124_U6 ( .A1(maj_124_n20), .A2(maj_124_n19), .ZN(maj_124_n24) );
  NAND2_X1 maj_124_U5 ( .A1(maj_124_n24), .A2(maj_124_n23), .ZN(maj_124_n25)
         );
  NAND2_X1 maj_124_U4 ( .A1(maj_124_n20), .A2(maj_124_n19), .ZN(maj_124_n26)
         );
  NAND2_X1 maj_124_U3 ( .A1(maj_124_n26), .A2(maj_124_n25), .ZN(maj_124_port_o) );
  XOR2_X1 maj_124_U2 ( .A(maj_124_n22), .B(maj_124_n21), .Z(maj_124_n23) );
  NAND2_X1 maj_125_U15 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_125_n18) );
  NAND2_X1 maj_125_U14 ( .A1(maj_125_n21), .A2(maj_125_n22), .ZN(maj_125_n17)
         );
  NAND2_X1 maj_125_U13 ( .A1(maj_125_n18), .A2(maj_125_n17), .ZN(maj_125_n19)
         );
  NAND2_X1 maj_125_U12 ( .A1(v_0_2[2]), .A2(maj_125_n16), .ZN(maj_125_n14) );
  NAND2_X1 maj_125_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_125_n15) );
  NAND2_X1 maj_125_U10 ( .A1(maj_125_n15), .A2(maj_125_n14), .ZN(maj_125_n20)
         );
  XOR2_X1 maj_125_U9 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_125_n22) );
  XOR2_X1 maj_125_U8 ( .A(v_0_2[2]), .B(maj_125_n16), .Z(maj_125_n21) );
  XOR2_X1 maj_125_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_125_n16) );
  OR2_X1 maj_125_U6 ( .A1(maj_125_n20), .A2(maj_125_n19), .ZN(maj_125_n24) );
  NAND2_X1 maj_125_U5 ( .A1(maj_125_n24), .A2(maj_125_n23), .ZN(maj_125_n25)
         );
  NAND2_X1 maj_125_U4 ( .A1(maj_125_n20), .A2(maj_125_n19), .ZN(maj_125_n26)
         );
  NAND2_X1 maj_125_U3 ( .A1(maj_125_n26), .A2(maj_125_n25), .ZN(maj_125_port_o) );
  XOR2_X1 maj_125_U2 ( .A(maj_125_n22), .B(maj_125_n21), .Z(maj_125_n23) );
  NAND2_X1 maj_126_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_126_n18) );
  NAND2_X1 maj_126_U14 ( .A1(maj_126_n21), .A2(maj_126_n22), .ZN(maj_126_n17)
         );
  NAND2_X1 maj_126_U13 ( .A1(maj_126_n18), .A2(maj_126_n17), .ZN(maj_126_n19)
         );
  NAND2_X1 maj_126_U12 ( .A1(u_1_0[2]), .A2(maj_126_n16), .ZN(maj_126_n14) );
  NAND2_X1 maj_126_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_126_n15) );
  NAND2_X1 maj_126_U10 ( .A1(maj_126_n15), .A2(maj_126_n14), .ZN(maj_126_n20)
         );
  XOR2_X1 maj_126_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_126_n22) );
  XOR2_X1 maj_126_U8 ( .A(u_1_0[2]), .B(maj_126_n16), .Z(maj_126_n21) );
  XOR2_X1 maj_126_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_126_n16) );
  OR2_X1 maj_126_U6 ( .A1(maj_126_n20), .A2(maj_126_n19), .ZN(maj_126_n24) );
  NAND2_X1 maj_126_U5 ( .A1(maj_126_n24), .A2(maj_126_n23), .ZN(maj_126_n25)
         );
  NAND2_X1 maj_126_U4 ( .A1(maj_126_n20), .A2(maj_126_n19), .ZN(maj_126_n26)
         );
  NAND2_X1 maj_126_U3 ( .A1(maj_126_n26), .A2(maj_126_n25), .ZN(maj_126_port_o) );
  XOR2_X1 maj_126_U2 ( .A(maj_126_n22), .B(maj_126_n21), .Z(maj_126_n23) );
  NAND2_X1 maj_127_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_127_n18) );
  NAND2_X1 maj_127_U14 ( .A1(maj_127_n21), .A2(maj_127_n22), .ZN(maj_127_n17)
         );
  NAND2_X1 maj_127_U13 ( .A1(maj_127_n18), .A2(maj_127_n17), .ZN(maj_127_n19)
         );
  NAND2_X1 maj_127_U12 ( .A1(v_1_0[2]), .A2(maj_127_n16), .ZN(maj_127_n14) );
  NAND2_X1 maj_127_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_127_n15) );
  NAND2_X1 maj_127_U10 ( .A1(maj_127_n15), .A2(maj_127_n14), .ZN(maj_127_n20)
         );
  XOR2_X1 maj_127_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_127_n22) );
  XOR2_X1 maj_127_U8 ( .A(v_1_0[2]), .B(maj_127_n16), .Z(maj_127_n21) );
  XOR2_X1 maj_127_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_127_n16) );
  OR2_X1 maj_127_U6 ( .A1(maj_127_n20), .A2(maj_127_n19), .ZN(maj_127_n24) );
  NAND2_X1 maj_127_U5 ( .A1(maj_127_n24), .A2(maj_127_n23), .ZN(maj_127_n25)
         );
  NAND2_X1 maj_127_U4 ( .A1(maj_127_n20), .A2(maj_127_n19), .ZN(maj_127_n26)
         );
  NAND2_X1 maj_127_U3 ( .A1(maj_127_n26), .A2(maj_127_n25), .ZN(maj_127_port_o) );
  XOR2_X1 maj_127_U2 ( .A(maj_127_n22), .B(maj_127_n21), .Z(maj_127_n23) );
  NAND2_X1 maj_128_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_128_n18) );
  NAND2_X1 maj_128_U14 ( .A1(maj_128_n21), .A2(maj_128_n22), .ZN(maj_128_n17)
         );
  NAND2_X1 maj_128_U13 ( .A1(maj_128_n18), .A2(maj_128_n17), .ZN(maj_128_n19)
         );
  NAND2_X1 maj_128_U12 ( .A1(u_1_1[2]), .A2(maj_128_n16), .ZN(maj_128_n14) );
  NAND2_X1 maj_128_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_128_n15) );
  NAND2_X1 maj_128_U10 ( .A1(maj_128_n15), .A2(maj_128_n14), .ZN(maj_128_n20)
         );
  XOR2_X1 maj_128_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_128_n22) );
  XOR2_X1 maj_128_U8 ( .A(u_1_1[2]), .B(maj_128_n16), .Z(maj_128_n21) );
  XOR2_X1 maj_128_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_128_n16) );
  OR2_X1 maj_128_U6 ( .A1(maj_128_n20), .A2(maj_128_n19), .ZN(maj_128_n24) );
  NAND2_X1 maj_128_U5 ( .A1(maj_128_n24), .A2(maj_128_n23), .ZN(maj_128_n25)
         );
  NAND2_X1 maj_128_U4 ( .A1(maj_128_n20), .A2(maj_128_n19), .ZN(maj_128_n26)
         );
  NAND2_X1 maj_128_U3 ( .A1(maj_128_n26), .A2(maj_128_n25), .ZN(maj_128_port_o) );
  XOR2_X1 maj_128_U2 ( .A(maj_128_n22), .B(maj_128_n21), .Z(maj_128_n23) );
  NAND2_X1 maj_129_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_129_n18) );
  NAND2_X1 maj_129_U14 ( .A1(maj_129_n21), .A2(maj_129_n22), .ZN(maj_129_n17)
         );
  NAND2_X1 maj_129_U13 ( .A1(maj_129_n18), .A2(maj_129_n17), .ZN(maj_129_n19)
         );
  NAND2_X1 maj_129_U12 ( .A1(v_1_1[2]), .A2(maj_129_n16), .ZN(maj_129_n14) );
  NAND2_X1 maj_129_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_129_n15) );
  NAND2_X1 maj_129_U10 ( .A1(maj_129_n15), .A2(maj_129_n14), .ZN(maj_129_n20)
         );
  XOR2_X1 maj_129_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_129_n22) );
  XOR2_X1 maj_129_U8 ( .A(v_1_1[2]), .B(maj_129_n16), .Z(maj_129_n21) );
  XOR2_X1 maj_129_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_129_n16) );
  OR2_X1 maj_129_U6 ( .A1(maj_129_n20), .A2(maj_129_n19), .ZN(maj_129_n24) );
  NAND2_X1 maj_129_U5 ( .A1(maj_129_n24), .A2(maj_129_n23), .ZN(maj_129_n25)
         );
  NAND2_X1 maj_129_U4 ( .A1(maj_129_n20), .A2(maj_129_n19), .ZN(maj_129_n26)
         );
  NAND2_X1 maj_129_U3 ( .A1(maj_129_n26), .A2(maj_129_n25), .ZN(maj_129_port_o) );
  XOR2_X1 maj_129_U2 ( .A(maj_129_n22), .B(maj_129_n21), .Z(maj_129_n23) );
  NAND2_X1 maj_130_U15 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_130_n18) );
  NAND2_X1 maj_130_U14 ( .A1(maj_130_n21), .A2(maj_130_n22), .ZN(maj_130_n17)
         );
  NAND2_X1 maj_130_U13 ( .A1(maj_130_n18), .A2(maj_130_n17), .ZN(maj_130_n19)
         );
  NAND2_X1 maj_130_U12 ( .A1(u_1_2[2]), .A2(maj_130_n16), .ZN(maj_130_n14) );
  NAND2_X1 maj_130_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_130_n15) );
  NAND2_X1 maj_130_U10 ( .A1(maj_130_n15), .A2(maj_130_n14), .ZN(maj_130_n20)
         );
  XOR2_X1 maj_130_U9 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_130_n22) );
  XOR2_X1 maj_130_U8 ( .A(u_1_2[2]), .B(maj_130_n16), .Z(maj_130_n21) );
  XOR2_X1 maj_130_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_130_n16) );
  OR2_X1 maj_130_U6 ( .A1(maj_130_n20), .A2(maj_130_n19), .ZN(maj_130_n24) );
  NAND2_X1 maj_130_U5 ( .A1(maj_130_n24), .A2(maj_130_n23), .ZN(maj_130_n25)
         );
  NAND2_X1 maj_130_U4 ( .A1(maj_130_n20), .A2(maj_130_n19), .ZN(maj_130_n26)
         );
  NAND2_X1 maj_130_U3 ( .A1(maj_130_n26), .A2(maj_130_n25), .ZN(maj_130_port_o) );
  XOR2_X1 maj_130_U2 ( .A(maj_130_n22), .B(maj_130_n21), .Z(maj_130_n23) );
  NAND2_X1 maj_131_U15 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_131_n18) );
  NAND2_X1 maj_131_U14 ( .A1(maj_131_n21), .A2(maj_131_n22), .ZN(maj_131_n17)
         );
  NAND2_X1 maj_131_U13 ( .A1(maj_131_n18), .A2(maj_131_n17), .ZN(maj_131_n19)
         );
  NAND2_X1 maj_131_U12 ( .A1(v_1_2[2]), .A2(maj_131_n16), .ZN(maj_131_n14) );
  NAND2_X1 maj_131_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_131_n15) );
  NAND2_X1 maj_131_U10 ( .A1(maj_131_n15), .A2(maj_131_n14), .ZN(maj_131_n20)
         );
  XOR2_X1 maj_131_U9 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_131_n22) );
  XOR2_X1 maj_131_U8 ( .A(v_1_2[2]), .B(maj_131_n16), .Z(maj_131_n21) );
  XOR2_X1 maj_131_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_131_n16) );
  OR2_X1 maj_131_U6 ( .A1(maj_131_n20), .A2(maj_131_n19), .ZN(maj_131_n24) );
  NAND2_X1 maj_131_U5 ( .A1(maj_131_n24), .A2(maj_131_n23), .ZN(maj_131_n25)
         );
  NAND2_X1 maj_131_U4 ( .A1(maj_131_n20), .A2(maj_131_n19), .ZN(maj_131_n26)
         );
  NAND2_X1 maj_131_U3 ( .A1(maj_131_n26), .A2(maj_131_n25), .ZN(maj_131_port_o) );
  XOR2_X1 maj_131_U2 ( .A(maj_131_n22), .B(maj_131_n21), .Z(maj_131_n23) );
  NAND2_X1 maj_132_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_132_n18) );
  NAND2_X1 maj_132_U14 ( .A1(maj_132_n21), .A2(maj_132_n22), .ZN(maj_132_n17)
         );
  NAND2_X1 maj_132_U13 ( .A1(maj_132_n18), .A2(maj_132_n17), .ZN(maj_132_n19)
         );
  NAND2_X1 maj_132_U12 ( .A1(u_2_0[2]), .A2(maj_132_n16), .ZN(maj_132_n14) );
  NAND2_X1 maj_132_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_132_n15) );
  NAND2_X1 maj_132_U10 ( .A1(maj_132_n15), .A2(maj_132_n14), .ZN(maj_132_n20)
         );
  XOR2_X1 maj_132_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_132_n22) );
  XOR2_X1 maj_132_U8 ( .A(u_2_0[2]), .B(maj_132_n16), .Z(maj_132_n21) );
  XOR2_X1 maj_132_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_132_n16) );
  OR2_X1 maj_132_U6 ( .A1(maj_132_n20), .A2(maj_132_n19), .ZN(maj_132_n24) );
  NAND2_X1 maj_132_U5 ( .A1(maj_132_n24), .A2(maj_132_n23), .ZN(maj_132_n25)
         );
  NAND2_X1 maj_132_U4 ( .A1(maj_132_n20), .A2(maj_132_n19), .ZN(maj_132_n26)
         );
  NAND2_X1 maj_132_U3 ( .A1(maj_132_n26), .A2(maj_132_n25), .ZN(maj_132_port_o) );
  XOR2_X1 maj_132_U2 ( .A(maj_132_n22), .B(maj_132_n21), .Z(maj_132_n23) );
  NAND2_X1 maj_133_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_133_n18) );
  NAND2_X1 maj_133_U14 ( .A1(maj_133_n21), .A2(maj_133_n22), .ZN(maj_133_n17)
         );
  NAND2_X1 maj_133_U13 ( .A1(maj_133_n18), .A2(maj_133_n17), .ZN(maj_133_n19)
         );
  NAND2_X1 maj_133_U12 ( .A1(v_2_0[2]), .A2(maj_133_n16), .ZN(maj_133_n14) );
  NAND2_X1 maj_133_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_133_n15) );
  NAND2_X1 maj_133_U10 ( .A1(maj_133_n15), .A2(maj_133_n14), .ZN(maj_133_n20)
         );
  XOR2_X1 maj_133_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_133_n22) );
  XOR2_X1 maj_133_U8 ( .A(v_2_0[2]), .B(maj_133_n16), .Z(maj_133_n21) );
  XOR2_X1 maj_133_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_133_n16) );
  OR2_X1 maj_133_U6 ( .A1(maj_133_n20), .A2(maj_133_n19), .ZN(maj_133_n24) );
  NAND2_X1 maj_133_U5 ( .A1(maj_133_n24), .A2(maj_133_n23), .ZN(maj_133_n25)
         );
  NAND2_X1 maj_133_U4 ( .A1(maj_133_n20), .A2(maj_133_n19), .ZN(maj_133_n26)
         );
  NAND2_X1 maj_133_U3 ( .A1(maj_133_n26), .A2(maj_133_n25), .ZN(maj_133_port_o) );
  XOR2_X1 maj_133_U2 ( .A(maj_133_n22), .B(maj_133_n21), .Z(maj_133_n23) );
  NAND2_X1 maj_134_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_134_n18) );
  NAND2_X1 maj_134_U14 ( .A1(maj_134_n21), .A2(maj_134_n22), .ZN(maj_134_n17)
         );
  NAND2_X1 maj_134_U13 ( .A1(maj_134_n18), .A2(maj_134_n17), .ZN(maj_134_n19)
         );
  NAND2_X1 maj_134_U12 ( .A1(u_2_1[2]), .A2(maj_134_n16), .ZN(maj_134_n14) );
  NAND2_X1 maj_134_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_134_n15) );
  NAND2_X1 maj_134_U10 ( .A1(maj_134_n15), .A2(maj_134_n14), .ZN(maj_134_n20)
         );
  XOR2_X1 maj_134_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_134_n22) );
  XOR2_X1 maj_134_U8 ( .A(u_2_1[2]), .B(maj_134_n16), .Z(maj_134_n21) );
  XOR2_X1 maj_134_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_134_n16) );
  OR2_X1 maj_134_U6 ( .A1(maj_134_n20), .A2(maj_134_n19), .ZN(maj_134_n24) );
  NAND2_X1 maj_134_U5 ( .A1(maj_134_n24), .A2(maj_134_n23), .ZN(maj_134_n25)
         );
  NAND2_X1 maj_134_U4 ( .A1(maj_134_n20), .A2(maj_134_n19), .ZN(maj_134_n26)
         );
  NAND2_X1 maj_134_U3 ( .A1(maj_134_n26), .A2(maj_134_n25), .ZN(maj_134_port_o) );
  XOR2_X1 maj_134_U2 ( .A(maj_134_n22), .B(maj_134_n21), .Z(maj_134_n23) );
  NAND2_X1 maj_135_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_135_n18) );
  NAND2_X1 maj_135_U14 ( .A1(maj_135_n21), .A2(maj_135_n22), .ZN(maj_135_n17)
         );
  NAND2_X1 maj_135_U13 ( .A1(maj_135_n18), .A2(maj_135_n17), .ZN(maj_135_n19)
         );
  NAND2_X1 maj_135_U12 ( .A1(v_2_1[2]), .A2(maj_135_n16), .ZN(maj_135_n14) );
  NAND2_X1 maj_135_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_135_n15) );
  NAND2_X1 maj_135_U10 ( .A1(maj_135_n15), .A2(maj_135_n14), .ZN(maj_135_n20)
         );
  XOR2_X1 maj_135_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_135_n22) );
  XOR2_X1 maj_135_U8 ( .A(v_2_1[2]), .B(maj_135_n16), .Z(maj_135_n21) );
  XOR2_X1 maj_135_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_135_n16) );
  OR2_X1 maj_135_U6 ( .A1(maj_135_n20), .A2(maj_135_n19), .ZN(maj_135_n24) );
  NAND2_X1 maj_135_U5 ( .A1(maj_135_n24), .A2(maj_135_n23), .ZN(maj_135_n25)
         );
  NAND2_X1 maj_135_U4 ( .A1(maj_135_n20), .A2(maj_135_n19), .ZN(maj_135_n26)
         );
  NAND2_X1 maj_135_U3 ( .A1(maj_135_n26), .A2(maj_135_n25), .ZN(maj_135_port_o) );
  XOR2_X1 maj_135_U2 ( .A(maj_135_n22), .B(maj_135_n21), .Z(maj_135_n23) );
  NAND2_X1 maj_136_U15 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_136_n18) );
  NAND2_X1 maj_136_U14 ( .A1(maj_136_n21), .A2(maj_136_n22), .ZN(maj_136_n17)
         );
  NAND2_X1 maj_136_U13 ( .A1(maj_136_n18), .A2(maj_136_n17), .ZN(maj_136_n19)
         );
  NAND2_X1 maj_136_U12 ( .A1(u_2_2[2]), .A2(maj_136_n16), .ZN(maj_136_n14) );
  NAND2_X1 maj_136_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_136_n15) );
  NAND2_X1 maj_136_U10 ( .A1(maj_136_n15), .A2(maj_136_n14), .ZN(maj_136_n20)
         );
  XOR2_X1 maj_136_U9 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_136_n22) );
  XOR2_X1 maj_136_U8 ( .A(u_2_2[2]), .B(maj_136_n16), .Z(maj_136_n21) );
  XOR2_X1 maj_136_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_136_n16) );
  OR2_X1 maj_136_U6 ( .A1(maj_136_n20), .A2(maj_136_n19), .ZN(maj_136_n24) );
  NAND2_X1 maj_136_U5 ( .A1(maj_136_n24), .A2(maj_136_n23), .ZN(maj_136_n25)
         );
  NAND2_X1 maj_136_U4 ( .A1(maj_136_n20), .A2(maj_136_n19), .ZN(maj_136_n26)
         );
  NAND2_X1 maj_136_U3 ( .A1(maj_136_n26), .A2(maj_136_n25), .ZN(maj_136_port_o) );
  XOR2_X1 maj_136_U2 ( .A(maj_136_n22), .B(maj_136_n21), .Z(maj_136_n23) );
  NAND2_X1 maj_137_U15 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_137_n18) );
  NAND2_X1 maj_137_U14 ( .A1(maj_137_n21), .A2(maj_137_n22), .ZN(maj_137_n17)
         );
  NAND2_X1 maj_137_U13 ( .A1(maj_137_n18), .A2(maj_137_n17), .ZN(maj_137_n19)
         );
  NAND2_X1 maj_137_U12 ( .A1(v_2_2[2]), .A2(maj_137_n16), .ZN(maj_137_n14) );
  NAND2_X1 maj_137_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_137_n15) );
  NAND2_X1 maj_137_U10 ( .A1(maj_137_n15), .A2(maj_137_n14), .ZN(maj_137_n20)
         );
  XOR2_X1 maj_137_U9 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_137_n22) );
  XOR2_X1 maj_137_U8 ( .A(v_2_2[2]), .B(maj_137_n16), .Z(maj_137_n21) );
  XOR2_X1 maj_137_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_137_n16) );
  OR2_X1 maj_137_U6 ( .A1(maj_137_n20), .A2(maj_137_n19), .ZN(maj_137_n24) );
  NAND2_X1 maj_137_U5 ( .A1(maj_137_n24), .A2(maj_137_n23), .ZN(maj_137_n25)
         );
  NAND2_X1 maj_137_U4 ( .A1(maj_137_n20), .A2(maj_137_n19), .ZN(maj_137_n26)
         );
  NAND2_X1 maj_137_U3 ( .A1(maj_137_n26), .A2(maj_137_n25), .ZN(maj_137_port_o) );
  XOR2_X1 maj_137_U2 ( .A(maj_137_n22), .B(maj_137_n21), .Z(maj_137_n23) );
  NAND2_X1 maj_138_U15 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_138_n18) );
  NAND2_X1 maj_138_U14 ( .A1(maj_138_n21), .A2(maj_138_n22), .ZN(maj_138_n17)
         );
  NAND2_X1 maj_138_U13 ( .A1(maj_138_n18), .A2(maj_138_n17), .ZN(maj_138_n19)
         );
  NAND2_X1 maj_138_U12 ( .A1(u_3_0[2]), .A2(maj_138_n16), .ZN(maj_138_n14) );
  NAND2_X1 maj_138_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_138_n15) );
  NAND2_X1 maj_138_U10 ( .A1(maj_138_n15), .A2(maj_138_n14), .ZN(maj_138_n20)
         );
  XOR2_X1 maj_138_U9 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_138_n22) );
  XOR2_X1 maj_138_U8 ( .A(u_3_0[2]), .B(maj_138_n16), .Z(maj_138_n21) );
  XOR2_X1 maj_138_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_138_n16) );
  OR2_X1 maj_138_U6 ( .A1(maj_138_n20), .A2(maj_138_n19), .ZN(maj_138_n24) );
  NAND2_X1 maj_138_U5 ( .A1(maj_138_n24), .A2(maj_138_n23), .ZN(maj_138_n25)
         );
  NAND2_X1 maj_138_U4 ( .A1(maj_138_n20), .A2(maj_138_n19), .ZN(maj_138_n26)
         );
  NAND2_X1 maj_138_U3 ( .A1(maj_138_n26), .A2(maj_138_n25), .ZN(maj_138_port_o) );
  XOR2_X1 maj_138_U2 ( .A(maj_138_n22), .B(maj_138_n21), .Z(maj_138_n23) );
  NAND2_X1 maj_139_U15 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_139_n18) );
  NAND2_X1 maj_139_U14 ( .A1(maj_139_n21), .A2(maj_139_n22), .ZN(maj_139_n17)
         );
  NAND2_X1 maj_139_U13 ( .A1(maj_139_n18), .A2(maj_139_n17), .ZN(maj_139_n19)
         );
  NAND2_X1 maj_139_U12 ( .A1(v_3_0[2]), .A2(maj_139_n16), .ZN(maj_139_n14) );
  NAND2_X1 maj_139_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_139_n15) );
  NAND2_X1 maj_139_U10 ( .A1(maj_139_n15), .A2(maj_139_n14), .ZN(maj_139_n20)
         );
  XOR2_X1 maj_139_U9 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_139_n22) );
  XOR2_X1 maj_139_U8 ( .A(v_3_0[2]), .B(maj_139_n16), .Z(maj_139_n21) );
  XOR2_X1 maj_139_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_139_n16) );
  OR2_X1 maj_139_U6 ( .A1(maj_139_n20), .A2(maj_139_n19), .ZN(maj_139_n24) );
  NAND2_X1 maj_139_U5 ( .A1(maj_139_n24), .A2(maj_139_n23), .ZN(maj_139_n25)
         );
  NAND2_X1 maj_139_U4 ( .A1(maj_139_n20), .A2(maj_139_n19), .ZN(maj_139_n26)
         );
  NAND2_X1 maj_139_U3 ( .A1(maj_139_n26), .A2(maj_139_n25), .ZN(maj_139_port_o) );
  XOR2_X1 maj_139_U2 ( .A(maj_139_n22), .B(maj_139_n21), .Z(maj_139_n23) );
  NAND2_X1 maj_140_U15 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_140_n18) );
  NAND2_X1 maj_140_U14 ( .A1(maj_140_n21), .A2(maj_140_n22), .ZN(maj_140_n17)
         );
  NAND2_X1 maj_140_U13 ( .A1(maj_140_n18), .A2(maj_140_n17), .ZN(maj_140_n19)
         );
  NAND2_X1 maj_140_U12 ( .A1(u_3_1[2]), .A2(maj_140_n16), .ZN(maj_140_n14) );
  NAND2_X1 maj_140_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_140_n15) );
  NAND2_X1 maj_140_U10 ( .A1(maj_140_n15), .A2(maj_140_n14), .ZN(maj_140_n20)
         );
  XOR2_X1 maj_140_U9 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_140_n22) );
  XOR2_X1 maj_140_U8 ( .A(u_3_1[2]), .B(maj_140_n16), .Z(maj_140_n21) );
  XOR2_X1 maj_140_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_140_n16) );
  OR2_X1 maj_140_U6 ( .A1(maj_140_n20), .A2(maj_140_n19), .ZN(maj_140_n24) );
  NAND2_X1 maj_140_U5 ( .A1(maj_140_n24), .A2(maj_140_n23), .ZN(maj_140_n25)
         );
  NAND2_X1 maj_140_U4 ( .A1(maj_140_n20), .A2(maj_140_n19), .ZN(maj_140_n26)
         );
  NAND2_X1 maj_140_U3 ( .A1(maj_140_n26), .A2(maj_140_n25), .ZN(maj_140_port_o) );
  XOR2_X1 maj_140_U2 ( .A(maj_140_n22), .B(maj_140_n21), .Z(maj_140_n23) );
  NAND2_X1 maj_141_U15 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_141_n18) );
  NAND2_X1 maj_141_U14 ( .A1(maj_141_n21), .A2(maj_141_n22), .ZN(maj_141_n17)
         );
  NAND2_X1 maj_141_U13 ( .A1(maj_141_n18), .A2(maj_141_n17), .ZN(maj_141_n19)
         );
  NAND2_X1 maj_141_U12 ( .A1(v_3_1[2]), .A2(maj_141_n16), .ZN(maj_141_n14) );
  NAND2_X1 maj_141_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_141_n15) );
  NAND2_X1 maj_141_U10 ( .A1(maj_141_n15), .A2(maj_141_n14), .ZN(maj_141_n20)
         );
  XOR2_X1 maj_141_U9 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_141_n22) );
  XOR2_X1 maj_141_U8 ( .A(v_3_1[2]), .B(maj_141_n16), .Z(maj_141_n21) );
  XOR2_X1 maj_141_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_141_n16) );
  OR2_X1 maj_141_U6 ( .A1(maj_141_n20), .A2(maj_141_n19), .ZN(maj_141_n24) );
  NAND2_X1 maj_141_U5 ( .A1(maj_141_n24), .A2(maj_141_n23), .ZN(maj_141_n25)
         );
  NAND2_X1 maj_141_U4 ( .A1(maj_141_n20), .A2(maj_141_n19), .ZN(maj_141_n26)
         );
  NAND2_X1 maj_141_U3 ( .A1(maj_141_n26), .A2(maj_141_n25), .ZN(maj_141_port_o) );
  XOR2_X1 maj_141_U2 ( .A(maj_141_n22), .B(maj_141_n21), .Z(maj_141_n23) );
  NAND2_X1 maj_142_U15 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_142_n18) );
  NAND2_X1 maj_142_U14 ( .A1(maj_142_n21), .A2(maj_142_n22), .ZN(maj_142_n17)
         );
  NAND2_X1 maj_142_U13 ( .A1(maj_142_n18), .A2(maj_142_n17), .ZN(maj_142_n19)
         );
  NAND2_X1 maj_142_U12 ( .A1(u_3_2[2]), .A2(maj_142_n16), .ZN(maj_142_n14) );
  NAND2_X1 maj_142_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_142_n15) );
  NAND2_X1 maj_142_U10 ( .A1(maj_142_n15), .A2(maj_142_n14), .ZN(maj_142_n20)
         );
  XOR2_X1 maj_142_U9 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_142_n22) );
  XOR2_X1 maj_142_U8 ( .A(u_3_2[2]), .B(maj_142_n16), .Z(maj_142_n21) );
  XOR2_X1 maj_142_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_142_n16) );
  OR2_X1 maj_142_U6 ( .A1(maj_142_n20), .A2(maj_142_n19), .ZN(maj_142_n24) );
  NAND2_X1 maj_142_U5 ( .A1(maj_142_n24), .A2(maj_142_n23), .ZN(maj_142_n25)
         );
  NAND2_X1 maj_142_U4 ( .A1(maj_142_n20), .A2(maj_142_n19), .ZN(maj_142_n26)
         );
  NAND2_X1 maj_142_U3 ( .A1(maj_142_n26), .A2(maj_142_n25), .ZN(maj_142_port_o) );
  XOR2_X1 maj_142_U2 ( .A(maj_142_n22), .B(maj_142_n21), .Z(maj_142_n23) );
  NAND2_X1 maj_143_U15 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_143_n18) );
  NAND2_X1 maj_143_U14 ( .A1(maj_143_n21), .A2(maj_143_n22), .ZN(maj_143_n17)
         );
  NAND2_X1 maj_143_U13 ( .A1(maj_143_n18), .A2(maj_143_n17), .ZN(maj_143_n19)
         );
  NAND2_X1 maj_143_U12 ( .A1(v_3_2[2]), .A2(maj_143_n16), .ZN(maj_143_n14) );
  NAND2_X1 maj_143_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_143_n15) );
  NAND2_X1 maj_143_U10 ( .A1(maj_143_n15), .A2(maj_143_n14), .ZN(maj_143_n20)
         );
  XOR2_X1 maj_143_U9 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_143_n22) );
  XOR2_X1 maj_143_U8 ( .A(v_3_2[2]), .B(maj_143_n16), .Z(maj_143_n21) );
  XOR2_X1 maj_143_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_143_n16) );
  OR2_X1 maj_143_U6 ( .A1(maj_143_n20), .A2(maj_143_n19), .ZN(maj_143_n24) );
  NAND2_X1 maj_143_U5 ( .A1(maj_143_n24), .A2(maj_143_n23), .ZN(maj_143_n25)
         );
  NAND2_X1 maj_143_U4 ( .A1(maj_143_n20), .A2(maj_143_n19), .ZN(maj_143_n26)
         );
  NAND2_X1 maj_143_U3 ( .A1(maj_143_n26), .A2(maj_143_n25), .ZN(maj_143_port_o) );
  XOR2_X1 maj_143_U2 ( .A(maj_143_n22), .B(maj_143_n21), .Z(maj_143_n23) );
  NAND2_X1 maj_144_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_144_n18) );
  NAND2_X1 maj_144_U14 ( .A1(maj_144_n21), .A2(maj_144_n22), .ZN(maj_144_n17)
         );
  NAND2_X1 maj_144_U13 ( .A1(maj_144_n18), .A2(maj_144_n17), .ZN(maj_144_n19)
         );
  NAND2_X1 maj_144_U12 ( .A1(u_0_0[2]), .A2(maj_144_n16), .ZN(maj_144_n14) );
  NAND2_X1 maj_144_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_144_n15) );
  NAND2_X1 maj_144_U10 ( .A1(maj_144_n15), .A2(maj_144_n14), .ZN(maj_144_n20)
         );
  XOR2_X1 maj_144_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_144_n22) );
  XOR2_X1 maj_144_U8 ( .A(u_0_0[2]), .B(maj_144_n16), .Z(maj_144_n21) );
  XOR2_X1 maj_144_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_144_n16) );
  OR2_X1 maj_144_U6 ( .A1(maj_144_n20), .A2(maj_144_n19), .ZN(maj_144_n24) );
  NAND2_X1 maj_144_U5 ( .A1(maj_144_n24), .A2(maj_144_n23), .ZN(maj_144_n25)
         );
  NAND2_X1 maj_144_U4 ( .A1(maj_144_n20), .A2(maj_144_n19), .ZN(maj_144_n26)
         );
  NAND2_X1 maj_144_U3 ( .A1(maj_144_n26), .A2(maj_144_n25), .ZN(maj_144_port_o) );
  XOR2_X1 maj_144_U2 ( .A(maj_144_n22), .B(maj_144_n21), .Z(maj_144_n23) );
  NAND2_X1 maj_145_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_145_n18) );
  NAND2_X1 maj_145_U14 ( .A1(maj_145_n21), .A2(maj_145_n22), .ZN(maj_145_n17)
         );
  NAND2_X1 maj_145_U13 ( .A1(maj_145_n18), .A2(maj_145_n17), .ZN(maj_145_n19)
         );
  NAND2_X1 maj_145_U12 ( .A1(v_0_0[2]), .A2(maj_145_n16), .ZN(maj_145_n14) );
  NAND2_X1 maj_145_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_145_n15) );
  NAND2_X1 maj_145_U10 ( .A1(maj_145_n15), .A2(maj_145_n14), .ZN(maj_145_n20)
         );
  XOR2_X1 maj_145_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_145_n22) );
  XOR2_X1 maj_145_U8 ( .A(v_0_0[2]), .B(maj_145_n16), .Z(maj_145_n21) );
  XOR2_X1 maj_145_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_145_n16) );
  OR2_X1 maj_145_U6 ( .A1(maj_145_n20), .A2(maj_145_n19), .ZN(maj_145_n24) );
  NAND2_X1 maj_145_U5 ( .A1(maj_145_n24), .A2(maj_145_n23), .ZN(maj_145_n25)
         );
  NAND2_X1 maj_145_U4 ( .A1(maj_145_n20), .A2(maj_145_n19), .ZN(maj_145_n26)
         );
  NAND2_X1 maj_145_U3 ( .A1(maj_145_n26), .A2(maj_145_n25), .ZN(maj_145_port_o) );
  XOR2_X1 maj_145_U2 ( .A(maj_145_n22), .B(maj_145_n21), .Z(maj_145_n23) );
  NAND2_X1 maj_146_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_146_n18) );
  NAND2_X1 maj_146_U14 ( .A1(maj_146_n21), .A2(maj_146_n22), .ZN(maj_146_n17)
         );
  NAND2_X1 maj_146_U13 ( .A1(maj_146_n18), .A2(maj_146_n17), .ZN(maj_146_n19)
         );
  NAND2_X1 maj_146_U12 ( .A1(u_0_1[2]), .A2(maj_146_n16), .ZN(maj_146_n14) );
  NAND2_X1 maj_146_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_146_n15) );
  NAND2_X1 maj_146_U10 ( .A1(maj_146_n15), .A2(maj_146_n14), .ZN(maj_146_n20)
         );
  XOR2_X1 maj_146_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_146_n22) );
  XOR2_X1 maj_146_U8 ( .A(u_0_1[2]), .B(maj_146_n16), .Z(maj_146_n21) );
  XOR2_X1 maj_146_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_146_n16) );
  OR2_X1 maj_146_U6 ( .A1(maj_146_n20), .A2(maj_146_n19), .ZN(maj_146_n24) );
  NAND2_X1 maj_146_U5 ( .A1(maj_146_n24), .A2(maj_146_n23), .ZN(maj_146_n25)
         );
  NAND2_X1 maj_146_U4 ( .A1(maj_146_n20), .A2(maj_146_n19), .ZN(maj_146_n26)
         );
  NAND2_X1 maj_146_U3 ( .A1(maj_146_n26), .A2(maj_146_n25), .ZN(maj_146_port_o) );
  XOR2_X1 maj_146_U2 ( .A(maj_146_n22), .B(maj_146_n21), .Z(maj_146_n23) );
  NAND2_X1 maj_147_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_147_n18) );
  NAND2_X1 maj_147_U14 ( .A1(maj_147_n21), .A2(maj_147_n22), .ZN(maj_147_n17)
         );
  NAND2_X1 maj_147_U13 ( .A1(maj_147_n18), .A2(maj_147_n17), .ZN(maj_147_n19)
         );
  NAND2_X1 maj_147_U12 ( .A1(v_0_1[2]), .A2(maj_147_n16), .ZN(maj_147_n14) );
  NAND2_X1 maj_147_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_147_n15) );
  NAND2_X1 maj_147_U10 ( .A1(maj_147_n15), .A2(maj_147_n14), .ZN(maj_147_n20)
         );
  XOR2_X1 maj_147_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_147_n22) );
  XOR2_X1 maj_147_U8 ( .A(v_0_1[2]), .B(maj_147_n16), .Z(maj_147_n21) );
  XOR2_X1 maj_147_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_147_n16) );
  OR2_X1 maj_147_U6 ( .A1(maj_147_n20), .A2(maj_147_n19), .ZN(maj_147_n24) );
  NAND2_X1 maj_147_U5 ( .A1(maj_147_n24), .A2(maj_147_n23), .ZN(maj_147_n25)
         );
  NAND2_X1 maj_147_U4 ( .A1(maj_147_n20), .A2(maj_147_n19), .ZN(maj_147_n26)
         );
  NAND2_X1 maj_147_U3 ( .A1(maj_147_n26), .A2(maj_147_n25), .ZN(maj_147_port_o) );
  XOR2_X1 maj_147_U2 ( .A(maj_147_n22), .B(maj_147_n21), .Z(maj_147_n23) );
  NAND2_X1 maj_148_U15 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_148_n18) );
  NAND2_X1 maj_148_U14 ( .A1(maj_148_n21), .A2(maj_148_n22), .ZN(maj_148_n17)
         );
  NAND2_X1 maj_148_U13 ( .A1(maj_148_n18), .A2(maj_148_n17), .ZN(maj_148_n19)
         );
  NAND2_X1 maj_148_U12 ( .A1(u_0_2[2]), .A2(maj_148_n16), .ZN(maj_148_n14) );
  NAND2_X1 maj_148_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_148_n15) );
  NAND2_X1 maj_148_U10 ( .A1(maj_148_n15), .A2(maj_148_n14), .ZN(maj_148_n20)
         );
  XOR2_X1 maj_148_U9 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_148_n22) );
  XOR2_X1 maj_148_U8 ( .A(u_0_2[2]), .B(maj_148_n16), .Z(maj_148_n21) );
  XOR2_X1 maj_148_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_148_n16) );
  OR2_X1 maj_148_U6 ( .A1(maj_148_n20), .A2(maj_148_n19), .ZN(maj_148_n24) );
  NAND2_X1 maj_148_U5 ( .A1(maj_148_n24), .A2(maj_148_n23), .ZN(maj_148_n25)
         );
  NAND2_X1 maj_148_U4 ( .A1(maj_148_n20), .A2(maj_148_n19), .ZN(maj_148_n26)
         );
  NAND2_X1 maj_148_U3 ( .A1(maj_148_n26), .A2(maj_148_n25), .ZN(maj_148_port_o) );
  XOR2_X1 maj_148_U2 ( .A(maj_148_n22), .B(maj_148_n21), .Z(maj_148_n23) );
  NAND2_X1 maj_149_U15 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_149_n18) );
  NAND2_X1 maj_149_U14 ( .A1(maj_149_n21), .A2(maj_149_n22), .ZN(maj_149_n17)
         );
  NAND2_X1 maj_149_U13 ( .A1(maj_149_n18), .A2(maj_149_n17), .ZN(maj_149_n19)
         );
  NAND2_X1 maj_149_U12 ( .A1(v_0_2[2]), .A2(maj_149_n16), .ZN(maj_149_n14) );
  NAND2_X1 maj_149_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_149_n15) );
  NAND2_X1 maj_149_U10 ( .A1(maj_149_n15), .A2(maj_149_n14), .ZN(maj_149_n20)
         );
  XOR2_X1 maj_149_U9 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_149_n22) );
  XOR2_X1 maj_149_U8 ( .A(v_0_2[2]), .B(maj_149_n16), .Z(maj_149_n21) );
  XOR2_X1 maj_149_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_149_n16) );
  OR2_X1 maj_149_U6 ( .A1(maj_149_n20), .A2(maj_149_n19), .ZN(maj_149_n24) );
  NAND2_X1 maj_149_U5 ( .A1(maj_149_n24), .A2(maj_149_n23), .ZN(maj_149_n25)
         );
  NAND2_X1 maj_149_U4 ( .A1(maj_149_n20), .A2(maj_149_n19), .ZN(maj_149_n26)
         );
  NAND2_X1 maj_149_U3 ( .A1(maj_149_n26), .A2(maj_149_n25), .ZN(maj_149_port_o) );
  XOR2_X1 maj_149_U2 ( .A(maj_149_n22), .B(maj_149_n21), .Z(maj_149_n23) );
  NAND2_X1 maj_150_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_150_n18) );
  NAND2_X1 maj_150_U14 ( .A1(maj_150_n21), .A2(maj_150_n22), .ZN(maj_150_n17)
         );
  NAND2_X1 maj_150_U13 ( .A1(maj_150_n18), .A2(maj_150_n17), .ZN(maj_150_n19)
         );
  NAND2_X1 maj_150_U12 ( .A1(u_1_0[2]), .A2(maj_150_n16), .ZN(maj_150_n14) );
  NAND2_X1 maj_150_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_150_n15) );
  NAND2_X1 maj_150_U10 ( .A1(maj_150_n15), .A2(maj_150_n14), .ZN(maj_150_n20)
         );
  XOR2_X1 maj_150_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_150_n22) );
  XOR2_X1 maj_150_U8 ( .A(u_1_0[2]), .B(maj_150_n16), .Z(maj_150_n21) );
  XOR2_X1 maj_150_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_150_n16) );
  OR2_X1 maj_150_U6 ( .A1(maj_150_n20), .A2(maj_150_n19), .ZN(maj_150_n24) );
  NAND2_X1 maj_150_U5 ( .A1(maj_150_n24), .A2(maj_150_n23), .ZN(maj_150_n25)
         );
  NAND2_X1 maj_150_U4 ( .A1(maj_150_n20), .A2(maj_150_n19), .ZN(maj_150_n26)
         );
  NAND2_X1 maj_150_U3 ( .A1(maj_150_n26), .A2(maj_150_n25), .ZN(maj_150_port_o) );
  XOR2_X1 maj_150_U2 ( .A(maj_150_n22), .B(maj_150_n21), .Z(maj_150_n23) );
  NAND2_X1 maj_151_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_151_n18) );
  NAND2_X1 maj_151_U14 ( .A1(maj_151_n21), .A2(maj_151_n22), .ZN(maj_151_n17)
         );
  NAND2_X1 maj_151_U13 ( .A1(maj_151_n18), .A2(maj_151_n17), .ZN(maj_151_n19)
         );
  NAND2_X1 maj_151_U12 ( .A1(v_1_0[2]), .A2(maj_151_n16), .ZN(maj_151_n14) );
  NAND2_X1 maj_151_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_151_n15) );
  NAND2_X1 maj_151_U10 ( .A1(maj_151_n15), .A2(maj_151_n14), .ZN(maj_151_n20)
         );
  XOR2_X1 maj_151_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_151_n22) );
  XOR2_X1 maj_151_U8 ( .A(v_1_0[2]), .B(maj_151_n16), .Z(maj_151_n21) );
  XOR2_X1 maj_151_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_151_n16) );
  OR2_X1 maj_151_U6 ( .A1(maj_151_n20), .A2(maj_151_n19), .ZN(maj_151_n24) );
  NAND2_X1 maj_151_U5 ( .A1(maj_151_n24), .A2(maj_151_n23), .ZN(maj_151_n25)
         );
  NAND2_X1 maj_151_U4 ( .A1(maj_151_n20), .A2(maj_151_n19), .ZN(maj_151_n26)
         );
  NAND2_X1 maj_151_U3 ( .A1(maj_151_n26), .A2(maj_151_n25), .ZN(maj_151_port_o) );
  XOR2_X1 maj_151_U2 ( .A(maj_151_n22), .B(maj_151_n21), .Z(maj_151_n23) );
  NAND2_X1 maj_152_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_152_n18) );
  NAND2_X1 maj_152_U14 ( .A1(maj_152_n21), .A2(maj_152_n22), .ZN(maj_152_n17)
         );
  NAND2_X1 maj_152_U13 ( .A1(maj_152_n18), .A2(maj_152_n17), .ZN(maj_152_n19)
         );
  NAND2_X1 maj_152_U12 ( .A1(u_1_1[2]), .A2(maj_152_n16), .ZN(maj_152_n14) );
  NAND2_X1 maj_152_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_152_n15) );
  NAND2_X1 maj_152_U10 ( .A1(maj_152_n15), .A2(maj_152_n14), .ZN(maj_152_n20)
         );
  XOR2_X1 maj_152_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_152_n22) );
  XOR2_X1 maj_152_U8 ( .A(u_1_1[2]), .B(maj_152_n16), .Z(maj_152_n21) );
  XOR2_X1 maj_152_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_152_n16) );
  OR2_X1 maj_152_U6 ( .A1(maj_152_n20), .A2(maj_152_n19), .ZN(maj_152_n24) );
  NAND2_X1 maj_152_U5 ( .A1(maj_152_n24), .A2(maj_152_n23), .ZN(maj_152_n25)
         );
  NAND2_X1 maj_152_U4 ( .A1(maj_152_n20), .A2(maj_152_n19), .ZN(maj_152_n26)
         );
  NAND2_X1 maj_152_U3 ( .A1(maj_152_n26), .A2(maj_152_n25), .ZN(maj_152_port_o) );
  XOR2_X1 maj_152_U2 ( .A(maj_152_n22), .B(maj_152_n21), .Z(maj_152_n23) );
  NAND2_X1 maj_153_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_153_n18) );
  NAND2_X1 maj_153_U14 ( .A1(maj_153_n21), .A2(maj_153_n22), .ZN(maj_153_n17)
         );
  NAND2_X1 maj_153_U13 ( .A1(maj_153_n18), .A2(maj_153_n17), .ZN(maj_153_n19)
         );
  NAND2_X1 maj_153_U12 ( .A1(v_1_1[2]), .A2(maj_153_n16), .ZN(maj_153_n14) );
  NAND2_X1 maj_153_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_153_n15) );
  NAND2_X1 maj_153_U10 ( .A1(maj_153_n15), .A2(maj_153_n14), .ZN(maj_153_n20)
         );
  XOR2_X1 maj_153_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_153_n22) );
  XOR2_X1 maj_153_U8 ( .A(v_1_1[2]), .B(maj_153_n16), .Z(maj_153_n21) );
  XOR2_X1 maj_153_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_153_n16) );
  OR2_X1 maj_153_U6 ( .A1(maj_153_n20), .A2(maj_153_n19), .ZN(maj_153_n24) );
  NAND2_X1 maj_153_U5 ( .A1(maj_153_n24), .A2(maj_153_n23), .ZN(maj_153_n25)
         );
  NAND2_X1 maj_153_U4 ( .A1(maj_153_n20), .A2(maj_153_n19), .ZN(maj_153_n26)
         );
  NAND2_X1 maj_153_U3 ( .A1(maj_153_n26), .A2(maj_153_n25), .ZN(maj_153_port_o) );
  XOR2_X1 maj_153_U2 ( .A(maj_153_n22), .B(maj_153_n21), .Z(maj_153_n23) );
  NAND2_X1 maj_154_U15 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_154_n18) );
  NAND2_X1 maj_154_U14 ( .A1(maj_154_n21), .A2(maj_154_n22), .ZN(maj_154_n17)
         );
  NAND2_X1 maj_154_U13 ( .A1(maj_154_n18), .A2(maj_154_n17), .ZN(maj_154_n19)
         );
  NAND2_X1 maj_154_U12 ( .A1(u_1_2[2]), .A2(maj_154_n16), .ZN(maj_154_n14) );
  NAND2_X1 maj_154_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_154_n15) );
  NAND2_X1 maj_154_U10 ( .A1(maj_154_n15), .A2(maj_154_n14), .ZN(maj_154_n20)
         );
  XOR2_X1 maj_154_U9 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_154_n22) );
  XOR2_X1 maj_154_U8 ( .A(u_1_2[2]), .B(maj_154_n16), .Z(maj_154_n21) );
  XOR2_X1 maj_154_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_154_n16) );
  OR2_X1 maj_154_U6 ( .A1(maj_154_n20), .A2(maj_154_n19), .ZN(maj_154_n24) );
  NAND2_X1 maj_154_U5 ( .A1(maj_154_n24), .A2(maj_154_n23), .ZN(maj_154_n25)
         );
  NAND2_X1 maj_154_U4 ( .A1(maj_154_n20), .A2(maj_154_n19), .ZN(maj_154_n26)
         );
  NAND2_X1 maj_154_U3 ( .A1(maj_154_n26), .A2(maj_154_n25), .ZN(maj_154_port_o) );
  XOR2_X1 maj_154_U2 ( .A(maj_154_n22), .B(maj_154_n21), .Z(maj_154_n23) );
  NAND2_X1 maj_155_U15 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_155_n18) );
  NAND2_X1 maj_155_U14 ( .A1(maj_155_n21), .A2(maj_155_n22), .ZN(maj_155_n17)
         );
  NAND2_X1 maj_155_U13 ( .A1(maj_155_n18), .A2(maj_155_n17), .ZN(maj_155_n19)
         );
  NAND2_X1 maj_155_U12 ( .A1(v_1_2[2]), .A2(maj_155_n16), .ZN(maj_155_n14) );
  NAND2_X1 maj_155_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_155_n15) );
  NAND2_X1 maj_155_U10 ( .A1(maj_155_n15), .A2(maj_155_n14), .ZN(maj_155_n20)
         );
  XOR2_X1 maj_155_U9 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_155_n22) );
  XOR2_X1 maj_155_U8 ( .A(v_1_2[2]), .B(maj_155_n16), .Z(maj_155_n21) );
  XOR2_X1 maj_155_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_155_n16) );
  OR2_X1 maj_155_U6 ( .A1(maj_155_n20), .A2(maj_155_n19), .ZN(maj_155_n24) );
  NAND2_X1 maj_155_U5 ( .A1(maj_155_n24), .A2(maj_155_n23), .ZN(maj_155_n25)
         );
  NAND2_X1 maj_155_U4 ( .A1(maj_155_n20), .A2(maj_155_n19), .ZN(maj_155_n26)
         );
  NAND2_X1 maj_155_U3 ( .A1(maj_155_n26), .A2(maj_155_n25), .ZN(maj_155_port_o) );
  XOR2_X1 maj_155_U2 ( .A(maj_155_n22), .B(maj_155_n21), .Z(maj_155_n23) );
  NAND2_X1 maj_156_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_156_n18) );
  NAND2_X1 maj_156_U14 ( .A1(maj_156_n21), .A2(maj_156_n22), .ZN(maj_156_n17)
         );
  NAND2_X1 maj_156_U13 ( .A1(maj_156_n18), .A2(maj_156_n17), .ZN(maj_156_n19)
         );
  NAND2_X1 maj_156_U12 ( .A1(u_2_0[2]), .A2(maj_156_n16), .ZN(maj_156_n14) );
  NAND2_X1 maj_156_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_156_n15) );
  NAND2_X1 maj_156_U10 ( .A1(maj_156_n15), .A2(maj_156_n14), .ZN(maj_156_n20)
         );
  XOR2_X1 maj_156_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_156_n22) );
  XOR2_X1 maj_156_U8 ( .A(u_2_0[2]), .B(maj_156_n16), .Z(maj_156_n21) );
  XOR2_X1 maj_156_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_156_n16) );
  OR2_X1 maj_156_U6 ( .A1(maj_156_n20), .A2(maj_156_n19), .ZN(maj_156_n24) );
  NAND2_X1 maj_156_U5 ( .A1(maj_156_n24), .A2(maj_156_n23), .ZN(maj_156_n25)
         );
  NAND2_X1 maj_156_U4 ( .A1(maj_156_n20), .A2(maj_156_n19), .ZN(maj_156_n26)
         );
  NAND2_X1 maj_156_U3 ( .A1(maj_156_n26), .A2(maj_156_n25), .ZN(maj_156_port_o) );
  XOR2_X1 maj_156_U2 ( .A(maj_156_n22), .B(maj_156_n21), .Z(maj_156_n23) );
  NAND2_X1 maj_157_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_157_n18) );
  NAND2_X1 maj_157_U14 ( .A1(maj_157_n21), .A2(maj_157_n22), .ZN(maj_157_n17)
         );
  NAND2_X1 maj_157_U13 ( .A1(maj_157_n18), .A2(maj_157_n17), .ZN(maj_157_n19)
         );
  NAND2_X1 maj_157_U12 ( .A1(v_2_0[2]), .A2(maj_157_n16), .ZN(maj_157_n14) );
  NAND2_X1 maj_157_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_157_n15) );
  NAND2_X1 maj_157_U10 ( .A1(maj_157_n15), .A2(maj_157_n14), .ZN(maj_157_n20)
         );
  XOR2_X1 maj_157_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_157_n22) );
  XOR2_X1 maj_157_U8 ( .A(v_2_0[2]), .B(maj_157_n16), .Z(maj_157_n21) );
  XOR2_X1 maj_157_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_157_n16) );
  OR2_X1 maj_157_U6 ( .A1(maj_157_n20), .A2(maj_157_n19), .ZN(maj_157_n24) );
  NAND2_X1 maj_157_U5 ( .A1(maj_157_n24), .A2(maj_157_n23), .ZN(maj_157_n25)
         );
  NAND2_X1 maj_157_U4 ( .A1(maj_157_n20), .A2(maj_157_n19), .ZN(maj_157_n26)
         );
  NAND2_X1 maj_157_U3 ( .A1(maj_157_n26), .A2(maj_157_n25), .ZN(maj_157_port_o) );
  XOR2_X1 maj_157_U2 ( .A(maj_157_n22), .B(maj_157_n21), .Z(maj_157_n23) );
  NAND2_X1 maj_158_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_158_n18) );
  NAND2_X1 maj_158_U14 ( .A1(maj_158_n21), .A2(maj_158_n22), .ZN(maj_158_n17)
         );
  NAND2_X1 maj_158_U13 ( .A1(maj_158_n18), .A2(maj_158_n17), .ZN(maj_158_n19)
         );
  NAND2_X1 maj_158_U12 ( .A1(u_2_1[2]), .A2(maj_158_n16), .ZN(maj_158_n14) );
  NAND2_X1 maj_158_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_158_n15) );
  NAND2_X1 maj_158_U10 ( .A1(maj_158_n15), .A2(maj_158_n14), .ZN(maj_158_n20)
         );
  XOR2_X1 maj_158_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_158_n22) );
  XOR2_X1 maj_158_U8 ( .A(u_2_1[2]), .B(maj_158_n16), .Z(maj_158_n21) );
  XOR2_X1 maj_158_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_158_n16) );
  OR2_X1 maj_158_U6 ( .A1(maj_158_n20), .A2(maj_158_n19), .ZN(maj_158_n24) );
  NAND2_X1 maj_158_U5 ( .A1(maj_158_n24), .A2(maj_158_n23), .ZN(maj_158_n25)
         );
  NAND2_X1 maj_158_U4 ( .A1(maj_158_n20), .A2(maj_158_n19), .ZN(maj_158_n26)
         );
  NAND2_X1 maj_158_U3 ( .A1(maj_158_n26), .A2(maj_158_n25), .ZN(maj_158_port_o) );
  XOR2_X1 maj_158_U2 ( .A(maj_158_n22), .B(maj_158_n21), .Z(maj_158_n23) );
  NAND2_X1 maj_159_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_159_n18) );
  NAND2_X1 maj_159_U14 ( .A1(maj_159_n21), .A2(maj_159_n22), .ZN(maj_159_n17)
         );
  NAND2_X1 maj_159_U13 ( .A1(maj_159_n18), .A2(maj_159_n17), .ZN(maj_159_n19)
         );
  NAND2_X1 maj_159_U12 ( .A1(v_2_1[2]), .A2(maj_159_n16), .ZN(maj_159_n14) );
  NAND2_X1 maj_159_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_159_n15) );
  NAND2_X1 maj_159_U10 ( .A1(maj_159_n15), .A2(maj_159_n14), .ZN(maj_159_n20)
         );
  XOR2_X1 maj_159_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_159_n22) );
  XOR2_X1 maj_159_U8 ( .A(v_2_1[2]), .B(maj_159_n16), .Z(maj_159_n21) );
  XOR2_X1 maj_159_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_159_n16) );
  OR2_X1 maj_159_U6 ( .A1(maj_159_n20), .A2(maj_159_n19), .ZN(maj_159_n24) );
  NAND2_X1 maj_159_U5 ( .A1(maj_159_n24), .A2(maj_159_n23), .ZN(maj_159_n25)
         );
  NAND2_X1 maj_159_U4 ( .A1(maj_159_n20), .A2(maj_159_n19), .ZN(maj_159_n26)
         );
  NAND2_X1 maj_159_U3 ( .A1(maj_159_n26), .A2(maj_159_n25), .ZN(maj_159_port_o) );
  XOR2_X1 maj_159_U2 ( .A(maj_159_n22), .B(maj_159_n21), .Z(maj_159_n23) );
  NAND2_X1 maj_160_U15 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_160_n18) );
  NAND2_X1 maj_160_U14 ( .A1(maj_160_n21), .A2(maj_160_n22), .ZN(maj_160_n17)
         );
  NAND2_X1 maj_160_U13 ( .A1(maj_160_n18), .A2(maj_160_n17), .ZN(maj_160_n19)
         );
  NAND2_X1 maj_160_U12 ( .A1(u_2_2[2]), .A2(maj_160_n16), .ZN(maj_160_n14) );
  NAND2_X1 maj_160_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_160_n15) );
  NAND2_X1 maj_160_U10 ( .A1(maj_160_n15), .A2(maj_160_n14), .ZN(maj_160_n20)
         );
  XOR2_X1 maj_160_U9 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_160_n22) );
  XOR2_X1 maj_160_U8 ( .A(u_2_2[2]), .B(maj_160_n16), .Z(maj_160_n21) );
  XOR2_X1 maj_160_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_160_n16) );
  OR2_X1 maj_160_U6 ( .A1(maj_160_n20), .A2(maj_160_n19), .ZN(maj_160_n24) );
  NAND2_X1 maj_160_U5 ( .A1(maj_160_n24), .A2(maj_160_n23), .ZN(maj_160_n25)
         );
  NAND2_X1 maj_160_U4 ( .A1(maj_160_n20), .A2(maj_160_n19), .ZN(maj_160_n26)
         );
  NAND2_X1 maj_160_U3 ( .A1(maj_160_n26), .A2(maj_160_n25), .ZN(maj_160_port_o) );
  XOR2_X1 maj_160_U2 ( .A(maj_160_n22), .B(maj_160_n21), .Z(maj_160_n23) );
  NAND2_X1 maj_161_U15 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_161_n18) );
  NAND2_X1 maj_161_U14 ( .A1(maj_161_n21), .A2(maj_161_n22), .ZN(maj_161_n17)
         );
  NAND2_X1 maj_161_U13 ( .A1(maj_161_n18), .A2(maj_161_n17), .ZN(maj_161_n19)
         );
  NAND2_X1 maj_161_U12 ( .A1(v_2_2[2]), .A2(maj_161_n16), .ZN(maj_161_n14) );
  NAND2_X1 maj_161_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_161_n15) );
  NAND2_X1 maj_161_U10 ( .A1(maj_161_n15), .A2(maj_161_n14), .ZN(maj_161_n20)
         );
  XOR2_X1 maj_161_U9 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_161_n22) );
  XOR2_X1 maj_161_U8 ( .A(v_2_2[2]), .B(maj_161_n16), .Z(maj_161_n21) );
  XOR2_X1 maj_161_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_161_n16) );
  OR2_X1 maj_161_U6 ( .A1(maj_161_n20), .A2(maj_161_n19), .ZN(maj_161_n24) );
  NAND2_X1 maj_161_U5 ( .A1(maj_161_n24), .A2(maj_161_n23), .ZN(maj_161_n25)
         );
  NAND2_X1 maj_161_U4 ( .A1(maj_161_n20), .A2(maj_161_n19), .ZN(maj_161_n26)
         );
  NAND2_X1 maj_161_U3 ( .A1(maj_161_n26), .A2(maj_161_n25), .ZN(maj_161_port_o) );
  XOR2_X1 maj_161_U2 ( .A(maj_161_n22), .B(maj_161_n21), .Z(maj_161_n23) );
  NAND2_X1 maj_162_U15 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_162_n18) );
  NAND2_X1 maj_162_U14 ( .A1(maj_162_n21), .A2(maj_162_n22), .ZN(maj_162_n17)
         );
  NAND2_X1 maj_162_U13 ( .A1(maj_162_n18), .A2(maj_162_n17), .ZN(maj_162_n19)
         );
  NAND2_X1 maj_162_U12 ( .A1(u_3_0[2]), .A2(maj_162_n16), .ZN(maj_162_n14) );
  NAND2_X1 maj_162_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_162_n15) );
  NAND2_X1 maj_162_U10 ( .A1(maj_162_n15), .A2(maj_162_n14), .ZN(maj_162_n20)
         );
  XOR2_X1 maj_162_U9 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_162_n22) );
  XOR2_X1 maj_162_U8 ( .A(u_3_0[2]), .B(maj_162_n16), .Z(maj_162_n21) );
  XOR2_X1 maj_162_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_162_n16) );
  OR2_X1 maj_162_U6 ( .A1(maj_162_n20), .A2(maj_162_n19), .ZN(maj_162_n24) );
  NAND2_X1 maj_162_U5 ( .A1(maj_162_n24), .A2(maj_162_n23), .ZN(maj_162_n25)
         );
  NAND2_X1 maj_162_U4 ( .A1(maj_162_n20), .A2(maj_162_n19), .ZN(maj_162_n26)
         );
  NAND2_X1 maj_162_U3 ( .A1(maj_162_n26), .A2(maj_162_n25), .ZN(maj_162_port_o) );
  XOR2_X1 maj_162_U2 ( .A(maj_162_n22), .B(maj_162_n21), .Z(maj_162_n23) );
  NAND2_X1 maj_163_U15 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_163_n18) );
  NAND2_X1 maj_163_U14 ( .A1(maj_163_n21), .A2(maj_163_n22), .ZN(maj_163_n17)
         );
  NAND2_X1 maj_163_U13 ( .A1(maj_163_n18), .A2(maj_163_n17), .ZN(maj_163_n19)
         );
  NAND2_X1 maj_163_U12 ( .A1(v_3_0[2]), .A2(maj_163_n16), .ZN(maj_163_n14) );
  NAND2_X1 maj_163_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_163_n15) );
  NAND2_X1 maj_163_U10 ( .A1(maj_163_n15), .A2(maj_163_n14), .ZN(maj_163_n20)
         );
  XOR2_X1 maj_163_U9 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_163_n22) );
  XOR2_X1 maj_163_U8 ( .A(v_3_0[2]), .B(maj_163_n16), .Z(maj_163_n21) );
  XOR2_X1 maj_163_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_163_n16) );
  OR2_X1 maj_163_U6 ( .A1(maj_163_n20), .A2(maj_163_n19), .ZN(maj_163_n24) );
  NAND2_X1 maj_163_U5 ( .A1(maj_163_n24), .A2(maj_163_n23), .ZN(maj_163_n25)
         );
  NAND2_X1 maj_163_U4 ( .A1(maj_163_n20), .A2(maj_163_n19), .ZN(maj_163_n26)
         );
  NAND2_X1 maj_163_U3 ( .A1(maj_163_n26), .A2(maj_163_n25), .ZN(maj_163_port_o) );
  XOR2_X1 maj_163_U2 ( .A(maj_163_n22), .B(maj_163_n21), .Z(maj_163_n23) );
  NAND2_X1 maj_164_U15 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_164_n18) );
  NAND2_X1 maj_164_U14 ( .A1(maj_164_n21), .A2(maj_164_n22), .ZN(maj_164_n17)
         );
  NAND2_X1 maj_164_U13 ( .A1(maj_164_n18), .A2(maj_164_n17), .ZN(maj_164_n19)
         );
  NAND2_X1 maj_164_U12 ( .A1(u_3_1[2]), .A2(maj_164_n16), .ZN(maj_164_n14) );
  NAND2_X1 maj_164_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_164_n15) );
  NAND2_X1 maj_164_U10 ( .A1(maj_164_n15), .A2(maj_164_n14), .ZN(maj_164_n20)
         );
  XOR2_X1 maj_164_U9 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_164_n22) );
  XOR2_X1 maj_164_U8 ( .A(u_3_1[2]), .B(maj_164_n16), .Z(maj_164_n21) );
  XOR2_X1 maj_164_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_164_n16) );
  OR2_X1 maj_164_U6 ( .A1(maj_164_n20), .A2(maj_164_n19), .ZN(maj_164_n24) );
  NAND2_X1 maj_164_U5 ( .A1(maj_164_n24), .A2(maj_164_n23), .ZN(maj_164_n25)
         );
  NAND2_X1 maj_164_U4 ( .A1(maj_164_n20), .A2(maj_164_n19), .ZN(maj_164_n26)
         );
  NAND2_X1 maj_164_U3 ( .A1(maj_164_n26), .A2(maj_164_n25), .ZN(maj_164_port_o) );
  XOR2_X1 maj_164_U2 ( .A(maj_164_n22), .B(maj_164_n21), .Z(maj_164_n23) );
  NAND2_X1 maj_165_U15 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_165_n18) );
  NAND2_X1 maj_165_U14 ( .A1(maj_165_n21), .A2(maj_165_n22), .ZN(maj_165_n17)
         );
  NAND2_X1 maj_165_U13 ( .A1(maj_165_n18), .A2(maj_165_n17), .ZN(maj_165_n19)
         );
  NAND2_X1 maj_165_U12 ( .A1(v_3_1[2]), .A2(maj_165_n16), .ZN(maj_165_n14) );
  NAND2_X1 maj_165_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_165_n15) );
  NAND2_X1 maj_165_U10 ( .A1(maj_165_n15), .A2(maj_165_n14), .ZN(maj_165_n20)
         );
  XOR2_X1 maj_165_U9 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_165_n22) );
  XOR2_X1 maj_165_U8 ( .A(v_3_1[2]), .B(maj_165_n16), .Z(maj_165_n21) );
  XOR2_X1 maj_165_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_165_n16) );
  OR2_X1 maj_165_U6 ( .A1(maj_165_n20), .A2(maj_165_n19), .ZN(maj_165_n24) );
  NAND2_X1 maj_165_U5 ( .A1(maj_165_n24), .A2(maj_165_n23), .ZN(maj_165_n25)
         );
  NAND2_X1 maj_165_U4 ( .A1(maj_165_n20), .A2(maj_165_n19), .ZN(maj_165_n26)
         );
  NAND2_X1 maj_165_U3 ( .A1(maj_165_n26), .A2(maj_165_n25), .ZN(maj_165_port_o) );
  XOR2_X1 maj_165_U2 ( .A(maj_165_n22), .B(maj_165_n21), .Z(maj_165_n23) );
  NAND2_X1 maj_166_U15 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_166_n18) );
  NAND2_X1 maj_166_U14 ( .A1(maj_166_n21), .A2(maj_166_n22), .ZN(maj_166_n17)
         );
  NAND2_X1 maj_166_U13 ( .A1(maj_166_n18), .A2(maj_166_n17), .ZN(maj_166_n19)
         );
  NAND2_X1 maj_166_U12 ( .A1(u_3_2[2]), .A2(maj_166_n16), .ZN(maj_166_n14) );
  NAND2_X1 maj_166_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_166_n15) );
  NAND2_X1 maj_166_U10 ( .A1(maj_166_n15), .A2(maj_166_n14), .ZN(maj_166_n20)
         );
  XOR2_X1 maj_166_U9 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_166_n22) );
  XOR2_X1 maj_166_U8 ( .A(u_3_2[2]), .B(maj_166_n16), .Z(maj_166_n21) );
  XOR2_X1 maj_166_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_166_n16) );
  OR2_X1 maj_166_U6 ( .A1(maj_166_n20), .A2(maj_166_n19), .ZN(maj_166_n24) );
  NAND2_X1 maj_166_U5 ( .A1(maj_166_n24), .A2(maj_166_n23), .ZN(maj_166_n25)
         );
  NAND2_X1 maj_166_U4 ( .A1(maj_166_n20), .A2(maj_166_n19), .ZN(maj_166_n26)
         );
  NAND2_X1 maj_166_U3 ( .A1(maj_166_n26), .A2(maj_166_n25), .ZN(maj_166_port_o) );
  XOR2_X1 maj_166_U2 ( .A(maj_166_n22), .B(maj_166_n21), .Z(maj_166_n23) );
  NAND2_X1 maj_167_U15 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_167_n18) );
  NAND2_X1 maj_167_U14 ( .A1(maj_167_n21), .A2(maj_167_n22), .ZN(maj_167_n17)
         );
  NAND2_X1 maj_167_U13 ( .A1(maj_167_n18), .A2(maj_167_n17), .ZN(maj_167_n19)
         );
  NAND2_X1 maj_167_U12 ( .A1(v_3_2[2]), .A2(maj_167_n16), .ZN(maj_167_n14) );
  NAND2_X1 maj_167_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_167_n15) );
  NAND2_X1 maj_167_U10 ( .A1(maj_167_n15), .A2(maj_167_n14), .ZN(maj_167_n20)
         );
  XOR2_X1 maj_167_U9 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_167_n22) );
  XOR2_X1 maj_167_U8 ( .A(v_3_2[2]), .B(maj_167_n16), .Z(maj_167_n21) );
  XOR2_X1 maj_167_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_167_n16) );
  OR2_X1 maj_167_U6 ( .A1(maj_167_n20), .A2(maj_167_n19), .ZN(maj_167_n24) );
  NAND2_X1 maj_167_U5 ( .A1(maj_167_n24), .A2(maj_167_n23), .ZN(maj_167_n25)
         );
  NAND2_X1 maj_167_U4 ( .A1(maj_167_n20), .A2(maj_167_n19), .ZN(maj_167_n26)
         );
  NAND2_X1 maj_167_U3 ( .A1(maj_167_n26), .A2(maj_167_n25), .ZN(maj_167_port_o) );
  XOR2_X1 maj_167_U2 ( .A(maj_167_n22), .B(maj_167_n21), .Z(maj_167_n23) );
  NAND2_X1 maj_168_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_168_n18) );
  NAND2_X1 maj_168_U14 ( .A1(maj_168_n21), .A2(maj_168_n22), .ZN(maj_168_n17)
         );
  NAND2_X1 maj_168_U13 ( .A1(maj_168_n18), .A2(maj_168_n17), .ZN(maj_168_n19)
         );
  NAND2_X1 maj_168_U12 ( .A1(u_0_0[2]), .A2(maj_168_n16), .ZN(maj_168_n14) );
  NAND2_X1 maj_168_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_168_n15) );
  NAND2_X1 maj_168_U10 ( .A1(maj_168_n15), .A2(maj_168_n14), .ZN(maj_168_n20)
         );
  XOR2_X1 maj_168_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_168_n22) );
  XOR2_X1 maj_168_U8 ( .A(u_0_0[2]), .B(maj_168_n16), .Z(maj_168_n21) );
  XOR2_X1 maj_168_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_168_n16) );
  OR2_X1 maj_168_U6 ( .A1(maj_168_n20), .A2(maj_168_n19), .ZN(maj_168_n24) );
  NAND2_X1 maj_168_U5 ( .A1(maj_168_n24), .A2(maj_168_n23), .ZN(maj_168_n25)
         );
  NAND2_X1 maj_168_U4 ( .A1(maj_168_n20), .A2(maj_168_n19), .ZN(maj_168_n26)
         );
  NAND2_X1 maj_168_U3 ( .A1(maj_168_n26), .A2(maj_168_n25), .ZN(maj_168_port_o) );
  XOR2_X1 maj_168_U2 ( .A(maj_168_n22), .B(maj_168_n21), .Z(maj_168_n23) );
  NAND2_X1 maj_169_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_169_n18) );
  NAND2_X1 maj_169_U14 ( .A1(maj_169_n21), .A2(maj_169_n22), .ZN(maj_169_n17)
         );
  NAND2_X1 maj_169_U13 ( .A1(maj_169_n18), .A2(maj_169_n17), .ZN(maj_169_n19)
         );
  NAND2_X1 maj_169_U12 ( .A1(v_0_0[2]), .A2(maj_169_n16), .ZN(maj_169_n14) );
  NAND2_X1 maj_169_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_169_n15) );
  NAND2_X1 maj_169_U10 ( .A1(maj_169_n15), .A2(maj_169_n14), .ZN(maj_169_n20)
         );
  XOR2_X1 maj_169_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_169_n22) );
  XOR2_X1 maj_169_U8 ( .A(v_0_0[2]), .B(maj_169_n16), .Z(maj_169_n21) );
  XOR2_X1 maj_169_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_169_n16) );
  OR2_X1 maj_169_U6 ( .A1(maj_169_n20), .A2(maj_169_n19), .ZN(maj_169_n24) );
  NAND2_X1 maj_169_U5 ( .A1(maj_169_n24), .A2(maj_169_n23), .ZN(maj_169_n25)
         );
  NAND2_X1 maj_169_U4 ( .A1(maj_169_n20), .A2(maj_169_n19), .ZN(maj_169_n26)
         );
  NAND2_X1 maj_169_U3 ( .A1(maj_169_n26), .A2(maj_169_n25), .ZN(maj_169_port_o) );
  XOR2_X1 maj_169_U2 ( .A(maj_169_n22), .B(maj_169_n21), .Z(maj_169_n23) );
  NAND2_X1 maj_170_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_170_n18) );
  NAND2_X1 maj_170_U14 ( .A1(maj_170_n21), .A2(maj_170_n22), .ZN(maj_170_n17)
         );
  NAND2_X1 maj_170_U13 ( .A1(maj_170_n18), .A2(maj_170_n17), .ZN(maj_170_n19)
         );
  NAND2_X1 maj_170_U12 ( .A1(u_0_1[2]), .A2(maj_170_n16), .ZN(maj_170_n14) );
  NAND2_X1 maj_170_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_170_n15) );
  NAND2_X1 maj_170_U10 ( .A1(maj_170_n15), .A2(maj_170_n14), .ZN(maj_170_n20)
         );
  XOR2_X1 maj_170_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_170_n22) );
  XOR2_X1 maj_170_U8 ( .A(u_0_1[2]), .B(maj_170_n16), .Z(maj_170_n21) );
  XOR2_X1 maj_170_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_170_n16) );
  OR2_X1 maj_170_U6 ( .A1(maj_170_n20), .A2(maj_170_n19), .ZN(maj_170_n24) );
  NAND2_X1 maj_170_U5 ( .A1(maj_170_n24), .A2(maj_170_n23), .ZN(maj_170_n25)
         );
  NAND2_X1 maj_170_U4 ( .A1(maj_170_n20), .A2(maj_170_n19), .ZN(maj_170_n26)
         );
  NAND2_X1 maj_170_U3 ( .A1(maj_170_n26), .A2(maj_170_n25), .ZN(maj_170_port_o) );
  XOR2_X1 maj_170_U2 ( .A(maj_170_n22), .B(maj_170_n21), .Z(maj_170_n23) );
  NAND2_X1 maj_171_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_171_n18) );
  NAND2_X1 maj_171_U14 ( .A1(maj_171_n21), .A2(maj_171_n22), .ZN(maj_171_n17)
         );
  NAND2_X1 maj_171_U13 ( .A1(maj_171_n18), .A2(maj_171_n17), .ZN(maj_171_n19)
         );
  NAND2_X1 maj_171_U12 ( .A1(v_0_1[2]), .A2(maj_171_n16), .ZN(maj_171_n14) );
  NAND2_X1 maj_171_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_171_n15) );
  NAND2_X1 maj_171_U10 ( .A1(maj_171_n15), .A2(maj_171_n14), .ZN(maj_171_n20)
         );
  XOR2_X1 maj_171_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_171_n22) );
  XOR2_X1 maj_171_U8 ( .A(v_0_1[2]), .B(maj_171_n16), .Z(maj_171_n21) );
  XOR2_X1 maj_171_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_171_n16) );
  OR2_X1 maj_171_U6 ( .A1(maj_171_n20), .A2(maj_171_n19), .ZN(maj_171_n24) );
  NAND2_X1 maj_171_U5 ( .A1(maj_171_n24), .A2(maj_171_n23), .ZN(maj_171_n25)
         );
  NAND2_X1 maj_171_U4 ( .A1(maj_171_n20), .A2(maj_171_n19), .ZN(maj_171_n26)
         );
  NAND2_X1 maj_171_U3 ( .A1(maj_171_n26), .A2(maj_171_n25), .ZN(maj_171_port_o) );
  XOR2_X1 maj_171_U2 ( .A(maj_171_n22), .B(maj_171_n21), .Z(maj_171_n23) );
  NAND2_X1 maj_172_U15 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_172_n18) );
  NAND2_X1 maj_172_U14 ( .A1(maj_172_n21), .A2(maj_172_n22), .ZN(maj_172_n17)
         );
  NAND2_X1 maj_172_U13 ( .A1(maj_172_n18), .A2(maj_172_n17), .ZN(maj_172_n19)
         );
  NAND2_X1 maj_172_U12 ( .A1(u_0_2[2]), .A2(maj_172_n16), .ZN(maj_172_n14) );
  NAND2_X1 maj_172_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_172_n15) );
  NAND2_X1 maj_172_U10 ( .A1(maj_172_n15), .A2(maj_172_n14), .ZN(maj_172_n20)
         );
  XOR2_X1 maj_172_U9 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_172_n22) );
  XOR2_X1 maj_172_U8 ( .A(u_0_2[2]), .B(maj_172_n16), .Z(maj_172_n21) );
  XOR2_X1 maj_172_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_172_n16) );
  OR2_X1 maj_172_U6 ( .A1(maj_172_n20), .A2(maj_172_n19), .ZN(maj_172_n24) );
  NAND2_X1 maj_172_U5 ( .A1(maj_172_n24), .A2(maj_172_n23), .ZN(maj_172_n25)
         );
  NAND2_X1 maj_172_U4 ( .A1(maj_172_n20), .A2(maj_172_n19), .ZN(maj_172_n26)
         );
  NAND2_X1 maj_172_U3 ( .A1(maj_172_n26), .A2(maj_172_n25), .ZN(maj_172_port_o) );
  XOR2_X1 maj_172_U2 ( .A(maj_172_n22), .B(maj_172_n21), .Z(maj_172_n23) );
  NAND2_X1 maj_173_U15 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_173_n18) );
  NAND2_X1 maj_173_U14 ( .A1(maj_173_n21), .A2(maj_173_n22), .ZN(maj_173_n17)
         );
  NAND2_X1 maj_173_U13 ( .A1(maj_173_n18), .A2(maj_173_n17), .ZN(maj_173_n19)
         );
  NAND2_X1 maj_173_U12 ( .A1(v_0_2[2]), .A2(maj_173_n16), .ZN(maj_173_n14) );
  NAND2_X1 maj_173_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_173_n15) );
  NAND2_X1 maj_173_U10 ( .A1(maj_173_n15), .A2(maj_173_n14), .ZN(maj_173_n20)
         );
  XOR2_X1 maj_173_U9 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_173_n22) );
  XOR2_X1 maj_173_U8 ( .A(v_0_2[2]), .B(maj_173_n16), .Z(maj_173_n21) );
  XOR2_X1 maj_173_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_173_n16) );
  OR2_X1 maj_173_U6 ( .A1(maj_173_n20), .A2(maj_173_n19), .ZN(maj_173_n24) );
  NAND2_X1 maj_173_U5 ( .A1(maj_173_n24), .A2(maj_173_n23), .ZN(maj_173_n25)
         );
  NAND2_X1 maj_173_U4 ( .A1(maj_173_n20), .A2(maj_173_n19), .ZN(maj_173_n26)
         );
  NAND2_X1 maj_173_U3 ( .A1(maj_173_n26), .A2(maj_173_n25), .ZN(maj_173_port_o) );
  XOR2_X1 maj_173_U2 ( .A(maj_173_n22), .B(maj_173_n21), .Z(maj_173_n23) );
  NAND2_X1 maj_174_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_174_n18) );
  NAND2_X1 maj_174_U14 ( .A1(maj_174_n21), .A2(maj_174_n22), .ZN(maj_174_n17)
         );
  NAND2_X1 maj_174_U13 ( .A1(maj_174_n18), .A2(maj_174_n17), .ZN(maj_174_n19)
         );
  NAND2_X1 maj_174_U12 ( .A1(u_1_0[2]), .A2(maj_174_n16), .ZN(maj_174_n14) );
  NAND2_X1 maj_174_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_174_n15) );
  NAND2_X1 maj_174_U10 ( .A1(maj_174_n15), .A2(maj_174_n14), .ZN(maj_174_n20)
         );
  XOR2_X1 maj_174_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_174_n22) );
  XOR2_X1 maj_174_U8 ( .A(u_1_0[2]), .B(maj_174_n16), .Z(maj_174_n21) );
  XOR2_X1 maj_174_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_174_n16) );
  OR2_X1 maj_174_U6 ( .A1(maj_174_n20), .A2(maj_174_n19), .ZN(maj_174_n24) );
  NAND2_X1 maj_174_U5 ( .A1(maj_174_n24), .A2(maj_174_n23), .ZN(maj_174_n25)
         );
  NAND2_X1 maj_174_U4 ( .A1(maj_174_n20), .A2(maj_174_n19), .ZN(maj_174_n26)
         );
  NAND2_X1 maj_174_U3 ( .A1(maj_174_n26), .A2(maj_174_n25), .ZN(maj_174_port_o) );
  XOR2_X1 maj_174_U2 ( .A(maj_174_n22), .B(maj_174_n21), .Z(maj_174_n23) );
  NAND2_X1 maj_175_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_175_n18) );
  NAND2_X1 maj_175_U14 ( .A1(maj_175_n21), .A2(maj_175_n22), .ZN(maj_175_n17)
         );
  NAND2_X1 maj_175_U13 ( .A1(maj_175_n18), .A2(maj_175_n17), .ZN(maj_175_n19)
         );
  NAND2_X1 maj_175_U12 ( .A1(v_1_0[2]), .A2(maj_175_n16), .ZN(maj_175_n14) );
  NAND2_X1 maj_175_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_175_n15) );
  NAND2_X1 maj_175_U10 ( .A1(maj_175_n15), .A2(maj_175_n14), .ZN(maj_175_n20)
         );
  XOR2_X1 maj_175_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_175_n22) );
  XOR2_X1 maj_175_U8 ( .A(v_1_0[2]), .B(maj_175_n16), .Z(maj_175_n21) );
  XOR2_X1 maj_175_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_175_n16) );
  OR2_X1 maj_175_U6 ( .A1(maj_175_n20), .A2(maj_175_n19), .ZN(maj_175_n24) );
  NAND2_X1 maj_175_U5 ( .A1(maj_175_n24), .A2(maj_175_n23), .ZN(maj_175_n25)
         );
  NAND2_X1 maj_175_U4 ( .A1(maj_175_n20), .A2(maj_175_n19), .ZN(maj_175_n26)
         );
  NAND2_X1 maj_175_U3 ( .A1(maj_175_n26), .A2(maj_175_n25), .ZN(maj_175_port_o) );
  XOR2_X1 maj_175_U2 ( .A(maj_175_n22), .B(maj_175_n21), .Z(maj_175_n23) );
  NAND2_X1 maj_176_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_176_n18) );
  NAND2_X1 maj_176_U14 ( .A1(maj_176_n21), .A2(maj_176_n22), .ZN(maj_176_n17)
         );
  NAND2_X1 maj_176_U13 ( .A1(maj_176_n18), .A2(maj_176_n17), .ZN(maj_176_n19)
         );
  NAND2_X1 maj_176_U12 ( .A1(u_1_1[2]), .A2(maj_176_n16), .ZN(maj_176_n14) );
  NAND2_X1 maj_176_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_176_n15) );
  NAND2_X1 maj_176_U10 ( .A1(maj_176_n15), .A2(maj_176_n14), .ZN(maj_176_n20)
         );
  XOR2_X1 maj_176_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_176_n22) );
  XOR2_X1 maj_176_U8 ( .A(u_1_1[2]), .B(maj_176_n16), .Z(maj_176_n21) );
  XOR2_X1 maj_176_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_176_n16) );
  OR2_X1 maj_176_U6 ( .A1(maj_176_n20), .A2(maj_176_n19), .ZN(maj_176_n24) );
  NAND2_X1 maj_176_U5 ( .A1(maj_176_n24), .A2(maj_176_n23), .ZN(maj_176_n25)
         );
  NAND2_X1 maj_176_U4 ( .A1(maj_176_n20), .A2(maj_176_n19), .ZN(maj_176_n26)
         );
  NAND2_X1 maj_176_U3 ( .A1(maj_176_n26), .A2(maj_176_n25), .ZN(maj_176_port_o) );
  XOR2_X1 maj_176_U2 ( .A(maj_176_n22), .B(maj_176_n21), .Z(maj_176_n23) );
  NAND2_X1 maj_177_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_177_n18) );
  NAND2_X1 maj_177_U14 ( .A1(maj_177_n21), .A2(maj_177_n22), .ZN(maj_177_n17)
         );
  NAND2_X1 maj_177_U13 ( .A1(maj_177_n18), .A2(maj_177_n17), .ZN(maj_177_n19)
         );
  NAND2_X1 maj_177_U12 ( .A1(v_1_1[2]), .A2(maj_177_n16), .ZN(maj_177_n14) );
  NAND2_X1 maj_177_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_177_n15) );
  NAND2_X1 maj_177_U10 ( .A1(maj_177_n15), .A2(maj_177_n14), .ZN(maj_177_n20)
         );
  XOR2_X1 maj_177_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_177_n22) );
  XOR2_X1 maj_177_U8 ( .A(v_1_1[2]), .B(maj_177_n16), .Z(maj_177_n21) );
  XOR2_X1 maj_177_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_177_n16) );
  OR2_X1 maj_177_U6 ( .A1(maj_177_n20), .A2(maj_177_n19), .ZN(maj_177_n24) );
  NAND2_X1 maj_177_U5 ( .A1(maj_177_n24), .A2(maj_177_n23), .ZN(maj_177_n25)
         );
  NAND2_X1 maj_177_U4 ( .A1(maj_177_n20), .A2(maj_177_n19), .ZN(maj_177_n26)
         );
  NAND2_X1 maj_177_U3 ( .A1(maj_177_n26), .A2(maj_177_n25), .ZN(maj_177_port_o) );
  XOR2_X1 maj_177_U2 ( .A(maj_177_n22), .B(maj_177_n21), .Z(maj_177_n23) );
  NAND2_X1 maj_178_U15 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_178_n18) );
  NAND2_X1 maj_178_U14 ( .A1(maj_178_n21), .A2(maj_178_n22), .ZN(maj_178_n17)
         );
  NAND2_X1 maj_178_U13 ( .A1(maj_178_n18), .A2(maj_178_n17), .ZN(maj_178_n19)
         );
  NAND2_X1 maj_178_U12 ( .A1(u_1_2[2]), .A2(maj_178_n16), .ZN(maj_178_n14) );
  NAND2_X1 maj_178_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_178_n15) );
  NAND2_X1 maj_178_U10 ( .A1(maj_178_n15), .A2(maj_178_n14), .ZN(maj_178_n20)
         );
  XOR2_X1 maj_178_U9 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_178_n22) );
  XOR2_X1 maj_178_U8 ( .A(u_1_2[2]), .B(maj_178_n16), .Z(maj_178_n21) );
  XOR2_X1 maj_178_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_178_n16) );
  OR2_X1 maj_178_U6 ( .A1(maj_178_n20), .A2(maj_178_n19), .ZN(maj_178_n24) );
  NAND2_X1 maj_178_U5 ( .A1(maj_178_n24), .A2(maj_178_n23), .ZN(maj_178_n25)
         );
  NAND2_X1 maj_178_U4 ( .A1(maj_178_n20), .A2(maj_178_n19), .ZN(maj_178_n26)
         );
  NAND2_X1 maj_178_U3 ( .A1(maj_178_n26), .A2(maj_178_n25), .ZN(maj_178_port_o) );
  XOR2_X1 maj_178_U2 ( .A(maj_178_n22), .B(maj_178_n21), .Z(maj_178_n23) );
  NAND2_X1 maj_179_U15 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_179_n18) );
  NAND2_X1 maj_179_U14 ( .A1(maj_179_n21), .A2(maj_179_n22), .ZN(maj_179_n17)
         );
  NAND2_X1 maj_179_U13 ( .A1(maj_179_n18), .A2(maj_179_n17), .ZN(maj_179_n19)
         );
  NAND2_X1 maj_179_U12 ( .A1(v_1_2[2]), .A2(maj_179_n16), .ZN(maj_179_n14) );
  NAND2_X1 maj_179_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_179_n15) );
  NAND2_X1 maj_179_U10 ( .A1(maj_179_n15), .A2(maj_179_n14), .ZN(maj_179_n20)
         );
  XOR2_X1 maj_179_U9 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_179_n22) );
  XOR2_X1 maj_179_U8 ( .A(v_1_2[2]), .B(maj_179_n16), .Z(maj_179_n21) );
  XOR2_X1 maj_179_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_179_n16) );
  OR2_X1 maj_179_U6 ( .A1(maj_179_n20), .A2(maj_179_n19), .ZN(maj_179_n24) );
  NAND2_X1 maj_179_U5 ( .A1(maj_179_n24), .A2(maj_179_n23), .ZN(maj_179_n25)
         );
  NAND2_X1 maj_179_U4 ( .A1(maj_179_n20), .A2(maj_179_n19), .ZN(maj_179_n26)
         );
  NAND2_X1 maj_179_U3 ( .A1(maj_179_n26), .A2(maj_179_n25), .ZN(maj_179_port_o) );
  XOR2_X1 maj_179_U2 ( .A(maj_179_n22), .B(maj_179_n21), .Z(maj_179_n23) );
  NAND2_X1 maj_180_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_180_n18) );
  NAND2_X1 maj_180_U14 ( .A1(maj_180_n21), .A2(maj_180_n22), .ZN(maj_180_n17)
         );
  NAND2_X1 maj_180_U13 ( .A1(maj_180_n18), .A2(maj_180_n17), .ZN(maj_180_n19)
         );
  NAND2_X1 maj_180_U12 ( .A1(u_2_0[2]), .A2(maj_180_n16), .ZN(maj_180_n14) );
  NAND2_X1 maj_180_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_180_n15) );
  NAND2_X1 maj_180_U10 ( .A1(maj_180_n15), .A2(maj_180_n14), .ZN(maj_180_n20)
         );
  XOR2_X1 maj_180_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_180_n22) );
  XOR2_X1 maj_180_U8 ( .A(u_2_0[2]), .B(maj_180_n16), .Z(maj_180_n21) );
  XOR2_X1 maj_180_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_180_n16) );
  OR2_X1 maj_180_U6 ( .A1(maj_180_n20), .A2(maj_180_n19), .ZN(maj_180_n24) );
  NAND2_X1 maj_180_U5 ( .A1(maj_180_n24), .A2(maj_180_n23), .ZN(maj_180_n25)
         );
  NAND2_X1 maj_180_U4 ( .A1(maj_180_n20), .A2(maj_180_n19), .ZN(maj_180_n26)
         );
  NAND2_X1 maj_180_U3 ( .A1(maj_180_n26), .A2(maj_180_n25), .ZN(maj_180_port_o) );
  XOR2_X1 maj_180_U2 ( .A(maj_180_n22), .B(maj_180_n21), .Z(maj_180_n23) );
  NAND2_X1 maj_181_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_181_n18) );
  NAND2_X1 maj_181_U14 ( .A1(maj_181_n21), .A2(maj_181_n22), .ZN(maj_181_n17)
         );
  NAND2_X1 maj_181_U13 ( .A1(maj_181_n18), .A2(maj_181_n17), .ZN(maj_181_n19)
         );
  NAND2_X1 maj_181_U12 ( .A1(v_2_0[2]), .A2(maj_181_n16), .ZN(maj_181_n14) );
  NAND2_X1 maj_181_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_181_n15) );
  NAND2_X1 maj_181_U10 ( .A1(maj_181_n15), .A2(maj_181_n14), .ZN(maj_181_n20)
         );
  XOR2_X1 maj_181_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_181_n22) );
  XOR2_X1 maj_181_U8 ( .A(v_2_0[2]), .B(maj_181_n16), .Z(maj_181_n21) );
  XOR2_X1 maj_181_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_181_n16) );
  OR2_X1 maj_181_U6 ( .A1(maj_181_n20), .A2(maj_181_n19), .ZN(maj_181_n24) );
  NAND2_X1 maj_181_U5 ( .A1(maj_181_n24), .A2(maj_181_n23), .ZN(maj_181_n25)
         );
  NAND2_X1 maj_181_U4 ( .A1(maj_181_n20), .A2(maj_181_n19), .ZN(maj_181_n26)
         );
  NAND2_X1 maj_181_U3 ( .A1(maj_181_n26), .A2(maj_181_n25), .ZN(maj_181_port_o) );
  XOR2_X1 maj_181_U2 ( .A(maj_181_n22), .B(maj_181_n21), .Z(maj_181_n23) );
  NAND2_X1 maj_182_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_182_n18) );
  NAND2_X1 maj_182_U14 ( .A1(maj_182_n21), .A2(maj_182_n22), .ZN(maj_182_n17)
         );
  NAND2_X1 maj_182_U13 ( .A1(maj_182_n18), .A2(maj_182_n17), .ZN(maj_182_n19)
         );
  NAND2_X1 maj_182_U12 ( .A1(u_2_1[2]), .A2(maj_182_n16), .ZN(maj_182_n14) );
  NAND2_X1 maj_182_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_182_n15) );
  NAND2_X1 maj_182_U10 ( .A1(maj_182_n15), .A2(maj_182_n14), .ZN(maj_182_n20)
         );
  XOR2_X1 maj_182_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_182_n22) );
  XOR2_X1 maj_182_U8 ( .A(u_2_1[2]), .B(maj_182_n16), .Z(maj_182_n21) );
  XOR2_X1 maj_182_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_182_n16) );
  OR2_X1 maj_182_U6 ( .A1(maj_182_n20), .A2(maj_182_n19), .ZN(maj_182_n24) );
  NAND2_X1 maj_182_U5 ( .A1(maj_182_n24), .A2(maj_182_n23), .ZN(maj_182_n25)
         );
  NAND2_X1 maj_182_U4 ( .A1(maj_182_n20), .A2(maj_182_n19), .ZN(maj_182_n26)
         );
  NAND2_X1 maj_182_U3 ( .A1(maj_182_n26), .A2(maj_182_n25), .ZN(maj_182_port_o) );
  XOR2_X1 maj_182_U2 ( .A(maj_182_n22), .B(maj_182_n21), .Z(maj_182_n23) );
  NAND2_X1 maj_183_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_183_n18) );
  NAND2_X1 maj_183_U14 ( .A1(maj_183_n21), .A2(maj_183_n22), .ZN(maj_183_n17)
         );
  NAND2_X1 maj_183_U13 ( .A1(maj_183_n18), .A2(maj_183_n17), .ZN(maj_183_n19)
         );
  NAND2_X1 maj_183_U12 ( .A1(v_2_1[2]), .A2(maj_183_n16), .ZN(maj_183_n14) );
  NAND2_X1 maj_183_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_183_n15) );
  NAND2_X1 maj_183_U10 ( .A1(maj_183_n15), .A2(maj_183_n14), .ZN(maj_183_n20)
         );
  XOR2_X1 maj_183_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_183_n22) );
  XOR2_X1 maj_183_U8 ( .A(v_2_1[2]), .B(maj_183_n16), .Z(maj_183_n21) );
  XOR2_X1 maj_183_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_183_n16) );
  OR2_X1 maj_183_U6 ( .A1(maj_183_n20), .A2(maj_183_n19), .ZN(maj_183_n24) );
  NAND2_X1 maj_183_U5 ( .A1(maj_183_n24), .A2(maj_183_n23), .ZN(maj_183_n25)
         );
  NAND2_X1 maj_183_U4 ( .A1(maj_183_n20), .A2(maj_183_n19), .ZN(maj_183_n26)
         );
  NAND2_X1 maj_183_U3 ( .A1(maj_183_n26), .A2(maj_183_n25), .ZN(maj_183_port_o) );
  XOR2_X1 maj_183_U2 ( .A(maj_183_n22), .B(maj_183_n21), .Z(maj_183_n23) );
  NAND2_X1 maj_184_U15 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_184_n18) );
  NAND2_X1 maj_184_U14 ( .A1(maj_184_n21), .A2(maj_184_n22), .ZN(maj_184_n17)
         );
  NAND2_X1 maj_184_U13 ( .A1(maj_184_n18), .A2(maj_184_n17), .ZN(maj_184_n19)
         );
  NAND2_X1 maj_184_U12 ( .A1(u_2_2[2]), .A2(maj_184_n16), .ZN(maj_184_n14) );
  NAND2_X1 maj_184_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_184_n15) );
  NAND2_X1 maj_184_U10 ( .A1(maj_184_n15), .A2(maj_184_n14), .ZN(maj_184_n20)
         );
  XOR2_X1 maj_184_U9 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_184_n22) );
  XOR2_X1 maj_184_U8 ( .A(u_2_2[2]), .B(maj_184_n16), .Z(maj_184_n21) );
  XOR2_X1 maj_184_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_184_n16) );
  OR2_X1 maj_184_U6 ( .A1(maj_184_n20), .A2(maj_184_n19), .ZN(maj_184_n24) );
  NAND2_X1 maj_184_U5 ( .A1(maj_184_n24), .A2(maj_184_n23), .ZN(maj_184_n25)
         );
  NAND2_X1 maj_184_U4 ( .A1(maj_184_n20), .A2(maj_184_n19), .ZN(maj_184_n26)
         );
  NAND2_X1 maj_184_U3 ( .A1(maj_184_n26), .A2(maj_184_n25), .ZN(maj_184_port_o) );
  XOR2_X1 maj_184_U2 ( .A(maj_184_n22), .B(maj_184_n21), .Z(maj_184_n23) );
  NAND2_X1 maj_185_U15 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_185_n18) );
  NAND2_X1 maj_185_U14 ( .A1(maj_185_n21), .A2(maj_185_n22), .ZN(maj_185_n17)
         );
  NAND2_X1 maj_185_U13 ( .A1(maj_185_n18), .A2(maj_185_n17), .ZN(maj_185_n19)
         );
  NAND2_X1 maj_185_U12 ( .A1(v_2_2[2]), .A2(maj_185_n16), .ZN(maj_185_n14) );
  NAND2_X1 maj_185_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_185_n15) );
  NAND2_X1 maj_185_U10 ( .A1(maj_185_n15), .A2(maj_185_n14), .ZN(maj_185_n20)
         );
  XOR2_X1 maj_185_U9 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_185_n22) );
  XOR2_X1 maj_185_U8 ( .A(v_2_2[2]), .B(maj_185_n16), .Z(maj_185_n21) );
  XOR2_X1 maj_185_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_185_n16) );
  OR2_X1 maj_185_U6 ( .A1(maj_185_n20), .A2(maj_185_n19), .ZN(maj_185_n24) );
  NAND2_X1 maj_185_U5 ( .A1(maj_185_n24), .A2(maj_185_n23), .ZN(maj_185_n25)
         );
  NAND2_X1 maj_185_U4 ( .A1(maj_185_n20), .A2(maj_185_n19), .ZN(maj_185_n26)
         );
  NAND2_X1 maj_185_U3 ( .A1(maj_185_n26), .A2(maj_185_n25), .ZN(maj_185_port_o) );
  XOR2_X1 maj_185_U2 ( .A(maj_185_n22), .B(maj_185_n21), .Z(maj_185_n23) );
  NAND2_X1 maj_186_U15 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_186_n18) );
  NAND2_X1 maj_186_U14 ( .A1(maj_186_n21), .A2(maj_186_n22), .ZN(maj_186_n17)
         );
  NAND2_X1 maj_186_U13 ( .A1(maj_186_n18), .A2(maj_186_n17), .ZN(maj_186_n19)
         );
  NAND2_X1 maj_186_U12 ( .A1(u_3_0[2]), .A2(maj_186_n16), .ZN(maj_186_n14) );
  NAND2_X1 maj_186_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_186_n15) );
  NAND2_X1 maj_186_U10 ( .A1(maj_186_n15), .A2(maj_186_n14), .ZN(maj_186_n20)
         );
  XOR2_X1 maj_186_U9 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_186_n22) );
  XOR2_X1 maj_186_U8 ( .A(u_3_0[2]), .B(maj_186_n16), .Z(maj_186_n21) );
  XOR2_X1 maj_186_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_186_n16) );
  OR2_X1 maj_186_U6 ( .A1(maj_186_n20), .A2(maj_186_n19), .ZN(maj_186_n24) );
  NAND2_X1 maj_186_U5 ( .A1(maj_186_n24), .A2(maj_186_n23), .ZN(maj_186_n25)
         );
  NAND2_X1 maj_186_U4 ( .A1(maj_186_n20), .A2(maj_186_n19), .ZN(maj_186_n26)
         );
  NAND2_X1 maj_186_U3 ( .A1(maj_186_n26), .A2(maj_186_n25), .ZN(maj_186_port_o) );
  XOR2_X1 maj_186_U2 ( .A(maj_186_n22), .B(maj_186_n21), .Z(maj_186_n23) );
  NAND2_X1 maj_187_U15 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_187_n18) );
  NAND2_X1 maj_187_U14 ( .A1(maj_187_n21), .A2(maj_187_n22), .ZN(maj_187_n17)
         );
  NAND2_X1 maj_187_U13 ( .A1(maj_187_n18), .A2(maj_187_n17), .ZN(maj_187_n19)
         );
  NAND2_X1 maj_187_U12 ( .A1(v_3_0[2]), .A2(maj_187_n16), .ZN(maj_187_n14) );
  NAND2_X1 maj_187_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_187_n15) );
  NAND2_X1 maj_187_U10 ( .A1(maj_187_n15), .A2(maj_187_n14), .ZN(maj_187_n20)
         );
  XOR2_X1 maj_187_U9 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_187_n22) );
  XOR2_X1 maj_187_U8 ( .A(v_3_0[2]), .B(maj_187_n16), .Z(maj_187_n21) );
  XOR2_X1 maj_187_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_187_n16) );
  OR2_X1 maj_187_U6 ( .A1(maj_187_n20), .A2(maj_187_n19), .ZN(maj_187_n24) );
  NAND2_X1 maj_187_U5 ( .A1(maj_187_n24), .A2(maj_187_n23), .ZN(maj_187_n25)
         );
  NAND2_X1 maj_187_U4 ( .A1(maj_187_n20), .A2(maj_187_n19), .ZN(maj_187_n26)
         );
  NAND2_X1 maj_187_U3 ( .A1(maj_187_n26), .A2(maj_187_n25), .ZN(maj_187_port_o) );
  XOR2_X1 maj_187_U2 ( .A(maj_187_n22), .B(maj_187_n21), .Z(maj_187_n23) );
  NAND2_X1 maj_188_U15 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_188_n18) );
  NAND2_X1 maj_188_U14 ( .A1(maj_188_n21), .A2(maj_188_n22), .ZN(maj_188_n17)
         );
  NAND2_X1 maj_188_U13 ( .A1(maj_188_n18), .A2(maj_188_n17), .ZN(maj_188_n19)
         );
  NAND2_X1 maj_188_U12 ( .A1(u_3_1[2]), .A2(maj_188_n16), .ZN(maj_188_n14) );
  NAND2_X1 maj_188_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_188_n15) );
  NAND2_X1 maj_188_U10 ( .A1(maj_188_n15), .A2(maj_188_n14), .ZN(maj_188_n20)
         );
  XOR2_X1 maj_188_U9 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_188_n22) );
  XOR2_X1 maj_188_U8 ( .A(u_3_1[2]), .B(maj_188_n16), .Z(maj_188_n21) );
  XOR2_X1 maj_188_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_188_n16) );
  OR2_X1 maj_188_U6 ( .A1(maj_188_n20), .A2(maj_188_n19), .ZN(maj_188_n24) );
  NAND2_X1 maj_188_U5 ( .A1(maj_188_n24), .A2(maj_188_n23), .ZN(maj_188_n25)
         );
  NAND2_X1 maj_188_U4 ( .A1(maj_188_n20), .A2(maj_188_n19), .ZN(maj_188_n26)
         );
  NAND2_X1 maj_188_U3 ( .A1(maj_188_n26), .A2(maj_188_n25), .ZN(maj_188_port_o) );
  XOR2_X1 maj_188_U2 ( .A(maj_188_n22), .B(maj_188_n21), .Z(maj_188_n23) );
  NAND2_X1 maj_189_U15 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_189_n18) );
  NAND2_X1 maj_189_U14 ( .A1(maj_189_n21), .A2(maj_189_n22), .ZN(maj_189_n17)
         );
  NAND2_X1 maj_189_U13 ( .A1(maj_189_n18), .A2(maj_189_n17), .ZN(maj_189_n19)
         );
  NAND2_X1 maj_189_U12 ( .A1(v_3_1[2]), .A2(maj_189_n16), .ZN(maj_189_n14) );
  NAND2_X1 maj_189_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_189_n15) );
  NAND2_X1 maj_189_U10 ( .A1(maj_189_n15), .A2(maj_189_n14), .ZN(maj_189_n20)
         );
  XOR2_X1 maj_189_U9 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_189_n22) );
  XOR2_X1 maj_189_U8 ( .A(v_3_1[2]), .B(maj_189_n16), .Z(maj_189_n21) );
  XOR2_X1 maj_189_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_189_n16) );
  OR2_X1 maj_189_U6 ( .A1(maj_189_n20), .A2(maj_189_n19), .ZN(maj_189_n24) );
  NAND2_X1 maj_189_U5 ( .A1(maj_189_n24), .A2(maj_189_n23), .ZN(maj_189_n25)
         );
  NAND2_X1 maj_189_U4 ( .A1(maj_189_n20), .A2(maj_189_n19), .ZN(maj_189_n26)
         );
  NAND2_X1 maj_189_U3 ( .A1(maj_189_n26), .A2(maj_189_n25), .ZN(maj_189_port_o) );
  XOR2_X1 maj_189_U2 ( .A(maj_189_n22), .B(maj_189_n21), .Z(maj_189_n23) );
  NAND2_X1 maj_190_U15 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_190_n18) );
  NAND2_X1 maj_190_U14 ( .A1(maj_190_n21), .A2(maj_190_n22), .ZN(maj_190_n17)
         );
  NAND2_X1 maj_190_U13 ( .A1(maj_190_n18), .A2(maj_190_n17), .ZN(maj_190_n19)
         );
  NAND2_X1 maj_190_U12 ( .A1(u_3_2[2]), .A2(maj_190_n16), .ZN(maj_190_n14) );
  NAND2_X1 maj_190_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_190_n15) );
  NAND2_X1 maj_190_U10 ( .A1(maj_190_n15), .A2(maj_190_n14), .ZN(maj_190_n20)
         );
  XOR2_X1 maj_190_U9 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_190_n22) );
  XOR2_X1 maj_190_U8 ( .A(u_3_2[2]), .B(maj_190_n16), .Z(maj_190_n21) );
  XOR2_X1 maj_190_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_190_n16) );
  OR2_X1 maj_190_U6 ( .A1(maj_190_n20), .A2(maj_190_n19), .ZN(maj_190_n24) );
  NAND2_X1 maj_190_U5 ( .A1(maj_190_n24), .A2(maj_190_n23), .ZN(maj_190_n25)
         );
  NAND2_X1 maj_190_U4 ( .A1(maj_190_n20), .A2(maj_190_n19), .ZN(maj_190_n26)
         );
  NAND2_X1 maj_190_U3 ( .A1(maj_190_n26), .A2(maj_190_n25), .ZN(maj_190_port_o) );
  XOR2_X1 maj_190_U2 ( .A(maj_190_n22), .B(maj_190_n21), .Z(maj_190_n23) );
  NAND2_X1 maj_191_U15 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_191_n18) );
  NAND2_X1 maj_191_U14 ( .A1(maj_191_n21), .A2(maj_191_n22), .ZN(maj_191_n17)
         );
  NAND2_X1 maj_191_U13 ( .A1(maj_191_n18), .A2(maj_191_n17), .ZN(maj_191_n19)
         );
  NAND2_X1 maj_191_U12 ( .A1(v_3_2[2]), .A2(maj_191_n16), .ZN(maj_191_n14) );
  NAND2_X1 maj_191_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_191_n15) );
  NAND2_X1 maj_191_U10 ( .A1(maj_191_n15), .A2(maj_191_n14), .ZN(maj_191_n20)
         );
  XOR2_X1 maj_191_U9 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_191_n22) );
  XOR2_X1 maj_191_U8 ( .A(v_3_2[2]), .B(maj_191_n16), .Z(maj_191_n21) );
  XOR2_X1 maj_191_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_191_n16) );
  OR2_X1 maj_191_U6 ( .A1(maj_191_n20), .A2(maj_191_n19), .ZN(maj_191_n24) );
  NAND2_X1 maj_191_U5 ( .A1(maj_191_n24), .A2(maj_191_n23), .ZN(maj_191_n25)
         );
  NAND2_X1 maj_191_U4 ( .A1(maj_191_n20), .A2(maj_191_n19), .ZN(maj_191_n26)
         );
  NAND2_X1 maj_191_U3 ( .A1(maj_191_n26), .A2(maj_191_n25), .ZN(maj_191_port_o) );
  XOR2_X1 maj_191_U2 ( .A(maj_191_n22), .B(maj_191_n21), .Z(maj_191_n23) );
  NAND2_X1 maj_192_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_192_n18) );
  NAND2_X1 maj_192_U14 ( .A1(maj_192_n21), .A2(maj_192_n22), .ZN(maj_192_n17)
         );
  NAND2_X1 maj_192_U13 ( .A1(maj_192_n18), .A2(maj_192_n17), .ZN(maj_192_n19)
         );
  NAND2_X1 maj_192_U12 ( .A1(u_0_0[2]), .A2(maj_192_n16), .ZN(maj_192_n14) );
  NAND2_X1 maj_192_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_192_n15) );
  NAND2_X1 maj_192_U10 ( .A1(maj_192_n15), .A2(maj_192_n14), .ZN(maj_192_n20)
         );
  XOR2_X1 maj_192_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_192_n22) );
  XOR2_X1 maj_192_U8 ( .A(u_0_0[2]), .B(maj_192_n16), .Z(maj_192_n21) );
  XOR2_X1 maj_192_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_192_n16) );
  OR2_X1 maj_192_U6 ( .A1(maj_192_n20), .A2(maj_192_n19), .ZN(maj_192_n24) );
  NAND2_X1 maj_192_U5 ( .A1(maj_192_n24), .A2(maj_192_n23), .ZN(maj_192_n25)
         );
  NAND2_X1 maj_192_U4 ( .A1(maj_192_n20), .A2(maj_192_n19), .ZN(maj_192_n26)
         );
  NAND2_X1 maj_192_U3 ( .A1(maj_192_n26), .A2(maj_192_n25), .ZN(maj_192_port_o) );
  XOR2_X1 maj_192_U2 ( .A(maj_192_n22), .B(maj_192_n21), .Z(maj_192_n23) );
  NAND2_X1 maj_193_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_193_n18) );
  NAND2_X1 maj_193_U14 ( .A1(maj_193_n21), .A2(maj_193_n22), .ZN(maj_193_n17)
         );
  NAND2_X1 maj_193_U13 ( .A1(maj_193_n18), .A2(maj_193_n17), .ZN(maj_193_n19)
         );
  NAND2_X1 maj_193_U12 ( .A1(v_0_0[2]), .A2(maj_193_n16), .ZN(maj_193_n14) );
  NAND2_X1 maj_193_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_193_n15) );
  NAND2_X1 maj_193_U10 ( .A1(maj_193_n15), .A2(maj_193_n14), .ZN(maj_193_n20)
         );
  XOR2_X1 maj_193_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_193_n22) );
  XOR2_X1 maj_193_U8 ( .A(v_0_0[2]), .B(maj_193_n16), .Z(maj_193_n21) );
  XOR2_X1 maj_193_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_193_n16) );
  OR2_X1 maj_193_U6 ( .A1(maj_193_n20), .A2(maj_193_n19), .ZN(maj_193_n24) );
  NAND2_X1 maj_193_U5 ( .A1(maj_193_n24), .A2(maj_193_n23), .ZN(maj_193_n25)
         );
  NAND2_X1 maj_193_U4 ( .A1(maj_193_n20), .A2(maj_193_n19), .ZN(maj_193_n26)
         );
  NAND2_X1 maj_193_U3 ( .A1(maj_193_n26), .A2(maj_193_n25), .ZN(maj_193_port_o) );
  XOR2_X1 maj_193_U2 ( .A(maj_193_n22), .B(maj_193_n21), .Z(maj_193_n23) );
  NAND2_X1 maj_194_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_194_n18) );
  NAND2_X1 maj_194_U14 ( .A1(maj_194_n21), .A2(maj_194_n22), .ZN(maj_194_n17)
         );
  NAND2_X1 maj_194_U13 ( .A1(maj_194_n18), .A2(maj_194_n17), .ZN(maj_194_n19)
         );
  NAND2_X1 maj_194_U12 ( .A1(u_0_1[2]), .A2(maj_194_n16), .ZN(maj_194_n14) );
  NAND2_X1 maj_194_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_194_n15) );
  NAND2_X1 maj_194_U10 ( .A1(maj_194_n15), .A2(maj_194_n14), .ZN(maj_194_n20)
         );
  XOR2_X1 maj_194_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_194_n22) );
  XOR2_X1 maj_194_U8 ( .A(u_0_1[2]), .B(maj_194_n16), .Z(maj_194_n21) );
  XOR2_X1 maj_194_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_194_n16) );
  OR2_X1 maj_194_U6 ( .A1(maj_194_n20), .A2(maj_194_n19), .ZN(maj_194_n24) );
  NAND2_X1 maj_194_U5 ( .A1(maj_194_n24), .A2(maj_194_n23), .ZN(maj_194_n25)
         );
  NAND2_X1 maj_194_U4 ( .A1(maj_194_n20), .A2(maj_194_n19), .ZN(maj_194_n26)
         );
  NAND2_X1 maj_194_U3 ( .A1(maj_194_n26), .A2(maj_194_n25), .ZN(maj_194_port_o) );
  XOR2_X1 maj_194_U2 ( .A(maj_194_n22), .B(maj_194_n21), .Z(maj_194_n23) );
  NAND2_X1 maj_195_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_195_n18) );
  NAND2_X1 maj_195_U14 ( .A1(maj_195_n21), .A2(maj_195_n22), .ZN(maj_195_n17)
         );
  NAND2_X1 maj_195_U13 ( .A1(maj_195_n18), .A2(maj_195_n17), .ZN(maj_195_n19)
         );
  NAND2_X1 maj_195_U12 ( .A1(v_0_1[2]), .A2(maj_195_n16), .ZN(maj_195_n14) );
  NAND2_X1 maj_195_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_195_n15) );
  NAND2_X1 maj_195_U10 ( .A1(maj_195_n15), .A2(maj_195_n14), .ZN(maj_195_n20)
         );
  XOR2_X1 maj_195_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_195_n22) );
  XOR2_X1 maj_195_U8 ( .A(v_0_1[2]), .B(maj_195_n16), .Z(maj_195_n21) );
  XOR2_X1 maj_195_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_195_n16) );
  OR2_X1 maj_195_U6 ( .A1(maj_195_n20), .A2(maj_195_n19), .ZN(maj_195_n24) );
  NAND2_X1 maj_195_U5 ( .A1(maj_195_n24), .A2(maj_195_n23), .ZN(maj_195_n25)
         );
  NAND2_X1 maj_195_U4 ( .A1(maj_195_n20), .A2(maj_195_n19), .ZN(maj_195_n26)
         );
  NAND2_X1 maj_195_U3 ( .A1(maj_195_n26), .A2(maj_195_n25), .ZN(maj_195_port_o) );
  XOR2_X1 maj_195_U2 ( .A(maj_195_n22), .B(maj_195_n21), .Z(maj_195_n23) );
  NAND2_X1 maj_196_U15 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_196_n18) );
  NAND2_X1 maj_196_U14 ( .A1(maj_196_n21), .A2(maj_196_n22), .ZN(maj_196_n17)
         );
  NAND2_X1 maj_196_U13 ( .A1(maj_196_n18), .A2(maj_196_n17), .ZN(maj_196_n19)
         );
  NAND2_X1 maj_196_U12 ( .A1(u_0_2[2]), .A2(maj_196_n16), .ZN(maj_196_n14) );
  NAND2_X1 maj_196_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_196_n15) );
  NAND2_X1 maj_196_U10 ( .A1(maj_196_n15), .A2(maj_196_n14), .ZN(maj_196_n20)
         );
  XOR2_X1 maj_196_U9 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_196_n22) );
  XOR2_X1 maj_196_U8 ( .A(u_0_2[2]), .B(maj_196_n16), .Z(maj_196_n21) );
  XOR2_X1 maj_196_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_196_n16) );
  OR2_X1 maj_196_U6 ( .A1(maj_196_n20), .A2(maj_196_n19), .ZN(maj_196_n24) );
  NAND2_X1 maj_196_U5 ( .A1(maj_196_n24), .A2(maj_196_n23), .ZN(maj_196_n25)
         );
  NAND2_X1 maj_196_U4 ( .A1(maj_196_n20), .A2(maj_196_n19), .ZN(maj_196_n26)
         );
  NAND2_X1 maj_196_U3 ( .A1(maj_196_n26), .A2(maj_196_n25), .ZN(maj_196_port_o) );
  XOR2_X1 maj_196_U2 ( .A(maj_196_n22), .B(maj_196_n21), .Z(maj_196_n23) );
  NAND2_X1 maj_197_U15 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_197_n18) );
  NAND2_X1 maj_197_U14 ( .A1(maj_197_n21), .A2(maj_197_n22), .ZN(maj_197_n17)
         );
  NAND2_X1 maj_197_U13 ( .A1(maj_197_n18), .A2(maj_197_n17), .ZN(maj_197_n19)
         );
  NAND2_X1 maj_197_U12 ( .A1(v_0_2[2]), .A2(maj_197_n16), .ZN(maj_197_n14) );
  NAND2_X1 maj_197_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_197_n15) );
  NAND2_X1 maj_197_U10 ( .A1(maj_197_n15), .A2(maj_197_n14), .ZN(maj_197_n20)
         );
  XOR2_X1 maj_197_U9 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_197_n22) );
  XOR2_X1 maj_197_U8 ( .A(v_0_2[2]), .B(maj_197_n16), .Z(maj_197_n21) );
  XOR2_X1 maj_197_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_197_n16) );
  OR2_X1 maj_197_U6 ( .A1(maj_197_n20), .A2(maj_197_n19), .ZN(maj_197_n24) );
  NAND2_X1 maj_197_U5 ( .A1(maj_197_n24), .A2(maj_197_n23), .ZN(maj_197_n25)
         );
  NAND2_X1 maj_197_U4 ( .A1(maj_197_n20), .A2(maj_197_n19), .ZN(maj_197_n26)
         );
  NAND2_X1 maj_197_U3 ( .A1(maj_197_n26), .A2(maj_197_n25), .ZN(maj_197_port_o) );
  XOR2_X1 maj_197_U2 ( .A(maj_197_n22), .B(maj_197_n21), .Z(maj_197_n23) );
  NAND2_X1 maj_198_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_198_n18) );
  NAND2_X1 maj_198_U14 ( .A1(maj_198_n21), .A2(maj_198_n22), .ZN(maj_198_n17)
         );
  NAND2_X1 maj_198_U13 ( .A1(maj_198_n18), .A2(maj_198_n17), .ZN(maj_198_n19)
         );
  NAND2_X1 maj_198_U12 ( .A1(u_1_0[2]), .A2(maj_198_n16), .ZN(maj_198_n14) );
  NAND2_X1 maj_198_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_198_n15) );
  NAND2_X1 maj_198_U10 ( .A1(maj_198_n15), .A2(maj_198_n14), .ZN(maj_198_n20)
         );
  XOR2_X1 maj_198_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_198_n22) );
  XOR2_X1 maj_198_U8 ( .A(u_1_0[2]), .B(maj_198_n16), .Z(maj_198_n21) );
  XOR2_X1 maj_198_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_198_n16) );
  OR2_X1 maj_198_U6 ( .A1(maj_198_n20), .A2(maj_198_n19), .ZN(maj_198_n24) );
  NAND2_X1 maj_198_U5 ( .A1(maj_198_n24), .A2(maj_198_n23), .ZN(maj_198_n25)
         );
  NAND2_X1 maj_198_U4 ( .A1(maj_198_n20), .A2(maj_198_n19), .ZN(maj_198_n26)
         );
  NAND2_X1 maj_198_U3 ( .A1(maj_198_n26), .A2(maj_198_n25), .ZN(maj_198_port_o) );
  XOR2_X1 maj_198_U2 ( .A(maj_198_n22), .B(maj_198_n21), .Z(maj_198_n23) );
  NAND2_X1 maj_199_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_199_n18) );
  NAND2_X1 maj_199_U14 ( .A1(maj_199_n21), .A2(maj_199_n22), .ZN(maj_199_n17)
         );
  NAND2_X1 maj_199_U13 ( .A1(maj_199_n18), .A2(maj_199_n17), .ZN(maj_199_n19)
         );
  NAND2_X1 maj_199_U12 ( .A1(v_1_0[2]), .A2(maj_199_n16), .ZN(maj_199_n14) );
  NAND2_X1 maj_199_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_199_n15) );
  NAND2_X1 maj_199_U10 ( .A1(maj_199_n15), .A2(maj_199_n14), .ZN(maj_199_n20)
         );
  XOR2_X1 maj_199_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_199_n22) );
  XOR2_X1 maj_199_U8 ( .A(v_1_0[2]), .B(maj_199_n16), .Z(maj_199_n21) );
  XOR2_X1 maj_199_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_199_n16) );
  OR2_X1 maj_199_U6 ( .A1(maj_199_n20), .A2(maj_199_n19), .ZN(maj_199_n24) );
  NAND2_X1 maj_199_U5 ( .A1(maj_199_n24), .A2(maj_199_n23), .ZN(maj_199_n25)
         );
  NAND2_X1 maj_199_U4 ( .A1(maj_199_n20), .A2(maj_199_n19), .ZN(maj_199_n26)
         );
  NAND2_X1 maj_199_U3 ( .A1(maj_199_n26), .A2(maj_199_n25), .ZN(maj_199_port_o) );
  XOR2_X1 maj_199_U2 ( .A(maj_199_n22), .B(maj_199_n21), .Z(maj_199_n23) );
  NAND2_X1 maj_200_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_200_n18) );
  NAND2_X1 maj_200_U14 ( .A1(maj_200_n21), .A2(maj_200_n22), .ZN(maj_200_n17)
         );
  NAND2_X1 maj_200_U13 ( .A1(maj_200_n18), .A2(maj_200_n17), .ZN(maj_200_n19)
         );
  NAND2_X1 maj_200_U12 ( .A1(u_1_1[2]), .A2(maj_200_n16), .ZN(maj_200_n14) );
  NAND2_X1 maj_200_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_200_n15) );
  NAND2_X1 maj_200_U10 ( .A1(maj_200_n15), .A2(maj_200_n14), .ZN(maj_200_n20)
         );
  XOR2_X1 maj_200_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_200_n22) );
  XOR2_X1 maj_200_U8 ( .A(u_1_1[2]), .B(maj_200_n16), .Z(maj_200_n21) );
  XOR2_X1 maj_200_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_200_n16) );
  OR2_X1 maj_200_U6 ( .A1(maj_200_n20), .A2(maj_200_n19), .ZN(maj_200_n24) );
  NAND2_X1 maj_200_U5 ( .A1(maj_200_n24), .A2(maj_200_n23), .ZN(maj_200_n25)
         );
  NAND2_X1 maj_200_U4 ( .A1(maj_200_n20), .A2(maj_200_n19), .ZN(maj_200_n26)
         );
  NAND2_X1 maj_200_U3 ( .A1(maj_200_n26), .A2(maj_200_n25), .ZN(maj_200_port_o) );
  XOR2_X1 maj_200_U2 ( .A(maj_200_n22), .B(maj_200_n21), .Z(maj_200_n23) );
  NAND2_X1 maj_201_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_201_n18) );
  NAND2_X1 maj_201_U14 ( .A1(maj_201_n21), .A2(maj_201_n22), .ZN(maj_201_n17)
         );
  NAND2_X1 maj_201_U13 ( .A1(maj_201_n18), .A2(maj_201_n17), .ZN(maj_201_n19)
         );
  NAND2_X1 maj_201_U12 ( .A1(v_1_1[2]), .A2(maj_201_n16), .ZN(maj_201_n14) );
  NAND2_X1 maj_201_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_201_n15) );
  NAND2_X1 maj_201_U10 ( .A1(maj_201_n15), .A2(maj_201_n14), .ZN(maj_201_n20)
         );
  XOR2_X1 maj_201_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_201_n22) );
  XOR2_X1 maj_201_U8 ( .A(v_1_1[2]), .B(maj_201_n16), .Z(maj_201_n21) );
  XOR2_X1 maj_201_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_201_n16) );
  OR2_X1 maj_201_U6 ( .A1(maj_201_n20), .A2(maj_201_n19), .ZN(maj_201_n24) );
  NAND2_X1 maj_201_U5 ( .A1(maj_201_n24), .A2(maj_201_n23), .ZN(maj_201_n25)
         );
  NAND2_X1 maj_201_U4 ( .A1(maj_201_n20), .A2(maj_201_n19), .ZN(maj_201_n26)
         );
  NAND2_X1 maj_201_U3 ( .A1(maj_201_n26), .A2(maj_201_n25), .ZN(maj_201_port_o) );
  XOR2_X1 maj_201_U2 ( .A(maj_201_n22), .B(maj_201_n21), .Z(maj_201_n23) );
  NAND2_X1 maj_202_U15 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_202_n18) );
  NAND2_X1 maj_202_U14 ( .A1(maj_202_n21), .A2(maj_202_n22), .ZN(maj_202_n17)
         );
  NAND2_X1 maj_202_U13 ( .A1(maj_202_n18), .A2(maj_202_n17), .ZN(maj_202_n19)
         );
  NAND2_X1 maj_202_U12 ( .A1(u_1_2[2]), .A2(maj_202_n16), .ZN(maj_202_n14) );
  NAND2_X1 maj_202_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_202_n15) );
  NAND2_X1 maj_202_U10 ( .A1(maj_202_n15), .A2(maj_202_n14), .ZN(maj_202_n20)
         );
  XOR2_X1 maj_202_U9 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_202_n22) );
  XOR2_X1 maj_202_U8 ( .A(u_1_2[2]), .B(maj_202_n16), .Z(maj_202_n21) );
  XOR2_X1 maj_202_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_202_n16) );
  OR2_X1 maj_202_U6 ( .A1(maj_202_n20), .A2(maj_202_n19), .ZN(maj_202_n24) );
  NAND2_X1 maj_202_U5 ( .A1(maj_202_n24), .A2(maj_202_n23), .ZN(maj_202_n25)
         );
  NAND2_X1 maj_202_U4 ( .A1(maj_202_n20), .A2(maj_202_n19), .ZN(maj_202_n26)
         );
  NAND2_X1 maj_202_U3 ( .A1(maj_202_n26), .A2(maj_202_n25), .ZN(maj_202_port_o) );
  XOR2_X1 maj_202_U2 ( .A(maj_202_n22), .B(maj_202_n21), .Z(maj_202_n23) );
  NAND2_X1 maj_203_U15 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_203_n18) );
  NAND2_X1 maj_203_U14 ( .A1(maj_203_n21), .A2(maj_203_n22), .ZN(maj_203_n17)
         );
  NAND2_X1 maj_203_U13 ( .A1(maj_203_n18), .A2(maj_203_n17), .ZN(maj_203_n19)
         );
  NAND2_X1 maj_203_U12 ( .A1(v_1_2[2]), .A2(maj_203_n16), .ZN(maj_203_n14) );
  NAND2_X1 maj_203_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_203_n15) );
  NAND2_X1 maj_203_U10 ( .A1(maj_203_n15), .A2(maj_203_n14), .ZN(maj_203_n20)
         );
  XOR2_X1 maj_203_U9 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_203_n22) );
  XOR2_X1 maj_203_U8 ( .A(v_1_2[2]), .B(maj_203_n16), .Z(maj_203_n21) );
  XOR2_X1 maj_203_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_203_n16) );
  OR2_X1 maj_203_U6 ( .A1(maj_203_n20), .A2(maj_203_n19), .ZN(maj_203_n24) );
  NAND2_X1 maj_203_U5 ( .A1(maj_203_n24), .A2(maj_203_n23), .ZN(maj_203_n25)
         );
  NAND2_X1 maj_203_U4 ( .A1(maj_203_n20), .A2(maj_203_n19), .ZN(maj_203_n26)
         );
  NAND2_X1 maj_203_U3 ( .A1(maj_203_n26), .A2(maj_203_n25), .ZN(maj_203_port_o) );
  XOR2_X1 maj_203_U2 ( .A(maj_203_n22), .B(maj_203_n21), .Z(maj_203_n23) );
  NAND2_X1 maj_204_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_204_n18) );
  NAND2_X1 maj_204_U14 ( .A1(maj_204_n21), .A2(maj_204_n22), .ZN(maj_204_n17)
         );
  NAND2_X1 maj_204_U13 ( .A1(maj_204_n18), .A2(maj_204_n17), .ZN(maj_204_n19)
         );
  NAND2_X1 maj_204_U12 ( .A1(u_2_0[2]), .A2(maj_204_n16), .ZN(maj_204_n14) );
  NAND2_X1 maj_204_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_204_n15) );
  NAND2_X1 maj_204_U10 ( .A1(maj_204_n15), .A2(maj_204_n14), .ZN(maj_204_n20)
         );
  XOR2_X1 maj_204_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_204_n22) );
  XOR2_X1 maj_204_U8 ( .A(u_2_0[2]), .B(maj_204_n16), .Z(maj_204_n21) );
  XOR2_X1 maj_204_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_204_n16) );
  OR2_X1 maj_204_U6 ( .A1(maj_204_n20), .A2(maj_204_n19), .ZN(maj_204_n24) );
  NAND2_X1 maj_204_U5 ( .A1(maj_204_n24), .A2(maj_204_n23), .ZN(maj_204_n25)
         );
  NAND2_X1 maj_204_U4 ( .A1(maj_204_n20), .A2(maj_204_n19), .ZN(maj_204_n26)
         );
  NAND2_X1 maj_204_U3 ( .A1(maj_204_n26), .A2(maj_204_n25), .ZN(maj_204_port_o) );
  XOR2_X1 maj_204_U2 ( .A(maj_204_n22), .B(maj_204_n21), .Z(maj_204_n23) );
  NAND2_X1 maj_205_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_205_n18) );
  NAND2_X1 maj_205_U14 ( .A1(maj_205_n21), .A2(maj_205_n22), .ZN(maj_205_n17)
         );
  NAND2_X1 maj_205_U13 ( .A1(maj_205_n18), .A2(maj_205_n17), .ZN(maj_205_n19)
         );
  NAND2_X1 maj_205_U12 ( .A1(v_2_0[2]), .A2(maj_205_n16), .ZN(maj_205_n14) );
  NAND2_X1 maj_205_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_205_n15) );
  NAND2_X1 maj_205_U10 ( .A1(maj_205_n15), .A2(maj_205_n14), .ZN(maj_205_n20)
         );
  XOR2_X1 maj_205_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_205_n22) );
  XOR2_X1 maj_205_U8 ( .A(v_2_0[2]), .B(maj_205_n16), .Z(maj_205_n21) );
  XOR2_X1 maj_205_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_205_n16) );
  OR2_X1 maj_205_U6 ( .A1(maj_205_n20), .A2(maj_205_n19), .ZN(maj_205_n24) );
  NAND2_X1 maj_205_U5 ( .A1(maj_205_n24), .A2(maj_205_n23), .ZN(maj_205_n25)
         );
  NAND2_X1 maj_205_U4 ( .A1(maj_205_n20), .A2(maj_205_n19), .ZN(maj_205_n26)
         );
  NAND2_X1 maj_205_U3 ( .A1(maj_205_n26), .A2(maj_205_n25), .ZN(maj_205_port_o) );
  XOR2_X1 maj_205_U2 ( .A(maj_205_n22), .B(maj_205_n21), .Z(maj_205_n23) );
  NAND2_X1 maj_206_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_206_n18) );
  NAND2_X1 maj_206_U14 ( .A1(maj_206_n21), .A2(maj_206_n22), .ZN(maj_206_n17)
         );
  NAND2_X1 maj_206_U13 ( .A1(maj_206_n18), .A2(maj_206_n17), .ZN(maj_206_n19)
         );
  NAND2_X1 maj_206_U12 ( .A1(u_2_1[2]), .A2(maj_206_n16), .ZN(maj_206_n14) );
  NAND2_X1 maj_206_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_206_n15) );
  NAND2_X1 maj_206_U10 ( .A1(maj_206_n15), .A2(maj_206_n14), .ZN(maj_206_n20)
         );
  XOR2_X1 maj_206_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_206_n22) );
  XOR2_X1 maj_206_U8 ( .A(u_2_1[2]), .B(maj_206_n16), .Z(maj_206_n21) );
  XOR2_X1 maj_206_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_206_n16) );
  OR2_X1 maj_206_U6 ( .A1(maj_206_n20), .A2(maj_206_n19), .ZN(maj_206_n24) );
  NAND2_X1 maj_206_U5 ( .A1(maj_206_n24), .A2(maj_206_n23), .ZN(maj_206_n25)
         );
  NAND2_X1 maj_206_U4 ( .A1(maj_206_n20), .A2(maj_206_n19), .ZN(maj_206_n26)
         );
  NAND2_X1 maj_206_U3 ( .A1(maj_206_n26), .A2(maj_206_n25), .ZN(maj_206_port_o) );
  XOR2_X1 maj_206_U2 ( .A(maj_206_n22), .B(maj_206_n21), .Z(maj_206_n23) );
  NAND2_X1 maj_207_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_207_n18) );
  NAND2_X1 maj_207_U14 ( .A1(maj_207_n21), .A2(maj_207_n22), .ZN(maj_207_n17)
         );
  NAND2_X1 maj_207_U13 ( .A1(maj_207_n18), .A2(maj_207_n17), .ZN(maj_207_n19)
         );
  NAND2_X1 maj_207_U12 ( .A1(v_2_1[2]), .A2(maj_207_n16), .ZN(maj_207_n14) );
  NAND2_X1 maj_207_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_207_n15) );
  NAND2_X1 maj_207_U10 ( .A1(maj_207_n15), .A2(maj_207_n14), .ZN(maj_207_n20)
         );
  XOR2_X1 maj_207_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_207_n22) );
  XOR2_X1 maj_207_U8 ( .A(v_2_1[2]), .B(maj_207_n16), .Z(maj_207_n21) );
  XOR2_X1 maj_207_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_207_n16) );
  OR2_X1 maj_207_U6 ( .A1(maj_207_n20), .A2(maj_207_n19), .ZN(maj_207_n24) );
  NAND2_X1 maj_207_U5 ( .A1(maj_207_n24), .A2(maj_207_n23), .ZN(maj_207_n25)
         );
  NAND2_X1 maj_207_U4 ( .A1(maj_207_n20), .A2(maj_207_n19), .ZN(maj_207_n26)
         );
  NAND2_X1 maj_207_U3 ( .A1(maj_207_n26), .A2(maj_207_n25), .ZN(maj_207_port_o) );
  XOR2_X1 maj_207_U2 ( .A(maj_207_n22), .B(maj_207_n21), .Z(maj_207_n23) );
  NAND2_X1 maj_208_U15 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_208_n18) );
  NAND2_X1 maj_208_U14 ( .A1(maj_208_n21), .A2(maj_208_n22), .ZN(maj_208_n17)
         );
  NAND2_X1 maj_208_U13 ( .A1(maj_208_n18), .A2(maj_208_n17), .ZN(maj_208_n19)
         );
  NAND2_X1 maj_208_U12 ( .A1(u_2_2[2]), .A2(maj_208_n16), .ZN(maj_208_n14) );
  NAND2_X1 maj_208_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_208_n15) );
  NAND2_X1 maj_208_U10 ( .A1(maj_208_n15), .A2(maj_208_n14), .ZN(maj_208_n20)
         );
  XOR2_X1 maj_208_U9 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_208_n22) );
  XOR2_X1 maj_208_U8 ( .A(u_2_2[2]), .B(maj_208_n16), .Z(maj_208_n21) );
  XOR2_X1 maj_208_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_208_n16) );
  OR2_X1 maj_208_U6 ( .A1(maj_208_n20), .A2(maj_208_n19), .ZN(maj_208_n24) );
  NAND2_X1 maj_208_U5 ( .A1(maj_208_n24), .A2(maj_208_n23), .ZN(maj_208_n25)
         );
  NAND2_X1 maj_208_U4 ( .A1(maj_208_n20), .A2(maj_208_n19), .ZN(maj_208_n26)
         );
  NAND2_X1 maj_208_U3 ( .A1(maj_208_n26), .A2(maj_208_n25), .ZN(maj_208_port_o) );
  XOR2_X1 maj_208_U2 ( .A(maj_208_n22), .B(maj_208_n21), .Z(maj_208_n23) );
  NAND2_X1 maj_209_U15 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_209_n18) );
  NAND2_X1 maj_209_U14 ( .A1(maj_209_n21), .A2(maj_209_n22), .ZN(maj_209_n17)
         );
  NAND2_X1 maj_209_U13 ( .A1(maj_209_n18), .A2(maj_209_n17), .ZN(maj_209_n19)
         );
  NAND2_X1 maj_209_U12 ( .A1(v_2_2[2]), .A2(maj_209_n16), .ZN(maj_209_n14) );
  NAND2_X1 maj_209_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_209_n15) );
  NAND2_X1 maj_209_U10 ( .A1(maj_209_n15), .A2(maj_209_n14), .ZN(maj_209_n20)
         );
  XOR2_X1 maj_209_U9 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_209_n22) );
  XOR2_X1 maj_209_U8 ( .A(v_2_2[2]), .B(maj_209_n16), .Z(maj_209_n21) );
  XOR2_X1 maj_209_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_209_n16) );
  OR2_X1 maj_209_U6 ( .A1(maj_209_n20), .A2(maj_209_n19), .ZN(maj_209_n24) );
  NAND2_X1 maj_209_U5 ( .A1(maj_209_n24), .A2(maj_209_n23), .ZN(maj_209_n25)
         );
  NAND2_X1 maj_209_U4 ( .A1(maj_209_n20), .A2(maj_209_n19), .ZN(maj_209_n26)
         );
  NAND2_X1 maj_209_U3 ( .A1(maj_209_n26), .A2(maj_209_n25), .ZN(maj_209_port_o) );
  XOR2_X1 maj_209_U2 ( .A(maj_209_n22), .B(maj_209_n21), .Z(maj_209_n23) );
  NAND2_X1 maj_210_U15 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_210_n18) );
  NAND2_X1 maj_210_U14 ( .A1(maj_210_n21), .A2(maj_210_n22), .ZN(maj_210_n17)
         );
  NAND2_X1 maj_210_U13 ( .A1(maj_210_n18), .A2(maj_210_n17), .ZN(maj_210_n19)
         );
  NAND2_X1 maj_210_U12 ( .A1(u_3_0[2]), .A2(maj_210_n16), .ZN(maj_210_n14) );
  NAND2_X1 maj_210_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_210_n15) );
  NAND2_X1 maj_210_U10 ( .A1(maj_210_n15), .A2(maj_210_n14), .ZN(maj_210_n20)
         );
  XOR2_X1 maj_210_U9 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_210_n22) );
  XOR2_X1 maj_210_U8 ( .A(u_3_0[2]), .B(maj_210_n16), .Z(maj_210_n21) );
  XOR2_X1 maj_210_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_210_n16) );
  OR2_X1 maj_210_U6 ( .A1(maj_210_n20), .A2(maj_210_n19), .ZN(maj_210_n24) );
  NAND2_X1 maj_210_U5 ( .A1(maj_210_n24), .A2(maj_210_n23), .ZN(maj_210_n25)
         );
  NAND2_X1 maj_210_U4 ( .A1(maj_210_n20), .A2(maj_210_n19), .ZN(maj_210_n26)
         );
  NAND2_X1 maj_210_U3 ( .A1(maj_210_n26), .A2(maj_210_n25), .ZN(maj_210_port_o) );
  XOR2_X1 maj_210_U2 ( .A(maj_210_n22), .B(maj_210_n21), .Z(maj_210_n23) );
  NAND2_X1 maj_211_U15 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_211_n18) );
  NAND2_X1 maj_211_U14 ( .A1(maj_211_n21), .A2(maj_211_n22), .ZN(maj_211_n17)
         );
  NAND2_X1 maj_211_U13 ( .A1(maj_211_n18), .A2(maj_211_n17), .ZN(maj_211_n19)
         );
  NAND2_X1 maj_211_U12 ( .A1(v_3_0[2]), .A2(maj_211_n16), .ZN(maj_211_n14) );
  NAND2_X1 maj_211_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_211_n15) );
  NAND2_X1 maj_211_U10 ( .A1(maj_211_n15), .A2(maj_211_n14), .ZN(maj_211_n20)
         );
  XOR2_X1 maj_211_U9 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_211_n22) );
  XOR2_X1 maj_211_U8 ( .A(v_3_0[2]), .B(maj_211_n16), .Z(maj_211_n21) );
  XOR2_X1 maj_211_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_211_n16) );
  OR2_X1 maj_211_U6 ( .A1(maj_211_n20), .A2(maj_211_n19), .ZN(maj_211_n24) );
  NAND2_X1 maj_211_U5 ( .A1(maj_211_n24), .A2(maj_211_n23), .ZN(maj_211_n25)
         );
  NAND2_X1 maj_211_U4 ( .A1(maj_211_n20), .A2(maj_211_n19), .ZN(maj_211_n26)
         );
  NAND2_X1 maj_211_U3 ( .A1(maj_211_n26), .A2(maj_211_n25), .ZN(maj_211_port_o) );
  XOR2_X1 maj_211_U2 ( .A(maj_211_n22), .B(maj_211_n21), .Z(maj_211_n23) );
  NAND2_X1 maj_212_U15 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_212_n18) );
  NAND2_X1 maj_212_U14 ( .A1(maj_212_n21), .A2(maj_212_n22), .ZN(maj_212_n17)
         );
  NAND2_X1 maj_212_U13 ( .A1(maj_212_n18), .A2(maj_212_n17), .ZN(maj_212_n19)
         );
  NAND2_X1 maj_212_U12 ( .A1(u_3_1[2]), .A2(maj_212_n16), .ZN(maj_212_n14) );
  NAND2_X1 maj_212_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_212_n15) );
  NAND2_X1 maj_212_U10 ( .A1(maj_212_n15), .A2(maj_212_n14), .ZN(maj_212_n20)
         );
  XOR2_X1 maj_212_U9 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_212_n22) );
  XOR2_X1 maj_212_U8 ( .A(u_3_1[2]), .B(maj_212_n16), .Z(maj_212_n21) );
  XOR2_X1 maj_212_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_212_n16) );
  OR2_X1 maj_212_U6 ( .A1(maj_212_n20), .A2(maj_212_n19), .ZN(maj_212_n24) );
  NAND2_X1 maj_212_U5 ( .A1(maj_212_n24), .A2(maj_212_n23), .ZN(maj_212_n25)
         );
  NAND2_X1 maj_212_U4 ( .A1(maj_212_n20), .A2(maj_212_n19), .ZN(maj_212_n26)
         );
  NAND2_X1 maj_212_U3 ( .A1(maj_212_n26), .A2(maj_212_n25), .ZN(maj_212_port_o) );
  XOR2_X1 maj_212_U2 ( .A(maj_212_n22), .B(maj_212_n21), .Z(maj_212_n23) );
  NAND2_X1 maj_213_U15 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_213_n18) );
  NAND2_X1 maj_213_U14 ( .A1(maj_213_n21), .A2(maj_213_n22), .ZN(maj_213_n17)
         );
  NAND2_X1 maj_213_U13 ( .A1(maj_213_n18), .A2(maj_213_n17), .ZN(maj_213_n19)
         );
  NAND2_X1 maj_213_U12 ( .A1(v_3_1[2]), .A2(maj_213_n16), .ZN(maj_213_n14) );
  NAND2_X1 maj_213_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_213_n15) );
  NAND2_X1 maj_213_U10 ( .A1(maj_213_n15), .A2(maj_213_n14), .ZN(maj_213_n20)
         );
  XOR2_X1 maj_213_U9 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_213_n22) );
  XOR2_X1 maj_213_U8 ( .A(v_3_1[2]), .B(maj_213_n16), .Z(maj_213_n21) );
  XOR2_X1 maj_213_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_213_n16) );
  OR2_X1 maj_213_U6 ( .A1(maj_213_n20), .A2(maj_213_n19), .ZN(maj_213_n24) );
  NAND2_X1 maj_213_U5 ( .A1(maj_213_n24), .A2(maj_213_n23), .ZN(maj_213_n25)
         );
  NAND2_X1 maj_213_U4 ( .A1(maj_213_n20), .A2(maj_213_n19), .ZN(maj_213_n26)
         );
  NAND2_X1 maj_213_U3 ( .A1(maj_213_n26), .A2(maj_213_n25), .ZN(maj_213_port_o) );
  XOR2_X1 maj_213_U2 ( .A(maj_213_n22), .B(maj_213_n21), .Z(maj_213_n23) );
  NAND2_X1 maj_214_U15 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_214_n18) );
  NAND2_X1 maj_214_U14 ( .A1(maj_214_n21), .A2(maj_214_n22), .ZN(maj_214_n17)
         );
  NAND2_X1 maj_214_U13 ( .A1(maj_214_n18), .A2(maj_214_n17), .ZN(maj_214_n19)
         );
  NAND2_X1 maj_214_U12 ( .A1(u_3_2[2]), .A2(maj_214_n16), .ZN(maj_214_n14) );
  NAND2_X1 maj_214_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_214_n15) );
  NAND2_X1 maj_214_U10 ( .A1(maj_214_n15), .A2(maj_214_n14), .ZN(maj_214_n20)
         );
  XOR2_X1 maj_214_U9 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_214_n22) );
  XOR2_X1 maj_214_U8 ( .A(u_3_2[2]), .B(maj_214_n16), .Z(maj_214_n21) );
  XOR2_X1 maj_214_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_214_n16) );
  OR2_X1 maj_214_U6 ( .A1(maj_214_n20), .A2(maj_214_n19), .ZN(maj_214_n24) );
  NAND2_X1 maj_214_U5 ( .A1(maj_214_n24), .A2(maj_214_n23), .ZN(maj_214_n25)
         );
  NAND2_X1 maj_214_U4 ( .A1(maj_214_n20), .A2(maj_214_n19), .ZN(maj_214_n26)
         );
  NAND2_X1 maj_214_U3 ( .A1(maj_214_n26), .A2(maj_214_n25), .ZN(maj_214_port_o) );
  XOR2_X1 maj_214_U2 ( .A(maj_214_n22), .B(maj_214_n21), .Z(maj_214_n23) );
  NAND2_X1 maj_215_U15 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_215_n18) );
  NAND2_X1 maj_215_U14 ( .A1(maj_215_n21), .A2(maj_215_n22), .ZN(maj_215_n17)
         );
  NAND2_X1 maj_215_U13 ( .A1(maj_215_n18), .A2(maj_215_n17), .ZN(maj_215_n19)
         );
  NAND2_X1 maj_215_U12 ( .A1(v_3_2[2]), .A2(maj_215_n16), .ZN(maj_215_n14) );
  NAND2_X1 maj_215_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_215_n15) );
  NAND2_X1 maj_215_U10 ( .A1(maj_215_n15), .A2(maj_215_n14), .ZN(maj_215_n20)
         );
  XOR2_X1 maj_215_U9 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_215_n22) );
  XOR2_X1 maj_215_U8 ( .A(v_3_2[2]), .B(maj_215_n16), .Z(maj_215_n21) );
  XOR2_X1 maj_215_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_215_n16) );
  OR2_X1 maj_215_U6 ( .A1(maj_215_n20), .A2(maj_215_n19), .ZN(maj_215_n24) );
  NAND2_X1 maj_215_U5 ( .A1(maj_215_n24), .A2(maj_215_n23), .ZN(maj_215_n25)
         );
  NAND2_X1 maj_215_U4 ( .A1(maj_215_n20), .A2(maj_215_n19), .ZN(maj_215_n26)
         );
  NAND2_X1 maj_215_U3 ( .A1(maj_215_n26), .A2(maj_215_n25), .ZN(maj_215_port_o) );
  XOR2_X1 maj_215_U2 ( .A(maj_215_n22), .B(maj_215_n21), .Z(maj_215_n23) );
  NAND2_X1 maj_216_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_216_n18) );
  NAND2_X1 maj_216_U14 ( .A1(maj_216_n21), .A2(maj_216_n22), .ZN(maj_216_n17)
         );
  NAND2_X1 maj_216_U13 ( .A1(maj_216_n18), .A2(maj_216_n17), .ZN(maj_216_n19)
         );
  NAND2_X1 maj_216_U12 ( .A1(u_0_0[2]), .A2(maj_216_n16), .ZN(maj_216_n14) );
  NAND2_X1 maj_216_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_216_n15) );
  NAND2_X1 maj_216_U10 ( .A1(maj_216_n15), .A2(maj_216_n14), .ZN(maj_216_n20)
         );
  XOR2_X1 maj_216_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_216_n22) );
  XOR2_X1 maj_216_U8 ( .A(u_0_0[2]), .B(maj_216_n16), .Z(maj_216_n21) );
  XOR2_X1 maj_216_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_216_n16) );
  OR2_X1 maj_216_U6 ( .A1(maj_216_n20), .A2(maj_216_n19), .ZN(maj_216_n24) );
  NAND2_X1 maj_216_U5 ( .A1(maj_216_n24), .A2(maj_216_n23), .ZN(maj_216_n25)
         );
  NAND2_X1 maj_216_U4 ( .A1(maj_216_n20), .A2(maj_216_n19), .ZN(maj_216_n26)
         );
  NAND2_X1 maj_216_U3 ( .A1(maj_216_n26), .A2(maj_216_n25), .ZN(maj_216_port_o) );
  XOR2_X1 maj_216_U2 ( .A(maj_216_n22), .B(maj_216_n21), .Z(maj_216_n23) );
  NAND2_X1 maj_217_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_217_n18) );
  NAND2_X1 maj_217_U14 ( .A1(maj_217_n21), .A2(maj_217_n22), .ZN(maj_217_n17)
         );
  NAND2_X1 maj_217_U13 ( .A1(maj_217_n18), .A2(maj_217_n17), .ZN(maj_217_n19)
         );
  NAND2_X1 maj_217_U12 ( .A1(v_0_0[2]), .A2(maj_217_n16), .ZN(maj_217_n14) );
  NAND2_X1 maj_217_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_217_n15) );
  NAND2_X1 maj_217_U10 ( .A1(maj_217_n15), .A2(maj_217_n14), .ZN(maj_217_n20)
         );
  XOR2_X1 maj_217_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_217_n22) );
  XOR2_X1 maj_217_U8 ( .A(v_0_0[2]), .B(maj_217_n16), .Z(maj_217_n21) );
  XOR2_X1 maj_217_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_217_n16) );
  OR2_X1 maj_217_U6 ( .A1(maj_217_n20), .A2(maj_217_n19), .ZN(maj_217_n24) );
  NAND2_X1 maj_217_U5 ( .A1(maj_217_n24), .A2(maj_217_n23), .ZN(maj_217_n25)
         );
  NAND2_X1 maj_217_U4 ( .A1(maj_217_n20), .A2(maj_217_n19), .ZN(maj_217_n26)
         );
  NAND2_X1 maj_217_U3 ( .A1(maj_217_n26), .A2(maj_217_n25), .ZN(maj_217_port_o) );
  XOR2_X1 maj_217_U2 ( .A(maj_217_n22), .B(maj_217_n21), .Z(maj_217_n23) );
  NAND2_X1 maj_218_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_218_n18) );
  NAND2_X1 maj_218_U14 ( .A1(maj_218_n21), .A2(maj_218_n22), .ZN(maj_218_n17)
         );
  NAND2_X1 maj_218_U13 ( .A1(maj_218_n18), .A2(maj_218_n17), .ZN(maj_218_n19)
         );
  NAND2_X1 maj_218_U12 ( .A1(u_0_1[2]), .A2(maj_218_n16), .ZN(maj_218_n14) );
  NAND2_X1 maj_218_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_218_n15) );
  NAND2_X1 maj_218_U10 ( .A1(maj_218_n15), .A2(maj_218_n14), .ZN(maj_218_n20)
         );
  XOR2_X1 maj_218_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_218_n22) );
  XOR2_X1 maj_218_U8 ( .A(u_0_1[2]), .B(maj_218_n16), .Z(maj_218_n21) );
  XOR2_X1 maj_218_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_218_n16) );
  OR2_X1 maj_218_U6 ( .A1(maj_218_n20), .A2(maj_218_n19), .ZN(maj_218_n24) );
  NAND2_X1 maj_218_U5 ( .A1(maj_218_n24), .A2(maj_218_n23), .ZN(maj_218_n25)
         );
  NAND2_X1 maj_218_U4 ( .A1(maj_218_n20), .A2(maj_218_n19), .ZN(maj_218_n26)
         );
  NAND2_X1 maj_218_U3 ( .A1(maj_218_n26), .A2(maj_218_n25), .ZN(maj_218_port_o) );
  XOR2_X1 maj_218_U2 ( .A(maj_218_n22), .B(maj_218_n21), .Z(maj_218_n23) );
  NAND2_X1 maj_219_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_219_n18) );
  NAND2_X1 maj_219_U14 ( .A1(maj_219_n21), .A2(maj_219_n22), .ZN(maj_219_n17)
         );
  NAND2_X1 maj_219_U13 ( .A1(maj_219_n18), .A2(maj_219_n17), .ZN(maj_219_n19)
         );
  NAND2_X1 maj_219_U12 ( .A1(v_0_1[2]), .A2(maj_219_n16), .ZN(maj_219_n14) );
  NAND2_X1 maj_219_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_219_n15) );
  NAND2_X1 maj_219_U10 ( .A1(maj_219_n15), .A2(maj_219_n14), .ZN(maj_219_n20)
         );
  XOR2_X1 maj_219_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_219_n22) );
  XOR2_X1 maj_219_U8 ( .A(v_0_1[2]), .B(maj_219_n16), .Z(maj_219_n21) );
  XOR2_X1 maj_219_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_219_n16) );
  OR2_X1 maj_219_U6 ( .A1(maj_219_n20), .A2(maj_219_n19), .ZN(maj_219_n24) );
  NAND2_X1 maj_219_U5 ( .A1(maj_219_n24), .A2(maj_219_n23), .ZN(maj_219_n25)
         );
  NAND2_X1 maj_219_U4 ( .A1(maj_219_n20), .A2(maj_219_n19), .ZN(maj_219_n26)
         );
  NAND2_X1 maj_219_U3 ( .A1(maj_219_n26), .A2(maj_219_n25), .ZN(maj_219_port_o) );
  XOR2_X1 maj_219_U2 ( .A(maj_219_n22), .B(maj_219_n21), .Z(maj_219_n23) );
  NAND2_X1 maj_220_U15 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_220_n18) );
  NAND2_X1 maj_220_U14 ( .A1(maj_220_n21), .A2(maj_220_n22), .ZN(maj_220_n17)
         );
  NAND2_X1 maj_220_U13 ( .A1(maj_220_n18), .A2(maj_220_n17), .ZN(maj_220_n19)
         );
  NAND2_X1 maj_220_U12 ( .A1(u_0_2[2]), .A2(maj_220_n16), .ZN(maj_220_n14) );
  NAND2_X1 maj_220_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_220_n15) );
  NAND2_X1 maj_220_U10 ( .A1(maj_220_n15), .A2(maj_220_n14), .ZN(maj_220_n20)
         );
  XOR2_X1 maj_220_U9 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_220_n22) );
  XOR2_X1 maj_220_U8 ( .A(u_0_2[2]), .B(maj_220_n16), .Z(maj_220_n21) );
  XOR2_X1 maj_220_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_220_n16) );
  OR2_X1 maj_220_U6 ( .A1(maj_220_n20), .A2(maj_220_n19), .ZN(maj_220_n24) );
  NAND2_X1 maj_220_U5 ( .A1(maj_220_n24), .A2(maj_220_n23), .ZN(maj_220_n25)
         );
  NAND2_X1 maj_220_U4 ( .A1(maj_220_n20), .A2(maj_220_n19), .ZN(maj_220_n26)
         );
  NAND2_X1 maj_220_U3 ( .A1(maj_220_n26), .A2(maj_220_n25), .ZN(maj_220_port_o) );
  XOR2_X1 maj_220_U2 ( .A(maj_220_n22), .B(maj_220_n21), .Z(maj_220_n23) );
  NAND2_X1 maj_221_U15 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_221_n18) );
  NAND2_X1 maj_221_U14 ( .A1(maj_221_n21), .A2(maj_221_n22), .ZN(maj_221_n17)
         );
  NAND2_X1 maj_221_U13 ( .A1(maj_221_n18), .A2(maj_221_n17), .ZN(maj_221_n19)
         );
  NAND2_X1 maj_221_U12 ( .A1(v_0_2[2]), .A2(maj_221_n16), .ZN(maj_221_n14) );
  NAND2_X1 maj_221_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_221_n15) );
  NAND2_X1 maj_221_U10 ( .A1(maj_221_n15), .A2(maj_221_n14), .ZN(maj_221_n20)
         );
  XOR2_X1 maj_221_U9 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_221_n22) );
  XOR2_X1 maj_221_U8 ( .A(v_0_2[2]), .B(maj_221_n16), .Z(maj_221_n21) );
  XOR2_X1 maj_221_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_221_n16) );
  OR2_X1 maj_221_U6 ( .A1(maj_221_n20), .A2(maj_221_n19), .ZN(maj_221_n24) );
  NAND2_X1 maj_221_U5 ( .A1(maj_221_n24), .A2(maj_221_n23), .ZN(maj_221_n25)
         );
  NAND2_X1 maj_221_U4 ( .A1(maj_221_n20), .A2(maj_221_n19), .ZN(maj_221_n26)
         );
  NAND2_X1 maj_221_U3 ( .A1(maj_221_n26), .A2(maj_221_n25), .ZN(maj_221_port_o) );
  XOR2_X1 maj_221_U2 ( .A(maj_221_n22), .B(maj_221_n21), .Z(maj_221_n23) );
  NAND2_X1 maj_222_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_222_n18) );
  NAND2_X1 maj_222_U14 ( .A1(maj_222_n21), .A2(maj_222_n22), .ZN(maj_222_n17)
         );
  NAND2_X1 maj_222_U13 ( .A1(maj_222_n18), .A2(maj_222_n17), .ZN(maj_222_n19)
         );
  NAND2_X1 maj_222_U12 ( .A1(u_1_0[2]), .A2(maj_222_n16), .ZN(maj_222_n14) );
  NAND2_X1 maj_222_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_222_n15) );
  NAND2_X1 maj_222_U10 ( .A1(maj_222_n15), .A2(maj_222_n14), .ZN(maj_222_n20)
         );
  XOR2_X1 maj_222_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_222_n22) );
  XOR2_X1 maj_222_U8 ( .A(u_1_0[2]), .B(maj_222_n16), .Z(maj_222_n21) );
  XOR2_X1 maj_222_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_222_n16) );
  OR2_X1 maj_222_U6 ( .A1(maj_222_n20), .A2(maj_222_n19), .ZN(maj_222_n24) );
  NAND2_X1 maj_222_U5 ( .A1(maj_222_n24), .A2(maj_222_n23), .ZN(maj_222_n25)
         );
  NAND2_X1 maj_222_U4 ( .A1(maj_222_n20), .A2(maj_222_n19), .ZN(maj_222_n26)
         );
  NAND2_X1 maj_222_U3 ( .A1(maj_222_n26), .A2(maj_222_n25), .ZN(maj_222_port_o) );
  XOR2_X1 maj_222_U2 ( .A(maj_222_n22), .B(maj_222_n21), .Z(maj_222_n23) );
  NAND2_X1 maj_223_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_223_n18) );
  NAND2_X1 maj_223_U14 ( .A1(maj_223_n21), .A2(maj_223_n22), .ZN(maj_223_n17)
         );
  NAND2_X1 maj_223_U13 ( .A1(maj_223_n18), .A2(maj_223_n17), .ZN(maj_223_n19)
         );
  NAND2_X1 maj_223_U12 ( .A1(v_1_0[2]), .A2(maj_223_n16), .ZN(maj_223_n14) );
  NAND2_X1 maj_223_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_223_n15) );
  NAND2_X1 maj_223_U10 ( .A1(maj_223_n15), .A2(maj_223_n14), .ZN(maj_223_n20)
         );
  XOR2_X1 maj_223_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_223_n22) );
  XOR2_X1 maj_223_U8 ( .A(v_1_0[2]), .B(maj_223_n16), .Z(maj_223_n21) );
  XOR2_X1 maj_223_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_223_n16) );
  OR2_X1 maj_223_U6 ( .A1(maj_223_n20), .A2(maj_223_n19), .ZN(maj_223_n24) );
  NAND2_X1 maj_223_U5 ( .A1(maj_223_n24), .A2(maj_223_n23), .ZN(maj_223_n25)
         );
  NAND2_X1 maj_223_U4 ( .A1(maj_223_n20), .A2(maj_223_n19), .ZN(maj_223_n26)
         );
  NAND2_X1 maj_223_U3 ( .A1(maj_223_n26), .A2(maj_223_n25), .ZN(maj_223_port_o) );
  XOR2_X1 maj_223_U2 ( .A(maj_223_n22), .B(maj_223_n21), .Z(maj_223_n23) );
  NAND2_X1 maj_224_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_224_n18) );
  NAND2_X1 maj_224_U14 ( .A1(maj_224_n21), .A2(maj_224_n22), .ZN(maj_224_n17)
         );
  NAND2_X1 maj_224_U13 ( .A1(maj_224_n18), .A2(maj_224_n17), .ZN(maj_224_n19)
         );
  NAND2_X1 maj_224_U12 ( .A1(u_1_1[2]), .A2(maj_224_n16), .ZN(maj_224_n14) );
  NAND2_X1 maj_224_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_224_n15) );
  NAND2_X1 maj_224_U10 ( .A1(maj_224_n15), .A2(maj_224_n14), .ZN(maj_224_n20)
         );
  XOR2_X1 maj_224_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_224_n22) );
  XOR2_X1 maj_224_U8 ( .A(u_1_1[2]), .B(maj_224_n16), .Z(maj_224_n21) );
  XOR2_X1 maj_224_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_224_n16) );
  OR2_X1 maj_224_U6 ( .A1(maj_224_n20), .A2(maj_224_n19), .ZN(maj_224_n24) );
  NAND2_X1 maj_224_U5 ( .A1(maj_224_n24), .A2(maj_224_n23), .ZN(maj_224_n25)
         );
  NAND2_X1 maj_224_U4 ( .A1(maj_224_n20), .A2(maj_224_n19), .ZN(maj_224_n26)
         );
  NAND2_X1 maj_224_U3 ( .A1(maj_224_n26), .A2(maj_224_n25), .ZN(maj_224_port_o) );
  XOR2_X1 maj_224_U2 ( .A(maj_224_n22), .B(maj_224_n21), .Z(maj_224_n23) );
  NAND2_X1 maj_225_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_225_n18) );
  NAND2_X1 maj_225_U14 ( .A1(maj_225_n21), .A2(maj_225_n22), .ZN(maj_225_n17)
         );
  NAND2_X1 maj_225_U13 ( .A1(maj_225_n18), .A2(maj_225_n17), .ZN(maj_225_n19)
         );
  NAND2_X1 maj_225_U12 ( .A1(v_1_1[2]), .A2(maj_225_n16), .ZN(maj_225_n14) );
  NAND2_X1 maj_225_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_225_n15) );
  NAND2_X1 maj_225_U10 ( .A1(maj_225_n15), .A2(maj_225_n14), .ZN(maj_225_n20)
         );
  XOR2_X1 maj_225_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_225_n22) );
  XOR2_X1 maj_225_U8 ( .A(v_1_1[2]), .B(maj_225_n16), .Z(maj_225_n21) );
  XOR2_X1 maj_225_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_225_n16) );
  OR2_X1 maj_225_U6 ( .A1(maj_225_n20), .A2(maj_225_n19), .ZN(maj_225_n24) );
  NAND2_X1 maj_225_U5 ( .A1(maj_225_n24), .A2(maj_225_n23), .ZN(maj_225_n25)
         );
  NAND2_X1 maj_225_U4 ( .A1(maj_225_n20), .A2(maj_225_n19), .ZN(maj_225_n26)
         );
  NAND2_X1 maj_225_U3 ( .A1(maj_225_n26), .A2(maj_225_n25), .ZN(maj_225_port_o) );
  XOR2_X1 maj_225_U2 ( .A(maj_225_n22), .B(maj_225_n21), .Z(maj_225_n23) );
  NAND2_X1 maj_226_U15 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_226_n18) );
  NAND2_X1 maj_226_U14 ( .A1(maj_226_n21), .A2(maj_226_n22), .ZN(maj_226_n17)
         );
  NAND2_X1 maj_226_U13 ( .A1(maj_226_n18), .A2(maj_226_n17), .ZN(maj_226_n19)
         );
  NAND2_X1 maj_226_U12 ( .A1(u_1_2[2]), .A2(maj_226_n16), .ZN(maj_226_n14) );
  NAND2_X1 maj_226_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_226_n15) );
  NAND2_X1 maj_226_U10 ( .A1(maj_226_n15), .A2(maj_226_n14), .ZN(maj_226_n20)
         );
  XOR2_X1 maj_226_U9 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_226_n22) );
  XOR2_X1 maj_226_U8 ( .A(u_1_2[2]), .B(maj_226_n16), .Z(maj_226_n21) );
  XOR2_X1 maj_226_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_226_n16) );
  OR2_X1 maj_226_U6 ( .A1(maj_226_n20), .A2(maj_226_n19), .ZN(maj_226_n24) );
  NAND2_X1 maj_226_U5 ( .A1(maj_226_n24), .A2(maj_226_n23), .ZN(maj_226_n25)
         );
  NAND2_X1 maj_226_U4 ( .A1(maj_226_n20), .A2(maj_226_n19), .ZN(maj_226_n26)
         );
  NAND2_X1 maj_226_U3 ( .A1(maj_226_n26), .A2(maj_226_n25), .ZN(maj_226_port_o) );
  XOR2_X1 maj_226_U2 ( .A(maj_226_n22), .B(maj_226_n21), .Z(maj_226_n23) );
  NAND2_X1 maj_227_U15 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_227_n18) );
  NAND2_X1 maj_227_U14 ( .A1(maj_227_n21), .A2(maj_227_n22), .ZN(maj_227_n17)
         );
  NAND2_X1 maj_227_U13 ( .A1(maj_227_n18), .A2(maj_227_n17), .ZN(maj_227_n19)
         );
  NAND2_X1 maj_227_U12 ( .A1(v_1_2[2]), .A2(maj_227_n16), .ZN(maj_227_n14) );
  NAND2_X1 maj_227_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_227_n15) );
  NAND2_X1 maj_227_U10 ( .A1(maj_227_n15), .A2(maj_227_n14), .ZN(maj_227_n20)
         );
  XOR2_X1 maj_227_U9 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_227_n22) );
  XOR2_X1 maj_227_U8 ( .A(v_1_2[2]), .B(maj_227_n16), .Z(maj_227_n21) );
  XOR2_X1 maj_227_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_227_n16) );
  OR2_X1 maj_227_U6 ( .A1(maj_227_n20), .A2(maj_227_n19), .ZN(maj_227_n24) );
  NAND2_X1 maj_227_U5 ( .A1(maj_227_n24), .A2(maj_227_n23), .ZN(maj_227_n25)
         );
  NAND2_X1 maj_227_U4 ( .A1(maj_227_n20), .A2(maj_227_n19), .ZN(maj_227_n26)
         );
  NAND2_X1 maj_227_U3 ( .A1(maj_227_n26), .A2(maj_227_n25), .ZN(maj_227_port_o) );
  XOR2_X1 maj_227_U2 ( .A(maj_227_n22), .B(maj_227_n21), .Z(maj_227_n23) );
  NAND2_X1 maj_228_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_228_n18) );
  NAND2_X1 maj_228_U14 ( .A1(maj_228_n21), .A2(maj_228_n22), .ZN(maj_228_n17)
         );
  NAND2_X1 maj_228_U13 ( .A1(maj_228_n18), .A2(maj_228_n17), .ZN(maj_228_n19)
         );
  NAND2_X1 maj_228_U12 ( .A1(u_2_0[2]), .A2(maj_228_n16), .ZN(maj_228_n14) );
  NAND2_X1 maj_228_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_228_n15) );
  NAND2_X1 maj_228_U10 ( .A1(maj_228_n15), .A2(maj_228_n14), .ZN(maj_228_n20)
         );
  XOR2_X1 maj_228_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_228_n22) );
  XOR2_X1 maj_228_U8 ( .A(u_2_0[2]), .B(maj_228_n16), .Z(maj_228_n21) );
  XOR2_X1 maj_228_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_228_n16) );
  OR2_X1 maj_228_U6 ( .A1(maj_228_n20), .A2(maj_228_n19), .ZN(maj_228_n24) );
  NAND2_X1 maj_228_U5 ( .A1(maj_228_n24), .A2(maj_228_n23), .ZN(maj_228_n25)
         );
  NAND2_X1 maj_228_U4 ( .A1(maj_228_n20), .A2(maj_228_n19), .ZN(maj_228_n26)
         );
  NAND2_X1 maj_228_U3 ( .A1(maj_228_n26), .A2(maj_228_n25), .ZN(maj_228_port_o) );
  XOR2_X1 maj_228_U2 ( .A(maj_228_n22), .B(maj_228_n21), .Z(maj_228_n23) );
  NAND2_X1 maj_229_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_229_n18) );
  NAND2_X1 maj_229_U14 ( .A1(maj_229_n21), .A2(maj_229_n22), .ZN(maj_229_n17)
         );
  NAND2_X1 maj_229_U13 ( .A1(maj_229_n18), .A2(maj_229_n17), .ZN(maj_229_n19)
         );
  NAND2_X1 maj_229_U12 ( .A1(v_2_0[2]), .A2(maj_229_n16), .ZN(maj_229_n14) );
  NAND2_X1 maj_229_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_229_n15) );
  NAND2_X1 maj_229_U10 ( .A1(maj_229_n15), .A2(maj_229_n14), .ZN(maj_229_n20)
         );
  XOR2_X1 maj_229_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_229_n22) );
  XOR2_X1 maj_229_U8 ( .A(v_2_0[2]), .B(maj_229_n16), .Z(maj_229_n21) );
  XOR2_X1 maj_229_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_229_n16) );
  OR2_X1 maj_229_U6 ( .A1(maj_229_n20), .A2(maj_229_n19), .ZN(maj_229_n24) );
  NAND2_X1 maj_229_U5 ( .A1(maj_229_n24), .A2(maj_229_n23), .ZN(maj_229_n25)
         );
  NAND2_X1 maj_229_U4 ( .A1(maj_229_n20), .A2(maj_229_n19), .ZN(maj_229_n26)
         );
  NAND2_X1 maj_229_U3 ( .A1(maj_229_n26), .A2(maj_229_n25), .ZN(maj_229_port_o) );
  XOR2_X1 maj_229_U2 ( .A(maj_229_n22), .B(maj_229_n21), .Z(maj_229_n23) );
  NAND2_X1 maj_230_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_230_n18) );
  NAND2_X1 maj_230_U14 ( .A1(maj_230_n21), .A2(maj_230_n22), .ZN(maj_230_n17)
         );
  NAND2_X1 maj_230_U13 ( .A1(maj_230_n18), .A2(maj_230_n17), .ZN(maj_230_n19)
         );
  NAND2_X1 maj_230_U12 ( .A1(u_2_1[2]), .A2(maj_230_n16), .ZN(maj_230_n14) );
  NAND2_X1 maj_230_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_230_n15) );
  NAND2_X1 maj_230_U10 ( .A1(maj_230_n15), .A2(maj_230_n14), .ZN(maj_230_n20)
         );
  XOR2_X1 maj_230_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_230_n22) );
  XOR2_X1 maj_230_U8 ( .A(u_2_1[2]), .B(maj_230_n16), .Z(maj_230_n21) );
  XOR2_X1 maj_230_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_230_n16) );
  OR2_X1 maj_230_U6 ( .A1(maj_230_n20), .A2(maj_230_n19), .ZN(maj_230_n24) );
  NAND2_X1 maj_230_U5 ( .A1(maj_230_n24), .A2(maj_230_n23), .ZN(maj_230_n25)
         );
  NAND2_X1 maj_230_U4 ( .A1(maj_230_n20), .A2(maj_230_n19), .ZN(maj_230_n26)
         );
  NAND2_X1 maj_230_U3 ( .A1(maj_230_n26), .A2(maj_230_n25), .ZN(maj_230_port_o) );
  XOR2_X1 maj_230_U2 ( .A(maj_230_n22), .B(maj_230_n21), .Z(maj_230_n23) );
  NAND2_X1 maj_231_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_231_n18) );
  NAND2_X1 maj_231_U14 ( .A1(maj_231_n21), .A2(maj_231_n22), .ZN(maj_231_n17)
         );
  NAND2_X1 maj_231_U13 ( .A1(maj_231_n18), .A2(maj_231_n17), .ZN(maj_231_n19)
         );
  NAND2_X1 maj_231_U12 ( .A1(v_2_1[2]), .A2(maj_231_n16), .ZN(maj_231_n14) );
  NAND2_X1 maj_231_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_231_n15) );
  NAND2_X1 maj_231_U10 ( .A1(maj_231_n15), .A2(maj_231_n14), .ZN(maj_231_n20)
         );
  XOR2_X1 maj_231_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_231_n22) );
  XOR2_X1 maj_231_U8 ( .A(v_2_1[2]), .B(maj_231_n16), .Z(maj_231_n21) );
  XOR2_X1 maj_231_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_231_n16) );
  OR2_X1 maj_231_U6 ( .A1(maj_231_n20), .A2(maj_231_n19), .ZN(maj_231_n24) );
  NAND2_X1 maj_231_U5 ( .A1(maj_231_n24), .A2(maj_231_n23), .ZN(maj_231_n25)
         );
  NAND2_X1 maj_231_U4 ( .A1(maj_231_n20), .A2(maj_231_n19), .ZN(maj_231_n26)
         );
  NAND2_X1 maj_231_U3 ( .A1(maj_231_n26), .A2(maj_231_n25), .ZN(maj_231_port_o) );
  XOR2_X1 maj_231_U2 ( .A(maj_231_n22), .B(maj_231_n21), .Z(maj_231_n23) );
  NAND2_X1 maj_232_U15 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_232_n18) );
  NAND2_X1 maj_232_U14 ( .A1(maj_232_n21), .A2(maj_232_n22), .ZN(maj_232_n17)
         );
  NAND2_X1 maj_232_U13 ( .A1(maj_232_n18), .A2(maj_232_n17), .ZN(maj_232_n19)
         );
  NAND2_X1 maj_232_U12 ( .A1(u_2_2[2]), .A2(maj_232_n16), .ZN(maj_232_n14) );
  NAND2_X1 maj_232_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_232_n15) );
  NAND2_X1 maj_232_U10 ( .A1(maj_232_n15), .A2(maj_232_n14), .ZN(maj_232_n20)
         );
  XOR2_X1 maj_232_U9 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_232_n22) );
  XOR2_X1 maj_232_U8 ( .A(u_2_2[2]), .B(maj_232_n16), .Z(maj_232_n21) );
  XOR2_X1 maj_232_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_232_n16) );
  OR2_X1 maj_232_U6 ( .A1(maj_232_n20), .A2(maj_232_n19), .ZN(maj_232_n24) );
  NAND2_X1 maj_232_U5 ( .A1(maj_232_n24), .A2(maj_232_n23), .ZN(maj_232_n25)
         );
  NAND2_X1 maj_232_U4 ( .A1(maj_232_n20), .A2(maj_232_n19), .ZN(maj_232_n26)
         );
  NAND2_X1 maj_232_U3 ( .A1(maj_232_n26), .A2(maj_232_n25), .ZN(maj_232_port_o) );
  XOR2_X1 maj_232_U2 ( .A(maj_232_n22), .B(maj_232_n21), .Z(maj_232_n23) );
  NAND2_X1 maj_233_U15 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_233_n18) );
  NAND2_X1 maj_233_U14 ( .A1(maj_233_n21), .A2(maj_233_n22), .ZN(maj_233_n17)
         );
  NAND2_X1 maj_233_U13 ( .A1(maj_233_n18), .A2(maj_233_n17), .ZN(maj_233_n19)
         );
  NAND2_X1 maj_233_U12 ( .A1(v_2_2[2]), .A2(maj_233_n16), .ZN(maj_233_n14) );
  NAND2_X1 maj_233_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_233_n15) );
  NAND2_X1 maj_233_U10 ( .A1(maj_233_n15), .A2(maj_233_n14), .ZN(maj_233_n20)
         );
  XOR2_X1 maj_233_U9 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_233_n22) );
  XOR2_X1 maj_233_U8 ( .A(v_2_2[2]), .B(maj_233_n16), .Z(maj_233_n21) );
  XOR2_X1 maj_233_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_233_n16) );
  OR2_X1 maj_233_U6 ( .A1(maj_233_n20), .A2(maj_233_n19), .ZN(maj_233_n24) );
  NAND2_X1 maj_233_U5 ( .A1(maj_233_n24), .A2(maj_233_n23), .ZN(maj_233_n25)
         );
  NAND2_X1 maj_233_U4 ( .A1(maj_233_n20), .A2(maj_233_n19), .ZN(maj_233_n26)
         );
  NAND2_X1 maj_233_U3 ( .A1(maj_233_n26), .A2(maj_233_n25), .ZN(maj_233_port_o) );
  XOR2_X1 maj_233_U2 ( .A(maj_233_n22), .B(maj_233_n21), .Z(maj_233_n23) );
  NAND2_X1 maj_234_U15 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_234_n18) );
  NAND2_X1 maj_234_U14 ( .A1(maj_234_n21), .A2(maj_234_n22), .ZN(maj_234_n17)
         );
  NAND2_X1 maj_234_U13 ( .A1(maj_234_n18), .A2(maj_234_n17), .ZN(maj_234_n19)
         );
  NAND2_X1 maj_234_U12 ( .A1(u_3_0[2]), .A2(maj_234_n16), .ZN(maj_234_n14) );
  NAND2_X1 maj_234_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_234_n15) );
  NAND2_X1 maj_234_U10 ( .A1(maj_234_n15), .A2(maj_234_n14), .ZN(maj_234_n20)
         );
  XOR2_X1 maj_234_U9 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_234_n22) );
  XOR2_X1 maj_234_U8 ( .A(u_3_0[2]), .B(maj_234_n16), .Z(maj_234_n21) );
  XOR2_X1 maj_234_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_234_n16) );
  OR2_X1 maj_234_U6 ( .A1(maj_234_n20), .A2(maj_234_n19), .ZN(maj_234_n24) );
  NAND2_X1 maj_234_U5 ( .A1(maj_234_n24), .A2(maj_234_n23), .ZN(maj_234_n25)
         );
  NAND2_X1 maj_234_U4 ( .A1(maj_234_n20), .A2(maj_234_n19), .ZN(maj_234_n26)
         );
  NAND2_X1 maj_234_U3 ( .A1(maj_234_n26), .A2(maj_234_n25), .ZN(maj_234_port_o) );
  XOR2_X1 maj_234_U2 ( .A(maj_234_n22), .B(maj_234_n21), .Z(maj_234_n23) );
  NAND2_X1 maj_235_U15 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_235_n18) );
  NAND2_X1 maj_235_U14 ( .A1(maj_235_n21), .A2(maj_235_n22), .ZN(maj_235_n17)
         );
  NAND2_X1 maj_235_U13 ( .A1(maj_235_n18), .A2(maj_235_n17), .ZN(maj_235_n19)
         );
  NAND2_X1 maj_235_U12 ( .A1(v_3_0[2]), .A2(maj_235_n16), .ZN(maj_235_n14) );
  NAND2_X1 maj_235_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_235_n15) );
  NAND2_X1 maj_235_U10 ( .A1(maj_235_n15), .A2(maj_235_n14), .ZN(maj_235_n20)
         );
  XOR2_X1 maj_235_U9 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_235_n22) );
  XOR2_X1 maj_235_U8 ( .A(v_3_0[2]), .B(maj_235_n16), .Z(maj_235_n21) );
  XOR2_X1 maj_235_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_235_n16) );
  OR2_X1 maj_235_U6 ( .A1(maj_235_n20), .A2(maj_235_n19), .ZN(maj_235_n24) );
  NAND2_X1 maj_235_U5 ( .A1(maj_235_n24), .A2(maj_235_n23), .ZN(maj_235_n25)
         );
  NAND2_X1 maj_235_U4 ( .A1(maj_235_n20), .A2(maj_235_n19), .ZN(maj_235_n26)
         );
  NAND2_X1 maj_235_U3 ( .A1(maj_235_n26), .A2(maj_235_n25), .ZN(maj_235_port_o) );
  XOR2_X1 maj_235_U2 ( .A(maj_235_n22), .B(maj_235_n21), .Z(maj_235_n23) );
  NAND2_X1 maj_236_U15 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_236_n18) );
  NAND2_X1 maj_236_U14 ( .A1(maj_236_n21), .A2(maj_236_n22), .ZN(maj_236_n17)
         );
  NAND2_X1 maj_236_U13 ( .A1(maj_236_n18), .A2(maj_236_n17), .ZN(maj_236_n19)
         );
  NAND2_X1 maj_236_U12 ( .A1(u_3_1[2]), .A2(maj_236_n16), .ZN(maj_236_n14) );
  NAND2_X1 maj_236_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_236_n15) );
  NAND2_X1 maj_236_U10 ( .A1(maj_236_n15), .A2(maj_236_n14), .ZN(maj_236_n20)
         );
  XOR2_X1 maj_236_U9 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_236_n22) );
  XOR2_X1 maj_236_U8 ( .A(u_3_1[2]), .B(maj_236_n16), .Z(maj_236_n21) );
  XOR2_X1 maj_236_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_236_n16) );
  OR2_X1 maj_236_U6 ( .A1(maj_236_n20), .A2(maj_236_n19), .ZN(maj_236_n24) );
  NAND2_X1 maj_236_U5 ( .A1(maj_236_n24), .A2(maj_236_n23), .ZN(maj_236_n25)
         );
  NAND2_X1 maj_236_U4 ( .A1(maj_236_n20), .A2(maj_236_n19), .ZN(maj_236_n26)
         );
  NAND2_X1 maj_236_U3 ( .A1(maj_236_n26), .A2(maj_236_n25), .ZN(maj_236_port_o) );
  XOR2_X1 maj_236_U2 ( .A(maj_236_n22), .B(maj_236_n21), .Z(maj_236_n23) );
  NAND2_X1 maj_237_U15 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_237_n18) );
  NAND2_X1 maj_237_U14 ( .A1(maj_237_n21), .A2(maj_237_n22), .ZN(maj_237_n17)
         );
  NAND2_X1 maj_237_U13 ( .A1(maj_237_n18), .A2(maj_237_n17), .ZN(maj_237_n19)
         );
  NAND2_X1 maj_237_U12 ( .A1(v_3_1[2]), .A2(maj_237_n16), .ZN(maj_237_n14) );
  NAND2_X1 maj_237_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_237_n15) );
  NAND2_X1 maj_237_U10 ( .A1(maj_237_n15), .A2(maj_237_n14), .ZN(maj_237_n20)
         );
  XOR2_X1 maj_237_U9 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_237_n22) );
  XOR2_X1 maj_237_U8 ( .A(v_3_1[2]), .B(maj_237_n16), .Z(maj_237_n21) );
  XOR2_X1 maj_237_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_237_n16) );
  OR2_X1 maj_237_U6 ( .A1(maj_237_n20), .A2(maj_237_n19), .ZN(maj_237_n24) );
  NAND2_X1 maj_237_U5 ( .A1(maj_237_n24), .A2(maj_237_n23), .ZN(maj_237_n25)
         );
  NAND2_X1 maj_237_U4 ( .A1(maj_237_n20), .A2(maj_237_n19), .ZN(maj_237_n26)
         );
  NAND2_X1 maj_237_U3 ( .A1(maj_237_n26), .A2(maj_237_n25), .ZN(maj_237_port_o) );
  XOR2_X1 maj_237_U2 ( .A(maj_237_n22), .B(maj_237_n21), .Z(maj_237_n23) );
  NAND2_X1 maj_238_U15 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_238_n18) );
  NAND2_X1 maj_238_U14 ( .A1(maj_238_n21), .A2(maj_238_n22), .ZN(maj_238_n17)
         );
  NAND2_X1 maj_238_U13 ( .A1(maj_238_n18), .A2(maj_238_n17), .ZN(maj_238_n19)
         );
  NAND2_X1 maj_238_U12 ( .A1(u_3_2[2]), .A2(maj_238_n16), .ZN(maj_238_n14) );
  NAND2_X1 maj_238_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_238_n15) );
  NAND2_X1 maj_238_U10 ( .A1(maj_238_n15), .A2(maj_238_n14), .ZN(maj_238_n20)
         );
  XOR2_X1 maj_238_U9 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_238_n22) );
  XOR2_X1 maj_238_U8 ( .A(u_3_2[2]), .B(maj_238_n16), .Z(maj_238_n21) );
  XOR2_X1 maj_238_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_238_n16) );
  OR2_X1 maj_238_U6 ( .A1(maj_238_n20), .A2(maj_238_n19), .ZN(maj_238_n24) );
  NAND2_X1 maj_238_U5 ( .A1(maj_238_n24), .A2(maj_238_n23), .ZN(maj_238_n25)
         );
  NAND2_X1 maj_238_U4 ( .A1(maj_238_n20), .A2(maj_238_n19), .ZN(maj_238_n26)
         );
  NAND2_X1 maj_238_U3 ( .A1(maj_238_n26), .A2(maj_238_n25), .ZN(maj_238_port_o) );
  XOR2_X1 maj_238_U2 ( .A(maj_238_n22), .B(maj_238_n21), .Z(maj_238_n23) );
  NAND2_X1 maj_239_U15 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_239_n18) );
  NAND2_X1 maj_239_U14 ( .A1(maj_239_n21), .A2(maj_239_n22), .ZN(maj_239_n17)
         );
  NAND2_X1 maj_239_U13 ( .A1(maj_239_n18), .A2(maj_239_n17), .ZN(maj_239_n19)
         );
  NAND2_X1 maj_239_U12 ( .A1(v_3_2[2]), .A2(maj_239_n16), .ZN(maj_239_n14) );
  NAND2_X1 maj_239_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_239_n15) );
  NAND2_X1 maj_239_U10 ( .A1(maj_239_n15), .A2(maj_239_n14), .ZN(maj_239_n20)
         );
  XOR2_X1 maj_239_U9 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_239_n22) );
  XOR2_X1 maj_239_U8 ( .A(v_3_2[2]), .B(maj_239_n16), .Z(maj_239_n21) );
  XOR2_X1 maj_239_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_239_n16) );
  OR2_X1 maj_239_U6 ( .A1(maj_239_n20), .A2(maj_239_n19), .ZN(maj_239_n24) );
  NAND2_X1 maj_239_U5 ( .A1(maj_239_n24), .A2(maj_239_n23), .ZN(maj_239_n25)
         );
  NAND2_X1 maj_239_U4 ( .A1(maj_239_n20), .A2(maj_239_n19), .ZN(maj_239_n26)
         );
  NAND2_X1 maj_239_U3 ( .A1(maj_239_n26), .A2(maj_239_n25), .ZN(maj_239_port_o) );
  XOR2_X1 maj_239_U2 ( .A(maj_239_n22), .B(maj_239_n21), .Z(maj_239_n23) );
endmodule

