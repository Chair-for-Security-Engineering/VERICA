
module And_gate ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, 
        io_i0_s4, io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, p_rand_0, 
        p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7, 
        p_rand_8, p_rand_9, io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4
 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i0_s2, io_i0_s3, io_i0_s4,
         io_i1_s0, io_i1_s1, io_i1_s2, io_i1_s3, io_i1_s4, p_rand_0, p_rand_1,
         p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7, p_rand_8,
         p_rand_9;
  output io_o0_s0, io_o0_s1, io_o0_s2, io_o0_s3, io_o0_s4;
  wire   n_hpc2_0_n140, n_hpc2_0_n139, n_hpc2_0_n138, n_hpc2_0_n137,
         n_hpc2_0_n136, n_hpc2_0_n135, n_hpc2_0_n134, n_hpc2_0_n133,
         n_hpc2_0_n132, n_hpc2_0_n131, n_hpc2_0_n130, n_hpc2_0_n129,
         n_hpc2_0_n128, n_hpc2_0_n127, n_hpc2_0_n126, n_hpc2_0_n125,
         n_hpc2_0_n124, n_hpc2_0_n123, n_hpc2_0_n122, n_hpc2_0_n121,
         n_hpc2_0_n120, n_hpc2_0_n119, n_hpc2_0_n118, n_hpc2_0_n117,
         n_hpc2_0_n116, n_hpc2_0_n115, n_hpc2_0_n114, n_hpc2_0_n113,
         n_hpc2_0_n112, n_hpc2_0_n111, n_hpc2_0_n110, n_hpc2_0_n109,
         n_hpc2_0_n108, n_hpc2_0_n107, n_hpc2_0_n106, n_hpc2_0_n105,
         n_hpc2_0_n104, n_hpc2_0_n103, n_hpc2_0_n102, n_hpc2_0_n101,
         n_hpc2_0_n100, n_hpc2_0_n99, n_hpc2_0_n98, n_hpc2_0_n97, n_hpc2_0_n96,
         n_hpc2_0_n95, n_hpc2_0_n94, n_hpc2_0_n93, n_hpc2_0_n92, n_hpc2_0_n91,
         n_hpc2_0_n90, n_hpc2_0_n89, n_hpc2_0_n88, n_hpc2_0_n87, n_hpc2_0_n86,
         n_hpc2_0_n85, n_hpc2_0_n84, n_hpc2_0_n83, n_hpc2_0_n82, n_hpc2_0_n81,
         n_hpc2_0_n80, n_hpc2_0_n79, n_hpc2_0_n78, n_hpc2_0_n77, n_hpc2_0_n76,
         n_hpc2_0_n75, n_hpc2_0_n74, n_hpc2_0_n73, n_hpc2_0_n72, n_hpc2_0_n71,
         n_hpc2_0_n70, n_hpc2_0_n69, n_hpc2_0_n68, n_hpc2_0_n67, n_hpc2_0_n66,
         n_hpc2_0_n65, n_hpc2_0_n64, n_hpc2_0_n63, n_hpc2_0_n62, n_hpc2_0_n61,
         n_hpc2_0_n60, n_hpc2_0_n59, n_hpc2_0_n58, n_hpc2_0_n57, n_hpc2_0_n56,
         n_hpc2_0_n55, n_hpc2_0_n54, n_hpc2_0_n53, n_hpc2_0_n52, n_hpc2_0_n51,
         n_hpc2_0_n50, n_hpc2_0_n49, n_hpc2_0_n48, n_hpc2_0_n47, n_hpc2_0_n46,
         n_hpc2_0_n45, n_hpc2_0_n44, n_hpc2_0_n43, n_hpc2_0_n42, n_hpc2_0_n41,
         n_hpc2_0_n40, n_hpc2_0_n39, n_hpc2_0_n38, n_hpc2_0_n37, n_hpc2_0_n36,
         n_hpc2_0_n35, n_hpc2_0_n34, n_hpc2_0_n33, n_hpc2_0_n32, n_hpc2_0_n31,
         n_hpc2_0_n30, n_hpc2_0_n29, n_hpc2_0_n28, n_hpc2_0_n27, n_hpc2_0_n26,
         n_hpc2_0_n25, n_hpc2_0_n24, n_hpc2_0_n23, n_hpc2_0_n22, n_hpc2_0_n21,
         n_hpc2_0_n20, n_hpc2_0_n19, n_hpc2_0_n18, n_hpc2_0_n17, n_hpc2_0_n16,
         n_hpc2_0_n15, n_hpc2_0_n14, n_hpc2_0_n13, n_hpc2_0_n12, n_hpc2_0_n11,
         n_hpc2_0_n10, n_hpc2_0_n9, n_hpc2_0_n8, n_hpc2_0_n7, n_hpc2_0_n6,
         n_hpc2_0_n5, n_hpc2_0_n4, n_hpc2_0_n3, n_hpc2_0_n2, n_hpc2_0_n1,
         n_hpc2_0_N69, n_hpc2_0_N68, n_hpc2_0_N67, n_hpc2_0_N66, n_hpc2_0_N65,
         n_hpc2_0_N64, n_hpc2_0_N63, n_hpc2_0_N62, n_hpc2_0_N61, n_hpc2_0_N60,
         n_hpc2_0_N59, n_hpc2_0_N58, n_hpc2_0_N57, n_hpc2_0_N56, n_hpc2_0_N55,
         n_hpc2_0_N54, n_hpc2_0_N53, n_hpc2_0_N52, n_hpc2_0_N51, n_hpc2_0_N50,
         n_hpc2_0_N49, n_hpc2_0_N48, n_hpc2_0_N47, n_hpc2_0_N46, n_hpc2_0_N45,
         n_hpc2_0_N44, n_hpc2_0_N43, n_hpc2_0_N42, n_hpc2_0_N41, n_hpc2_0_N40,
         n_hpc2_0_N39, n_hpc2_0_N38, n_hpc2_0_N37, n_hpc2_0_N36, n_hpc2_0_N35,
         n_hpc2_0_N34, n_hpc2_0_N33, n_hpc2_0_N32, n_hpc2_0_N31, n_hpc2_0_N30,
         n_hpc2_0_N29, n_hpc2_0_N28, n_hpc2_0_N27, n_hpc2_0_N26, n_hpc2_0_N25,
         n_hpc2_0_N24, n_hpc2_0_N23, n_hpc2_0_N22, n_hpc2_0_N21, n_hpc2_0_N20,
         n_hpc2_0_N19, n_hpc2_0_N18, n_hpc2_0_N17, n_hpc2_0_N16, n_hpc2_0_N15,
         n_hpc2_0_N14, n_hpc2_0_N13, n_hpc2_0_N12, n_hpc2_0_N11, n_hpc2_0_N10,
         n_hpc2_0_N9, n_hpc2_0_N8, n_hpc2_0_N7, n_hpc2_0_N6, n_hpc2_0_N5,
         n_hpc2_0__hpc_u43, n_hpc2_0__hpc_u34, n_hpc2_0__hpc_u24,
         n_hpc2_0__hpc_u14, n_hpc2_0__hpc_u04;

  NOR2_X1 u_hpc2_0_U112 ( .A1(n_hpc2_0_n140), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N10) );
  NOR2_X1 u_hpc2_0_U111 ( .A1(n_hpc2_0_n139), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N11) );
  NOR2_X1 u_hpc2_0_U110 ( .A1(n_hpc2_0_n138), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N12) );
  NOR2_X1 u_hpc2_0_U109 ( .A1(n_hpc2_0_n137), .A2(n_hpc2_0_n10), .ZN(
        n_hpc2_0_N13) );
  NOR2_X1 u_hpc2_0_U108 ( .A1(n_hpc2_0_n136), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N14) );
  NOR2_X1 u_hpc2_0_U107 ( .A1(n_hpc2_0_n135), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N15) );
  NOR2_X1 u_hpc2_0_U106 ( .A1(n_hpc2_0_n134), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N16) );
  NOR2_X1 u_hpc2_0_U105 ( .A1(n_hpc2_0_n133), .A2(n_hpc2_0_n9), .ZN(
        n_hpc2_0_N17) );
  NOR2_X1 u_hpc2_0_U104 ( .A1(n_hpc2_0_n132), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N18) );
  NOR2_X1 u_hpc2_0_U103 ( .A1(n_hpc2_0_n131), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N19) );
  NOR2_X1 u_hpc2_0_U102 ( .A1(n_hpc2_0_n130), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N20) );
  NOR2_X1 u_hpc2_0_U101 ( .A1(n_hpc2_0_n129), .A2(n_hpc2_0_n8), .ZN(
        n_hpc2_0_N21) );
  NOR2_X1 u_hpc2_0_U100 ( .A1(n_hpc2_0_n128), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N22) );
  NOR2_X1 u_hpc2_0_U99 ( .A1(n_hpc2_0_n127), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N23) );
  NOR2_X1 u_hpc2_0_U98 ( .A1(n_hpc2_0_n126), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N24) );
  NOR2_X1 u_hpc2_0_U97 ( .A1(n_hpc2_0_n125), .A2(n_hpc2_0_n7), .ZN(
        n_hpc2_0_N25) );
  NOR2_X1 u_hpc2_0_U96 ( .A1(n_hpc2_0_n124), .A2(n_hpc2_0_n6), .ZN(
        n_hpc2_0_N26) );
  NOR2_X1 u_hpc2_0_U95 ( .A1(n_hpc2_0_n123), .A2(n_hpc2_0_n6), .ZN(
        n_hpc2_0_N27) );
  NOR2_X1 u_hpc2_0_U94 ( .A1(n_hpc2_0_n122), .A2(n_hpc2_0_n6), .ZN(
        n_hpc2_0_N28) );
  NOR2_X1 u_hpc2_0_U93 ( .A1(n_hpc2_0_n121), .A2(n_hpc2_0_n6), .ZN(
        n_hpc2_0_N29) );
  NOR2_X1 u_hpc2_0_U92 ( .A1(n_hpc2_0_n119), .A2(n_hpc2_0_n120), .ZN(
        n_hpc2_0_N30) );
  NOR2_X1 u_hpc2_0_U91 ( .A1(n_hpc2_0_n117), .A2(n_hpc2_0_n118), .ZN(
        n_hpc2_0_N31) );
  NOR2_X1 u_hpc2_0_U90 ( .A1(n_hpc2_0_n115), .A2(n_hpc2_0_n116), .ZN(
        n_hpc2_0_N32) );
  NOR2_X1 u_hpc2_0_U89 ( .A1(n_hpc2_0_n113), .A2(n_hpc2_0_n114), .ZN(
        n_hpc2_0_N33) );
  NOR2_X1 u_hpc2_0_U88 ( .A1(n_hpc2_0_n119), .A2(n_hpc2_0_n112), .ZN(
        n_hpc2_0_N34) );
  NOR2_X1 u_hpc2_0_U87 ( .A1(n_hpc2_0_n110), .A2(n_hpc2_0_n111), .ZN(
        n_hpc2_0_N35) );
  NOR2_X1 u_hpc2_0_U86 ( .A1(n_hpc2_0_n108), .A2(n_hpc2_0_n109), .ZN(
        n_hpc2_0_N36) );
  NOR2_X1 u_hpc2_0_U85 ( .A1(n_hpc2_0_n106), .A2(n_hpc2_0_n107), .ZN(
        n_hpc2_0_N37) );
  NOR2_X1 u_hpc2_0_U84 ( .A1(n_hpc2_0_n117), .A2(n_hpc2_0_n105), .ZN(
        n_hpc2_0_N38) );
  NOR2_X1 u_hpc2_0_U83 ( .A1(n_hpc2_0_n110), .A2(n_hpc2_0_n104), .ZN(
        n_hpc2_0_N39) );
  NOR2_X1 u_hpc2_0_U82 ( .A1(n_hpc2_0_n102), .A2(n_hpc2_0_n103), .ZN(
        n_hpc2_0_N40) );
  NOR2_X1 u_hpc2_0_U81 ( .A1(n_hpc2_0_n100), .A2(n_hpc2_0_n101), .ZN(
        n_hpc2_0_N41) );
  NOR2_X1 u_hpc2_0_U80 ( .A1(n_hpc2_0_n115), .A2(n_hpc2_0_n99), .ZN(
        n_hpc2_0_N42) );
  NOR2_X1 u_hpc2_0_U79 ( .A1(n_hpc2_0_n108), .A2(n_hpc2_0_n98), .ZN(
        n_hpc2_0_N43) );
  NOR2_X1 u_hpc2_0_U78 ( .A1(n_hpc2_0_n102), .A2(n_hpc2_0_n97), .ZN(
        n_hpc2_0_N44) );
  NOR2_X1 u_hpc2_0_U77 ( .A1(n_hpc2_0_n95), .A2(n_hpc2_0_n96), .ZN(
        n_hpc2_0_N45) );
  NOR2_X1 u_hpc2_0_U76 ( .A1(n_hpc2_0_n113), .A2(n_hpc2_0_n94), .ZN(
        n_hpc2_0_N46) );
  NOR2_X1 u_hpc2_0_U75 ( .A1(n_hpc2_0_n106), .A2(n_hpc2_0_n93), .ZN(
        n_hpc2_0_N47) );
  NOR2_X1 u_hpc2_0_U74 ( .A1(n_hpc2_0_n100), .A2(n_hpc2_0_n92), .ZN(
        n_hpc2_0_N48) );
  NOR2_X1 u_hpc2_0_U73 ( .A1(n_hpc2_0_n95), .A2(n_hpc2_0_n91), .ZN(
        n_hpc2_0_N49) );
  NOR2_X1 u_hpc2_0_U72 ( .A1(n_hpc2_0_n90), .A2(n_hpc2_0_n10), .ZN(n_hpc2_0_N5) );
  XOR2_X1 u_hpc2_0_U71 ( .A(io_i1_s1), .B(p_rand_0), .Z(n_hpc2_0_N50) );
  XOR2_X1 u_hpc2_0_U70 ( .A(io_i1_s2), .B(p_rand_1), .Z(n_hpc2_0_N51) );
  XOR2_X1 u_hpc2_0_U69 ( .A(io_i1_s3), .B(p_rand_2), .Z(n_hpc2_0_N52) );
  XOR2_X1 u_hpc2_0_U68 ( .A(io_i1_s4), .B(p_rand_3), .Z(n_hpc2_0_N53) );
  XOR2_X1 u_hpc2_0_U67 ( .A(io_i1_s0), .B(p_rand_0), .Z(n_hpc2_0_N54) );
  XOR2_X1 u_hpc2_0_U66 ( .A(io_i1_s2), .B(p_rand_4), .Z(n_hpc2_0_N55) );
  XOR2_X1 u_hpc2_0_U65 ( .A(io_i1_s3), .B(p_rand_5), .Z(n_hpc2_0_N56) );
  XOR2_X1 u_hpc2_0_U64 ( .A(io_i1_s4), .B(p_rand_6), .Z(n_hpc2_0_N57) );
  XOR2_X1 u_hpc2_0_U63 ( .A(io_i1_s0), .B(p_rand_1), .Z(n_hpc2_0_N58) );
  XOR2_X1 u_hpc2_0_U62 ( .A(io_i1_s1), .B(p_rand_4), .Z(n_hpc2_0_N59) );
  NOR2_X1 u_hpc2_0_U61 ( .A1(n_hpc2_0_n89), .A2(n_hpc2_0_n9), .ZN(n_hpc2_0_N6)
         );
  XOR2_X1 u_hpc2_0_U60 ( .A(io_i1_s3), .B(p_rand_7), .Z(n_hpc2_0_N60) );
  XOR2_X1 u_hpc2_0_U59 ( .A(io_i1_s4), .B(p_rand_8), .Z(n_hpc2_0_N61) );
  XOR2_X1 u_hpc2_0_U58 ( .A(io_i1_s0), .B(p_rand_2), .Z(n_hpc2_0_N62) );
  XOR2_X1 u_hpc2_0_U57 ( .A(io_i1_s1), .B(p_rand_5), .Z(n_hpc2_0_N63) );
  XOR2_X1 u_hpc2_0_U56 ( .A(io_i1_s2), .B(p_rand_7), .Z(n_hpc2_0_N64) );
  XOR2_X1 u_hpc2_0_U55 ( .A(io_i1_s4), .B(p_rand_9), .Z(n_hpc2_0_N65) );
  XOR2_X1 u_hpc2_0_U54 ( .A(io_i1_s0), .B(p_rand_3), .Z(n_hpc2_0_N66) );
  XOR2_X1 u_hpc2_0_U53 ( .A(io_i1_s1), .B(p_rand_6), .Z(n_hpc2_0_N67) );
  XOR2_X1 u_hpc2_0_U52 ( .A(io_i1_s2), .B(p_rand_8), .Z(n_hpc2_0_N68) );
  XOR2_X1 u_hpc2_0_U51 ( .A(io_i1_s3), .B(p_rand_9), .Z(n_hpc2_0_N69) );
  NOR2_X1 u_hpc2_0_U50 ( .A1(n_hpc2_0_n88), .A2(n_hpc2_0_n8), .ZN(n_hpc2_0_N7)
         );
  NOR2_X1 u_hpc2_0_U49 ( .A1(n_hpc2_0_n87), .A2(n_hpc2_0_n7), .ZN(n_hpc2_0_N8)
         );
  NOR2_X1 u_hpc2_0_U48 ( .A1(n_hpc2_0_n86), .A2(n_hpc2_0_n6), .ZN(n_hpc2_0_N9)
         );
  INV_X1 u_hpc2_0_U47 ( .A(io_i0_s0), .ZN(n_hpc2_0_n1) );
  INV_X1 u_hpc2_0_U46 ( .A(io_i0_s1), .ZN(n_hpc2_0_n2) );
  INV_X1 u_hpc2_0_U45 ( .A(io_i0_s2), .ZN(n_hpc2_0_n3) );
  INV_X1 u_hpc2_0_U44 ( .A(io_i0_s3), .ZN(n_hpc2_0_n4) );
  INV_X1 u_hpc2_0_U43 ( .A(io_i0_s4), .ZN(n_hpc2_0_n5) );
  XOR2_X1 u_hpc2_0_U42 ( .A(n_hpc2_0__hpc_u04), .B(n_hpc2_0_n85), .Z(
        n_hpc2_0_n44) );
  XOR2_X1 u_hpc2_0_U41 ( .A(n_hpc2_0_n83), .B(n_hpc2_0_n84), .Z(n_hpc2_0_n45)
         );
  XOR2_X1 u_hpc2_0_U40 ( .A(n_hpc2_0_n44), .B(n_hpc2_0_n45), .Z(n_hpc2_0_n40)
         );
  XOR2_X1 u_hpc2_0_U39 ( .A(n_hpc2_0_n79), .B(n_hpc2_0_n80), .Z(n_hpc2_0_n42)
         );
  XOR2_X1 u_hpc2_0_U38 ( .A(n_hpc2_0_n81), .B(n_hpc2_0_n82), .Z(n_hpc2_0_n43)
         );
  XOR2_X1 u_hpc2_0_U37 ( .A(n_hpc2_0_n42), .B(n_hpc2_0_n43), .Z(n_hpc2_0_n41)
         );
  XOR2_X1 u_hpc2_0_U36 ( .A(n_hpc2_0_n40), .B(n_hpc2_0_n41), .Z(n_hpc2_0_n39)
         );
  XOR2_X1 u_hpc2_0_U35 ( .A(n_hpc2_0_n39), .B(n_hpc2_0_n78), .Z(io_o0_s0) );
  XOR2_X1 u_hpc2_0_U34 ( .A(n_hpc2_0__hpc_u14), .B(n_hpc2_0_n77), .Z(
        n_hpc2_0_n37) );
  XOR2_X1 u_hpc2_0_U33 ( .A(n_hpc2_0_n75), .B(n_hpc2_0_n76), .Z(n_hpc2_0_n38)
         );
  XOR2_X1 u_hpc2_0_U32 ( .A(n_hpc2_0_n37), .B(n_hpc2_0_n38), .Z(n_hpc2_0_n33)
         );
  XOR2_X1 u_hpc2_0_U31 ( .A(n_hpc2_0_n71), .B(n_hpc2_0_n72), .Z(n_hpc2_0_n35)
         );
  XOR2_X1 u_hpc2_0_U30 ( .A(n_hpc2_0_n73), .B(n_hpc2_0_n74), .Z(n_hpc2_0_n36)
         );
  XOR2_X1 u_hpc2_0_U29 ( .A(n_hpc2_0_n35), .B(n_hpc2_0_n36), .Z(n_hpc2_0_n34)
         );
  XOR2_X1 u_hpc2_0_U28 ( .A(n_hpc2_0_n33), .B(n_hpc2_0_n34), .Z(n_hpc2_0_n32)
         );
  XOR2_X1 u_hpc2_0_U27 ( .A(n_hpc2_0_n32), .B(n_hpc2_0_n70), .Z(io_o0_s1) );
  XOR2_X1 u_hpc2_0_U26 ( .A(n_hpc2_0__hpc_u24), .B(n_hpc2_0_n69), .Z(
        n_hpc2_0_n30) );
  XOR2_X1 u_hpc2_0_U25 ( .A(n_hpc2_0_n67), .B(n_hpc2_0_n68), .Z(n_hpc2_0_n31)
         );
  XOR2_X1 u_hpc2_0_U24 ( .A(n_hpc2_0_n30), .B(n_hpc2_0_n31), .Z(n_hpc2_0_n26)
         );
  XOR2_X1 u_hpc2_0_U23 ( .A(n_hpc2_0_n63), .B(n_hpc2_0_n64), .Z(n_hpc2_0_n28)
         );
  XOR2_X1 u_hpc2_0_U22 ( .A(n_hpc2_0_n65), .B(n_hpc2_0_n66), .Z(n_hpc2_0_n29)
         );
  XOR2_X1 u_hpc2_0_U21 ( .A(n_hpc2_0_n28), .B(n_hpc2_0_n29), .Z(n_hpc2_0_n27)
         );
  XOR2_X1 u_hpc2_0_U20 ( .A(n_hpc2_0_n26), .B(n_hpc2_0_n27), .Z(n_hpc2_0_n25)
         );
  XOR2_X1 u_hpc2_0_U19 ( .A(n_hpc2_0_n25), .B(n_hpc2_0_n62), .Z(io_o0_s2) );
  XOR2_X1 u_hpc2_0_U18 ( .A(n_hpc2_0__hpc_u34), .B(n_hpc2_0_n61), .Z(
        n_hpc2_0_n23) );
  XOR2_X1 u_hpc2_0_U17 ( .A(n_hpc2_0_n59), .B(n_hpc2_0_n60), .Z(n_hpc2_0_n24)
         );
  XOR2_X1 u_hpc2_0_U16 ( .A(n_hpc2_0_n23), .B(n_hpc2_0_n24), .Z(n_hpc2_0_n19)
         );
  XOR2_X1 u_hpc2_0_U15 ( .A(n_hpc2_0_n55), .B(n_hpc2_0_n56), .Z(n_hpc2_0_n21)
         );
  XOR2_X1 u_hpc2_0_U14 ( .A(n_hpc2_0_n57), .B(n_hpc2_0_n58), .Z(n_hpc2_0_n22)
         );
  XOR2_X1 u_hpc2_0_U13 ( .A(n_hpc2_0_n21), .B(n_hpc2_0_n22), .Z(n_hpc2_0_n20)
         );
  XOR2_X1 u_hpc2_0_U12 ( .A(n_hpc2_0_n19), .B(n_hpc2_0_n20), .Z(n_hpc2_0_n18)
         );
  XOR2_X1 u_hpc2_0_U11 ( .A(n_hpc2_0_n18), .B(n_hpc2_0_n54), .Z(io_o0_s3) );
  XOR2_X1 u_hpc2_0_U10 ( .A(n_hpc2_0__hpc_u43), .B(n_hpc2_0_n53), .Z(
        n_hpc2_0_n16) );
  XOR2_X1 u_hpc2_0_U9 ( .A(n_hpc2_0_n51), .B(n_hpc2_0_n52), .Z(n_hpc2_0_n17)
         );
  XOR2_X1 u_hpc2_0_U8 ( .A(n_hpc2_0_n16), .B(n_hpc2_0_n17), .Z(n_hpc2_0_n12)
         );
  XOR2_X1 u_hpc2_0_U7 ( .A(n_hpc2_0_n47), .B(n_hpc2_0_n48), .Z(n_hpc2_0_n14)
         );
  XOR2_X1 u_hpc2_0_U6 ( .A(n_hpc2_0_n49), .B(n_hpc2_0_n50), .Z(n_hpc2_0_n15)
         );
  XOR2_X1 u_hpc2_0_U5 ( .A(n_hpc2_0_n14), .B(n_hpc2_0_n15), .Z(n_hpc2_0_n13)
         );
  XOR2_X1 u_hpc2_0_U4 ( .A(n_hpc2_0_n12), .B(n_hpc2_0_n13), .Z(n_hpc2_0_n11)
         );
  XOR2_X1 u_hpc2_0_U3 ( .A(n_hpc2_0_n11), .B(n_hpc2_0_n46), .Z(io_o0_s4) );
  DFF_X1 u_hpc2_0__hpc_av32_reg ( .D(n_hpc2_0_N24), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n58) );
  DFF_X1 u_hpc2_0__hpc_v32_reg ( .D(n_hpc2_0_N64), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n126) );
  DFF_X1 u_hpc2_0__hpc_av31_reg ( .D(n_hpc2_0_N23), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n57) );
  DFF_X1 u_hpc2_0__hpc_v31_reg ( .D(n_hpc2_0_N63), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n127) );
  DFF_X1 u_hpc2_0__hpc_av30_reg ( .D(n_hpc2_0_N22), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n56) );
  DFF_X1 u_hpc2_0__hpc_v30_reg ( .D(n_hpc2_0_N62), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n128) );
  DFF_X1 u_hpc2_0__hpc_av24_reg ( .D(n_hpc2_0_N21), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n67) );
  DFF_X1 u_hpc2_0__hpc_v24_reg ( .D(n_hpc2_0_N61), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n129) );
  DFF_X1 u_hpc2_0__hpc_av23_reg ( .D(n_hpc2_0_N20), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n66) );
  DFF_X1 u_hpc2_0__hpc_v23_reg ( .D(n_hpc2_0_N60), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n130) );
  DFF_X1 u_hpc2_0__hpc_av21_reg ( .D(n_hpc2_0_N19), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n65) );
  DFF_X1 u_hpc2_0__hpc_v21_reg ( .D(n_hpc2_0_N59), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n131) );
  DFF_X1 u_hpc2_0__hpc_av20_reg ( .D(n_hpc2_0_N18), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n64) );
  DFF_X1 u_hpc2_0__hpc_v20_reg ( .D(n_hpc2_0_N58), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n132) );
  DFF_X1 u_hpc2_0__hpc_av14_reg ( .D(n_hpc2_0_N17), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n75) );
  DFF_X1 u_hpc2_0__hpc_v14_reg ( .D(n_hpc2_0_N57), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n133) );
  DFF_X1 u_hpc2_0__hpc_av13_reg ( .D(n_hpc2_0_N16), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n74) );
  DFF_X1 u_hpc2_0__hpc_v13_reg ( .D(n_hpc2_0_N56), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n134) );
  DFF_X1 u_hpc2_0__hpc_av12_reg ( .D(n_hpc2_0_N15), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n73) );
  DFF_X1 u_hpc2_0__hpc_v12_reg ( .D(n_hpc2_0_N55), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n135) );
  DFF_X1 u_hpc2_0__hpc_av10_reg ( .D(n_hpc2_0_N14), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n72) );
  DFF_X1 u_hpc2_0__hpc_v10_reg ( .D(n_hpc2_0_N54), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n136) );
  DFF_X1 u_hpc2_0__hpc_av04_reg ( .D(n_hpc2_0_N13), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n83) );
  DFF_X1 u_hpc2_0__hpc_v04_reg ( .D(n_hpc2_0_N53), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n137) );
  DFF_X1 u_hpc2_0__hpc_av03_reg ( .D(n_hpc2_0_N12), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n82) );
  DFF_X1 u_hpc2_0__hpc_v03_reg ( .D(n_hpc2_0_N52), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n138) );
  DFF_X1 u_hpc2_0__hpc_av02_reg ( .D(n_hpc2_0_N11), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n81) );
  DFF_X1 u_hpc2_0__hpc_v02_reg ( .D(n_hpc2_0_N51), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n139) );
  DFF_X1 u_hpc2_0__hpc_av01_reg ( .D(n_hpc2_0_N10), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n80) );
  DFF_X1 u_hpc2_0__hpc_v01_reg ( .D(n_hpc2_0_N50), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n140) );
  DFF_X1 u_hpc2_0__hpc_u43_reg ( .D(n_hpc2_0_N49), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u43), .QN() );
  DFF_X1 u_hpc2_0__hpc_u42_reg ( .D(n_hpc2_0_N48), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n53) );
  DFF_X1 u_hpc2_0__hpc_u41_reg ( .D(n_hpc2_0_N47), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n52) );
  DFF_X1 u_hpc2_0__hpc_u40_reg ( .D(n_hpc2_0_N46), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n46) );
  DFF_X1 u_hpc2_0__hpc_u34_reg ( .D(n_hpc2_0_N45), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u34), .QN() );
  DFF_X1 u_hpc2_0__hpc_u32_reg ( .D(n_hpc2_0_N44), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n61) );
  DFF_X1 u_hpc2_0__hpc_u31_reg ( .D(n_hpc2_0_N43), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n60) );
  DFF_X1 u_hpc2_0__hpc_u30_reg ( .D(n_hpc2_0_N42), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n54) );
  DFF_X1 u_hpc2_0__hpc_u24_reg ( .D(n_hpc2_0_N41), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u24), .QN() );
  DFF_X1 u_hpc2_0__hpc_u23_reg ( .D(n_hpc2_0_N40), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n69) );
  DFF_X1 u_hpc2_0__hpc_u21_reg ( .D(n_hpc2_0_N39), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n68) );
  DFF_X1 u_hpc2_0__hpc_u20_reg ( .D(n_hpc2_0_N38), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n62) );
  DFF_X1 u_hpc2_0__hpc_u14_reg ( .D(n_hpc2_0_N37), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u14), .QN() );
  DFF_X1 u_hpc2_0__hpc_u13_reg ( .D(n_hpc2_0_N36), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n77) );
  DFF_X1 u_hpc2_0__hpc_u12_reg ( .D(n_hpc2_0_N35), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n76) );
  DFF_X1 u_hpc2_0__hpc_u10_reg ( .D(n_hpc2_0_N34), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n70) );
  DFF_X1 u_hpc2_0__hpc_u04_reg ( .D(n_hpc2_0_N33), .CK(clock_0), .Q(
        n_hpc2_0__hpc_u04), .QN() );
  DFF_X1 u_hpc2_0__hpc_u03_reg ( .D(n_hpc2_0_N32), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n85) );
  DFF_X1 u_hpc2_0__hpc_u02_reg ( .D(n_hpc2_0_N31), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n84) );
  DFF_X1 u_hpc2_0__hpc_u01_reg ( .D(n_hpc2_0_N30), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n78) );
  DFF_X1 u_hpc2_0__hpc_ab4_reg ( .D(n_hpc2_0_N9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n47) );
  DFF_X1 u_hpc2_0__hpc_b4_reg ( .D(io_i1_s4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n86) );
  DFF_X1 u_hpc2_0__hpc_ab3_reg ( .D(n_hpc2_0_N8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n55) );
  DFF_X1 u_hpc2_0__hpc_b3_reg ( .D(io_i1_s3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n87) );
  DFF_X1 u_hpc2_0__hpc_ab2_reg ( .D(n_hpc2_0_N7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n63) );
  DFF_X1 u_hpc2_0__hpc_b2_reg ( .D(io_i1_s2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n88) );
  DFF_X1 u_hpc2_0__hpc_ab1_reg ( .D(n_hpc2_0_N6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n71) );
  DFF_X1 u_hpc2_0__hpc_b1_reg ( .D(io_i1_s1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n89) );
  DFF_X1 u_hpc2_0__hpc_ab0_reg ( .D(n_hpc2_0_N5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n79) );
  DFF_X1 u_hpc2_0__hpc_b0_reg ( .D(io_i1_s0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n90) );
  DFF_X1 u_hpc2_0__hpc_av43_reg ( .D(n_hpc2_0_N29), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n51) );
  DFF_X1 u_hpc2_0__hpc_av42_reg ( .D(n_hpc2_0_N28), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n50) );
  DFF_X1 u_hpc2_0__hpc_av41_reg ( .D(n_hpc2_0_N27), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n49) );
  DFF_X1 u_hpc2_0__hpc_av40_reg ( .D(n_hpc2_0_N26), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n48) );
  DFF_X1 u_hpc2_0__hpc_av34_reg ( .D(n_hpc2_0_N25), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n59) );
  DFF_X1 u_hpc2_0_reg_pipeline_13_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n111) );
  DFF_X1 u_hpc2_0_reg_pipeline_15_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n114) );
  DFF_X1 u_hpc2_0_reg_pipeline_2_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n94) );
  DFF_X1 u_hpc2_0_reg_pipeline_19_reg ( .D(io_i0_s0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n10) );
  DFF_X1 u_hpc2_0_reg_pipeline_20_reg ( .D(io_i0_s1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n9) );
  DFF_X1 u_hpc2_0_reg_pipeline_17_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n118) );
  DFF_X1 u_hpc2_0_reg_pipeline_12_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n109) );
  DFF_X1 u_hpc2_0_reg_pipeline_16_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n116) );
  DFF_X1 u_hpc2_0_reg_pipeline_18_reg ( .D(n_hpc2_0_n1), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n120) );
  DFF_X1 u_hpc2_0_reg_pipeline_14_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n112) );
  DFF_X1 u_hpc2_0_reg_pipeline_5_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n98) );
  DFF_X1 u_hpc2_0_reg_pipeline_6_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n99) );
  DFF_X1 u_hpc2_0_reg_pipeline_9_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n104) );
  DFF_X1 u_hpc2_0_reg_pipeline_7_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n101) );
  DFF_X1 u_hpc2_0__hpc_r9_reg ( .D(p_rand_9), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n95) );
  DFF_X1 u_hpc2_0__hpc_r7_reg ( .D(p_rand_7), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n102) );
  DFF_X1 u_hpc2_0_reg_pipeline_8_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n103) );
  DFF_X1 u_hpc2_0__hpc_r8_reg ( .D(p_rand_8), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n100) );
  DFF_X1 u_hpc2_0__hpc_r6_reg ( .D(p_rand_6), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n106) );
  DFF_X1 u_hpc2_0__hpc_r5_reg ( .D(p_rand_5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n108) );
  DFF_X1 u_hpc2_0_reg_pipeline_11_reg ( .D(n_hpc2_0_n2), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n107) );
  DFF_X1 u_hpc2_0_reg_pipeline_10_reg ( .D(n_hpc2_0_n3), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n105) );
  DFF_X1 u_hpc2_0_reg_pipeline_1_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n93) );
  DFF_X1 u_hpc2_0_reg_pipeline_0_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n92) );
  DFF_X1 u_hpc2_0_reg_pipeline_reg ( .D(n_hpc2_0_n5), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n91) );
  DFF_X1 u_hpc2_0__hpc_v43_reg ( .D(n_hpc2_0_N69), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n121) );
  DFF_X1 u_hpc2_0__hpc_v42_reg ( .D(n_hpc2_0_N68), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n122) );
  DFF_X1 u_hpc2_0__hpc_v41_reg ( .D(n_hpc2_0_N67), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n123) );
  DFF_X1 u_hpc2_0__hpc_v40_reg ( .D(n_hpc2_0_N66), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n124) );
  DFF_X1 u_hpc2_0__hpc_v34_reg ( .D(n_hpc2_0_N65), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n125) );
  DFF_X1 u_hpc2_0_reg_pipeline_4_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n97) );
  DFF_X1 u_hpc2_0_reg_pipeline_21_reg ( .D(io_i0_s2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n8) );
  DFF_X1 u_hpc2_0_reg_pipeline_22_reg ( .D(io_i0_s3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n7) );
  DFF_X1 u_hpc2_0_reg_pipeline_23_reg ( .D(io_i0_s4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n6) );
  DFF_X1 u_hpc2_0_reg_pipeline_3_reg ( .D(n_hpc2_0_n4), .CK(clock_0), .Q(), 
        .QN(n_hpc2_0_n96) );
  DFF_X1 u_hpc2_0__hpc_r4_reg ( .D(p_rand_4), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n110) );
  DFF_X1 u_hpc2_0__hpc_r3_reg ( .D(p_rand_3), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n113) );
  DFF_X1 u_hpc2_0__hpc_r2_reg ( .D(p_rand_2), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n115) );
  DFF_X1 u_hpc2_0__hpc_r1_reg ( .D(p_rand_1), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n117) );
  DFF_X1 u_hpc2_0__hpc_r0_reg ( .D(p_rand_0), .CK(clock_0), .Q(), .QN(
        n_hpc2_0_n119) );
endmodule

