
module keccak_b25_r10_i2_o1 ( clock, reset, io_block_i0, io_block_i1, 
        io_block_o0 );
  input [9:0] io_block_i0;
  input [9:0] io_block_i1;
  output [9:0] io_block_o0;
  input clock, reset;
  wire   f0_io_state_out_0_0, f0_io_state_out_0_1, f0_io_state_out_1_0,
         f0_io_state_out_1_1, f0_io_state_out_2_0, f0_io_state_out_2_1,
         f0_io_state_out_3_0, f0_io_state_out_3_1, f0_io_state_out_4_0,
         f0_io_state_out_4_1, abs1_io_state_out_0_0, abs1_io_state_out_0_1,
         abs1_io_state_out_0_2, abs1_io_state_out_0_3, abs1_io_state_out_0_4,
         abs1_io_state_out_1_0, abs1_io_state_out_1_1, abs1_io_state_out_1_2,
         abs1_io_state_out_1_3, abs1_io_state_out_1_4, abs1_io_state_out_2_0,
         abs1_io_state_out_2_1, abs1_io_state_out_2_2, abs1_io_state_out_2_3,
         abs1_io_state_out_2_4, abs1_io_state_out_3_0, abs1_io_state_out_3_1,
         abs1_io_state_out_3_2, abs1_io_state_out_3_3, abs1_io_state_out_3_4,
         abs1_io_state_out_4_0, abs1_io_state_out_4_1, abs1_io_state_out_4_2,
         abs1_io_state_out_4_3, abs1_io_state_out_4_4,
         f0_round_9_io_state_out_4_4, f0_round_9_io_state_out_4_3,
         f0_round_9_io_state_out_4_2, f0_round_9_io_state_out_4_1,
         f0_round_9_io_state_out_4_0, f0_round_9_io_state_out_3_4,
         f0_round_9_io_state_out_3_3, f0_round_9_io_state_out_3_2,
         f0_round_9_io_state_out_3_1, f0_round_9_io_state_out_3_0,
         f0_round_9_io_state_out_2_4, f0_round_9_io_state_out_2_3,
         f0_round_9_io_state_out_2_2, f0_round_9_io_state_out_2_1,
         f0_round_9_io_state_out_2_0, f0_round_9_io_state_out_1_4,
         f0_round_9_io_state_out_1_3, f0_round_9_io_state_out_1_2,
         f0_round_9_io_state_out_1_1, f0_round_9_io_state_out_1_0,
         f0_round_9_io_state_out_0_4, f0_round_9_io_state_out_0_3,
         f0_round_9_io_state_out_0_2, f0_round_9_io_state_out_0_1,
         f0_round_9_io_state_out_0_0, f0_round_8_io_state_out_4_4,
         f0_round_8_io_state_out_4_3, f0_round_8_io_state_out_4_2,
         f0_round_8_io_state_out_4_1, f0_round_8_io_state_out_4_0,
         f0_round_8_io_state_out_3_4, f0_round_8_io_state_out_3_3,
         f0_round_8_io_state_out_3_2, f0_round_8_io_state_out_3_1,
         f0_round_8_io_state_out_3_0, f0_round_8_io_state_out_2_4,
         f0_round_8_io_state_out_2_3, f0_round_8_io_state_out_2_2,
         f0_round_8_io_state_out_2_1, f0_round_8_io_state_out_2_0,
         f0_round_8_io_state_out_1_4, f0_round_8_io_state_out_1_3,
         f0_round_8_io_state_out_1_2, f0_round_8_io_state_out_1_1,
         f0_round_8_io_state_out_1_0, f0_round_8_io_state_out_0_4,
         f0_round_8_io_state_out_0_3, f0_round_8_io_state_out_0_2,
         f0_round_8_io_state_out_0_1, f0_round_8_io_state_out_0_0,
         f0_round_7_io_state_out_4_4, f0_round_7_io_state_out_4_3,
         f0_round_7_io_state_out_4_2, f0_round_7_io_state_out_4_1,
         f0_round_7_io_state_out_4_0, f0_round_7_io_state_out_3_4,
         f0_round_7_io_state_out_3_3, f0_round_7_io_state_out_3_2,
         f0_round_7_io_state_out_3_1, f0_round_7_io_state_out_3_0,
         f0_round_7_io_state_out_2_4, f0_round_7_io_state_out_2_3,
         f0_round_7_io_state_out_2_2, f0_round_7_io_state_out_2_1,
         f0_round_7_io_state_out_2_0, f0_round_7_io_state_out_1_4,
         f0_round_7_io_state_out_1_3, f0_round_7_io_state_out_1_2,
         f0_round_7_io_state_out_1_1, f0_round_7_io_state_out_1_0,
         f0_round_7_io_state_out_0_4, f0_round_7_io_state_out_0_3,
         f0_round_7_io_state_out_0_2, f0_round_7_io_state_out_0_1,
         f0_round_7_io_state_out_0_0, f0_round_6_io_state_out_4_4,
         f0_round_6_io_state_out_4_3, f0_round_6_io_state_out_4_2,
         f0_round_6_io_state_out_4_1, f0_round_6_io_state_out_4_0,
         f0_round_6_io_state_out_3_4, f0_round_6_io_state_out_3_3,
         f0_round_6_io_state_out_3_2, f0_round_6_io_state_out_3_1,
         f0_round_6_io_state_out_3_0, f0_round_6_io_state_out_2_4,
         f0_round_6_io_state_out_2_3, f0_round_6_io_state_out_2_2,
         f0_round_6_io_state_out_2_1, f0_round_6_io_state_out_2_0,
         f0_round_6_io_state_out_1_4, f0_round_6_io_state_out_1_3,
         f0_round_6_io_state_out_1_2, f0_round_6_io_state_out_1_1,
         f0_round_6_io_state_out_1_0, f0_round_6_io_state_out_0_4,
         f0_round_6_io_state_out_0_3, f0_round_6_io_state_out_0_2,
         f0_round_6_io_state_out_0_1, f0_round_6_io_state_out_0_0,
         f0_round_5_io_state_out_4_4, f0_round_5_io_state_out_4_3,
         f0_round_5_io_state_out_4_2, f0_round_5_io_state_out_4_1,
         f0_round_5_io_state_out_4_0, f0_round_5_io_state_out_3_4,
         f0_round_5_io_state_out_3_3, f0_round_5_io_state_out_3_2,
         f0_round_5_io_state_out_3_1, f0_round_5_io_state_out_3_0,
         f0_round_5_io_state_out_2_4, f0_round_5_io_state_out_2_3,
         f0_round_5_io_state_out_2_2, f0_round_5_io_state_out_2_1,
         f0_round_5_io_state_out_2_0, f0_round_5_io_state_out_1_4,
         f0_round_5_io_state_out_1_3, f0_round_5_io_state_out_1_2,
         f0_round_5_io_state_out_1_1, f0_round_5_io_state_out_1_0,
         f0_round_5_io_state_out_0_4, f0_round_5_io_state_out_0_3,
         f0_round_5_io_state_out_0_2, f0_round_5_io_state_out_0_1,
         f0_round_5_io_state_out_0_0, f0_round_4_io_state_out_4_4,
         f0_round_4_io_state_out_4_3, f0_round_4_io_state_out_4_2,
         f0_round_4_io_state_out_4_1, f0_round_4_io_state_out_4_0,
         f0_round_4_io_state_out_3_4, f0_round_4_io_state_out_3_3,
         f0_round_4_io_state_out_3_2, f0_round_4_io_state_out_3_1,
         f0_round_4_io_state_out_3_0, f0_round_4_io_state_out_2_4,
         f0_round_4_io_state_out_2_3, f0_round_4_io_state_out_2_2,
         f0_round_4_io_state_out_2_1, f0_round_4_io_state_out_2_0,
         f0_round_4_io_state_out_1_4, f0_round_4_io_state_out_1_3,
         f0_round_4_io_state_out_1_2, f0_round_4_io_state_out_1_1,
         f0_round_4_io_state_out_1_0, f0_round_4_io_state_out_0_4,
         f0_round_4_io_state_out_0_3, f0_round_4_io_state_out_0_2,
         f0_round_4_io_state_out_0_1, f0_round_4_io_state_out_0_0,
         f0_round_3_io_state_out_4_4, f0_round_3_io_state_out_4_3,
         f0_round_3_io_state_out_4_2, f0_round_3_io_state_out_4_1,
         f0_round_3_io_state_out_4_0, f0_round_3_io_state_out_3_4,
         f0_round_3_io_state_out_3_3, f0_round_3_io_state_out_3_2,
         f0_round_3_io_state_out_3_1, f0_round_3_io_state_out_3_0,
         f0_round_3_io_state_out_2_4, f0_round_3_io_state_out_2_3,
         f0_round_3_io_state_out_2_2, f0_round_3_io_state_out_2_1,
         f0_round_3_io_state_out_2_0, f0_round_3_io_state_out_1_4,
         f0_round_3_io_state_out_1_3, f0_round_3_io_state_out_1_2,
         f0_round_3_io_state_out_1_1, f0_round_3_io_state_out_1_0,
         f0_round_3_io_state_out_0_4, f0_round_3_io_state_out_0_3,
         f0_round_3_io_state_out_0_2, f0_round_3_io_state_out_0_1,
         f0_round_3_io_state_out_0_0, f0_round_2_io_state_out_4_4,
         f0_round_2_io_state_out_4_3, f0_round_2_io_state_out_4_2,
         f0_round_2_io_state_out_4_1, f0_round_2_io_state_out_4_0,
         f0_round_2_io_state_out_3_4, f0_round_2_io_state_out_3_3,
         f0_round_2_io_state_out_3_2, f0_round_2_io_state_out_3_1,
         f0_round_2_io_state_out_3_0, f0_round_2_io_state_out_2_4,
         f0_round_2_io_state_out_2_3, f0_round_2_io_state_out_2_2,
         f0_round_2_io_state_out_2_1, f0_round_2_io_state_out_2_0,
         f0_round_2_io_state_out_1_4, f0_round_2_io_state_out_1_3,
         f0_round_2_io_state_out_1_2, f0_round_2_io_state_out_1_1,
         f0_round_2_io_state_out_1_0, f0_round_2_io_state_out_0_4,
         f0_round_2_io_state_out_0_3, f0_round_2_io_state_out_0_2,
         f0_round_2_io_state_out_0_1, f0_round_2_io_state_out_0_0,
         f0_round_1_io_state_out_4_4, f0_round_1_io_state_out_4_3,
         f0_round_1_io_state_out_4_2, f0_round_1_io_state_out_4_1,
         f0_round_1_io_state_out_4_0, f0_round_1_io_state_out_3_4,
         f0_round_1_io_state_out_3_3, f0_round_1_io_state_out_3_2,
         f0_round_1_io_state_out_3_1, f0_round_1_io_state_out_3_0,
         f0_round_1_io_state_out_2_4, f0_round_1_io_state_out_2_3,
         f0_round_1_io_state_out_2_2, f0_round_1_io_state_out_2_1,
         f0_round_1_io_state_out_2_0, f0_round_1_io_state_out_1_4,
         f0_round_1_io_state_out_1_3, f0_round_1_io_state_out_1_2,
         f0_round_1_io_state_out_1_1, f0_round_1_io_state_out_1_0,
         f0_round_1_io_state_out_0_4, f0_round_1_io_state_out_0_3,
         f0_round_1_io_state_out_0_2, f0_round_1_io_state_out_0_1,
         f0_round_1_io_state_out_0_0, f0_round_io_state_out_4_4,
         f0_round_io_state_out_4_3, f0_round_io_state_out_4_2,
         f0_round_io_state_out_4_1, f0_round_io_state_out_4_0,
         f0_round_io_state_out_3_4, f0_round_io_state_out_3_3,
         f0_round_io_state_out_3_2, f0_round_io_state_out_3_1,
         f0_round_io_state_out_3_0, f0_round_io_state_out_2_4,
         f0_round_io_state_out_2_3, f0_round_io_state_out_2_2,
         f0_round_io_state_out_2_1, f0_round_io_state_out_2_0,
         f0_round_io_state_out_1_4, f0_round_io_state_out_1_3,
         f0_round_io_state_out_1_2, f0_round_io_state_out_1_1,
         f0_round_io_state_out_1_0, f0_round_io_state_out_0_4,
         f0_round_io_state_out_0_3, f0_round_io_state_out_0_2,
         f0_round_io_state_out_0_1, f0_round_io_state_out_0_0,
         f0_round0_io_state_out_4_4, f0_round0_io_state_out_4_3,
         f0_round0_io_state_out_4_2, f0_round0_io_state_out_4_1,
         f0_round0_io_state_out_4_0, f0_round0_io_state_out_3_4,
         f0_round0_io_state_out_3_3, f0_round0_io_state_out_3_2,
         f0_round0_io_state_out_3_1, f0_round0_io_state_out_3_0,
         f0_round0_io_state_out_2_4, f0_round0_io_state_out_2_3,
         f0_round0_io_state_out_2_2, f0_round0_io_state_out_2_1,
         f0_round0_io_state_out_2_0, f0_round0_io_state_out_1_4,
         f0_round0_io_state_out_1_3, f0_round0_io_state_out_1_2,
         f0_round0_io_state_out_1_1, f0_round0_io_state_out_1_0,
         f0_round0_io_state_out_0_4, f0_round0_io_state_out_0_3,
         f0_round0_io_state_out_0_2, f0_round0_io_state_out_0_1,
         f0_round0_io_state_out_0_0, f0_round0_c_io_state_out_0_0,
         f0_round0_p_io_state_out_2_4, f0_round0_p_io_state_out_2_3,
         f0_round0_p_io_state_out_2_2, f0_round0_p_io_state_out_2_1,
         f0_round0_p_io_state_out_2_0, f0_round0_p_io_state_out_1_4,
         f0_round0_p_io_state_out_1_3, f0_round0_p_io_state_out_1_2,
         f0_round0_p_io_state_out_1_1, f0_round0_p_io_state_out_1_0,
         f0_round0_p_io_state_out_0_4, f0_round0_p_io_state_out_0_3,
         f0_round0_p_io_state_out_0_2, f0_round0_p_io_state_out_0_1,
         f0_round0_p_io_state_out_0_0, f0_round0_t_n5, f0_round0_t_n4,
         f0_round0_t_n3, f0_round0_t_n2, f0_round0_t_n1, f0_round0_c_n25,
         f0_round0_c_n24, f0_round0_c_n23, f0_round0_c_n22, f0_round0_c_n21,
         f0_round0_c_n20, f0_round0_c_n19, f0_round0_c_n18, f0_round0_c_n17,
         f0_round0_c_n16, f0_round0_c_n15, f0_round0_c_n14, f0_round0_c_n13,
         f0_round0_c_n12, f0_round0_c_n11, f0_round0_c_n10, f0_round0_c_n9,
         f0_round0_c_n8, f0_round0_c_n7, f0_round0_c_n6, f0_round0_c_n5,
         f0_round0_c_n4, f0_round0_c_n3, f0_round0_c_n2, f0_round0_c_n1,
         f0_round_p_io_state_out_4_4, f0_round_p_io_state_out_4_3,
         f0_round_p_io_state_out_4_2, f0_round_p_io_state_out_4_1,
         f0_round_p_io_state_out_4_0, f0_round_p_io_state_out_3_4,
         f0_round_p_io_state_out_3_3, f0_round_p_io_state_out_3_2,
         f0_round_p_io_state_out_3_1, f0_round_p_io_state_out_3_0,
         f0_round_p_io_state_out_2_4, f0_round_p_io_state_out_2_3,
         f0_round_p_io_state_out_2_2, f0_round_p_io_state_out_2_1,
         f0_round_p_io_state_out_2_0, f0_round_p_io_state_out_1_4,
         f0_round_p_io_state_out_1_3, f0_round_p_io_state_out_1_2,
         f0_round_p_io_state_out_1_1, f0_round_p_io_state_out_1_0,
         f0_round_p_io_state_out_0_4, f0_round_p_io_state_out_0_3,
         f0_round_p_io_state_out_0_2, f0_round_p_io_state_out_0_1,
         f0_round_p_io_state_out_0_0, f0_round_t_n25, f0_round_t_n24,
         f0_round_t_n23, f0_round_t_n22, f0_round_t_n21, f0_round_t_n20,
         f0_round_t_n19, f0_round_t_n18, f0_round_t_n17, f0_round_t_n16,
         f0_round_t_n15, f0_round_t_n14, f0_round_t_n13, f0_round_t_n12,
         f0_round_t_n11, f0_round_t_n10, f0_round_t_n9, f0_round_t_n8,
         f0_round_t_n7, f0_round_t_n6, f0_round_t_n5, f0_round_t_n4,
         f0_round_t_n3, f0_round_t_n2, f0_round_t_n1, f0_round_c_n25,
         f0_round_c_n24, f0_round_c_n23, f0_round_c_n22, f0_round_c_n21,
         f0_round_c_n20, f0_round_c_n19, f0_round_c_n18, f0_round_c_n17,
         f0_round_c_n16, f0_round_c_n15, f0_round_c_n14, f0_round_c_n13,
         f0_round_c_n12, f0_round_c_n11, f0_round_c_n10, f0_round_c_n9,
         f0_round_c_n8, f0_round_c_n7, f0_round_c_n6, f0_round_c_n5,
         f0_round_c_n4, f0_round_c_n3, f0_round_c_n2, f0_round_c_n1,
         f0_round_1_p_io_state_out_4_4, f0_round_1_p_io_state_out_4_3,
         f0_round_1_p_io_state_out_4_2, f0_round_1_p_io_state_out_4_1,
         f0_round_1_p_io_state_out_4_0, f0_round_1_p_io_state_out_3_4,
         f0_round_1_p_io_state_out_3_3, f0_round_1_p_io_state_out_3_2,
         f0_round_1_p_io_state_out_3_1, f0_round_1_p_io_state_out_3_0,
         f0_round_1_p_io_state_out_2_4, f0_round_1_p_io_state_out_2_3,
         f0_round_1_p_io_state_out_2_2, f0_round_1_p_io_state_out_2_1,
         f0_round_1_p_io_state_out_2_0, f0_round_1_p_io_state_out_1_4,
         f0_round_1_p_io_state_out_1_3, f0_round_1_p_io_state_out_1_2,
         f0_round_1_p_io_state_out_1_1, f0_round_1_p_io_state_out_1_0,
         f0_round_1_p_io_state_out_0_4, f0_round_1_p_io_state_out_0_3,
         f0_round_1_p_io_state_out_0_2, f0_round_1_p_io_state_out_0_1,
         f0_round_1_p_io_state_out_0_0, f0_round_1_t_n25, f0_round_1_t_n24,
         f0_round_1_t_n23, f0_round_1_t_n22, f0_round_1_t_n21,
         f0_round_1_t_n20, f0_round_1_t_n19, f0_round_1_t_n18,
         f0_round_1_t_n17, f0_round_1_t_n16, f0_round_1_t_n15,
         f0_round_1_t_n14, f0_round_1_t_n13, f0_round_1_t_n12,
         f0_round_1_t_n11, f0_round_1_t_n10, f0_round_1_t_n9, f0_round_1_t_n8,
         f0_round_1_t_n7, f0_round_1_t_n6, f0_round_1_t_n5, f0_round_1_t_n4,
         f0_round_1_t_n3, f0_round_1_t_n2, f0_round_1_t_n1, f0_round_1_c_n25,
         f0_round_1_c_n24, f0_round_1_c_n23, f0_round_1_c_n22,
         f0_round_1_c_n21, f0_round_1_c_n20, f0_round_1_c_n19,
         f0_round_1_c_n18, f0_round_1_c_n17, f0_round_1_c_n16,
         f0_round_1_c_n15, f0_round_1_c_n14, f0_round_1_c_n13,
         f0_round_1_c_n12, f0_round_1_c_n11, f0_round_1_c_n10, f0_round_1_c_n9,
         f0_round_1_c_n8, f0_round_1_c_n7, f0_round_1_c_n6, f0_round_1_c_n5,
         f0_round_1_c_n4, f0_round_1_c_n3, f0_round_1_c_n2, f0_round_1_c_n1,
         f0_round_2_p_io_state_out_4_4, f0_round_2_p_io_state_out_4_3,
         f0_round_2_p_io_state_out_4_2, f0_round_2_p_io_state_out_4_1,
         f0_round_2_p_io_state_out_4_0, f0_round_2_p_io_state_out_3_4,
         f0_round_2_p_io_state_out_3_3, f0_round_2_p_io_state_out_3_2,
         f0_round_2_p_io_state_out_3_1, f0_round_2_p_io_state_out_3_0,
         f0_round_2_p_io_state_out_2_4, f0_round_2_p_io_state_out_2_3,
         f0_round_2_p_io_state_out_2_2, f0_round_2_p_io_state_out_2_1,
         f0_round_2_p_io_state_out_2_0, f0_round_2_p_io_state_out_1_4,
         f0_round_2_p_io_state_out_1_3, f0_round_2_p_io_state_out_1_2,
         f0_round_2_p_io_state_out_1_1, f0_round_2_p_io_state_out_1_0,
         f0_round_2_p_io_state_out_0_4, f0_round_2_p_io_state_out_0_3,
         f0_round_2_p_io_state_out_0_2, f0_round_2_p_io_state_out_0_1,
         f0_round_2_p_io_state_out_0_0, f0_round_2_t_n25, f0_round_2_t_n24,
         f0_round_2_t_n23, f0_round_2_t_n22, f0_round_2_t_n21,
         f0_round_2_t_n20, f0_round_2_t_n19, f0_round_2_t_n18,
         f0_round_2_t_n17, f0_round_2_t_n16, f0_round_2_t_n15,
         f0_round_2_t_n14, f0_round_2_t_n13, f0_round_2_t_n12,
         f0_round_2_t_n11, f0_round_2_t_n10, f0_round_2_t_n9, f0_round_2_t_n8,
         f0_round_2_t_n7, f0_round_2_t_n6, f0_round_2_t_n5, f0_round_2_t_n4,
         f0_round_2_t_n3, f0_round_2_t_n2, f0_round_2_t_n1, f0_round_2_c_n25,
         f0_round_2_c_n24, f0_round_2_c_n23, f0_round_2_c_n22,
         f0_round_2_c_n21, f0_round_2_c_n20, f0_round_2_c_n19,
         f0_round_2_c_n18, f0_round_2_c_n17, f0_round_2_c_n16,
         f0_round_2_c_n15, f0_round_2_c_n14, f0_round_2_c_n13,
         f0_round_2_c_n12, f0_round_2_c_n11, f0_round_2_c_n10, f0_round_2_c_n9,
         f0_round_2_c_n8, f0_round_2_c_n7, f0_round_2_c_n6, f0_round_2_c_n5,
         f0_round_2_c_n4, f0_round_2_c_n3, f0_round_2_c_n2, f0_round_2_c_n1,
         f0_round_3_c_io_state_out_0_0, f0_round_3_p_io_state_out_4_4,
         f0_round_3_p_io_state_out_4_3, f0_round_3_p_io_state_out_4_2,
         f0_round_3_p_io_state_out_4_1, f0_round_3_p_io_state_out_4_0,
         f0_round_3_p_io_state_out_3_4, f0_round_3_p_io_state_out_3_3,
         f0_round_3_p_io_state_out_3_2, f0_round_3_p_io_state_out_3_1,
         f0_round_3_p_io_state_out_3_0, f0_round_3_p_io_state_out_2_4,
         f0_round_3_p_io_state_out_2_3, f0_round_3_p_io_state_out_2_2,
         f0_round_3_p_io_state_out_2_1, f0_round_3_p_io_state_out_2_0,
         f0_round_3_p_io_state_out_1_4, f0_round_3_p_io_state_out_1_3,
         f0_round_3_p_io_state_out_1_2, f0_round_3_p_io_state_out_1_1,
         f0_round_3_p_io_state_out_1_0, f0_round_3_p_io_state_out_0_4,
         f0_round_3_p_io_state_out_0_3, f0_round_3_p_io_state_out_0_2,
         f0_round_3_p_io_state_out_0_1, f0_round_3_p_io_state_out_0_0,
         f0_round_3_t_n25, f0_round_3_t_n24, f0_round_3_t_n23,
         f0_round_3_t_n22, f0_round_3_t_n21, f0_round_3_t_n20,
         f0_round_3_t_n19, f0_round_3_t_n18, f0_round_3_t_n17,
         f0_round_3_t_n16, f0_round_3_t_n15, f0_round_3_t_n14,
         f0_round_3_t_n13, f0_round_3_t_n12, f0_round_3_t_n11,
         f0_round_3_t_n10, f0_round_3_t_n9, f0_round_3_t_n8, f0_round_3_t_n7,
         f0_round_3_t_n6, f0_round_3_t_n5, f0_round_3_t_n4, f0_round_3_t_n3,
         f0_round_3_t_n2, f0_round_3_t_n1, f0_round_3_c_n25, f0_round_3_c_n24,
         f0_round_3_c_n23, f0_round_3_c_n22, f0_round_3_c_n21,
         f0_round_3_c_n20, f0_round_3_c_n19, f0_round_3_c_n18,
         f0_round_3_c_n17, f0_round_3_c_n16, f0_round_3_c_n15,
         f0_round_3_c_n14, f0_round_3_c_n13, f0_round_3_c_n12,
         f0_round_3_c_n11, f0_round_3_c_n10, f0_round_3_c_n9, f0_round_3_c_n8,
         f0_round_3_c_n7, f0_round_3_c_n6, f0_round_3_c_n5, f0_round_3_c_n4,
         f0_round_3_c_n3, f0_round_3_c_n2, f0_round_3_c_n1,
         f0_round_4_c_io_state_out_0_0, f0_round_4_p_io_state_out_4_4,
         f0_round_4_p_io_state_out_4_3, f0_round_4_p_io_state_out_4_2,
         f0_round_4_p_io_state_out_4_1, f0_round_4_p_io_state_out_4_0,
         f0_round_4_p_io_state_out_3_4, f0_round_4_p_io_state_out_3_3,
         f0_round_4_p_io_state_out_3_2, f0_round_4_p_io_state_out_3_1,
         f0_round_4_p_io_state_out_3_0, f0_round_4_p_io_state_out_2_4,
         f0_round_4_p_io_state_out_2_3, f0_round_4_p_io_state_out_2_2,
         f0_round_4_p_io_state_out_2_1, f0_round_4_p_io_state_out_2_0,
         f0_round_4_p_io_state_out_1_4, f0_round_4_p_io_state_out_1_3,
         f0_round_4_p_io_state_out_1_2, f0_round_4_p_io_state_out_1_1,
         f0_round_4_p_io_state_out_1_0, f0_round_4_p_io_state_out_0_4,
         f0_round_4_p_io_state_out_0_3, f0_round_4_p_io_state_out_0_2,
         f0_round_4_p_io_state_out_0_1, f0_round_4_p_io_state_out_0_0,
         f0_round_4_t_n25, f0_round_4_t_n24, f0_round_4_t_n23,
         f0_round_4_t_n22, f0_round_4_t_n21, f0_round_4_t_n20,
         f0_round_4_t_n19, f0_round_4_t_n18, f0_round_4_t_n17,
         f0_round_4_t_n16, f0_round_4_t_n15, f0_round_4_t_n14,
         f0_round_4_t_n13, f0_round_4_t_n12, f0_round_4_t_n11,
         f0_round_4_t_n10, f0_round_4_t_n9, f0_round_4_t_n8, f0_round_4_t_n7,
         f0_round_4_t_n6, f0_round_4_t_n5, f0_round_4_t_n4, f0_round_4_t_n3,
         f0_round_4_t_n2, f0_round_4_t_n1, f0_round_4_c_n25, f0_round_4_c_n24,
         f0_round_4_c_n23, f0_round_4_c_n22, f0_round_4_c_n21,
         f0_round_4_c_n20, f0_round_4_c_n19, f0_round_4_c_n18,
         f0_round_4_c_n17, f0_round_4_c_n16, f0_round_4_c_n15,
         f0_round_4_c_n14, f0_round_4_c_n13, f0_round_4_c_n12,
         f0_round_4_c_n11, f0_round_4_c_n10, f0_round_4_c_n9, f0_round_4_c_n8,
         f0_round_4_c_n7, f0_round_4_c_n6, f0_round_4_c_n5, f0_round_4_c_n4,
         f0_round_4_c_n3, f0_round_4_c_n2, f0_round_4_c_n1,
         f0_round_5_c_io_state_out_0_0, f0_round_5_p_io_state_out_4_4,
         f0_round_5_p_io_state_out_4_3, f0_round_5_p_io_state_out_4_2,
         f0_round_5_p_io_state_out_4_1, f0_round_5_p_io_state_out_4_0,
         f0_round_5_p_io_state_out_3_4, f0_round_5_p_io_state_out_3_3,
         f0_round_5_p_io_state_out_3_2, f0_round_5_p_io_state_out_3_1,
         f0_round_5_p_io_state_out_3_0, f0_round_5_p_io_state_out_2_4,
         f0_round_5_p_io_state_out_2_3, f0_round_5_p_io_state_out_2_2,
         f0_round_5_p_io_state_out_2_1, f0_round_5_p_io_state_out_2_0,
         f0_round_5_p_io_state_out_1_4, f0_round_5_p_io_state_out_1_3,
         f0_round_5_p_io_state_out_1_2, f0_round_5_p_io_state_out_1_1,
         f0_round_5_p_io_state_out_1_0, f0_round_5_p_io_state_out_0_4,
         f0_round_5_p_io_state_out_0_3, f0_round_5_p_io_state_out_0_2,
         f0_round_5_p_io_state_out_0_1, f0_round_5_p_io_state_out_0_0,
         f0_round_5_t_n25, f0_round_5_t_n24, f0_round_5_t_n23,
         f0_round_5_t_n22, f0_round_5_t_n21, f0_round_5_t_n20,
         f0_round_5_t_n19, f0_round_5_t_n18, f0_round_5_t_n17,
         f0_round_5_t_n16, f0_round_5_t_n15, f0_round_5_t_n14,
         f0_round_5_t_n13, f0_round_5_t_n12, f0_round_5_t_n11,
         f0_round_5_t_n10, f0_round_5_t_n9, f0_round_5_t_n8, f0_round_5_t_n7,
         f0_round_5_t_n6, f0_round_5_t_n5, f0_round_5_t_n4, f0_round_5_t_n3,
         f0_round_5_t_n2, f0_round_5_t_n1, f0_round_5_c_n25, f0_round_5_c_n24,
         f0_round_5_c_n23, f0_round_5_c_n22, f0_round_5_c_n21,
         f0_round_5_c_n20, f0_round_5_c_n19, f0_round_5_c_n18,
         f0_round_5_c_n17, f0_round_5_c_n16, f0_round_5_c_n15,
         f0_round_5_c_n14, f0_round_5_c_n13, f0_round_5_c_n12,
         f0_round_5_c_n11, f0_round_5_c_n10, f0_round_5_c_n9, f0_round_5_c_n8,
         f0_round_5_c_n7, f0_round_5_c_n6, f0_round_5_c_n5, f0_round_5_c_n4,
         f0_round_5_c_n3, f0_round_5_c_n2, f0_round_5_c_n1,
         f0_round_6_c_io_state_out_0_0, f0_round_6_p_io_state_out_4_4,
         f0_round_6_p_io_state_out_4_3, f0_round_6_p_io_state_out_4_2,
         f0_round_6_p_io_state_out_4_1, f0_round_6_p_io_state_out_4_0,
         f0_round_6_p_io_state_out_3_4, f0_round_6_p_io_state_out_3_3,
         f0_round_6_p_io_state_out_3_2, f0_round_6_p_io_state_out_3_1,
         f0_round_6_p_io_state_out_3_0, f0_round_6_p_io_state_out_2_4,
         f0_round_6_p_io_state_out_2_3, f0_round_6_p_io_state_out_2_2,
         f0_round_6_p_io_state_out_2_1, f0_round_6_p_io_state_out_2_0,
         f0_round_6_p_io_state_out_1_4, f0_round_6_p_io_state_out_1_3,
         f0_round_6_p_io_state_out_1_2, f0_round_6_p_io_state_out_1_1,
         f0_round_6_p_io_state_out_1_0, f0_round_6_p_io_state_out_0_4,
         f0_round_6_p_io_state_out_0_3, f0_round_6_p_io_state_out_0_2,
         f0_round_6_p_io_state_out_0_1, f0_round_6_p_io_state_out_0_0,
         f0_round_6_t_n25, f0_round_6_t_n24, f0_round_6_t_n23,
         f0_round_6_t_n22, f0_round_6_t_n21, f0_round_6_t_n20,
         f0_round_6_t_n19, f0_round_6_t_n18, f0_round_6_t_n17,
         f0_round_6_t_n16, f0_round_6_t_n15, f0_round_6_t_n14,
         f0_round_6_t_n13, f0_round_6_t_n12, f0_round_6_t_n11,
         f0_round_6_t_n10, f0_round_6_t_n9, f0_round_6_t_n8, f0_round_6_t_n7,
         f0_round_6_t_n6, f0_round_6_t_n5, f0_round_6_t_n4, f0_round_6_t_n3,
         f0_round_6_t_n2, f0_round_6_t_n1, f0_round_6_c_n25, f0_round_6_c_n24,
         f0_round_6_c_n23, f0_round_6_c_n22, f0_round_6_c_n21,
         f0_round_6_c_n20, f0_round_6_c_n19, f0_round_6_c_n18,
         f0_round_6_c_n17, f0_round_6_c_n16, f0_round_6_c_n15,
         f0_round_6_c_n14, f0_round_6_c_n13, f0_round_6_c_n12,
         f0_round_6_c_n11, f0_round_6_c_n10, f0_round_6_c_n9, f0_round_6_c_n8,
         f0_round_6_c_n7, f0_round_6_c_n6, f0_round_6_c_n5, f0_round_6_c_n4,
         f0_round_6_c_n3, f0_round_6_c_n2, f0_round_6_c_n1,
         f0_round_7_p_io_state_out_4_4, f0_round_7_p_io_state_out_4_3,
         f0_round_7_p_io_state_out_4_2, f0_round_7_p_io_state_out_4_1,
         f0_round_7_p_io_state_out_4_0, f0_round_7_p_io_state_out_3_4,
         f0_round_7_p_io_state_out_3_3, f0_round_7_p_io_state_out_3_2,
         f0_round_7_p_io_state_out_3_1, f0_round_7_p_io_state_out_3_0,
         f0_round_7_p_io_state_out_2_4, f0_round_7_p_io_state_out_2_3,
         f0_round_7_p_io_state_out_2_2, f0_round_7_p_io_state_out_2_1,
         f0_round_7_p_io_state_out_2_0, f0_round_7_p_io_state_out_1_4,
         f0_round_7_p_io_state_out_1_3, f0_round_7_p_io_state_out_1_2,
         f0_round_7_p_io_state_out_1_1, f0_round_7_p_io_state_out_1_0,
         f0_round_7_p_io_state_out_0_4, f0_round_7_p_io_state_out_0_3,
         f0_round_7_p_io_state_out_0_2, f0_round_7_p_io_state_out_0_1,
         f0_round_7_p_io_state_out_0_0, f0_round_7_t_n25, f0_round_7_t_n24,
         f0_round_7_t_n23, f0_round_7_t_n22, f0_round_7_t_n21,
         f0_round_7_t_n20, f0_round_7_t_n19, f0_round_7_t_n18,
         f0_round_7_t_n17, f0_round_7_t_n16, f0_round_7_t_n15,
         f0_round_7_t_n14, f0_round_7_t_n13, f0_round_7_t_n12,
         f0_round_7_t_n11, f0_round_7_t_n10, f0_round_7_t_n9, f0_round_7_t_n8,
         f0_round_7_t_n7, f0_round_7_t_n6, f0_round_7_t_n5, f0_round_7_t_n4,
         f0_round_7_t_n3, f0_round_7_t_n2, f0_round_7_t_n1, f0_round_7_c_n25,
         f0_round_7_c_n24, f0_round_7_c_n23, f0_round_7_c_n22,
         f0_round_7_c_n21, f0_round_7_c_n20, f0_round_7_c_n19,
         f0_round_7_c_n18, f0_round_7_c_n17, f0_round_7_c_n16,
         f0_round_7_c_n15, f0_round_7_c_n14, f0_round_7_c_n13,
         f0_round_7_c_n12, f0_round_7_c_n11, f0_round_7_c_n10, f0_round_7_c_n9,
         f0_round_7_c_n8, f0_round_7_c_n7, f0_round_7_c_n6, f0_round_7_c_n5,
         f0_round_7_c_n4, f0_round_7_c_n3, f0_round_7_c_n2, f0_round_7_c_n1,
         f0_round_8_p_io_state_out_4_4, f0_round_8_p_io_state_out_4_3,
         f0_round_8_p_io_state_out_4_2, f0_round_8_p_io_state_out_4_1,
         f0_round_8_p_io_state_out_4_0, f0_round_8_p_io_state_out_3_4,
         f0_round_8_p_io_state_out_3_3, f0_round_8_p_io_state_out_3_2,
         f0_round_8_p_io_state_out_3_1, f0_round_8_p_io_state_out_3_0,
         f0_round_8_p_io_state_out_2_4, f0_round_8_p_io_state_out_2_3,
         f0_round_8_p_io_state_out_2_2, f0_round_8_p_io_state_out_2_1,
         f0_round_8_p_io_state_out_2_0, f0_round_8_p_io_state_out_1_4,
         f0_round_8_p_io_state_out_1_3, f0_round_8_p_io_state_out_1_2,
         f0_round_8_p_io_state_out_1_1, f0_round_8_p_io_state_out_1_0,
         f0_round_8_p_io_state_out_0_4, f0_round_8_p_io_state_out_0_3,
         f0_round_8_p_io_state_out_0_2, f0_round_8_p_io_state_out_0_1,
         f0_round_8_p_io_state_out_0_0, f0_round_8_t_n25, f0_round_8_t_n24,
         f0_round_8_t_n23, f0_round_8_t_n22, f0_round_8_t_n21,
         f0_round_8_t_n20, f0_round_8_t_n19, f0_round_8_t_n18,
         f0_round_8_t_n17, f0_round_8_t_n16, f0_round_8_t_n15,
         f0_round_8_t_n14, f0_round_8_t_n13, f0_round_8_t_n12,
         f0_round_8_t_n11, f0_round_8_t_n10, f0_round_8_t_n9, f0_round_8_t_n8,
         f0_round_8_t_n7, f0_round_8_t_n6, f0_round_8_t_n5, f0_round_8_t_n4,
         f0_round_8_t_n3, f0_round_8_t_n2, f0_round_8_t_n1, f0_round_8_c_n25,
         f0_round_8_c_n24, f0_round_8_c_n23, f0_round_8_c_n22,
         f0_round_8_c_n21, f0_round_8_c_n20, f0_round_8_c_n19,
         f0_round_8_c_n18, f0_round_8_c_n17, f0_round_8_c_n16,
         f0_round_8_c_n15, f0_round_8_c_n14, f0_round_8_c_n13,
         f0_round_8_c_n12, f0_round_8_c_n11, f0_round_8_c_n10, f0_round_8_c_n9,
         f0_round_8_c_n8, f0_round_8_c_n7, f0_round_8_c_n6, f0_round_8_c_n5,
         f0_round_8_c_n4, f0_round_8_c_n3, f0_round_8_c_n2, f0_round_8_c_n1,
         f0_round_9_c_io_state_out_0_0, f0_round_9_p_io_state_out_4_4,
         f0_round_9_p_io_state_out_4_3, f0_round_9_p_io_state_out_4_2,
         f0_round_9_p_io_state_out_4_1, f0_round_9_p_io_state_out_4_0,
         f0_round_9_p_io_state_out_3_4, f0_round_9_p_io_state_out_3_3,
         f0_round_9_p_io_state_out_3_2, f0_round_9_p_io_state_out_3_1,
         f0_round_9_p_io_state_out_3_0, f0_round_9_p_io_state_out_2_4,
         f0_round_9_p_io_state_out_2_3, f0_round_9_p_io_state_out_2_2,
         f0_round_9_p_io_state_out_2_1, f0_round_9_p_io_state_out_2_0,
         f0_round_9_p_io_state_out_1_4, f0_round_9_p_io_state_out_1_3,
         f0_round_9_p_io_state_out_1_2, f0_round_9_p_io_state_out_1_1,
         f0_round_9_p_io_state_out_1_0, f0_round_9_p_io_state_out_0_4,
         f0_round_9_p_io_state_out_0_3, f0_round_9_p_io_state_out_0_2,
         f0_round_9_p_io_state_out_0_1, f0_round_9_p_io_state_out_0_0,
         f0_round_9_t_n25, f0_round_9_t_n24, f0_round_9_t_n23,
         f0_round_9_t_n22, f0_round_9_t_n21, f0_round_9_t_n20,
         f0_round_9_t_n19, f0_round_9_t_n18, f0_round_9_t_n17,
         f0_round_9_t_n16, f0_round_9_t_n15, f0_round_9_t_n14,
         f0_round_9_t_n13, f0_round_9_t_n12, f0_round_9_t_n11,
         f0_round_9_t_n10, f0_round_9_t_n9, f0_round_9_t_n8, f0_round_9_t_n7,
         f0_round_9_t_n6, f0_round_9_t_n5, f0_round_9_t_n4, f0_round_9_t_n3,
         f0_round_9_t_n2, f0_round_9_t_n1, f0_round_9_c_n25, f0_round_9_c_n24,
         f0_round_9_c_n23, f0_round_9_c_n22, f0_round_9_c_n21,
         f0_round_9_c_n20, f0_round_9_c_n19, f0_round_9_c_n18,
         f0_round_9_c_n17, f0_round_9_c_n16, f0_round_9_c_n15,
         f0_round_9_c_n14, f0_round_9_c_n13, f0_round_9_c_n12,
         f0_round_9_c_n11, f0_round_9_c_n10, f0_round_9_c_n9, f0_round_9_c_n8,
         f0_round_9_c_n7, f0_round_9_c_n6, f0_round_9_c_n5, f0_round_9_c_n4,
         f0_round_9_c_n3, f0_round_9_c_n2, f0_round_9_c_n1,
         f0_round_10_p_io_state_out_4_4, f0_round_10_p_io_state_out_4_3,
         f0_round_10_p_io_state_out_4_2, f0_round_10_p_io_state_out_4_1,
         f0_round_10_p_io_state_out_4_0, f0_round_10_p_io_state_out_3_4,
         f0_round_10_p_io_state_out_3_3, f0_round_10_p_io_state_out_3_2,
         f0_round_10_p_io_state_out_3_1, f0_round_10_p_io_state_out_3_0,
         f0_round_10_p_io_state_out_2_4, f0_round_10_p_io_state_out_2_3,
         f0_round_10_p_io_state_out_2_2, f0_round_10_p_io_state_out_2_1,
         f0_round_10_p_io_state_out_2_0, f0_round_10_p_io_state_out_1_4,
         f0_round_10_p_io_state_out_1_3, f0_round_10_p_io_state_out_1_2,
         f0_round_10_p_io_state_out_1_1, f0_round_10_p_io_state_out_1_0,
         f0_round_10_p_io_state_out_0_4, f0_round_10_p_io_state_out_0_3,
         f0_round_10_p_io_state_out_0_2, f0_round_10_p_io_state_out_0_1,
         f0_round_10_p_io_state_out_0_0, f0_round_10_t_n25, f0_round_10_t_n24,
         f0_round_10_t_n23, f0_round_10_t_n22, f0_round_10_t_n21,
         f0_round_10_t_n20, f0_round_10_t_n19, f0_round_10_t_n18,
         f0_round_10_t_n17, f0_round_10_t_n16, f0_round_10_t_n15,
         f0_round_10_t_n14, f0_round_10_t_n13, f0_round_10_t_n12,
         f0_round_10_t_n11, f0_round_10_t_n10, f0_round_10_t_n9,
         f0_round_10_t_n8, f0_round_10_t_n7, f0_round_10_t_n6,
         f0_round_10_t_n5, f0_round_10_t_n4, f0_round_10_t_n3,
         f0_round_10_t_n2, f0_round_10_t_n1, f0_round_10_c_n25,
         f0_round_10_c_n24, f0_round_10_c_n23, f0_round_10_c_n22,
         f0_round_10_c_n21, f0_round_10_c_n20, f0_round_10_c_n19,
         f0_round_10_c_n18, f0_round_10_c_n17, f0_round_10_c_n16,
         f0_round_10_c_n15, f0_round_10_c_n14, f0_round_10_c_n13,
         f0_round_10_c_n12, f0_round_10_c_n11, f0_round_10_c_n10,
         f0_round_10_c_n9, f0_round_10_c_n8, f0_round_10_c_n7,
         f0_round_10_c_n6, f0_round_10_c_n5, f0_round_10_c_n4,
         f0_round_10_c_n3, f0_round_10_c_n2, f0_round_10_c_n1,
         f1_round_10_io_state_out_4_4, f1_round_10_io_state_out_4_3,
         f1_round_10_io_state_out_4_2, f1_round_10_io_state_out_4_1,
         f1_round_10_io_state_out_4_0, f1_round_10_io_state_out_3_4,
         f1_round_10_io_state_out_3_3, f1_round_10_io_state_out_3_2,
         f1_round_10_io_state_out_3_1, f1_round_10_io_state_out_3_0,
         f1_round_10_io_state_out_2_4, f1_round_10_io_state_out_2_3,
         f1_round_10_io_state_out_2_2, f1_round_10_io_state_out_2_1,
         f1_round_10_io_state_out_2_0, f1_round_10_io_state_out_1_4,
         f1_round_10_io_state_out_1_3, f1_round_10_io_state_out_1_2,
         f1_round_10_io_state_out_1_1, f1_round_10_io_state_out_1_0,
         f1_round_10_io_state_out_0_4, f1_round_10_io_state_out_0_3,
         f1_round_10_io_state_out_0_2, f1_round_10_io_state_out_0_1,
         f1_round_10_io_state_out_0_0, f1_round_9_io_state_out_4_4,
         f1_round_9_io_state_out_4_3, f1_round_9_io_state_out_4_2,
         f1_round_9_io_state_out_4_1, f1_round_9_io_state_out_4_0,
         f1_round_9_io_state_out_3_4, f1_round_9_io_state_out_3_3,
         f1_round_9_io_state_out_3_2, f1_round_9_io_state_out_3_1,
         f1_round_9_io_state_out_3_0, f1_round_9_io_state_out_2_4,
         f1_round_9_io_state_out_2_3, f1_round_9_io_state_out_2_2,
         f1_round_9_io_state_out_2_1, f1_round_9_io_state_out_2_0,
         f1_round_9_io_state_out_1_4, f1_round_9_io_state_out_1_3,
         f1_round_9_io_state_out_1_2, f1_round_9_io_state_out_1_1,
         f1_round_9_io_state_out_1_0, f1_round_9_io_state_out_0_4,
         f1_round_9_io_state_out_0_3, f1_round_9_io_state_out_0_2,
         f1_round_9_io_state_out_0_1, f1_round_9_io_state_out_0_0,
         f1_round_8_io_state_out_4_4, f1_round_8_io_state_out_4_3,
         f1_round_8_io_state_out_4_2, f1_round_8_io_state_out_4_1,
         f1_round_8_io_state_out_4_0, f1_round_8_io_state_out_3_4,
         f1_round_8_io_state_out_3_3, f1_round_8_io_state_out_3_2,
         f1_round_8_io_state_out_3_1, f1_round_8_io_state_out_3_0,
         f1_round_8_io_state_out_2_4, f1_round_8_io_state_out_2_3,
         f1_round_8_io_state_out_2_2, f1_round_8_io_state_out_2_1,
         f1_round_8_io_state_out_2_0, f1_round_8_io_state_out_1_4,
         f1_round_8_io_state_out_1_3, f1_round_8_io_state_out_1_2,
         f1_round_8_io_state_out_1_1, f1_round_8_io_state_out_1_0,
         f1_round_8_io_state_out_0_4, f1_round_8_io_state_out_0_3,
         f1_round_8_io_state_out_0_2, f1_round_8_io_state_out_0_1,
         f1_round_8_io_state_out_0_0, f1_round_7_io_state_out_4_4,
         f1_round_7_io_state_out_4_3, f1_round_7_io_state_out_4_2,
         f1_round_7_io_state_out_4_1, f1_round_7_io_state_out_4_0,
         f1_round_7_io_state_out_3_4, f1_round_7_io_state_out_3_3,
         f1_round_7_io_state_out_3_2, f1_round_7_io_state_out_3_1,
         f1_round_7_io_state_out_3_0, f1_round_7_io_state_out_2_4,
         f1_round_7_io_state_out_2_3, f1_round_7_io_state_out_2_2,
         f1_round_7_io_state_out_2_1, f1_round_7_io_state_out_2_0,
         f1_round_7_io_state_out_1_4, f1_round_7_io_state_out_1_3,
         f1_round_7_io_state_out_1_2, f1_round_7_io_state_out_1_1,
         f1_round_7_io_state_out_1_0, f1_round_7_io_state_out_0_4,
         f1_round_7_io_state_out_0_3, f1_round_7_io_state_out_0_2,
         f1_round_7_io_state_out_0_1, f1_round_7_io_state_out_0_0,
         f1_round_6_io_state_out_4_4, f1_round_6_io_state_out_4_3,
         f1_round_6_io_state_out_4_2, f1_round_6_io_state_out_4_1,
         f1_round_6_io_state_out_4_0, f1_round_6_io_state_out_3_4,
         f1_round_6_io_state_out_3_3, f1_round_6_io_state_out_3_2,
         f1_round_6_io_state_out_3_1, f1_round_6_io_state_out_3_0,
         f1_round_6_io_state_out_2_4, f1_round_6_io_state_out_2_3,
         f1_round_6_io_state_out_2_2, f1_round_6_io_state_out_2_1,
         f1_round_6_io_state_out_2_0, f1_round_6_io_state_out_1_4,
         f1_round_6_io_state_out_1_3, f1_round_6_io_state_out_1_2,
         f1_round_6_io_state_out_1_1, f1_round_6_io_state_out_1_0,
         f1_round_6_io_state_out_0_4, f1_round_6_io_state_out_0_3,
         f1_round_6_io_state_out_0_2, f1_round_6_io_state_out_0_1,
         f1_round_6_io_state_out_0_0, f1_round_5_io_state_out_4_4,
         f1_round_5_io_state_out_4_3, f1_round_5_io_state_out_4_2,
         f1_round_5_io_state_out_4_1, f1_round_5_io_state_out_4_0,
         f1_round_5_io_state_out_3_4, f1_round_5_io_state_out_3_3,
         f1_round_5_io_state_out_3_2, f1_round_5_io_state_out_3_1,
         f1_round_5_io_state_out_3_0, f1_round_5_io_state_out_2_4,
         f1_round_5_io_state_out_2_3, f1_round_5_io_state_out_2_2,
         f1_round_5_io_state_out_2_1, f1_round_5_io_state_out_2_0,
         f1_round_5_io_state_out_1_4, f1_round_5_io_state_out_1_3,
         f1_round_5_io_state_out_1_2, f1_round_5_io_state_out_1_1,
         f1_round_5_io_state_out_1_0, f1_round_5_io_state_out_0_4,
         f1_round_5_io_state_out_0_3, f1_round_5_io_state_out_0_2,
         f1_round_5_io_state_out_0_1, f1_round_5_io_state_out_0_0,
         f1_round_4_io_state_out_4_4, f1_round_4_io_state_out_4_3,
         f1_round_4_io_state_out_4_2, f1_round_4_io_state_out_4_1,
         f1_round_4_io_state_out_4_0, f1_round_4_io_state_out_3_4,
         f1_round_4_io_state_out_3_3, f1_round_4_io_state_out_3_2,
         f1_round_4_io_state_out_3_1, f1_round_4_io_state_out_3_0,
         f1_round_4_io_state_out_2_4, f1_round_4_io_state_out_2_3,
         f1_round_4_io_state_out_2_2, f1_round_4_io_state_out_2_1,
         f1_round_4_io_state_out_2_0, f1_round_4_io_state_out_1_4,
         f1_round_4_io_state_out_1_3, f1_round_4_io_state_out_1_2,
         f1_round_4_io_state_out_1_1, f1_round_4_io_state_out_1_0,
         f1_round_4_io_state_out_0_4, f1_round_4_io_state_out_0_3,
         f1_round_4_io_state_out_0_2, f1_round_4_io_state_out_0_1,
         f1_round_4_io_state_out_0_0, f1_round_3_io_state_out_4_4,
         f1_round_3_io_state_out_4_3, f1_round_3_io_state_out_4_2,
         f1_round_3_io_state_out_4_1, f1_round_3_io_state_out_4_0,
         f1_round_3_io_state_out_3_4, f1_round_3_io_state_out_3_3,
         f1_round_3_io_state_out_3_2, f1_round_3_io_state_out_3_1,
         f1_round_3_io_state_out_3_0, f1_round_3_io_state_out_2_4,
         f1_round_3_io_state_out_2_3, f1_round_3_io_state_out_2_2,
         f1_round_3_io_state_out_2_1, f1_round_3_io_state_out_2_0,
         f1_round_3_io_state_out_1_4, f1_round_3_io_state_out_1_3,
         f1_round_3_io_state_out_1_2, f1_round_3_io_state_out_1_1,
         f1_round_3_io_state_out_1_0, f1_round_3_io_state_out_0_4,
         f1_round_3_io_state_out_0_3, f1_round_3_io_state_out_0_2,
         f1_round_3_io_state_out_0_1, f1_round_3_io_state_out_0_0,
         f1_round_2_io_state_out_4_4, f1_round_2_io_state_out_4_3,
         f1_round_2_io_state_out_4_2, f1_round_2_io_state_out_4_1,
         f1_round_2_io_state_out_4_0, f1_round_2_io_state_out_3_4,
         f1_round_2_io_state_out_3_3, f1_round_2_io_state_out_3_2,
         f1_round_2_io_state_out_3_1, f1_round_2_io_state_out_3_0,
         f1_round_2_io_state_out_2_4, f1_round_2_io_state_out_2_3,
         f1_round_2_io_state_out_2_2, f1_round_2_io_state_out_2_1,
         f1_round_2_io_state_out_2_0, f1_round_2_io_state_out_1_4,
         f1_round_2_io_state_out_1_3, f1_round_2_io_state_out_1_2,
         f1_round_2_io_state_out_1_1, f1_round_2_io_state_out_1_0,
         f1_round_2_io_state_out_0_4, f1_round_2_io_state_out_0_3,
         f1_round_2_io_state_out_0_2, f1_round_2_io_state_out_0_1,
         f1_round_2_io_state_out_0_0, f1_round_1_io_state_out_4_4,
         f1_round_1_io_state_out_4_3, f1_round_1_io_state_out_4_2,
         f1_round_1_io_state_out_4_1, f1_round_1_io_state_out_4_0,
         f1_round_1_io_state_out_3_4, f1_round_1_io_state_out_3_3,
         f1_round_1_io_state_out_3_2, f1_round_1_io_state_out_3_1,
         f1_round_1_io_state_out_3_0, f1_round_1_io_state_out_2_4,
         f1_round_1_io_state_out_2_3, f1_round_1_io_state_out_2_2,
         f1_round_1_io_state_out_2_1, f1_round_1_io_state_out_2_0,
         f1_round_1_io_state_out_1_4, f1_round_1_io_state_out_1_3,
         f1_round_1_io_state_out_1_2, f1_round_1_io_state_out_1_1,
         f1_round_1_io_state_out_1_0, f1_round_1_io_state_out_0_4,
         f1_round_1_io_state_out_0_3, f1_round_1_io_state_out_0_2,
         f1_round_1_io_state_out_0_1, f1_round_1_io_state_out_0_0,
         f1_round_io_state_out_4_4, f1_round_io_state_out_4_3,
         f1_round_io_state_out_4_2, f1_round_io_state_out_4_1,
         f1_round_io_state_out_4_0, f1_round_io_state_out_3_4,
         f1_round_io_state_out_3_3, f1_round_io_state_out_3_2,
         f1_round_io_state_out_3_1, f1_round_io_state_out_3_0,
         f1_round_io_state_out_2_4, f1_round_io_state_out_2_3,
         f1_round_io_state_out_2_2, f1_round_io_state_out_2_1,
         f1_round_io_state_out_2_0, f1_round_io_state_out_1_4,
         f1_round_io_state_out_1_3, f1_round_io_state_out_1_2,
         f1_round_io_state_out_1_1, f1_round_io_state_out_1_0,
         f1_round_io_state_out_0_4, f1_round_io_state_out_0_3,
         f1_round_io_state_out_0_2, f1_round_io_state_out_0_1,
         f1_round_io_state_out_0_0, f1_round_c_io_state_out_0_0,
         f1_round_p_io_state_out_4_4, f1_round_p_io_state_out_4_3,
         f1_round_p_io_state_out_4_2, f1_round_p_io_state_out_4_1,
         f1_round_p_io_state_out_4_0, f1_round_p_io_state_out_3_4,
         f1_round_p_io_state_out_3_3, f1_round_p_io_state_out_3_2,
         f1_round_p_io_state_out_3_1, f1_round_p_io_state_out_3_0,
         f1_round_p_io_state_out_2_4, f1_round_p_io_state_out_2_3,
         f1_round_p_io_state_out_2_2, f1_round_p_io_state_out_2_1,
         f1_round_p_io_state_out_2_0, f1_round_p_io_state_out_1_4,
         f1_round_p_io_state_out_1_3, f1_round_p_io_state_out_1_2,
         f1_round_p_io_state_out_1_1, f1_round_p_io_state_out_1_0,
         f1_round_p_io_state_out_0_4, f1_round_p_io_state_out_0_3,
         f1_round_p_io_state_out_0_2, f1_round_p_io_state_out_0_1,
         f1_round_p_io_state_out_0_0, f1_round_t_n25, f1_round_t_n24,
         f1_round_t_n23, f1_round_t_n22, f1_round_t_n21, f1_round_t_n20,
         f1_round_t_n19, f1_round_t_n18, f1_round_t_n17, f1_round_t_n16,
         f1_round_t_n15, f1_round_t_n14, f1_round_t_n13, f1_round_t_n12,
         f1_round_t_n11, f1_round_t_n10, f1_round_t_n9, f1_round_t_n8,
         f1_round_t_n7, f1_round_t_n6, f1_round_t_n5, f1_round_t_n4,
         f1_round_t_n3, f1_round_t_n2, f1_round_t_n1, f1_round_c_n25,
         f1_round_c_n24, f1_round_c_n23, f1_round_c_n22, f1_round_c_n21,
         f1_round_c_n20, f1_round_c_n19, f1_round_c_n18, f1_round_c_n17,
         f1_round_c_n16, f1_round_c_n15, f1_round_c_n14, f1_round_c_n13,
         f1_round_c_n12, f1_round_c_n11, f1_round_c_n10, f1_round_c_n9,
         f1_round_c_n8, f1_round_c_n7, f1_round_c_n6, f1_round_c_n5,
         f1_round_c_n4, f1_round_c_n3, f1_round_c_n2, f1_round_c_n1,
         f1_round_1_p_io_state_out_4_4, f1_round_1_p_io_state_out_4_3,
         f1_round_1_p_io_state_out_4_2, f1_round_1_p_io_state_out_4_1,
         f1_round_1_p_io_state_out_4_0, f1_round_1_p_io_state_out_3_4,
         f1_round_1_p_io_state_out_3_3, f1_round_1_p_io_state_out_3_2,
         f1_round_1_p_io_state_out_3_1, f1_round_1_p_io_state_out_3_0,
         f1_round_1_p_io_state_out_2_4, f1_round_1_p_io_state_out_2_3,
         f1_round_1_p_io_state_out_2_2, f1_round_1_p_io_state_out_2_1,
         f1_round_1_p_io_state_out_2_0, f1_round_1_p_io_state_out_1_4,
         f1_round_1_p_io_state_out_1_3, f1_round_1_p_io_state_out_1_2,
         f1_round_1_p_io_state_out_1_1, f1_round_1_p_io_state_out_1_0,
         f1_round_1_p_io_state_out_0_4, f1_round_1_p_io_state_out_0_3,
         f1_round_1_p_io_state_out_0_2, f1_round_1_p_io_state_out_0_1,
         f1_round_1_p_io_state_out_0_0, f1_round_1_t_n25, f1_round_1_t_n24,
         f1_round_1_t_n23, f1_round_1_t_n22, f1_round_1_t_n21,
         f1_round_1_t_n20, f1_round_1_t_n19, f1_round_1_t_n18,
         f1_round_1_t_n17, f1_round_1_t_n16, f1_round_1_t_n15,
         f1_round_1_t_n14, f1_round_1_t_n13, f1_round_1_t_n12,
         f1_round_1_t_n11, f1_round_1_t_n10, f1_round_1_t_n9, f1_round_1_t_n8,
         f1_round_1_t_n7, f1_round_1_t_n6, f1_round_1_t_n5, f1_round_1_t_n4,
         f1_round_1_t_n3, f1_round_1_t_n2, f1_round_1_t_n1, f1_round_1_c_n25,
         f1_round_1_c_n24, f1_round_1_c_n23, f1_round_1_c_n22,
         f1_round_1_c_n21, f1_round_1_c_n20, f1_round_1_c_n19,
         f1_round_1_c_n18, f1_round_1_c_n17, f1_round_1_c_n16,
         f1_round_1_c_n15, f1_round_1_c_n14, f1_round_1_c_n13,
         f1_round_1_c_n12, f1_round_1_c_n11, f1_round_1_c_n10, f1_round_1_c_n9,
         f1_round_1_c_n8, f1_round_1_c_n7, f1_round_1_c_n6, f1_round_1_c_n5,
         f1_round_1_c_n4, f1_round_1_c_n3, f1_round_1_c_n2, f1_round_1_c_n1,
         f1_round_2_p_io_state_out_4_4, f1_round_2_p_io_state_out_4_3,
         f1_round_2_p_io_state_out_4_2, f1_round_2_p_io_state_out_4_1,
         f1_round_2_p_io_state_out_4_0, f1_round_2_p_io_state_out_3_4,
         f1_round_2_p_io_state_out_3_3, f1_round_2_p_io_state_out_3_2,
         f1_round_2_p_io_state_out_3_1, f1_round_2_p_io_state_out_3_0,
         f1_round_2_p_io_state_out_2_4, f1_round_2_p_io_state_out_2_3,
         f1_round_2_p_io_state_out_2_2, f1_round_2_p_io_state_out_2_1,
         f1_round_2_p_io_state_out_2_0, f1_round_2_p_io_state_out_1_4,
         f1_round_2_p_io_state_out_1_3, f1_round_2_p_io_state_out_1_2,
         f1_round_2_p_io_state_out_1_1, f1_round_2_p_io_state_out_1_0,
         f1_round_2_p_io_state_out_0_4, f1_round_2_p_io_state_out_0_3,
         f1_round_2_p_io_state_out_0_2, f1_round_2_p_io_state_out_0_1,
         f1_round_2_p_io_state_out_0_0, f1_round_2_t_n25, f1_round_2_t_n24,
         f1_round_2_t_n23, f1_round_2_t_n22, f1_round_2_t_n21,
         f1_round_2_t_n20, f1_round_2_t_n19, f1_round_2_t_n18,
         f1_round_2_t_n17, f1_round_2_t_n16, f1_round_2_t_n15,
         f1_round_2_t_n14, f1_round_2_t_n13, f1_round_2_t_n12,
         f1_round_2_t_n11, f1_round_2_t_n10, f1_round_2_t_n9, f1_round_2_t_n8,
         f1_round_2_t_n7, f1_round_2_t_n6, f1_round_2_t_n5, f1_round_2_t_n4,
         f1_round_2_t_n3, f1_round_2_t_n2, f1_round_2_t_n1, f1_round_2_c_n25,
         f1_round_2_c_n24, f1_round_2_c_n23, f1_round_2_c_n22,
         f1_round_2_c_n21, f1_round_2_c_n20, f1_round_2_c_n19,
         f1_round_2_c_n18, f1_round_2_c_n17, f1_round_2_c_n16,
         f1_round_2_c_n15, f1_round_2_c_n14, f1_round_2_c_n13,
         f1_round_2_c_n12, f1_round_2_c_n11, f1_round_2_c_n10, f1_round_2_c_n9,
         f1_round_2_c_n8, f1_round_2_c_n7, f1_round_2_c_n6, f1_round_2_c_n5,
         f1_round_2_c_n4, f1_round_2_c_n3, f1_round_2_c_n2, f1_round_2_c_n1,
         f1_round_3_p_io_state_out_4_4, f1_round_3_p_io_state_out_4_3,
         f1_round_3_p_io_state_out_4_2, f1_round_3_p_io_state_out_4_1,
         f1_round_3_p_io_state_out_4_0, f1_round_3_p_io_state_out_3_4,
         f1_round_3_p_io_state_out_3_3, f1_round_3_p_io_state_out_3_2,
         f1_round_3_p_io_state_out_3_1, f1_round_3_p_io_state_out_3_0,
         f1_round_3_p_io_state_out_2_4, f1_round_3_p_io_state_out_2_3,
         f1_round_3_p_io_state_out_2_2, f1_round_3_p_io_state_out_2_1,
         f1_round_3_p_io_state_out_2_0, f1_round_3_p_io_state_out_1_4,
         f1_round_3_p_io_state_out_1_3, f1_round_3_p_io_state_out_1_2,
         f1_round_3_p_io_state_out_1_1, f1_round_3_p_io_state_out_1_0,
         f1_round_3_p_io_state_out_0_4, f1_round_3_p_io_state_out_0_3,
         f1_round_3_p_io_state_out_0_2, f1_round_3_p_io_state_out_0_1,
         f1_round_3_p_io_state_out_0_0, f1_round_3_t_n25, f1_round_3_t_n24,
         f1_round_3_t_n23, f1_round_3_t_n22, f1_round_3_t_n21,
         f1_round_3_t_n20, f1_round_3_t_n19, f1_round_3_t_n18,
         f1_round_3_t_n17, f1_round_3_t_n16, f1_round_3_t_n15,
         f1_round_3_t_n14, f1_round_3_t_n13, f1_round_3_t_n12,
         f1_round_3_t_n11, f1_round_3_t_n10, f1_round_3_t_n9, f1_round_3_t_n8,
         f1_round_3_t_n7, f1_round_3_t_n6, f1_round_3_t_n5, f1_round_3_t_n4,
         f1_round_3_t_n3, f1_round_3_t_n2, f1_round_3_t_n1, f1_round_3_c_n25,
         f1_round_3_c_n24, f1_round_3_c_n23, f1_round_3_c_n22,
         f1_round_3_c_n21, f1_round_3_c_n20, f1_round_3_c_n19,
         f1_round_3_c_n18, f1_round_3_c_n17, f1_round_3_c_n16,
         f1_round_3_c_n15, f1_round_3_c_n14, f1_round_3_c_n13,
         f1_round_3_c_n12, f1_round_3_c_n11, f1_round_3_c_n10, f1_round_3_c_n9,
         f1_round_3_c_n8, f1_round_3_c_n7, f1_round_3_c_n6, f1_round_3_c_n5,
         f1_round_3_c_n4, f1_round_3_c_n3, f1_round_3_c_n2, f1_round_3_c_n1,
         f1_round_4_c_io_state_out_0_0, f1_round_4_p_io_state_out_4_4,
         f1_round_4_p_io_state_out_4_3, f1_round_4_p_io_state_out_4_2,
         f1_round_4_p_io_state_out_4_1, f1_round_4_p_io_state_out_4_0,
         f1_round_4_p_io_state_out_3_4, f1_round_4_p_io_state_out_3_3,
         f1_round_4_p_io_state_out_3_2, f1_round_4_p_io_state_out_3_1,
         f1_round_4_p_io_state_out_3_0, f1_round_4_p_io_state_out_2_4,
         f1_round_4_p_io_state_out_2_3, f1_round_4_p_io_state_out_2_2,
         f1_round_4_p_io_state_out_2_1, f1_round_4_p_io_state_out_2_0,
         f1_round_4_p_io_state_out_1_4, f1_round_4_p_io_state_out_1_3,
         f1_round_4_p_io_state_out_1_2, f1_round_4_p_io_state_out_1_1,
         f1_round_4_p_io_state_out_1_0, f1_round_4_p_io_state_out_0_4,
         f1_round_4_p_io_state_out_0_3, f1_round_4_p_io_state_out_0_2,
         f1_round_4_p_io_state_out_0_1, f1_round_4_p_io_state_out_0_0,
         f1_round_4_t_n25, f1_round_4_t_n24, f1_round_4_t_n23,
         f1_round_4_t_n22, f1_round_4_t_n21, f1_round_4_t_n20,
         f1_round_4_t_n19, f1_round_4_t_n18, f1_round_4_t_n17,
         f1_round_4_t_n16, f1_round_4_t_n15, f1_round_4_t_n14,
         f1_round_4_t_n13, f1_round_4_t_n12, f1_round_4_t_n11,
         f1_round_4_t_n10, f1_round_4_t_n9, f1_round_4_t_n8, f1_round_4_t_n7,
         f1_round_4_t_n6, f1_round_4_t_n5, f1_round_4_t_n4, f1_round_4_t_n3,
         f1_round_4_t_n2, f1_round_4_t_n1, f1_round_4_c_n25, f1_round_4_c_n24,
         f1_round_4_c_n23, f1_round_4_c_n22, f1_round_4_c_n21,
         f1_round_4_c_n20, f1_round_4_c_n19, f1_round_4_c_n18,
         f1_round_4_c_n17, f1_round_4_c_n16, f1_round_4_c_n15,
         f1_round_4_c_n14, f1_round_4_c_n13, f1_round_4_c_n12,
         f1_round_4_c_n11, f1_round_4_c_n10, f1_round_4_c_n9, f1_round_4_c_n8,
         f1_round_4_c_n7, f1_round_4_c_n6, f1_round_4_c_n5, f1_round_4_c_n4,
         f1_round_4_c_n3, f1_round_4_c_n2, f1_round_4_c_n1,
         f1_round_5_c_io_state_out_0_0, f1_round_5_p_io_state_out_4_4,
         f1_round_5_p_io_state_out_4_3, f1_round_5_p_io_state_out_4_2,
         f1_round_5_p_io_state_out_4_1, f1_round_5_p_io_state_out_4_0,
         f1_round_5_p_io_state_out_3_4, f1_round_5_p_io_state_out_3_3,
         f1_round_5_p_io_state_out_3_2, f1_round_5_p_io_state_out_3_1,
         f1_round_5_p_io_state_out_3_0, f1_round_5_p_io_state_out_2_4,
         f1_round_5_p_io_state_out_2_3, f1_round_5_p_io_state_out_2_2,
         f1_round_5_p_io_state_out_2_1, f1_round_5_p_io_state_out_2_0,
         f1_round_5_p_io_state_out_1_4, f1_round_5_p_io_state_out_1_3,
         f1_round_5_p_io_state_out_1_2, f1_round_5_p_io_state_out_1_1,
         f1_round_5_p_io_state_out_1_0, f1_round_5_p_io_state_out_0_4,
         f1_round_5_p_io_state_out_0_3, f1_round_5_p_io_state_out_0_2,
         f1_round_5_p_io_state_out_0_1, f1_round_5_p_io_state_out_0_0,
         f1_round_5_t_n25, f1_round_5_t_n24, f1_round_5_t_n23,
         f1_round_5_t_n22, f1_round_5_t_n21, f1_round_5_t_n20,
         f1_round_5_t_n19, f1_round_5_t_n18, f1_round_5_t_n17,
         f1_round_5_t_n16, f1_round_5_t_n15, f1_round_5_t_n14,
         f1_round_5_t_n13, f1_round_5_t_n12, f1_round_5_t_n11,
         f1_round_5_t_n10, f1_round_5_t_n9, f1_round_5_t_n8, f1_round_5_t_n7,
         f1_round_5_t_n6, f1_round_5_t_n5, f1_round_5_t_n4, f1_round_5_t_n3,
         f1_round_5_t_n2, f1_round_5_t_n1, f1_round_5_c_n25, f1_round_5_c_n24,
         f1_round_5_c_n23, f1_round_5_c_n22, f1_round_5_c_n21,
         f1_round_5_c_n20, f1_round_5_c_n19, f1_round_5_c_n18,
         f1_round_5_c_n17, f1_round_5_c_n16, f1_round_5_c_n15,
         f1_round_5_c_n14, f1_round_5_c_n13, f1_round_5_c_n12,
         f1_round_5_c_n11, f1_round_5_c_n10, f1_round_5_c_n9, f1_round_5_c_n8,
         f1_round_5_c_n7, f1_round_5_c_n6, f1_round_5_c_n5, f1_round_5_c_n4,
         f1_round_5_c_n3, f1_round_5_c_n2, f1_round_5_c_n1,
         f1_round_6_c_io_state_out_0_0, f1_round_6_p_io_state_out_4_4,
         f1_round_6_p_io_state_out_4_3, f1_round_6_p_io_state_out_4_2,
         f1_round_6_p_io_state_out_4_1, f1_round_6_p_io_state_out_4_0,
         f1_round_6_p_io_state_out_3_4, f1_round_6_p_io_state_out_3_3,
         f1_round_6_p_io_state_out_3_2, f1_round_6_p_io_state_out_3_1,
         f1_round_6_p_io_state_out_3_0, f1_round_6_p_io_state_out_2_4,
         f1_round_6_p_io_state_out_2_3, f1_round_6_p_io_state_out_2_2,
         f1_round_6_p_io_state_out_2_1, f1_round_6_p_io_state_out_2_0,
         f1_round_6_p_io_state_out_1_4, f1_round_6_p_io_state_out_1_3,
         f1_round_6_p_io_state_out_1_2, f1_round_6_p_io_state_out_1_1,
         f1_round_6_p_io_state_out_1_0, f1_round_6_p_io_state_out_0_4,
         f1_round_6_p_io_state_out_0_3, f1_round_6_p_io_state_out_0_2,
         f1_round_6_p_io_state_out_0_1, f1_round_6_p_io_state_out_0_0,
         f1_round_6_t_n25, f1_round_6_t_n24, f1_round_6_t_n23,
         f1_round_6_t_n22, f1_round_6_t_n21, f1_round_6_t_n20,
         f1_round_6_t_n19, f1_round_6_t_n18, f1_round_6_t_n17,
         f1_round_6_t_n16, f1_round_6_t_n15, f1_round_6_t_n14,
         f1_round_6_t_n13, f1_round_6_t_n12, f1_round_6_t_n11,
         f1_round_6_t_n10, f1_round_6_t_n9, f1_round_6_t_n8, f1_round_6_t_n7,
         f1_round_6_t_n6, f1_round_6_t_n5, f1_round_6_t_n4, f1_round_6_t_n3,
         f1_round_6_t_n2, f1_round_6_t_n1, f1_round_6_c_n25, f1_round_6_c_n24,
         f1_round_6_c_n23, f1_round_6_c_n22, f1_round_6_c_n21,
         f1_round_6_c_n20, f1_round_6_c_n19, f1_round_6_c_n18,
         f1_round_6_c_n17, f1_round_6_c_n16, f1_round_6_c_n15,
         f1_round_6_c_n14, f1_round_6_c_n13, f1_round_6_c_n12,
         f1_round_6_c_n11, f1_round_6_c_n10, f1_round_6_c_n9, f1_round_6_c_n8,
         f1_round_6_c_n7, f1_round_6_c_n6, f1_round_6_c_n5, f1_round_6_c_n4,
         f1_round_6_c_n3, f1_round_6_c_n2, f1_round_6_c_n1,
         f1_round_7_c_io_state_out_0_0, f1_round_7_p_io_state_out_4_4,
         f1_round_7_p_io_state_out_4_3, f1_round_7_p_io_state_out_4_2,
         f1_round_7_p_io_state_out_4_1, f1_round_7_p_io_state_out_4_0,
         f1_round_7_p_io_state_out_3_4, f1_round_7_p_io_state_out_3_3,
         f1_round_7_p_io_state_out_3_2, f1_round_7_p_io_state_out_3_1,
         f1_round_7_p_io_state_out_3_0, f1_round_7_p_io_state_out_2_4,
         f1_round_7_p_io_state_out_2_3, f1_round_7_p_io_state_out_2_2,
         f1_round_7_p_io_state_out_2_1, f1_round_7_p_io_state_out_2_0,
         f1_round_7_p_io_state_out_1_4, f1_round_7_p_io_state_out_1_3,
         f1_round_7_p_io_state_out_1_2, f1_round_7_p_io_state_out_1_1,
         f1_round_7_p_io_state_out_1_0, f1_round_7_p_io_state_out_0_4,
         f1_round_7_p_io_state_out_0_3, f1_round_7_p_io_state_out_0_2,
         f1_round_7_p_io_state_out_0_1, f1_round_7_p_io_state_out_0_0,
         f1_round_7_t_n25, f1_round_7_t_n24, f1_round_7_t_n23,
         f1_round_7_t_n22, f1_round_7_t_n21, f1_round_7_t_n20,
         f1_round_7_t_n19, f1_round_7_t_n18, f1_round_7_t_n17,
         f1_round_7_t_n16, f1_round_7_t_n15, f1_round_7_t_n14,
         f1_round_7_t_n13, f1_round_7_t_n12, f1_round_7_t_n11,
         f1_round_7_t_n10, f1_round_7_t_n9, f1_round_7_t_n8, f1_round_7_t_n7,
         f1_round_7_t_n6, f1_round_7_t_n5, f1_round_7_t_n4, f1_round_7_t_n3,
         f1_round_7_t_n2, f1_round_7_t_n1, f1_round_7_c_n25, f1_round_7_c_n24,
         f1_round_7_c_n23, f1_round_7_c_n22, f1_round_7_c_n21,
         f1_round_7_c_n20, f1_round_7_c_n19, f1_round_7_c_n18,
         f1_round_7_c_n17, f1_round_7_c_n16, f1_round_7_c_n15,
         f1_round_7_c_n14, f1_round_7_c_n13, f1_round_7_c_n12,
         f1_round_7_c_n11, f1_round_7_c_n10, f1_round_7_c_n9, f1_round_7_c_n8,
         f1_round_7_c_n7, f1_round_7_c_n6, f1_round_7_c_n5, f1_round_7_c_n4,
         f1_round_7_c_n3, f1_round_7_c_n2, f1_round_7_c_n1,
         f1_round_8_p_io_state_out_4_4, f1_round_8_p_io_state_out_4_3,
         f1_round_8_p_io_state_out_4_2, f1_round_8_p_io_state_out_4_1,
         f1_round_8_p_io_state_out_4_0, f1_round_8_p_io_state_out_3_4,
         f1_round_8_p_io_state_out_3_3, f1_round_8_p_io_state_out_3_2,
         f1_round_8_p_io_state_out_3_1, f1_round_8_p_io_state_out_3_0,
         f1_round_8_p_io_state_out_2_4, f1_round_8_p_io_state_out_2_3,
         f1_round_8_p_io_state_out_2_2, f1_round_8_p_io_state_out_2_1,
         f1_round_8_p_io_state_out_2_0, f1_round_8_p_io_state_out_1_4,
         f1_round_8_p_io_state_out_1_3, f1_round_8_p_io_state_out_1_2,
         f1_round_8_p_io_state_out_1_1, f1_round_8_p_io_state_out_1_0,
         f1_round_8_p_io_state_out_0_4, f1_round_8_p_io_state_out_0_3,
         f1_round_8_p_io_state_out_0_2, f1_round_8_p_io_state_out_0_1,
         f1_round_8_p_io_state_out_0_0, f1_round_8_t_n25, f1_round_8_t_n24,
         f1_round_8_t_n23, f1_round_8_t_n22, f1_round_8_t_n21,
         f1_round_8_t_n20, f1_round_8_t_n19, f1_round_8_t_n18,
         f1_round_8_t_n17, f1_round_8_t_n16, f1_round_8_t_n15,
         f1_round_8_t_n14, f1_round_8_t_n13, f1_round_8_t_n12,
         f1_round_8_t_n11, f1_round_8_t_n10, f1_round_8_t_n9, f1_round_8_t_n8,
         f1_round_8_t_n7, f1_round_8_t_n6, f1_round_8_t_n5, f1_round_8_t_n4,
         f1_round_8_t_n3, f1_round_8_t_n2, f1_round_8_t_n1, f1_round_8_c_n25,
         f1_round_8_c_n24, f1_round_8_c_n23, f1_round_8_c_n22,
         f1_round_8_c_n21, f1_round_8_c_n20, f1_round_8_c_n19,
         f1_round_8_c_n18, f1_round_8_c_n17, f1_round_8_c_n16,
         f1_round_8_c_n15, f1_round_8_c_n14, f1_round_8_c_n13,
         f1_round_8_c_n12, f1_round_8_c_n11, f1_round_8_c_n10, f1_round_8_c_n9,
         f1_round_8_c_n8, f1_round_8_c_n7, f1_round_8_c_n6, f1_round_8_c_n5,
         f1_round_8_c_n4, f1_round_8_c_n3, f1_round_8_c_n2, f1_round_8_c_n1,
         f1_round_9_p_io_state_out_4_4, f1_round_9_p_io_state_out_4_3,
         f1_round_9_p_io_state_out_4_2, f1_round_9_p_io_state_out_4_1,
         f1_round_9_p_io_state_out_4_0, f1_round_9_p_io_state_out_3_4,
         f1_round_9_p_io_state_out_3_3, f1_round_9_p_io_state_out_3_2,
         f1_round_9_p_io_state_out_3_1, f1_round_9_p_io_state_out_3_0,
         f1_round_9_p_io_state_out_2_4, f1_round_9_p_io_state_out_2_3,
         f1_round_9_p_io_state_out_2_2, f1_round_9_p_io_state_out_2_1,
         f1_round_9_p_io_state_out_2_0, f1_round_9_p_io_state_out_1_4,
         f1_round_9_p_io_state_out_1_3, f1_round_9_p_io_state_out_1_2,
         f1_round_9_p_io_state_out_1_1, f1_round_9_p_io_state_out_1_0,
         f1_round_9_p_io_state_out_0_4, f1_round_9_p_io_state_out_0_3,
         f1_round_9_p_io_state_out_0_2, f1_round_9_p_io_state_out_0_1,
         f1_round_9_p_io_state_out_0_0, f1_round_9_t_n25, f1_round_9_t_n24,
         f1_round_9_t_n23, f1_round_9_t_n22, f1_round_9_t_n21,
         f1_round_9_t_n20, f1_round_9_t_n19, f1_round_9_t_n18,
         f1_round_9_t_n17, f1_round_9_t_n16, f1_round_9_t_n15,
         f1_round_9_t_n14, f1_round_9_t_n13, f1_round_9_t_n12,
         f1_round_9_t_n11, f1_round_9_t_n10, f1_round_9_t_n9, f1_round_9_t_n8,
         f1_round_9_t_n7, f1_round_9_t_n6, f1_round_9_t_n5, f1_round_9_t_n4,
         f1_round_9_t_n3, f1_round_9_t_n2, f1_round_9_t_n1, f1_round_9_c_n25,
         f1_round_9_c_n24, f1_round_9_c_n23, f1_round_9_c_n22,
         f1_round_9_c_n21, f1_round_9_c_n20, f1_round_9_c_n19,
         f1_round_9_c_n18, f1_round_9_c_n17, f1_round_9_c_n16,
         f1_round_9_c_n15, f1_round_9_c_n14, f1_round_9_c_n13,
         f1_round_9_c_n12, f1_round_9_c_n11, f1_round_9_c_n10, f1_round_9_c_n9,
         f1_round_9_c_n8, f1_round_9_c_n7, f1_round_9_c_n6, f1_round_9_c_n5,
         f1_round_9_c_n4, f1_round_9_c_n3, f1_round_9_c_n2, f1_round_9_c_n1,
         f1_round_10_c_io_state_out_0_0, f1_round_10_p_io_state_out_4_4,
         f1_round_10_p_io_state_out_4_3, f1_round_10_p_io_state_out_4_2,
         f1_round_10_p_io_state_out_4_1, f1_round_10_p_io_state_out_4_0,
         f1_round_10_p_io_state_out_3_4, f1_round_10_p_io_state_out_3_3,
         f1_round_10_p_io_state_out_3_2, f1_round_10_p_io_state_out_3_1,
         f1_round_10_p_io_state_out_3_0, f1_round_10_p_io_state_out_2_4,
         f1_round_10_p_io_state_out_2_3, f1_round_10_p_io_state_out_2_2,
         f1_round_10_p_io_state_out_2_1, f1_round_10_p_io_state_out_2_0,
         f1_round_10_p_io_state_out_1_4, f1_round_10_p_io_state_out_1_3,
         f1_round_10_p_io_state_out_1_2, f1_round_10_p_io_state_out_1_1,
         f1_round_10_p_io_state_out_1_0, f1_round_10_p_io_state_out_0_4,
         f1_round_10_p_io_state_out_0_3, f1_round_10_p_io_state_out_0_2,
         f1_round_10_p_io_state_out_0_1, f1_round_10_p_io_state_out_0_0,
         f1_round_10_t_n25, f1_round_10_t_n24, f1_round_10_t_n23,
         f1_round_10_t_n22, f1_round_10_t_n21, f1_round_10_t_n20,
         f1_round_10_t_n19, f1_round_10_t_n18, f1_round_10_t_n17,
         f1_round_10_t_n16, f1_round_10_t_n15, f1_round_10_t_n14,
         f1_round_10_t_n13, f1_round_10_t_n12, f1_round_10_t_n11,
         f1_round_10_t_n10, f1_round_10_t_n9, f1_round_10_t_n8,
         f1_round_10_t_n7, f1_round_10_t_n6, f1_round_10_t_n5,
         f1_round_10_t_n4, f1_round_10_t_n3, f1_round_10_t_n2,
         f1_round_10_t_n1, f1_round_10_c_n25, f1_round_10_c_n24,
         f1_round_10_c_n23, f1_round_10_c_n22, f1_round_10_c_n21,
         f1_round_10_c_n20, f1_round_10_c_n19, f1_round_10_c_n18,
         f1_round_10_c_n17, f1_round_10_c_n16, f1_round_10_c_n15,
         f1_round_10_c_n14, f1_round_10_c_n13, f1_round_10_c_n12,
         f1_round_10_c_n11, f1_round_10_c_n10, f1_round_10_c_n9,
         f1_round_10_c_n8, f1_round_10_c_n7, f1_round_10_c_n6,
         f1_round_10_c_n5, f1_round_10_c_n4, f1_round_10_c_n3,
         f1_round_10_c_n2, f1_round_10_c_n1, f1_round_11_c_io_state_out_4_4,
         f1_round_11_c_io_state_out_4_3, f1_round_11_c_io_state_out_4_2,
         f1_round_11_c_io_state_out_3_4, f1_round_11_c_io_state_out_3_3,
         f1_round_11_c_io_state_out_3_2, f1_round_11_c_io_state_out_2_4,
         f1_round_11_c_io_state_out_2_3, f1_round_11_c_io_state_out_2_2,
         f1_round_11_c_io_state_out_1_4, f1_round_11_c_io_state_out_1_3,
         f1_round_11_c_io_state_out_1_2, f1_round_11_c_io_state_out_0_4,
         f1_round_11_c_io_state_out_0_3, f1_round_11_c_io_state_out_0_2,
         f1_round_11_p_io_state_out_4_4, f1_round_11_p_io_state_out_4_3,
         f1_round_11_p_io_state_out_4_2, f1_round_11_p_io_state_out_4_1,
         f1_round_11_p_io_state_out_4_0, f1_round_11_p_io_state_out_3_4,
         f1_round_11_p_io_state_out_3_3, f1_round_11_p_io_state_out_3_2,
         f1_round_11_p_io_state_out_3_1, f1_round_11_p_io_state_out_3_0,
         f1_round_11_p_io_state_out_2_4, f1_round_11_p_io_state_out_2_3,
         f1_round_11_p_io_state_out_2_2, f1_round_11_p_io_state_out_2_1,
         f1_round_11_p_io_state_out_2_0, f1_round_11_p_io_state_out_1_4,
         f1_round_11_p_io_state_out_1_3, f1_round_11_p_io_state_out_1_2,
         f1_round_11_p_io_state_out_1_1, f1_round_11_p_io_state_out_1_0,
         f1_round_11_p_io_state_out_0_4, f1_round_11_p_io_state_out_0_3,
         f1_round_11_p_io_state_out_0_2, f1_round_11_p_io_state_out_0_1,
         f1_round_11_p_io_state_out_0_0, f1_round_11_t_n25, f1_round_11_t_n24,
         f1_round_11_t_n23, f1_round_11_t_n22, f1_round_11_t_n21,
         f1_round_11_t_n20, f1_round_11_t_n19, f1_round_11_t_n18,
         f1_round_11_t_n17, f1_round_11_t_n16, f1_round_11_t_n15,
         f1_round_11_t_n14, f1_round_11_t_n13, f1_round_11_t_n12,
         f1_round_11_t_n11, f1_round_11_t_n10, f1_round_11_t_n9,
         f1_round_11_t_n8, f1_round_11_t_n7, f1_round_11_t_n6,
         f1_round_11_t_n5, f1_round_11_t_n4, f1_round_11_t_n3,
         f1_round_11_t_n2, f1_round_11_t_n1, f1_round_11_c_n25,
         f1_round_11_c_n24, f1_round_11_c_n23, f1_round_11_c_n22,
         f1_round_11_c_n21, f1_round_11_c_n20, f1_round_11_c_n19,
         f1_round_11_c_n18, f1_round_11_c_n17, f1_round_11_c_n16,
         f1_round_11_c_n15, f1_round_11_c_n14, f1_round_11_c_n13,
         f1_round_11_c_n12, f1_round_11_c_n11, f1_round_11_c_n10,
         f1_round_11_c_n9, f1_round_11_c_n8, f1_round_11_c_n7,
         f1_round_11_c_n6, f1_round_11_c_n5, f1_round_11_c_n4,
         f1_round_11_c_n3, f1_round_11_c_n2, f1_round_11_c_n1;

  XNOR2_X1 f0_round0_t_U20 ( .A(io_block_i0[1]), .B(io_block_i0[6]), .ZN(
        f0_round0_t_n5) );
  XOR2_X1 f0_round0_t_U19 ( .A(io_block_i0[4]), .B(io_block_i0[9]), .Z(
        f0_round0_t_n3) );
  XOR2_X1 f0_round0_t_U18 ( .A(io_block_i0[0]), .B(
        f0_round0_p_io_state_out_2_1), .Z(f0_round0_p_io_state_out_0_0) );
  XOR2_X1 f0_round0_t_U17 ( .A(io_block_i0[5]), .B(
        f0_round0_p_io_state_out_2_1), .Z(f0_round0_p_io_state_out_1_3) );
  XOR2_X1 f0_round0_t_U16 ( .A(io_block_i0[2]), .B(io_block_i0[7]), .Z(
        f0_round0_t_n4) );
  XOR2_X1 f0_round0_t_U15 ( .A(io_block_i0[0]), .B(io_block_i0[5]), .Z(
        f0_round0_t_n1) );
  XOR2_X1 f0_round0_t_U14 ( .A(io_block_i0[1]), .B(
        f0_round0_p_io_state_out_2_3), .Z(f0_round0_p_io_state_out_0_2) );
  XOR2_X1 f0_round0_t_U13 ( .A(io_block_i0[6]), .B(
        f0_round0_p_io_state_out_2_3), .Z(f0_round0_p_io_state_out_1_0) );
  XOR2_X1 f0_round0_t_U12 ( .A(io_block_i0[3]), .B(io_block_i0[8]), .Z(
        f0_round0_t_n2) );
  XOR2_X1 f0_round0_t_U11 ( .A(io_block_i0[2]), .B(
        f0_round0_p_io_state_out_2_0), .Z(f0_round0_p_io_state_out_0_4) );
  XOR2_X1 f0_round0_t_U10 ( .A(io_block_i0[7]), .B(
        f0_round0_p_io_state_out_2_0), .Z(f0_round0_p_io_state_out_1_2) );
  XOR2_X1 f0_round0_t_U9 ( .A(io_block_i0[3]), .B(f0_round0_p_io_state_out_2_2), .Z(f0_round0_p_io_state_out_0_1) );
  XOR2_X1 f0_round0_t_U8 ( .A(io_block_i0[8]), .B(f0_round0_p_io_state_out_2_2), .Z(f0_round0_p_io_state_out_1_4) );
  XOR2_X1 f0_round0_t_U7 ( .A(io_block_i0[4]), .B(f0_round0_p_io_state_out_2_4), .Z(f0_round0_p_io_state_out_0_3) );
  XOR2_X1 f0_round0_t_U6 ( .A(io_block_i0[9]), .B(f0_round0_p_io_state_out_2_4), .Z(f0_round0_p_io_state_out_1_1) );
  XOR2_X2 f0_round0_t_U5 ( .A(f0_round0_t_n1), .B(f0_round0_t_n2), .Z(
        f0_round0_p_io_state_out_2_4) );
  XOR2_X2 f0_round0_t_U4 ( .A(f0_round0_t_n3), .B(f0_round0_t_n4), .Z(
        f0_round0_p_io_state_out_2_2) );
  XOR2_X2 f0_round0_t_U3 ( .A(f0_round0_t_n4), .B(f0_round0_t_n1), .Z(
        f0_round0_p_io_state_out_2_3) );
  XNOR2_X2 f0_round0_t_U2 ( .A(f0_round0_t_n5), .B(f0_round0_t_n3), .ZN(
        f0_round0_p_io_state_out_2_1) );
  XNOR2_X2 f0_round0_t_U1 ( .A(f0_round0_t_n5), .B(f0_round0_t_n2), .ZN(
        f0_round0_p_io_state_out_2_0) );
  NAND2_X1 f0_round0_c_U50 ( .A1(f0_round0_p_io_state_out_2_0), .A2(
        f0_round0_p_io_state_out_1_0), .ZN(f0_round0_c_n25) );
  XOR2_X1 f0_round0_c_U49 ( .A(f0_round0_c_n25), .B(
        f0_round0_p_io_state_out_0_0), .Z(f0_round0_c_io_state_out_0_0) );
  NAND2_X1 f0_round0_c_U48 ( .A1(f0_round0_p_io_state_out_2_1), .A2(
        f0_round0_p_io_state_out_1_1), .ZN(f0_round0_c_n24) );
  XOR2_X1 f0_round0_c_U47 ( .A(f0_round0_c_n24), .B(
        f0_round0_p_io_state_out_0_1), .Z(f0_round0_io_state_out_0_1) );
  NAND2_X1 f0_round0_c_U46 ( .A1(f0_round0_p_io_state_out_2_2), .A2(
        f0_round0_p_io_state_out_1_2), .ZN(f0_round0_c_n23) );
  XOR2_X1 f0_round0_c_U45 ( .A(f0_round0_c_n23), .B(
        f0_round0_p_io_state_out_0_2), .Z(f0_round0_io_state_out_0_2) );
  NAND2_X1 f0_round0_c_U44 ( .A1(f0_round0_p_io_state_out_2_3), .A2(
        f0_round0_p_io_state_out_1_3), .ZN(f0_round0_c_n22) );
  XOR2_X1 f0_round0_c_U43 ( .A(f0_round0_c_n22), .B(
        f0_round0_p_io_state_out_0_3), .Z(f0_round0_io_state_out_0_3) );
  NAND2_X1 f0_round0_c_U42 ( .A1(f0_round0_p_io_state_out_2_4), .A2(
        f0_round0_p_io_state_out_1_4), .ZN(f0_round0_c_n21) );
  XOR2_X1 f0_round0_c_U41 ( .A(f0_round0_c_n21), .B(
        f0_round0_p_io_state_out_0_4), .Z(f0_round0_io_state_out_0_4) );
  NAND2_X1 f0_round0_c_U40 ( .A1(f0_round0_p_io_state_out_2_0), .A2(
        f0_round0_p_io_state_out_2_2), .ZN(f0_round0_c_n20) );
  XOR2_X1 f0_round0_c_U39 ( .A(f0_round0_c_n20), .B(
        f0_round0_p_io_state_out_1_0), .Z(f0_round0_io_state_out_1_0) );
  NAND2_X1 f0_round0_c_U38 ( .A1(f0_round0_p_io_state_out_2_1), .A2(
        f0_round0_p_io_state_out_2_3), .ZN(f0_round0_c_n19) );
  XOR2_X1 f0_round0_c_U37 ( .A(f0_round0_c_n19), .B(
        f0_round0_p_io_state_out_1_1), .Z(f0_round0_io_state_out_1_1) );
  NAND2_X1 f0_round0_c_U36 ( .A1(f0_round0_p_io_state_out_2_2), .A2(
        f0_round0_p_io_state_out_2_4), .ZN(f0_round0_c_n18) );
  XOR2_X1 f0_round0_c_U35 ( .A(f0_round0_c_n18), .B(
        f0_round0_p_io_state_out_1_2), .Z(f0_round0_io_state_out_1_2) );
  NAND2_X1 f0_round0_c_U34 ( .A1(f0_round0_p_io_state_out_2_3), .A2(
        f0_round0_p_io_state_out_2_0), .ZN(f0_round0_c_n17) );
  XOR2_X1 f0_round0_c_U33 ( .A(f0_round0_c_n17), .B(
        f0_round0_p_io_state_out_1_3), .Z(f0_round0_io_state_out_1_3) );
  NAND2_X1 f0_round0_c_U32 ( .A1(f0_round0_p_io_state_out_2_4), .A2(
        f0_round0_p_io_state_out_2_1), .ZN(f0_round0_c_n16) );
  XOR2_X1 f0_round0_c_U31 ( .A(f0_round0_c_n16), .B(
        f0_round0_p_io_state_out_1_4), .Z(f0_round0_io_state_out_1_4) );
  NAND2_X1 f0_round0_c_U30 ( .A1(f0_round0_p_io_state_out_2_2), .A2(
        f0_round0_p_io_state_out_2_4), .ZN(f0_round0_c_n15) );
  XOR2_X1 f0_round0_c_U29 ( .A(f0_round0_c_n15), .B(
        f0_round0_p_io_state_out_2_0), .Z(f0_round0_io_state_out_2_0) );
  NAND2_X1 f0_round0_c_U28 ( .A1(f0_round0_p_io_state_out_2_3), .A2(
        f0_round0_p_io_state_out_2_0), .ZN(f0_round0_c_n14) );
  XOR2_X1 f0_round0_c_U27 ( .A(f0_round0_c_n14), .B(
        f0_round0_p_io_state_out_2_1), .Z(f0_round0_io_state_out_2_1) );
  NAND2_X1 f0_round0_c_U26 ( .A1(f0_round0_p_io_state_out_2_4), .A2(
        f0_round0_p_io_state_out_2_1), .ZN(f0_round0_c_n13) );
  XOR2_X1 f0_round0_c_U25 ( .A(f0_round0_c_n13), .B(
        f0_round0_p_io_state_out_2_2), .Z(f0_round0_io_state_out_2_2) );
  NAND2_X1 f0_round0_c_U24 ( .A1(f0_round0_p_io_state_out_2_0), .A2(
        f0_round0_p_io_state_out_2_2), .ZN(f0_round0_c_n12) );
  XOR2_X1 f0_round0_c_U23 ( .A(f0_round0_c_n12), .B(
        f0_round0_p_io_state_out_2_3), .Z(f0_round0_io_state_out_2_3) );
  NAND2_X1 f0_round0_c_U22 ( .A1(f0_round0_p_io_state_out_2_1), .A2(
        f0_round0_p_io_state_out_2_3), .ZN(f0_round0_c_n11) );
  XOR2_X1 f0_round0_c_U21 ( .A(f0_round0_c_n11), .B(
        f0_round0_p_io_state_out_2_4), .Z(f0_round0_io_state_out_2_4) );
  NAND2_X1 f0_round0_c_U20 ( .A1(f0_round0_p_io_state_out_2_4), .A2(
        f0_round0_p_io_state_out_0_0), .ZN(f0_round0_c_n10) );
  XOR2_X1 f0_round0_c_U19 ( .A(f0_round0_c_n10), .B(
        f0_round0_p_io_state_out_2_2), .Z(f0_round0_io_state_out_3_0) );
  NAND2_X1 f0_round0_c_U18 ( .A1(f0_round0_p_io_state_out_2_0), .A2(
        f0_round0_p_io_state_out_0_1), .ZN(f0_round0_c_n9) );
  XOR2_X1 f0_round0_c_U17 ( .A(f0_round0_c_n9), .B(
        f0_round0_p_io_state_out_2_3), .Z(f0_round0_io_state_out_3_1) );
  NAND2_X1 f0_round0_c_U16 ( .A1(f0_round0_p_io_state_out_2_1), .A2(
        f0_round0_p_io_state_out_0_2), .ZN(f0_round0_c_n8) );
  XOR2_X1 f0_round0_c_U15 ( .A(f0_round0_c_n8), .B(
        f0_round0_p_io_state_out_2_4), .Z(f0_round0_io_state_out_3_2) );
  NAND2_X1 f0_round0_c_U14 ( .A1(f0_round0_p_io_state_out_2_2), .A2(
        f0_round0_p_io_state_out_0_3), .ZN(f0_round0_c_n7) );
  XOR2_X1 f0_round0_c_U13 ( .A(f0_round0_c_n7), .B(
        f0_round0_p_io_state_out_2_0), .Z(f0_round0_io_state_out_3_3) );
  NAND2_X1 f0_round0_c_U12 ( .A1(f0_round0_p_io_state_out_2_3), .A2(
        f0_round0_p_io_state_out_0_4), .ZN(f0_round0_c_n6) );
  XOR2_X1 f0_round0_c_U11 ( .A(f0_round0_c_n6), .B(
        f0_round0_p_io_state_out_2_1), .Z(f0_round0_io_state_out_3_4) );
  NAND2_X1 f0_round0_c_U10 ( .A1(f0_round0_p_io_state_out_1_0), .A2(
        f0_round0_p_io_state_out_0_0), .ZN(f0_round0_c_n5) );
  XOR2_X1 f0_round0_c_U9 ( .A(f0_round0_c_n5), .B(f0_round0_p_io_state_out_2_4), .Z(f0_round0_io_state_out_4_0) );
  NAND2_X1 f0_round0_c_U8 ( .A1(f0_round0_p_io_state_out_1_1), .A2(
        f0_round0_p_io_state_out_0_1), .ZN(f0_round0_c_n4) );
  XOR2_X1 f0_round0_c_U7 ( .A(f0_round0_c_n4), .B(f0_round0_p_io_state_out_2_0), .Z(f0_round0_io_state_out_4_1) );
  NAND2_X1 f0_round0_c_U6 ( .A1(f0_round0_p_io_state_out_1_2), .A2(
        f0_round0_p_io_state_out_0_2), .ZN(f0_round0_c_n3) );
  XOR2_X1 f0_round0_c_U5 ( .A(f0_round0_c_n3), .B(f0_round0_p_io_state_out_2_1), .Z(f0_round0_io_state_out_4_2) );
  NAND2_X1 f0_round0_c_U4 ( .A1(f0_round0_p_io_state_out_1_3), .A2(
        f0_round0_p_io_state_out_0_3), .ZN(f0_round0_c_n2) );
  XOR2_X1 f0_round0_c_U3 ( .A(f0_round0_c_n2), .B(f0_round0_p_io_state_out_2_2), .Z(f0_round0_io_state_out_4_3) );
  NAND2_X1 f0_round0_c_U2 ( .A1(f0_round0_p_io_state_out_1_4), .A2(
        f0_round0_p_io_state_out_0_4), .ZN(f0_round0_c_n1) );
  XOR2_X1 f0_round0_c_U1 ( .A(f0_round0_c_n1), .B(f0_round0_p_io_state_out_2_3), .Z(f0_round0_io_state_out_4_4) );
  INV_X1 f0_round0_i_U1 ( .A(f0_round0_c_io_state_out_0_0), .ZN(
        f0_round0_io_state_out_0_0) );
  XOR2_X1 f0_round_t_U50 ( .A(f0_round0_io_state_out_1_4), .B(
        f0_round0_io_state_out_1_3), .Z(f0_round_t_n25) );
  XNOR2_X1 f0_round_t_U49 ( .A(f0_round0_io_state_out_1_2), .B(f0_round_t_n25), 
        .ZN(f0_round_t_n23) );
  XOR2_X1 f0_round_t_U48 ( .A(f0_round0_io_state_out_1_1), .B(
        f0_round0_io_state_out_1_0), .Z(f0_round_t_n24) );
  XOR2_X1 f0_round_t_U47 ( .A(f0_round_t_n23), .B(f0_round_t_n24), .Z(
        f0_round_t_n8) );
  XOR2_X1 f0_round_t_U46 ( .A(f0_round0_io_state_out_4_4), .B(
        f0_round0_io_state_out_4_3), .Z(f0_round_t_n22) );
  XNOR2_X1 f0_round_t_U45 ( .A(f0_round0_io_state_out_4_2), .B(f0_round_t_n22), 
        .ZN(f0_round_t_n20) );
  XOR2_X1 f0_round_t_U44 ( .A(f0_round0_io_state_out_4_1), .B(
        f0_round0_io_state_out_4_0), .Z(f0_round_t_n21) );
  XNOR2_X1 f0_round_t_U43 ( .A(f0_round_t_n20), .B(f0_round_t_n21), .ZN(
        f0_round_t_n5) );
  XNOR2_X1 f0_round_t_U42 ( .A(f0_round_t_n8), .B(f0_round_t_n5), .ZN(
        f0_round_t_n19) );
  XOR2_X1 f0_round_t_U41 ( .A(f0_round0_io_state_out_0_0), .B(f0_round_t_n19), 
        .Z(f0_round_p_io_state_out_0_0) );
  XOR2_X1 f0_round_t_U40 ( .A(f0_round0_io_state_out_0_1), .B(f0_round_t_n19), 
        .Z(f0_round_p_io_state_out_1_3) );
  XOR2_X1 f0_round_t_U39 ( .A(f0_round0_io_state_out_0_2), .B(f0_round_t_n19), 
        .Z(f0_round_p_io_state_out_2_1) );
  XOR2_X1 f0_round_t_U38 ( .A(f0_round0_io_state_out_0_3), .B(f0_round_t_n19), 
        .Z(f0_round_p_io_state_out_3_4) );
  XOR2_X1 f0_round_t_U37 ( .A(f0_round0_io_state_out_0_4), .B(f0_round_t_n19), 
        .Z(f0_round_p_io_state_out_4_2) );
  XOR2_X1 f0_round_t_U36 ( .A(f0_round0_io_state_out_2_4), .B(
        f0_round0_io_state_out_2_3), .Z(f0_round_t_n18) );
  XNOR2_X1 f0_round_t_U35 ( .A(f0_round0_io_state_out_2_2), .B(f0_round_t_n18), 
        .ZN(f0_round_t_n16) );
  XOR2_X1 f0_round_t_U34 ( .A(f0_round0_io_state_out_2_1), .B(
        f0_round0_io_state_out_2_0), .Z(f0_round_t_n17) );
  XNOR2_X1 f0_round_t_U33 ( .A(f0_round_t_n16), .B(f0_round_t_n17), .ZN(
        f0_round_t_n6) );
  XOR2_X1 f0_round_t_U32 ( .A(f0_round0_io_state_out_0_4), .B(
        f0_round0_io_state_out_0_3), .Z(f0_round_t_n15) );
  XNOR2_X1 f0_round_t_U31 ( .A(f0_round0_io_state_out_0_2), .B(f0_round_t_n15), 
        .ZN(f0_round_t_n13) );
  XOR2_X1 f0_round_t_U30 ( .A(f0_round0_io_state_out_0_1), .B(
        f0_round0_io_state_out_0_0), .Z(f0_round_t_n14) );
  XNOR2_X1 f0_round_t_U29 ( .A(f0_round_t_n13), .B(f0_round_t_n14), .ZN(
        f0_round_t_n2) );
  XOR2_X1 f0_round_t_U28 ( .A(f0_round_t_n6), .B(f0_round_t_n2), .Z(
        f0_round_t_n12) );
  XOR2_X1 f0_round_t_U27 ( .A(f0_round0_io_state_out_1_0), .B(f0_round_t_n12), 
        .Z(f0_round_p_io_state_out_0_2) );
  XOR2_X1 f0_round_t_U26 ( .A(f0_round0_io_state_out_1_1), .B(f0_round_t_n12), 
        .Z(f0_round_p_io_state_out_1_0) );
  XOR2_X1 f0_round_t_U25 ( .A(f0_round0_io_state_out_1_2), .B(f0_round_t_n12), 
        .Z(f0_round_p_io_state_out_2_3) );
  XOR2_X1 f0_round_t_U24 ( .A(f0_round0_io_state_out_1_3), .B(f0_round_t_n12), 
        .Z(f0_round_p_io_state_out_3_1) );
  XOR2_X1 f0_round_t_U23 ( .A(f0_round0_io_state_out_1_4), .B(f0_round_t_n12), 
        .Z(f0_round_p_io_state_out_4_4) );
  XOR2_X1 f0_round_t_U22 ( .A(f0_round0_io_state_out_3_4), .B(
        f0_round0_io_state_out_3_3), .Z(f0_round_t_n11) );
  XNOR2_X1 f0_round_t_U21 ( .A(f0_round0_io_state_out_3_2), .B(f0_round_t_n11), 
        .ZN(f0_round_t_n9) );
  XOR2_X1 f0_round_t_U20 ( .A(f0_round0_io_state_out_3_1), .B(
        f0_round0_io_state_out_3_0), .Z(f0_round_t_n10) );
  XNOR2_X1 f0_round_t_U19 ( .A(f0_round_t_n9), .B(f0_round_t_n10), .ZN(
        f0_round_t_n3) );
  XNOR2_X1 f0_round_t_U18 ( .A(f0_round_t_n8), .B(f0_round_t_n3), .ZN(
        f0_round_t_n7) );
  XOR2_X1 f0_round_t_U17 ( .A(f0_round0_io_state_out_2_0), .B(f0_round_t_n7), 
        .Z(f0_round_p_io_state_out_0_4) );
  XOR2_X1 f0_round_t_U16 ( .A(f0_round0_io_state_out_2_1), .B(f0_round_t_n7), 
        .Z(f0_round_p_io_state_out_1_2) );
  XOR2_X1 f0_round_t_U15 ( .A(f0_round0_io_state_out_2_2), .B(f0_round_t_n7), 
        .Z(f0_round_p_io_state_out_2_0) );
  XOR2_X1 f0_round_t_U14 ( .A(f0_round0_io_state_out_2_3), .B(f0_round_t_n7), 
        .Z(f0_round_p_io_state_out_3_3) );
  XOR2_X1 f0_round_t_U13 ( .A(f0_round0_io_state_out_2_4), .B(f0_round_t_n7), 
        .Z(f0_round_p_io_state_out_4_1) );
  XOR2_X1 f0_round_t_U12 ( .A(f0_round_t_n5), .B(f0_round_t_n6), .Z(
        f0_round_t_n4) );
  XOR2_X1 f0_round_t_U11 ( .A(f0_round0_io_state_out_3_0), .B(f0_round_t_n4), 
        .Z(f0_round_p_io_state_out_0_1) );
  XOR2_X1 f0_round_t_U10 ( .A(f0_round0_io_state_out_3_1), .B(f0_round_t_n4), 
        .Z(f0_round_p_io_state_out_1_4) );
  XOR2_X1 f0_round_t_U9 ( .A(f0_round0_io_state_out_3_2), .B(f0_round_t_n4), 
        .Z(f0_round_p_io_state_out_2_2) );
  XOR2_X1 f0_round_t_U8 ( .A(f0_round0_io_state_out_3_3), .B(f0_round_t_n4), 
        .Z(f0_round_p_io_state_out_3_0) );
  XOR2_X1 f0_round_t_U7 ( .A(f0_round0_io_state_out_3_4), .B(f0_round_t_n4), 
        .Z(f0_round_p_io_state_out_4_3) );
  XOR2_X1 f0_round_t_U6 ( .A(f0_round_t_n2), .B(f0_round_t_n3), .Z(
        f0_round_t_n1) );
  XOR2_X1 f0_round_t_U5 ( .A(f0_round0_io_state_out_4_0), .B(f0_round_t_n1), 
        .Z(f0_round_p_io_state_out_0_3) );
  XOR2_X1 f0_round_t_U4 ( .A(f0_round0_io_state_out_4_1), .B(f0_round_t_n1), 
        .Z(f0_round_p_io_state_out_1_1) );
  XOR2_X1 f0_round_t_U3 ( .A(f0_round0_io_state_out_4_2), .B(f0_round_t_n1), 
        .Z(f0_round_p_io_state_out_2_4) );
  XOR2_X1 f0_round_t_U2 ( .A(f0_round0_io_state_out_4_3), .B(f0_round_t_n1), 
        .Z(f0_round_p_io_state_out_3_2) );
  XOR2_X1 f0_round_t_U1 ( .A(f0_round0_io_state_out_4_4), .B(f0_round_t_n1), 
        .Z(f0_round_p_io_state_out_4_0) );
  NAND2_X1 f0_round_c_U50 ( .A1(f0_round_p_io_state_out_2_0), .A2(
        f0_round_p_io_state_out_1_0), .ZN(f0_round_c_n25) );
  XOR2_X1 f0_round_c_U49 ( .A(f0_round_c_n25), .B(f0_round_p_io_state_out_0_0), 
        .Z(f0_round_io_state_out_0_0) );
  NAND2_X1 f0_round_c_U48 ( .A1(f0_round_p_io_state_out_2_1), .A2(
        f0_round_p_io_state_out_1_1), .ZN(f0_round_c_n24) );
  XOR2_X1 f0_round_c_U47 ( .A(f0_round_c_n24), .B(f0_round_p_io_state_out_0_1), 
        .Z(f0_round_io_state_out_0_1) );
  NAND2_X1 f0_round_c_U46 ( .A1(f0_round_p_io_state_out_2_2), .A2(
        f0_round_p_io_state_out_1_2), .ZN(f0_round_c_n23) );
  XOR2_X1 f0_round_c_U45 ( .A(f0_round_c_n23), .B(f0_round_p_io_state_out_0_2), 
        .Z(f0_round_io_state_out_0_2) );
  NAND2_X1 f0_round_c_U44 ( .A1(f0_round_p_io_state_out_2_3), .A2(
        f0_round_p_io_state_out_1_3), .ZN(f0_round_c_n22) );
  XOR2_X1 f0_round_c_U43 ( .A(f0_round_c_n22), .B(f0_round_p_io_state_out_0_3), 
        .Z(f0_round_io_state_out_0_3) );
  NAND2_X1 f0_round_c_U42 ( .A1(f0_round_p_io_state_out_2_4), .A2(
        f0_round_p_io_state_out_1_4), .ZN(f0_round_c_n21) );
  XOR2_X1 f0_round_c_U41 ( .A(f0_round_c_n21), .B(f0_round_p_io_state_out_0_4), 
        .Z(f0_round_io_state_out_0_4) );
  NAND2_X1 f0_round_c_U40 ( .A1(f0_round_p_io_state_out_2_0), .A2(
        f0_round_p_io_state_out_3_0), .ZN(f0_round_c_n20) );
  XOR2_X1 f0_round_c_U39 ( .A(f0_round_c_n20), .B(f0_round_p_io_state_out_1_0), 
        .Z(f0_round_io_state_out_1_0) );
  NAND2_X1 f0_round_c_U38 ( .A1(f0_round_p_io_state_out_2_1), .A2(
        f0_round_p_io_state_out_3_1), .ZN(f0_round_c_n19) );
  XOR2_X1 f0_round_c_U37 ( .A(f0_round_c_n19), .B(f0_round_p_io_state_out_1_1), 
        .Z(f0_round_io_state_out_1_1) );
  NAND2_X1 f0_round_c_U36 ( .A1(f0_round_p_io_state_out_2_2), .A2(
        f0_round_p_io_state_out_3_2), .ZN(f0_round_c_n18) );
  XOR2_X1 f0_round_c_U35 ( .A(f0_round_c_n18), .B(f0_round_p_io_state_out_1_2), 
        .Z(f0_round_io_state_out_1_2) );
  NAND2_X1 f0_round_c_U34 ( .A1(f0_round_p_io_state_out_2_3), .A2(
        f0_round_p_io_state_out_3_3), .ZN(f0_round_c_n17) );
  XOR2_X1 f0_round_c_U33 ( .A(f0_round_c_n17), .B(f0_round_p_io_state_out_1_3), 
        .Z(f0_round_io_state_out_1_3) );
  NAND2_X1 f0_round_c_U32 ( .A1(f0_round_p_io_state_out_2_4), .A2(
        f0_round_p_io_state_out_3_4), .ZN(f0_round_c_n16) );
  XOR2_X1 f0_round_c_U31 ( .A(f0_round_c_n16), .B(f0_round_p_io_state_out_1_4), 
        .Z(f0_round_io_state_out_1_4) );
  NAND2_X1 f0_round_c_U30 ( .A1(f0_round_p_io_state_out_3_0), .A2(
        f0_round_p_io_state_out_4_0), .ZN(f0_round_c_n15) );
  XOR2_X1 f0_round_c_U29 ( .A(f0_round_c_n15), .B(f0_round_p_io_state_out_2_0), 
        .Z(f0_round_io_state_out_2_0) );
  NAND2_X1 f0_round_c_U28 ( .A1(f0_round_p_io_state_out_3_1), .A2(
        f0_round_p_io_state_out_4_1), .ZN(f0_round_c_n14) );
  XOR2_X1 f0_round_c_U27 ( .A(f0_round_c_n14), .B(f0_round_p_io_state_out_2_1), 
        .Z(f0_round_io_state_out_2_1) );
  NAND2_X1 f0_round_c_U26 ( .A1(f0_round_p_io_state_out_3_2), .A2(
        f0_round_p_io_state_out_4_2), .ZN(f0_round_c_n13) );
  XOR2_X1 f0_round_c_U25 ( .A(f0_round_c_n13), .B(f0_round_p_io_state_out_2_2), 
        .Z(f0_round_io_state_out_2_2) );
  NAND2_X1 f0_round_c_U24 ( .A1(f0_round_p_io_state_out_3_3), .A2(
        f0_round_p_io_state_out_4_3), .ZN(f0_round_c_n12) );
  XOR2_X1 f0_round_c_U23 ( .A(f0_round_c_n12), .B(f0_round_p_io_state_out_2_3), 
        .Z(f0_round_io_state_out_2_3) );
  NAND2_X1 f0_round_c_U22 ( .A1(f0_round_p_io_state_out_3_4), .A2(
        f0_round_p_io_state_out_4_4), .ZN(f0_round_c_n11) );
  XOR2_X1 f0_round_c_U21 ( .A(f0_round_c_n11), .B(f0_round_p_io_state_out_2_4), 
        .Z(f0_round_io_state_out_2_4) );
  NAND2_X1 f0_round_c_U20 ( .A1(f0_round_p_io_state_out_4_0), .A2(
        f0_round_p_io_state_out_0_0), .ZN(f0_round_c_n10) );
  XOR2_X1 f0_round_c_U19 ( .A(f0_round_c_n10), .B(f0_round_p_io_state_out_3_0), 
        .Z(f0_round_io_state_out_3_0) );
  NAND2_X1 f0_round_c_U18 ( .A1(f0_round_p_io_state_out_4_1), .A2(
        f0_round_p_io_state_out_0_1), .ZN(f0_round_c_n9) );
  XOR2_X1 f0_round_c_U17 ( .A(f0_round_c_n9), .B(f0_round_p_io_state_out_3_1), 
        .Z(f0_round_io_state_out_3_1) );
  NAND2_X1 f0_round_c_U16 ( .A1(f0_round_p_io_state_out_4_2), .A2(
        f0_round_p_io_state_out_0_2), .ZN(f0_round_c_n8) );
  XOR2_X1 f0_round_c_U15 ( .A(f0_round_c_n8), .B(f0_round_p_io_state_out_3_2), 
        .Z(f0_round_io_state_out_3_2) );
  NAND2_X1 f0_round_c_U14 ( .A1(f0_round_p_io_state_out_4_3), .A2(
        f0_round_p_io_state_out_0_3), .ZN(f0_round_c_n7) );
  XOR2_X1 f0_round_c_U13 ( .A(f0_round_c_n7), .B(f0_round_p_io_state_out_3_3), 
        .Z(f0_round_io_state_out_3_3) );
  NAND2_X1 f0_round_c_U12 ( .A1(f0_round_p_io_state_out_4_4), .A2(
        f0_round_p_io_state_out_0_4), .ZN(f0_round_c_n6) );
  XOR2_X1 f0_round_c_U11 ( .A(f0_round_c_n6), .B(f0_round_p_io_state_out_3_4), 
        .Z(f0_round_io_state_out_3_4) );
  NAND2_X1 f0_round_c_U10 ( .A1(f0_round_p_io_state_out_1_0), .A2(
        f0_round_p_io_state_out_0_0), .ZN(f0_round_c_n5) );
  XOR2_X1 f0_round_c_U9 ( .A(f0_round_c_n5), .B(f0_round_p_io_state_out_4_0), 
        .Z(f0_round_io_state_out_4_0) );
  NAND2_X1 f0_round_c_U8 ( .A1(f0_round_p_io_state_out_1_1), .A2(
        f0_round_p_io_state_out_0_1), .ZN(f0_round_c_n4) );
  XOR2_X1 f0_round_c_U7 ( .A(f0_round_c_n4), .B(f0_round_p_io_state_out_4_1), 
        .Z(f0_round_io_state_out_4_1) );
  NAND2_X1 f0_round_c_U6 ( .A1(f0_round_p_io_state_out_1_2), .A2(
        f0_round_p_io_state_out_0_2), .ZN(f0_round_c_n3) );
  XOR2_X1 f0_round_c_U5 ( .A(f0_round_c_n3), .B(f0_round_p_io_state_out_4_2), 
        .Z(f0_round_io_state_out_4_2) );
  NAND2_X1 f0_round_c_U4 ( .A1(f0_round_p_io_state_out_1_3), .A2(
        f0_round_p_io_state_out_0_3), .ZN(f0_round_c_n2) );
  XOR2_X1 f0_round_c_U3 ( .A(f0_round_c_n2), .B(f0_round_p_io_state_out_4_3), 
        .Z(f0_round_io_state_out_4_3) );
  NAND2_X1 f0_round_c_U2 ( .A1(f0_round_p_io_state_out_1_4), .A2(
        f0_round_p_io_state_out_0_4), .ZN(f0_round_c_n1) );
  XOR2_X1 f0_round_c_U1 ( .A(f0_round_c_n1), .B(f0_round_p_io_state_out_4_4), 
        .Z(f0_round_io_state_out_4_4) );
  XOR2_X1 f0_round_1_t_U50 ( .A(f0_round_io_state_out_1_4), .B(
        f0_round_io_state_out_1_3), .Z(f0_round_1_t_n25) );
  XNOR2_X1 f0_round_1_t_U49 ( .A(f0_round_io_state_out_1_2), .B(
        f0_round_1_t_n25), .ZN(f0_round_1_t_n23) );
  XOR2_X1 f0_round_1_t_U48 ( .A(f0_round_io_state_out_1_1), .B(
        f0_round_io_state_out_1_0), .Z(f0_round_1_t_n24) );
  XOR2_X1 f0_round_1_t_U47 ( .A(f0_round_1_t_n23), .B(f0_round_1_t_n24), .Z(
        f0_round_1_t_n8) );
  XOR2_X1 f0_round_1_t_U46 ( .A(f0_round_io_state_out_4_4), .B(
        f0_round_io_state_out_4_3), .Z(f0_round_1_t_n22) );
  XNOR2_X1 f0_round_1_t_U45 ( .A(f0_round_io_state_out_4_2), .B(
        f0_round_1_t_n22), .ZN(f0_round_1_t_n20) );
  XOR2_X1 f0_round_1_t_U44 ( .A(f0_round_io_state_out_4_1), .B(
        f0_round_io_state_out_4_0), .Z(f0_round_1_t_n21) );
  XNOR2_X1 f0_round_1_t_U43 ( .A(f0_round_1_t_n20), .B(f0_round_1_t_n21), .ZN(
        f0_round_1_t_n5) );
  XNOR2_X1 f0_round_1_t_U42 ( .A(f0_round_1_t_n8), .B(f0_round_1_t_n5), .ZN(
        f0_round_1_t_n19) );
  XOR2_X1 f0_round_1_t_U41 ( .A(f0_round_io_state_out_0_0), .B(
        f0_round_1_t_n19), .Z(f0_round_1_p_io_state_out_0_0) );
  XOR2_X1 f0_round_1_t_U40 ( .A(f0_round_io_state_out_0_1), .B(
        f0_round_1_t_n19), .Z(f0_round_1_p_io_state_out_1_3) );
  XOR2_X1 f0_round_1_t_U39 ( .A(f0_round_io_state_out_0_2), .B(
        f0_round_1_t_n19), .Z(f0_round_1_p_io_state_out_2_1) );
  XOR2_X1 f0_round_1_t_U38 ( .A(f0_round_io_state_out_0_3), .B(
        f0_round_1_t_n19), .Z(f0_round_1_p_io_state_out_3_4) );
  XOR2_X1 f0_round_1_t_U37 ( .A(f0_round_io_state_out_0_4), .B(
        f0_round_1_t_n19), .Z(f0_round_1_p_io_state_out_4_2) );
  XOR2_X1 f0_round_1_t_U36 ( .A(f0_round_io_state_out_2_4), .B(
        f0_round_io_state_out_2_3), .Z(f0_round_1_t_n18) );
  XNOR2_X1 f0_round_1_t_U35 ( .A(f0_round_io_state_out_2_2), .B(
        f0_round_1_t_n18), .ZN(f0_round_1_t_n16) );
  XOR2_X1 f0_round_1_t_U34 ( .A(f0_round_io_state_out_2_1), .B(
        f0_round_io_state_out_2_0), .Z(f0_round_1_t_n17) );
  XNOR2_X1 f0_round_1_t_U33 ( .A(f0_round_1_t_n16), .B(f0_round_1_t_n17), .ZN(
        f0_round_1_t_n6) );
  XOR2_X1 f0_round_1_t_U32 ( .A(f0_round_io_state_out_0_4), .B(
        f0_round_io_state_out_0_3), .Z(f0_round_1_t_n15) );
  XNOR2_X1 f0_round_1_t_U31 ( .A(f0_round_io_state_out_0_2), .B(
        f0_round_1_t_n15), .ZN(f0_round_1_t_n13) );
  XOR2_X1 f0_round_1_t_U30 ( .A(f0_round_io_state_out_0_1), .B(
        f0_round_io_state_out_0_0), .Z(f0_round_1_t_n14) );
  XNOR2_X1 f0_round_1_t_U29 ( .A(f0_round_1_t_n13), .B(f0_round_1_t_n14), .ZN(
        f0_round_1_t_n2) );
  XOR2_X1 f0_round_1_t_U28 ( .A(f0_round_1_t_n6), .B(f0_round_1_t_n2), .Z(
        f0_round_1_t_n12) );
  XOR2_X1 f0_round_1_t_U27 ( .A(f0_round_io_state_out_1_0), .B(
        f0_round_1_t_n12), .Z(f0_round_1_p_io_state_out_0_2) );
  XOR2_X1 f0_round_1_t_U26 ( .A(f0_round_io_state_out_1_1), .B(
        f0_round_1_t_n12), .Z(f0_round_1_p_io_state_out_1_0) );
  XOR2_X1 f0_round_1_t_U25 ( .A(f0_round_io_state_out_1_2), .B(
        f0_round_1_t_n12), .Z(f0_round_1_p_io_state_out_2_3) );
  XOR2_X1 f0_round_1_t_U24 ( .A(f0_round_io_state_out_1_3), .B(
        f0_round_1_t_n12), .Z(f0_round_1_p_io_state_out_3_1) );
  XOR2_X1 f0_round_1_t_U23 ( .A(f0_round_io_state_out_1_4), .B(
        f0_round_1_t_n12), .Z(f0_round_1_p_io_state_out_4_4) );
  XOR2_X1 f0_round_1_t_U22 ( .A(f0_round_io_state_out_3_4), .B(
        f0_round_io_state_out_3_3), .Z(f0_round_1_t_n11) );
  XNOR2_X1 f0_round_1_t_U21 ( .A(f0_round_io_state_out_3_2), .B(
        f0_round_1_t_n11), .ZN(f0_round_1_t_n9) );
  XOR2_X1 f0_round_1_t_U20 ( .A(f0_round_io_state_out_3_1), .B(
        f0_round_io_state_out_3_0), .Z(f0_round_1_t_n10) );
  XNOR2_X1 f0_round_1_t_U19 ( .A(f0_round_1_t_n9), .B(f0_round_1_t_n10), .ZN(
        f0_round_1_t_n3) );
  XNOR2_X1 f0_round_1_t_U18 ( .A(f0_round_1_t_n8), .B(f0_round_1_t_n3), .ZN(
        f0_round_1_t_n7) );
  XOR2_X1 f0_round_1_t_U17 ( .A(f0_round_io_state_out_2_0), .B(f0_round_1_t_n7), .Z(f0_round_1_p_io_state_out_0_4) );
  XOR2_X1 f0_round_1_t_U16 ( .A(f0_round_io_state_out_2_1), .B(f0_round_1_t_n7), .Z(f0_round_1_p_io_state_out_1_2) );
  XOR2_X1 f0_round_1_t_U15 ( .A(f0_round_io_state_out_2_2), .B(f0_round_1_t_n7), .Z(f0_round_1_p_io_state_out_2_0) );
  XOR2_X1 f0_round_1_t_U14 ( .A(f0_round_io_state_out_2_3), .B(f0_round_1_t_n7), .Z(f0_round_1_p_io_state_out_3_3) );
  XOR2_X1 f0_round_1_t_U13 ( .A(f0_round_io_state_out_2_4), .B(f0_round_1_t_n7), .Z(f0_round_1_p_io_state_out_4_1) );
  XOR2_X1 f0_round_1_t_U12 ( .A(f0_round_1_t_n5), .B(f0_round_1_t_n6), .Z(
        f0_round_1_t_n4) );
  XOR2_X1 f0_round_1_t_U11 ( .A(f0_round_io_state_out_3_0), .B(f0_round_1_t_n4), .Z(f0_round_1_p_io_state_out_0_1) );
  XOR2_X1 f0_round_1_t_U10 ( .A(f0_round_io_state_out_3_1), .B(f0_round_1_t_n4), .Z(f0_round_1_p_io_state_out_1_4) );
  XOR2_X1 f0_round_1_t_U9 ( .A(f0_round_io_state_out_3_2), .B(f0_round_1_t_n4), 
        .Z(f0_round_1_p_io_state_out_2_2) );
  XOR2_X1 f0_round_1_t_U8 ( .A(f0_round_io_state_out_3_3), .B(f0_round_1_t_n4), 
        .Z(f0_round_1_p_io_state_out_3_0) );
  XOR2_X1 f0_round_1_t_U7 ( .A(f0_round_io_state_out_3_4), .B(f0_round_1_t_n4), 
        .Z(f0_round_1_p_io_state_out_4_3) );
  XOR2_X1 f0_round_1_t_U6 ( .A(f0_round_1_t_n2), .B(f0_round_1_t_n3), .Z(
        f0_round_1_t_n1) );
  XOR2_X1 f0_round_1_t_U5 ( .A(f0_round_io_state_out_4_0), .B(f0_round_1_t_n1), 
        .Z(f0_round_1_p_io_state_out_0_3) );
  XOR2_X1 f0_round_1_t_U4 ( .A(f0_round_io_state_out_4_1), .B(f0_round_1_t_n1), 
        .Z(f0_round_1_p_io_state_out_1_1) );
  XOR2_X1 f0_round_1_t_U3 ( .A(f0_round_io_state_out_4_2), .B(f0_round_1_t_n1), 
        .Z(f0_round_1_p_io_state_out_2_4) );
  XOR2_X1 f0_round_1_t_U2 ( .A(f0_round_io_state_out_4_3), .B(f0_round_1_t_n1), 
        .Z(f0_round_1_p_io_state_out_3_2) );
  XOR2_X1 f0_round_1_t_U1 ( .A(f0_round_io_state_out_4_4), .B(f0_round_1_t_n1), 
        .Z(f0_round_1_p_io_state_out_4_0) );
  NAND2_X1 f0_round_1_c_U50 ( .A1(f0_round_1_p_io_state_out_2_0), .A2(
        f0_round_1_p_io_state_out_1_0), .ZN(f0_round_1_c_n25) );
  XOR2_X1 f0_round_1_c_U49 ( .A(f0_round_1_c_n25), .B(
        f0_round_1_p_io_state_out_0_0), .Z(f0_round_1_io_state_out_0_0) );
  NAND2_X1 f0_round_1_c_U48 ( .A1(f0_round_1_p_io_state_out_2_1), .A2(
        f0_round_1_p_io_state_out_1_1), .ZN(f0_round_1_c_n24) );
  XOR2_X1 f0_round_1_c_U47 ( .A(f0_round_1_c_n24), .B(
        f0_round_1_p_io_state_out_0_1), .Z(f0_round_1_io_state_out_0_1) );
  NAND2_X1 f0_round_1_c_U46 ( .A1(f0_round_1_p_io_state_out_2_2), .A2(
        f0_round_1_p_io_state_out_1_2), .ZN(f0_round_1_c_n23) );
  XOR2_X1 f0_round_1_c_U45 ( .A(f0_round_1_c_n23), .B(
        f0_round_1_p_io_state_out_0_2), .Z(f0_round_1_io_state_out_0_2) );
  NAND2_X1 f0_round_1_c_U44 ( .A1(f0_round_1_p_io_state_out_2_3), .A2(
        f0_round_1_p_io_state_out_1_3), .ZN(f0_round_1_c_n22) );
  XOR2_X1 f0_round_1_c_U43 ( .A(f0_round_1_c_n22), .B(
        f0_round_1_p_io_state_out_0_3), .Z(f0_round_1_io_state_out_0_3) );
  NAND2_X1 f0_round_1_c_U42 ( .A1(f0_round_1_p_io_state_out_2_4), .A2(
        f0_round_1_p_io_state_out_1_4), .ZN(f0_round_1_c_n21) );
  XOR2_X1 f0_round_1_c_U41 ( .A(f0_round_1_c_n21), .B(
        f0_round_1_p_io_state_out_0_4), .Z(f0_round_1_io_state_out_0_4) );
  NAND2_X1 f0_round_1_c_U40 ( .A1(f0_round_1_p_io_state_out_2_0), .A2(
        f0_round_1_p_io_state_out_3_0), .ZN(f0_round_1_c_n20) );
  XOR2_X1 f0_round_1_c_U39 ( .A(f0_round_1_c_n20), .B(
        f0_round_1_p_io_state_out_1_0), .Z(f0_round_1_io_state_out_1_0) );
  NAND2_X1 f0_round_1_c_U38 ( .A1(f0_round_1_p_io_state_out_2_1), .A2(
        f0_round_1_p_io_state_out_3_1), .ZN(f0_round_1_c_n19) );
  XOR2_X1 f0_round_1_c_U37 ( .A(f0_round_1_c_n19), .B(
        f0_round_1_p_io_state_out_1_1), .Z(f0_round_1_io_state_out_1_1) );
  NAND2_X1 f0_round_1_c_U36 ( .A1(f0_round_1_p_io_state_out_2_2), .A2(
        f0_round_1_p_io_state_out_3_2), .ZN(f0_round_1_c_n18) );
  XOR2_X1 f0_round_1_c_U35 ( .A(f0_round_1_c_n18), .B(
        f0_round_1_p_io_state_out_1_2), .Z(f0_round_1_io_state_out_1_2) );
  NAND2_X1 f0_round_1_c_U34 ( .A1(f0_round_1_p_io_state_out_2_3), .A2(
        f0_round_1_p_io_state_out_3_3), .ZN(f0_round_1_c_n17) );
  XOR2_X1 f0_round_1_c_U33 ( .A(f0_round_1_c_n17), .B(
        f0_round_1_p_io_state_out_1_3), .Z(f0_round_1_io_state_out_1_3) );
  NAND2_X1 f0_round_1_c_U32 ( .A1(f0_round_1_p_io_state_out_2_4), .A2(
        f0_round_1_p_io_state_out_3_4), .ZN(f0_round_1_c_n16) );
  XOR2_X1 f0_round_1_c_U31 ( .A(f0_round_1_c_n16), .B(
        f0_round_1_p_io_state_out_1_4), .Z(f0_round_1_io_state_out_1_4) );
  NAND2_X1 f0_round_1_c_U30 ( .A1(f0_round_1_p_io_state_out_3_0), .A2(
        f0_round_1_p_io_state_out_4_0), .ZN(f0_round_1_c_n15) );
  XOR2_X1 f0_round_1_c_U29 ( .A(f0_round_1_c_n15), .B(
        f0_round_1_p_io_state_out_2_0), .Z(f0_round_1_io_state_out_2_0) );
  NAND2_X1 f0_round_1_c_U28 ( .A1(f0_round_1_p_io_state_out_3_1), .A2(
        f0_round_1_p_io_state_out_4_1), .ZN(f0_round_1_c_n14) );
  XOR2_X1 f0_round_1_c_U27 ( .A(f0_round_1_c_n14), .B(
        f0_round_1_p_io_state_out_2_1), .Z(f0_round_1_io_state_out_2_1) );
  NAND2_X1 f0_round_1_c_U26 ( .A1(f0_round_1_p_io_state_out_3_2), .A2(
        f0_round_1_p_io_state_out_4_2), .ZN(f0_round_1_c_n13) );
  XOR2_X1 f0_round_1_c_U25 ( .A(f0_round_1_c_n13), .B(
        f0_round_1_p_io_state_out_2_2), .Z(f0_round_1_io_state_out_2_2) );
  NAND2_X1 f0_round_1_c_U24 ( .A1(f0_round_1_p_io_state_out_3_3), .A2(
        f0_round_1_p_io_state_out_4_3), .ZN(f0_round_1_c_n12) );
  XOR2_X1 f0_round_1_c_U23 ( .A(f0_round_1_c_n12), .B(
        f0_round_1_p_io_state_out_2_3), .Z(f0_round_1_io_state_out_2_3) );
  NAND2_X1 f0_round_1_c_U22 ( .A1(f0_round_1_p_io_state_out_3_4), .A2(
        f0_round_1_p_io_state_out_4_4), .ZN(f0_round_1_c_n11) );
  XOR2_X1 f0_round_1_c_U21 ( .A(f0_round_1_c_n11), .B(
        f0_round_1_p_io_state_out_2_4), .Z(f0_round_1_io_state_out_2_4) );
  NAND2_X1 f0_round_1_c_U20 ( .A1(f0_round_1_p_io_state_out_4_0), .A2(
        f0_round_1_p_io_state_out_0_0), .ZN(f0_round_1_c_n10) );
  XOR2_X1 f0_round_1_c_U19 ( .A(f0_round_1_c_n10), .B(
        f0_round_1_p_io_state_out_3_0), .Z(f0_round_1_io_state_out_3_0) );
  NAND2_X1 f0_round_1_c_U18 ( .A1(f0_round_1_p_io_state_out_4_1), .A2(
        f0_round_1_p_io_state_out_0_1), .ZN(f0_round_1_c_n9) );
  XOR2_X1 f0_round_1_c_U17 ( .A(f0_round_1_c_n9), .B(
        f0_round_1_p_io_state_out_3_1), .Z(f0_round_1_io_state_out_3_1) );
  NAND2_X1 f0_round_1_c_U16 ( .A1(f0_round_1_p_io_state_out_4_2), .A2(
        f0_round_1_p_io_state_out_0_2), .ZN(f0_round_1_c_n8) );
  XOR2_X1 f0_round_1_c_U15 ( .A(f0_round_1_c_n8), .B(
        f0_round_1_p_io_state_out_3_2), .Z(f0_round_1_io_state_out_3_2) );
  NAND2_X1 f0_round_1_c_U14 ( .A1(f0_round_1_p_io_state_out_4_3), .A2(
        f0_round_1_p_io_state_out_0_3), .ZN(f0_round_1_c_n7) );
  XOR2_X1 f0_round_1_c_U13 ( .A(f0_round_1_c_n7), .B(
        f0_round_1_p_io_state_out_3_3), .Z(f0_round_1_io_state_out_3_3) );
  NAND2_X1 f0_round_1_c_U12 ( .A1(f0_round_1_p_io_state_out_4_4), .A2(
        f0_round_1_p_io_state_out_0_4), .ZN(f0_round_1_c_n6) );
  XOR2_X1 f0_round_1_c_U11 ( .A(f0_round_1_c_n6), .B(
        f0_round_1_p_io_state_out_3_4), .Z(f0_round_1_io_state_out_3_4) );
  NAND2_X1 f0_round_1_c_U10 ( .A1(f0_round_1_p_io_state_out_1_0), .A2(
        f0_round_1_p_io_state_out_0_0), .ZN(f0_round_1_c_n5) );
  XOR2_X1 f0_round_1_c_U9 ( .A(f0_round_1_c_n5), .B(
        f0_round_1_p_io_state_out_4_0), .Z(f0_round_1_io_state_out_4_0) );
  NAND2_X1 f0_round_1_c_U8 ( .A1(f0_round_1_p_io_state_out_1_1), .A2(
        f0_round_1_p_io_state_out_0_1), .ZN(f0_round_1_c_n4) );
  XOR2_X1 f0_round_1_c_U7 ( .A(f0_round_1_c_n4), .B(
        f0_round_1_p_io_state_out_4_1), .Z(f0_round_1_io_state_out_4_1) );
  NAND2_X1 f0_round_1_c_U6 ( .A1(f0_round_1_p_io_state_out_1_2), .A2(
        f0_round_1_p_io_state_out_0_2), .ZN(f0_round_1_c_n3) );
  XOR2_X1 f0_round_1_c_U5 ( .A(f0_round_1_c_n3), .B(
        f0_round_1_p_io_state_out_4_2), .Z(f0_round_1_io_state_out_4_2) );
  NAND2_X1 f0_round_1_c_U4 ( .A1(f0_round_1_p_io_state_out_1_3), .A2(
        f0_round_1_p_io_state_out_0_3), .ZN(f0_round_1_c_n2) );
  XOR2_X1 f0_round_1_c_U3 ( .A(f0_round_1_c_n2), .B(
        f0_round_1_p_io_state_out_4_3), .Z(f0_round_1_io_state_out_4_3) );
  NAND2_X1 f0_round_1_c_U2 ( .A1(f0_round_1_p_io_state_out_1_4), .A2(
        f0_round_1_p_io_state_out_0_4), .ZN(f0_round_1_c_n1) );
  XOR2_X1 f0_round_1_c_U1 ( .A(f0_round_1_c_n1), .B(
        f0_round_1_p_io_state_out_4_4), .Z(f0_round_1_io_state_out_4_4) );
  XOR2_X1 f0_round_2_t_U50 ( .A(f0_round_1_io_state_out_1_4), .B(
        f0_round_1_io_state_out_1_3), .Z(f0_round_2_t_n25) );
  XNOR2_X1 f0_round_2_t_U49 ( .A(f0_round_1_io_state_out_1_2), .B(
        f0_round_2_t_n25), .ZN(f0_round_2_t_n23) );
  XOR2_X1 f0_round_2_t_U48 ( .A(f0_round_1_io_state_out_1_1), .B(
        f0_round_1_io_state_out_1_0), .Z(f0_round_2_t_n24) );
  XOR2_X1 f0_round_2_t_U47 ( .A(f0_round_2_t_n23), .B(f0_round_2_t_n24), .Z(
        f0_round_2_t_n8) );
  XOR2_X1 f0_round_2_t_U46 ( .A(f0_round_1_io_state_out_4_4), .B(
        f0_round_1_io_state_out_4_3), .Z(f0_round_2_t_n22) );
  XNOR2_X1 f0_round_2_t_U45 ( .A(f0_round_1_io_state_out_4_2), .B(
        f0_round_2_t_n22), .ZN(f0_round_2_t_n20) );
  XOR2_X1 f0_round_2_t_U44 ( .A(f0_round_1_io_state_out_4_1), .B(
        f0_round_1_io_state_out_4_0), .Z(f0_round_2_t_n21) );
  XNOR2_X1 f0_round_2_t_U43 ( .A(f0_round_2_t_n20), .B(f0_round_2_t_n21), .ZN(
        f0_round_2_t_n5) );
  XNOR2_X1 f0_round_2_t_U42 ( .A(f0_round_2_t_n8), .B(f0_round_2_t_n5), .ZN(
        f0_round_2_t_n19) );
  XOR2_X1 f0_round_2_t_U41 ( .A(f0_round_1_io_state_out_0_0), .B(
        f0_round_2_t_n19), .Z(f0_round_2_p_io_state_out_0_0) );
  XOR2_X1 f0_round_2_t_U40 ( .A(f0_round_1_io_state_out_0_1), .B(
        f0_round_2_t_n19), .Z(f0_round_2_p_io_state_out_1_3) );
  XOR2_X1 f0_round_2_t_U39 ( .A(f0_round_1_io_state_out_0_2), .B(
        f0_round_2_t_n19), .Z(f0_round_2_p_io_state_out_2_1) );
  XOR2_X1 f0_round_2_t_U38 ( .A(f0_round_1_io_state_out_0_3), .B(
        f0_round_2_t_n19), .Z(f0_round_2_p_io_state_out_3_4) );
  XOR2_X1 f0_round_2_t_U37 ( .A(f0_round_1_io_state_out_0_4), .B(
        f0_round_2_t_n19), .Z(f0_round_2_p_io_state_out_4_2) );
  XOR2_X1 f0_round_2_t_U36 ( .A(f0_round_1_io_state_out_2_4), .B(
        f0_round_1_io_state_out_2_3), .Z(f0_round_2_t_n18) );
  XNOR2_X1 f0_round_2_t_U35 ( .A(f0_round_1_io_state_out_2_2), .B(
        f0_round_2_t_n18), .ZN(f0_round_2_t_n16) );
  XOR2_X1 f0_round_2_t_U34 ( .A(f0_round_1_io_state_out_2_1), .B(
        f0_round_1_io_state_out_2_0), .Z(f0_round_2_t_n17) );
  XNOR2_X1 f0_round_2_t_U33 ( .A(f0_round_2_t_n16), .B(f0_round_2_t_n17), .ZN(
        f0_round_2_t_n6) );
  XOR2_X1 f0_round_2_t_U32 ( .A(f0_round_1_io_state_out_0_4), .B(
        f0_round_1_io_state_out_0_3), .Z(f0_round_2_t_n15) );
  XNOR2_X1 f0_round_2_t_U31 ( .A(f0_round_1_io_state_out_0_2), .B(
        f0_round_2_t_n15), .ZN(f0_round_2_t_n13) );
  XOR2_X1 f0_round_2_t_U30 ( .A(f0_round_1_io_state_out_0_1), .B(
        f0_round_1_io_state_out_0_0), .Z(f0_round_2_t_n14) );
  XNOR2_X1 f0_round_2_t_U29 ( .A(f0_round_2_t_n13), .B(f0_round_2_t_n14), .ZN(
        f0_round_2_t_n2) );
  XOR2_X1 f0_round_2_t_U28 ( .A(f0_round_2_t_n6), .B(f0_round_2_t_n2), .Z(
        f0_round_2_t_n12) );
  XOR2_X1 f0_round_2_t_U27 ( .A(f0_round_1_io_state_out_1_0), .B(
        f0_round_2_t_n12), .Z(f0_round_2_p_io_state_out_0_2) );
  XOR2_X1 f0_round_2_t_U26 ( .A(f0_round_1_io_state_out_1_1), .B(
        f0_round_2_t_n12), .Z(f0_round_2_p_io_state_out_1_0) );
  XOR2_X1 f0_round_2_t_U25 ( .A(f0_round_1_io_state_out_1_2), .B(
        f0_round_2_t_n12), .Z(f0_round_2_p_io_state_out_2_3) );
  XOR2_X1 f0_round_2_t_U24 ( .A(f0_round_1_io_state_out_1_3), .B(
        f0_round_2_t_n12), .Z(f0_round_2_p_io_state_out_3_1) );
  XOR2_X1 f0_round_2_t_U23 ( .A(f0_round_1_io_state_out_1_4), .B(
        f0_round_2_t_n12), .Z(f0_round_2_p_io_state_out_4_4) );
  XOR2_X1 f0_round_2_t_U22 ( .A(f0_round_1_io_state_out_3_4), .B(
        f0_round_1_io_state_out_3_3), .Z(f0_round_2_t_n11) );
  XNOR2_X1 f0_round_2_t_U21 ( .A(f0_round_1_io_state_out_3_2), .B(
        f0_round_2_t_n11), .ZN(f0_round_2_t_n9) );
  XOR2_X1 f0_round_2_t_U20 ( .A(f0_round_1_io_state_out_3_1), .B(
        f0_round_1_io_state_out_3_0), .Z(f0_round_2_t_n10) );
  XNOR2_X1 f0_round_2_t_U19 ( .A(f0_round_2_t_n9), .B(f0_round_2_t_n10), .ZN(
        f0_round_2_t_n3) );
  XNOR2_X1 f0_round_2_t_U18 ( .A(f0_round_2_t_n8), .B(f0_round_2_t_n3), .ZN(
        f0_round_2_t_n7) );
  XOR2_X1 f0_round_2_t_U17 ( .A(f0_round_1_io_state_out_2_0), .B(
        f0_round_2_t_n7), .Z(f0_round_2_p_io_state_out_0_4) );
  XOR2_X1 f0_round_2_t_U16 ( .A(f0_round_1_io_state_out_2_1), .B(
        f0_round_2_t_n7), .Z(f0_round_2_p_io_state_out_1_2) );
  XOR2_X1 f0_round_2_t_U15 ( .A(f0_round_1_io_state_out_2_2), .B(
        f0_round_2_t_n7), .Z(f0_round_2_p_io_state_out_2_0) );
  XOR2_X1 f0_round_2_t_U14 ( .A(f0_round_1_io_state_out_2_3), .B(
        f0_round_2_t_n7), .Z(f0_round_2_p_io_state_out_3_3) );
  XOR2_X1 f0_round_2_t_U13 ( .A(f0_round_1_io_state_out_2_4), .B(
        f0_round_2_t_n7), .Z(f0_round_2_p_io_state_out_4_1) );
  XOR2_X1 f0_round_2_t_U12 ( .A(f0_round_2_t_n5), .B(f0_round_2_t_n6), .Z(
        f0_round_2_t_n4) );
  XOR2_X1 f0_round_2_t_U11 ( .A(f0_round_1_io_state_out_3_0), .B(
        f0_round_2_t_n4), .Z(f0_round_2_p_io_state_out_0_1) );
  XOR2_X1 f0_round_2_t_U10 ( .A(f0_round_1_io_state_out_3_1), .B(
        f0_round_2_t_n4), .Z(f0_round_2_p_io_state_out_1_4) );
  XOR2_X1 f0_round_2_t_U9 ( .A(f0_round_1_io_state_out_3_2), .B(
        f0_round_2_t_n4), .Z(f0_round_2_p_io_state_out_2_2) );
  XOR2_X1 f0_round_2_t_U8 ( .A(f0_round_1_io_state_out_3_3), .B(
        f0_round_2_t_n4), .Z(f0_round_2_p_io_state_out_3_0) );
  XOR2_X1 f0_round_2_t_U7 ( .A(f0_round_1_io_state_out_3_4), .B(
        f0_round_2_t_n4), .Z(f0_round_2_p_io_state_out_4_3) );
  XOR2_X1 f0_round_2_t_U6 ( .A(f0_round_2_t_n2), .B(f0_round_2_t_n3), .Z(
        f0_round_2_t_n1) );
  XOR2_X1 f0_round_2_t_U5 ( .A(f0_round_1_io_state_out_4_0), .B(
        f0_round_2_t_n1), .Z(f0_round_2_p_io_state_out_0_3) );
  XOR2_X1 f0_round_2_t_U4 ( .A(f0_round_1_io_state_out_4_1), .B(
        f0_round_2_t_n1), .Z(f0_round_2_p_io_state_out_1_1) );
  XOR2_X1 f0_round_2_t_U3 ( .A(f0_round_1_io_state_out_4_2), .B(
        f0_round_2_t_n1), .Z(f0_round_2_p_io_state_out_2_4) );
  XOR2_X1 f0_round_2_t_U2 ( .A(f0_round_1_io_state_out_4_3), .B(
        f0_round_2_t_n1), .Z(f0_round_2_p_io_state_out_3_2) );
  XOR2_X1 f0_round_2_t_U1 ( .A(f0_round_1_io_state_out_4_4), .B(
        f0_round_2_t_n1), .Z(f0_round_2_p_io_state_out_4_0) );
  NAND2_X1 f0_round_2_c_U50 ( .A1(f0_round_2_p_io_state_out_2_0), .A2(
        f0_round_2_p_io_state_out_1_0), .ZN(f0_round_2_c_n25) );
  XOR2_X1 f0_round_2_c_U49 ( .A(f0_round_2_c_n25), .B(
        f0_round_2_p_io_state_out_0_0), .Z(f0_round_2_io_state_out_0_0) );
  NAND2_X1 f0_round_2_c_U48 ( .A1(f0_round_2_p_io_state_out_2_1), .A2(
        f0_round_2_p_io_state_out_1_1), .ZN(f0_round_2_c_n24) );
  XOR2_X1 f0_round_2_c_U47 ( .A(f0_round_2_c_n24), .B(
        f0_round_2_p_io_state_out_0_1), .Z(f0_round_2_io_state_out_0_1) );
  NAND2_X1 f0_round_2_c_U46 ( .A1(f0_round_2_p_io_state_out_2_2), .A2(
        f0_round_2_p_io_state_out_1_2), .ZN(f0_round_2_c_n23) );
  XOR2_X1 f0_round_2_c_U45 ( .A(f0_round_2_c_n23), .B(
        f0_round_2_p_io_state_out_0_2), .Z(f0_round_2_io_state_out_0_2) );
  NAND2_X1 f0_round_2_c_U44 ( .A1(f0_round_2_p_io_state_out_2_3), .A2(
        f0_round_2_p_io_state_out_1_3), .ZN(f0_round_2_c_n22) );
  XOR2_X1 f0_round_2_c_U43 ( .A(f0_round_2_c_n22), .B(
        f0_round_2_p_io_state_out_0_3), .Z(f0_round_2_io_state_out_0_3) );
  NAND2_X1 f0_round_2_c_U42 ( .A1(f0_round_2_p_io_state_out_2_4), .A2(
        f0_round_2_p_io_state_out_1_4), .ZN(f0_round_2_c_n21) );
  XOR2_X1 f0_round_2_c_U41 ( .A(f0_round_2_c_n21), .B(
        f0_round_2_p_io_state_out_0_4), .Z(f0_round_2_io_state_out_0_4) );
  NAND2_X1 f0_round_2_c_U40 ( .A1(f0_round_2_p_io_state_out_2_0), .A2(
        f0_round_2_p_io_state_out_3_0), .ZN(f0_round_2_c_n20) );
  XOR2_X1 f0_round_2_c_U39 ( .A(f0_round_2_c_n20), .B(
        f0_round_2_p_io_state_out_1_0), .Z(f0_round_2_io_state_out_1_0) );
  NAND2_X1 f0_round_2_c_U38 ( .A1(f0_round_2_p_io_state_out_2_1), .A2(
        f0_round_2_p_io_state_out_3_1), .ZN(f0_round_2_c_n19) );
  XOR2_X1 f0_round_2_c_U37 ( .A(f0_round_2_c_n19), .B(
        f0_round_2_p_io_state_out_1_1), .Z(f0_round_2_io_state_out_1_1) );
  NAND2_X1 f0_round_2_c_U36 ( .A1(f0_round_2_p_io_state_out_2_2), .A2(
        f0_round_2_p_io_state_out_3_2), .ZN(f0_round_2_c_n18) );
  XOR2_X1 f0_round_2_c_U35 ( .A(f0_round_2_c_n18), .B(
        f0_round_2_p_io_state_out_1_2), .Z(f0_round_2_io_state_out_1_2) );
  NAND2_X1 f0_round_2_c_U34 ( .A1(f0_round_2_p_io_state_out_2_3), .A2(
        f0_round_2_p_io_state_out_3_3), .ZN(f0_round_2_c_n17) );
  XOR2_X1 f0_round_2_c_U33 ( .A(f0_round_2_c_n17), .B(
        f0_round_2_p_io_state_out_1_3), .Z(f0_round_2_io_state_out_1_3) );
  NAND2_X1 f0_round_2_c_U32 ( .A1(f0_round_2_p_io_state_out_2_4), .A2(
        f0_round_2_p_io_state_out_3_4), .ZN(f0_round_2_c_n16) );
  XOR2_X1 f0_round_2_c_U31 ( .A(f0_round_2_c_n16), .B(
        f0_round_2_p_io_state_out_1_4), .Z(f0_round_2_io_state_out_1_4) );
  NAND2_X1 f0_round_2_c_U30 ( .A1(f0_round_2_p_io_state_out_3_0), .A2(
        f0_round_2_p_io_state_out_4_0), .ZN(f0_round_2_c_n15) );
  XOR2_X1 f0_round_2_c_U29 ( .A(f0_round_2_c_n15), .B(
        f0_round_2_p_io_state_out_2_0), .Z(f0_round_2_io_state_out_2_0) );
  NAND2_X1 f0_round_2_c_U28 ( .A1(f0_round_2_p_io_state_out_3_1), .A2(
        f0_round_2_p_io_state_out_4_1), .ZN(f0_round_2_c_n14) );
  XOR2_X1 f0_round_2_c_U27 ( .A(f0_round_2_c_n14), .B(
        f0_round_2_p_io_state_out_2_1), .Z(f0_round_2_io_state_out_2_1) );
  NAND2_X1 f0_round_2_c_U26 ( .A1(f0_round_2_p_io_state_out_3_2), .A2(
        f0_round_2_p_io_state_out_4_2), .ZN(f0_round_2_c_n13) );
  XOR2_X1 f0_round_2_c_U25 ( .A(f0_round_2_c_n13), .B(
        f0_round_2_p_io_state_out_2_2), .Z(f0_round_2_io_state_out_2_2) );
  NAND2_X1 f0_round_2_c_U24 ( .A1(f0_round_2_p_io_state_out_3_3), .A2(
        f0_round_2_p_io_state_out_4_3), .ZN(f0_round_2_c_n12) );
  XOR2_X1 f0_round_2_c_U23 ( .A(f0_round_2_c_n12), .B(
        f0_round_2_p_io_state_out_2_3), .Z(f0_round_2_io_state_out_2_3) );
  NAND2_X1 f0_round_2_c_U22 ( .A1(f0_round_2_p_io_state_out_3_4), .A2(
        f0_round_2_p_io_state_out_4_4), .ZN(f0_round_2_c_n11) );
  XOR2_X1 f0_round_2_c_U21 ( .A(f0_round_2_c_n11), .B(
        f0_round_2_p_io_state_out_2_4), .Z(f0_round_2_io_state_out_2_4) );
  NAND2_X1 f0_round_2_c_U20 ( .A1(f0_round_2_p_io_state_out_4_0), .A2(
        f0_round_2_p_io_state_out_0_0), .ZN(f0_round_2_c_n10) );
  XOR2_X1 f0_round_2_c_U19 ( .A(f0_round_2_c_n10), .B(
        f0_round_2_p_io_state_out_3_0), .Z(f0_round_2_io_state_out_3_0) );
  NAND2_X1 f0_round_2_c_U18 ( .A1(f0_round_2_p_io_state_out_4_1), .A2(
        f0_round_2_p_io_state_out_0_1), .ZN(f0_round_2_c_n9) );
  XOR2_X1 f0_round_2_c_U17 ( .A(f0_round_2_c_n9), .B(
        f0_round_2_p_io_state_out_3_1), .Z(f0_round_2_io_state_out_3_1) );
  NAND2_X1 f0_round_2_c_U16 ( .A1(f0_round_2_p_io_state_out_4_2), .A2(
        f0_round_2_p_io_state_out_0_2), .ZN(f0_round_2_c_n8) );
  XOR2_X1 f0_round_2_c_U15 ( .A(f0_round_2_c_n8), .B(
        f0_round_2_p_io_state_out_3_2), .Z(f0_round_2_io_state_out_3_2) );
  NAND2_X1 f0_round_2_c_U14 ( .A1(f0_round_2_p_io_state_out_4_3), .A2(
        f0_round_2_p_io_state_out_0_3), .ZN(f0_round_2_c_n7) );
  XOR2_X1 f0_round_2_c_U13 ( .A(f0_round_2_c_n7), .B(
        f0_round_2_p_io_state_out_3_3), .Z(f0_round_2_io_state_out_3_3) );
  NAND2_X1 f0_round_2_c_U12 ( .A1(f0_round_2_p_io_state_out_4_4), .A2(
        f0_round_2_p_io_state_out_0_4), .ZN(f0_round_2_c_n6) );
  XOR2_X1 f0_round_2_c_U11 ( .A(f0_round_2_c_n6), .B(
        f0_round_2_p_io_state_out_3_4), .Z(f0_round_2_io_state_out_3_4) );
  NAND2_X1 f0_round_2_c_U10 ( .A1(f0_round_2_p_io_state_out_1_0), .A2(
        f0_round_2_p_io_state_out_0_0), .ZN(f0_round_2_c_n5) );
  XOR2_X1 f0_round_2_c_U9 ( .A(f0_round_2_c_n5), .B(
        f0_round_2_p_io_state_out_4_0), .Z(f0_round_2_io_state_out_4_0) );
  NAND2_X1 f0_round_2_c_U8 ( .A1(f0_round_2_p_io_state_out_1_1), .A2(
        f0_round_2_p_io_state_out_0_1), .ZN(f0_round_2_c_n4) );
  XOR2_X1 f0_round_2_c_U7 ( .A(f0_round_2_c_n4), .B(
        f0_round_2_p_io_state_out_4_1), .Z(f0_round_2_io_state_out_4_1) );
  NAND2_X1 f0_round_2_c_U6 ( .A1(f0_round_2_p_io_state_out_1_2), .A2(
        f0_round_2_p_io_state_out_0_2), .ZN(f0_round_2_c_n3) );
  XOR2_X1 f0_round_2_c_U5 ( .A(f0_round_2_c_n3), .B(
        f0_round_2_p_io_state_out_4_2), .Z(f0_round_2_io_state_out_4_2) );
  NAND2_X1 f0_round_2_c_U4 ( .A1(f0_round_2_p_io_state_out_1_3), .A2(
        f0_round_2_p_io_state_out_0_3), .ZN(f0_round_2_c_n2) );
  XOR2_X1 f0_round_2_c_U3 ( .A(f0_round_2_c_n2), .B(
        f0_round_2_p_io_state_out_4_3), .Z(f0_round_2_io_state_out_4_3) );
  NAND2_X1 f0_round_2_c_U2 ( .A1(f0_round_2_p_io_state_out_1_4), .A2(
        f0_round_2_p_io_state_out_0_4), .ZN(f0_round_2_c_n1) );
  XOR2_X1 f0_round_2_c_U1 ( .A(f0_round_2_c_n1), .B(
        f0_round_2_p_io_state_out_4_4), .Z(f0_round_2_io_state_out_4_4) );
  XOR2_X1 f0_round_3_t_U50 ( .A(f0_round_2_io_state_out_1_4), .B(
        f0_round_2_io_state_out_1_3), .Z(f0_round_3_t_n25) );
  XNOR2_X1 f0_round_3_t_U49 ( .A(f0_round_2_io_state_out_1_2), .B(
        f0_round_3_t_n25), .ZN(f0_round_3_t_n23) );
  XOR2_X1 f0_round_3_t_U48 ( .A(f0_round_2_io_state_out_1_1), .B(
        f0_round_2_io_state_out_1_0), .Z(f0_round_3_t_n24) );
  XOR2_X1 f0_round_3_t_U47 ( .A(f0_round_3_t_n23), .B(f0_round_3_t_n24), .Z(
        f0_round_3_t_n8) );
  XOR2_X1 f0_round_3_t_U46 ( .A(f0_round_2_io_state_out_4_4), .B(
        f0_round_2_io_state_out_4_3), .Z(f0_round_3_t_n22) );
  XNOR2_X1 f0_round_3_t_U45 ( .A(f0_round_2_io_state_out_4_2), .B(
        f0_round_3_t_n22), .ZN(f0_round_3_t_n20) );
  XOR2_X1 f0_round_3_t_U44 ( .A(f0_round_2_io_state_out_4_1), .B(
        f0_round_2_io_state_out_4_0), .Z(f0_round_3_t_n21) );
  XNOR2_X1 f0_round_3_t_U43 ( .A(f0_round_3_t_n20), .B(f0_round_3_t_n21), .ZN(
        f0_round_3_t_n5) );
  XNOR2_X1 f0_round_3_t_U42 ( .A(f0_round_3_t_n8), .B(f0_round_3_t_n5), .ZN(
        f0_round_3_t_n19) );
  XOR2_X1 f0_round_3_t_U41 ( .A(f0_round_2_io_state_out_0_0), .B(
        f0_round_3_t_n19), .Z(f0_round_3_p_io_state_out_0_0) );
  XOR2_X1 f0_round_3_t_U40 ( .A(f0_round_2_io_state_out_0_1), .B(
        f0_round_3_t_n19), .Z(f0_round_3_p_io_state_out_1_3) );
  XOR2_X1 f0_round_3_t_U39 ( .A(f0_round_2_io_state_out_0_2), .B(
        f0_round_3_t_n19), .Z(f0_round_3_p_io_state_out_2_1) );
  XOR2_X1 f0_round_3_t_U38 ( .A(f0_round_2_io_state_out_0_3), .B(
        f0_round_3_t_n19), .Z(f0_round_3_p_io_state_out_3_4) );
  XOR2_X1 f0_round_3_t_U37 ( .A(f0_round_2_io_state_out_0_4), .B(
        f0_round_3_t_n19), .Z(f0_round_3_p_io_state_out_4_2) );
  XOR2_X1 f0_round_3_t_U36 ( .A(f0_round_2_io_state_out_2_4), .B(
        f0_round_2_io_state_out_2_3), .Z(f0_round_3_t_n18) );
  XNOR2_X1 f0_round_3_t_U35 ( .A(f0_round_2_io_state_out_2_2), .B(
        f0_round_3_t_n18), .ZN(f0_round_3_t_n16) );
  XOR2_X1 f0_round_3_t_U34 ( .A(f0_round_2_io_state_out_2_1), .B(
        f0_round_2_io_state_out_2_0), .Z(f0_round_3_t_n17) );
  XNOR2_X1 f0_round_3_t_U33 ( .A(f0_round_3_t_n16), .B(f0_round_3_t_n17), .ZN(
        f0_round_3_t_n6) );
  XOR2_X1 f0_round_3_t_U32 ( .A(f0_round_2_io_state_out_0_4), .B(
        f0_round_2_io_state_out_0_3), .Z(f0_round_3_t_n15) );
  XNOR2_X1 f0_round_3_t_U31 ( .A(f0_round_2_io_state_out_0_2), .B(
        f0_round_3_t_n15), .ZN(f0_round_3_t_n13) );
  XOR2_X1 f0_round_3_t_U30 ( .A(f0_round_2_io_state_out_0_1), .B(
        f0_round_2_io_state_out_0_0), .Z(f0_round_3_t_n14) );
  XNOR2_X1 f0_round_3_t_U29 ( .A(f0_round_3_t_n13), .B(f0_round_3_t_n14), .ZN(
        f0_round_3_t_n2) );
  XOR2_X1 f0_round_3_t_U28 ( .A(f0_round_3_t_n6), .B(f0_round_3_t_n2), .Z(
        f0_round_3_t_n12) );
  XOR2_X1 f0_round_3_t_U27 ( .A(f0_round_2_io_state_out_1_0), .B(
        f0_round_3_t_n12), .Z(f0_round_3_p_io_state_out_0_2) );
  XOR2_X1 f0_round_3_t_U26 ( .A(f0_round_2_io_state_out_1_1), .B(
        f0_round_3_t_n12), .Z(f0_round_3_p_io_state_out_1_0) );
  XOR2_X1 f0_round_3_t_U25 ( .A(f0_round_2_io_state_out_1_2), .B(
        f0_round_3_t_n12), .Z(f0_round_3_p_io_state_out_2_3) );
  XOR2_X1 f0_round_3_t_U24 ( .A(f0_round_2_io_state_out_1_3), .B(
        f0_round_3_t_n12), .Z(f0_round_3_p_io_state_out_3_1) );
  XOR2_X1 f0_round_3_t_U23 ( .A(f0_round_2_io_state_out_1_4), .B(
        f0_round_3_t_n12), .Z(f0_round_3_p_io_state_out_4_4) );
  XOR2_X1 f0_round_3_t_U22 ( .A(f0_round_2_io_state_out_3_4), .B(
        f0_round_2_io_state_out_3_3), .Z(f0_round_3_t_n11) );
  XNOR2_X1 f0_round_3_t_U21 ( .A(f0_round_2_io_state_out_3_2), .B(
        f0_round_3_t_n11), .ZN(f0_round_3_t_n9) );
  XOR2_X1 f0_round_3_t_U20 ( .A(f0_round_2_io_state_out_3_1), .B(
        f0_round_2_io_state_out_3_0), .Z(f0_round_3_t_n10) );
  XNOR2_X1 f0_round_3_t_U19 ( .A(f0_round_3_t_n9), .B(f0_round_3_t_n10), .ZN(
        f0_round_3_t_n3) );
  XNOR2_X1 f0_round_3_t_U18 ( .A(f0_round_3_t_n8), .B(f0_round_3_t_n3), .ZN(
        f0_round_3_t_n7) );
  XOR2_X1 f0_round_3_t_U17 ( .A(f0_round_2_io_state_out_2_0), .B(
        f0_round_3_t_n7), .Z(f0_round_3_p_io_state_out_0_4) );
  XOR2_X1 f0_round_3_t_U16 ( .A(f0_round_2_io_state_out_2_1), .B(
        f0_round_3_t_n7), .Z(f0_round_3_p_io_state_out_1_2) );
  XOR2_X1 f0_round_3_t_U15 ( .A(f0_round_2_io_state_out_2_2), .B(
        f0_round_3_t_n7), .Z(f0_round_3_p_io_state_out_2_0) );
  XOR2_X1 f0_round_3_t_U14 ( .A(f0_round_2_io_state_out_2_3), .B(
        f0_round_3_t_n7), .Z(f0_round_3_p_io_state_out_3_3) );
  XOR2_X1 f0_round_3_t_U13 ( .A(f0_round_2_io_state_out_2_4), .B(
        f0_round_3_t_n7), .Z(f0_round_3_p_io_state_out_4_1) );
  XOR2_X1 f0_round_3_t_U12 ( .A(f0_round_3_t_n5), .B(f0_round_3_t_n6), .Z(
        f0_round_3_t_n4) );
  XOR2_X1 f0_round_3_t_U11 ( .A(f0_round_2_io_state_out_3_0), .B(
        f0_round_3_t_n4), .Z(f0_round_3_p_io_state_out_0_1) );
  XOR2_X1 f0_round_3_t_U10 ( .A(f0_round_2_io_state_out_3_1), .B(
        f0_round_3_t_n4), .Z(f0_round_3_p_io_state_out_1_4) );
  XOR2_X1 f0_round_3_t_U9 ( .A(f0_round_2_io_state_out_3_2), .B(
        f0_round_3_t_n4), .Z(f0_round_3_p_io_state_out_2_2) );
  XOR2_X1 f0_round_3_t_U8 ( .A(f0_round_2_io_state_out_3_3), .B(
        f0_round_3_t_n4), .Z(f0_round_3_p_io_state_out_3_0) );
  XOR2_X1 f0_round_3_t_U7 ( .A(f0_round_2_io_state_out_3_4), .B(
        f0_round_3_t_n4), .Z(f0_round_3_p_io_state_out_4_3) );
  XOR2_X1 f0_round_3_t_U6 ( .A(f0_round_3_t_n2), .B(f0_round_3_t_n3), .Z(
        f0_round_3_t_n1) );
  XOR2_X1 f0_round_3_t_U5 ( .A(f0_round_2_io_state_out_4_0), .B(
        f0_round_3_t_n1), .Z(f0_round_3_p_io_state_out_0_3) );
  XOR2_X1 f0_round_3_t_U4 ( .A(f0_round_2_io_state_out_4_1), .B(
        f0_round_3_t_n1), .Z(f0_round_3_p_io_state_out_1_1) );
  XOR2_X1 f0_round_3_t_U3 ( .A(f0_round_2_io_state_out_4_2), .B(
        f0_round_3_t_n1), .Z(f0_round_3_p_io_state_out_2_4) );
  XOR2_X1 f0_round_3_t_U2 ( .A(f0_round_2_io_state_out_4_3), .B(
        f0_round_3_t_n1), .Z(f0_round_3_p_io_state_out_3_2) );
  XOR2_X1 f0_round_3_t_U1 ( .A(f0_round_2_io_state_out_4_4), .B(
        f0_round_3_t_n1), .Z(f0_round_3_p_io_state_out_4_0) );
  NAND2_X1 f0_round_3_c_U50 ( .A1(f0_round_3_p_io_state_out_2_0), .A2(
        f0_round_3_p_io_state_out_1_0), .ZN(f0_round_3_c_n25) );
  XOR2_X1 f0_round_3_c_U49 ( .A(f0_round_3_c_n25), .B(
        f0_round_3_p_io_state_out_0_0), .Z(f0_round_3_c_io_state_out_0_0) );
  NAND2_X1 f0_round_3_c_U48 ( .A1(f0_round_3_p_io_state_out_2_1), .A2(
        f0_round_3_p_io_state_out_1_1), .ZN(f0_round_3_c_n24) );
  XOR2_X1 f0_round_3_c_U47 ( .A(f0_round_3_c_n24), .B(
        f0_round_3_p_io_state_out_0_1), .Z(f0_round_3_io_state_out_0_1) );
  NAND2_X1 f0_round_3_c_U46 ( .A1(f0_round_3_p_io_state_out_2_2), .A2(
        f0_round_3_p_io_state_out_1_2), .ZN(f0_round_3_c_n23) );
  XOR2_X1 f0_round_3_c_U45 ( .A(f0_round_3_c_n23), .B(
        f0_round_3_p_io_state_out_0_2), .Z(f0_round_3_io_state_out_0_2) );
  NAND2_X1 f0_round_3_c_U44 ( .A1(f0_round_3_p_io_state_out_2_3), .A2(
        f0_round_3_p_io_state_out_1_3), .ZN(f0_round_3_c_n22) );
  XOR2_X1 f0_round_3_c_U43 ( .A(f0_round_3_c_n22), .B(
        f0_round_3_p_io_state_out_0_3), .Z(f0_round_3_io_state_out_0_3) );
  NAND2_X1 f0_round_3_c_U42 ( .A1(f0_round_3_p_io_state_out_2_4), .A2(
        f0_round_3_p_io_state_out_1_4), .ZN(f0_round_3_c_n21) );
  XOR2_X1 f0_round_3_c_U41 ( .A(f0_round_3_c_n21), .B(
        f0_round_3_p_io_state_out_0_4), .Z(f0_round_3_io_state_out_0_4) );
  NAND2_X1 f0_round_3_c_U40 ( .A1(f0_round_3_p_io_state_out_2_0), .A2(
        f0_round_3_p_io_state_out_3_0), .ZN(f0_round_3_c_n20) );
  XOR2_X1 f0_round_3_c_U39 ( .A(f0_round_3_c_n20), .B(
        f0_round_3_p_io_state_out_1_0), .Z(f0_round_3_io_state_out_1_0) );
  NAND2_X1 f0_round_3_c_U38 ( .A1(f0_round_3_p_io_state_out_2_1), .A2(
        f0_round_3_p_io_state_out_3_1), .ZN(f0_round_3_c_n19) );
  XOR2_X1 f0_round_3_c_U37 ( .A(f0_round_3_c_n19), .B(
        f0_round_3_p_io_state_out_1_1), .Z(f0_round_3_io_state_out_1_1) );
  NAND2_X1 f0_round_3_c_U36 ( .A1(f0_round_3_p_io_state_out_2_2), .A2(
        f0_round_3_p_io_state_out_3_2), .ZN(f0_round_3_c_n18) );
  XOR2_X1 f0_round_3_c_U35 ( .A(f0_round_3_c_n18), .B(
        f0_round_3_p_io_state_out_1_2), .Z(f0_round_3_io_state_out_1_2) );
  NAND2_X1 f0_round_3_c_U34 ( .A1(f0_round_3_p_io_state_out_2_3), .A2(
        f0_round_3_p_io_state_out_3_3), .ZN(f0_round_3_c_n17) );
  XOR2_X1 f0_round_3_c_U33 ( .A(f0_round_3_c_n17), .B(
        f0_round_3_p_io_state_out_1_3), .Z(f0_round_3_io_state_out_1_3) );
  NAND2_X1 f0_round_3_c_U32 ( .A1(f0_round_3_p_io_state_out_2_4), .A2(
        f0_round_3_p_io_state_out_3_4), .ZN(f0_round_3_c_n16) );
  XOR2_X1 f0_round_3_c_U31 ( .A(f0_round_3_c_n16), .B(
        f0_round_3_p_io_state_out_1_4), .Z(f0_round_3_io_state_out_1_4) );
  NAND2_X1 f0_round_3_c_U30 ( .A1(f0_round_3_p_io_state_out_3_0), .A2(
        f0_round_3_p_io_state_out_4_0), .ZN(f0_round_3_c_n15) );
  XOR2_X1 f0_round_3_c_U29 ( .A(f0_round_3_c_n15), .B(
        f0_round_3_p_io_state_out_2_0), .Z(f0_round_3_io_state_out_2_0) );
  NAND2_X1 f0_round_3_c_U28 ( .A1(f0_round_3_p_io_state_out_3_1), .A2(
        f0_round_3_p_io_state_out_4_1), .ZN(f0_round_3_c_n14) );
  XOR2_X1 f0_round_3_c_U27 ( .A(f0_round_3_c_n14), .B(
        f0_round_3_p_io_state_out_2_1), .Z(f0_round_3_io_state_out_2_1) );
  NAND2_X1 f0_round_3_c_U26 ( .A1(f0_round_3_p_io_state_out_3_2), .A2(
        f0_round_3_p_io_state_out_4_2), .ZN(f0_round_3_c_n13) );
  XOR2_X1 f0_round_3_c_U25 ( .A(f0_round_3_c_n13), .B(
        f0_round_3_p_io_state_out_2_2), .Z(f0_round_3_io_state_out_2_2) );
  NAND2_X1 f0_round_3_c_U24 ( .A1(f0_round_3_p_io_state_out_3_3), .A2(
        f0_round_3_p_io_state_out_4_3), .ZN(f0_round_3_c_n12) );
  XOR2_X1 f0_round_3_c_U23 ( .A(f0_round_3_c_n12), .B(
        f0_round_3_p_io_state_out_2_3), .Z(f0_round_3_io_state_out_2_3) );
  NAND2_X1 f0_round_3_c_U22 ( .A1(f0_round_3_p_io_state_out_3_4), .A2(
        f0_round_3_p_io_state_out_4_4), .ZN(f0_round_3_c_n11) );
  XOR2_X1 f0_round_3_c_U21 ( .A(f0_round_3_c_n11), .B(
        f0_round_3_p_io_state_out_2_4), .Z(f0_round_3_io_state_out_2_4) );
  NAND2_X1 f0_round_3_c_U20 ( .A1(f0_round_3_p_io_state_out_4_0), .A2(
        f0_round_3_p_io_state_out_0_0), .ZN(f0_round_3_c_n10) );
  XOR2_X1 f0_round_3_c_U19 ( .A(f0_round_3_c_n10), .B(
        f0_round_3_p_io_state_out_3_0), .Z(f0_round_3_io_state_out_3_0) );
  NAND2_X1 f0_round_3_c_U18 ( .A1(f0_round_3_p_io_state_out_4_1), .A2(
        f0_round_3_p_io_state_out_0_1), .ZN(f0_round_3_c_n9) );
  XOR2_X1 f0_round_3_c_U17 ( .A(f0_round_3_c_n9), .B(
        f0_round_3_p_io_state_out_3_1), .Z(f0_round_3_io_state_out_3_1) );
  NAND2_X1 f0_round_3_c_U16 ( .A1(f0_round_3_p_io_state_out_4_2), .A2(
        f0_round_3_p_io_state_out_0_2), .ZN(f0_round_3_c_n8) );
  XOR2_X1 f0_round_3_c_U15 ( .A(f0_round_3_c_n8), .B(
        f0_round_3_p_io_state_out_3_2), .Z(f0_round_3_io_state_out_3_2) );
  NAND2_X1 f0_round_3_c_U14 ( .A1(f0_round_3_p_io_state_out_4_3), .A2(
        f0_round_3_p_io_state_out_0_3), .ZN(f0_round_3_c_n7) );
  XOR2_X1 f0_round_3_c_U13 ( .A(f0_round_3_c_n7), .B(
        f0_round_3_p_io_state_out_3_3), .Z(f0_round_3_io_state_out_3_3) );
  NAND2_X1 f0_round_3_c_U12 ( .A1(f0_round_3_p_io_state_out_4_4), .A2(
        f0_round_3_p_io_state_out_0_4), .ZN(f0_round_3_c_n6) );
  XOR2_X1 f0_round_3_c_U11 ( .A(f0_round_3_c_n6), .B(
        f0_round_3_p_io_state_out_3_4), .Z(f0_round_3_io_state_out_3_4) );
  NAND2_X1 f0_round_3_c_U10 ( .A1(f0_round_3_p_io_state_out_1_0), .A2(
        f0_round_3_p_io_state_out_0_0), .ZN(f0_round_3_c_n5) );
  XOR2_X1 f0_round_3_c_U9 ( .A(f0_round_3_c_n5), .B(
        f0_round_3_p_io_state_out_4_0), .Z(f0_round_3_io_state_out_4_0) );
  NAND2_X1 f0_round_3_c_U8 ( .A1(f0_round_3_p_io_state_out_1_1), .A2(
        f0_round_3_p_io_state_out_0_1), .ZN(f0_round_3_c_n4) );
  XOR2_X1 f0_round_3_c_U7 ( .A(f0_round_3_c_n4), .B(
        f0_round_3_p_io_state_out_4_1), .Z(f0_round_3_io_state_out_4_1) );
  NAND2_X1 f0_round_3_c_U6 ( .A1(f0_round_3_p_io_state_out_1_2), .A2(
        f0_round_3_p_io_state_out_0_2), .ZN(f0_round_3_c_n3) );
  XOR2_X1 f0_round_3_c_U5 ( .A(f0_round_3_c_n3), .B(
        f0_round_3_p_io_state_out_4_2), .Z(f0_round_3_io_state_out_4_2) );
  NAND2_X1 f0_round_3_c_U4 ( .A1(f0_round_3_p_io_state_out_1_3), .A2(
        f0_round_3_p_io_state_out_0_3), .ZN(f0_round_3_c_n2) );
  XOR2_X1 f0_round_3_c_U3 ( .A(f0_round_3_c_n2), .B(
        f0_round_3_p_io_state_out_4_3), .Z(f0_round_3_io_state_out_4_3) );
  NAND2_X1 f0_round_3_c_U2 ( .A1(f0_round_3_p_io_state_out_1_4), .A2(
        f0_round_3_p_io_state_out_0_4), .ZN(f0_round_3_c_n1) );
  XOR2_X1 f0_round_3_c_U1 ( .A(f0_round_3_c_n1), .B(
        f0_round_3_p_io_state_out_4_4), .Z(f0_round_3_io_state_out_4_4) );
  INV_X1 f0_round_3_i_U1 ( .A(f0_round_3_c_io_state_out_0_0), .ZN(
        f0_round_3_io_state_out_0_0) );
  XOR2_X1 f0_round_4_t_U50 ( .A(f0_round_3_io_state_out_1_4), .B(
        f0_round_3_io_state_out_1_3), .Z(f0_round_4_t_n25) );
  XNOR2_X1 f0_round_4_t_U49 ( .A(f0_round_3_io_state_out_1_2), .B(
        f0_round_4_t_n25), .ZN(f0_round_4_t_n23) );
  XOR2_X1 f0_round_4_t_U48 ( .A(f0_round_3_io_state_out_1_1), .B(
        f0_round_3_io_state_out_1_0), .Z(f0_round_4_t_n24) );
  XOR2_X1 f0_round_4_t_U47 ( .A(f0_round_4_t_n23), .B(f0_round_4_t_n24), .Z(
        f0_round_4_t_n8) );
  XOR2_X1 f0_round_4_t_U46 ( .A(f0_round_3_io_state_out_4_4), .B(
        f0_round_3_io_state_out_4_3), .Z(f0_round_4_t_n22) );
  XNOR2_X1 f0_round_4_t_U45 ( .A(f0_round_3_io_state_out_4_2), .B(
        f0_round_4_t_n22), .ZN(f0_round_4_t_n20) );
  XOR2_X1 f0_round_4_t_U44 ( .A(f0_round_3_io_state_out_4_1), .B(
        f0_round_3_io_state_out_4_0), .Z(f0_round_4_t_n21) );
  XNOR2_X1 f0_round_4_t_U43 ( .A(f0_round_4_t_n20), .B(f0_round_4_t_n21), .ZN(
        f0_round_4_t_n5) );
  XNOR2_X1 f0_round_4_t_U42 ( .A(f0_round_4_t_n8), .B(f0_round_4_t_n5), .ZN(
        f0_round_4_t_n19) );
  XOR2_X1 f0_round_4_t_U41 ( .A(f0_round_3_io_state_out_0_0), .B(
        f0_round_4_t_n19), .Z(f0_round_4_p_io_state_out_0_0) );
  XOR2_X1 f0_round_4_t_U40 ( .A(f0_round_3_io_state_out_0_1), .B(
        f0_round_4_t_n19), .Z(f0_round_4_p_io_state_out_1_3) );
  XOR2_X1 f0_round_4_t_U39 ( .A(f0_round_3_io_state_out_0_2), .B(
        f0_round_4_t_n19), .Z(f0_round_4_p_io_state_out_2_1) );
  XOR2_X1 f0_round_4_t_U38 ( .A(f0_round_3_io_state_out_0_3), .B(
        f0_round_4_t_n19), .Z(f0_round_4_p_io_state_out_3_4) );
  XOR2_X1 f0_round_4_t_U37 ( .A(f0_round_3_io_state_out_0_4), .B(
        f0_round_4_t_n19), .Z(f0_round_4_p_io_state_out_4_2) );
  XOR2_X1 f0_round_4_t_U36 ( .A(f0_round_3_io_state_out_2_4), .B(
        f0_round_3_io_state_out_2_3), .Z(f0_round_4_t_n18) );
  XNOR2_X1 f0_round_4_t_U35 ( .A(f0_round_3_io_state_out_2_2), .B(
        f0_round_4_t_n18), .ZN(f0_round_4_t_n16) );
  XOR2_X1 f0_round_4_t_U34 ( .A(f0_round_3_io_state_out_2_1), .B(
        f0_round_3_io_state_out_2_0), .Z(f0_round_4_t_n17) );
  XNOR2_X1 f0_round_4_t_U33 ( .A(f0_round_4_t_n16), .B(f0_round_4_t_n17), .ZN(
        f0_round_4_t_n6) );
  XOR2_X1 f0_round_4_t_U32 ( .A(f0_round_3_io_state_out_0_4), .B(
        f0_round_3_io_state_out_0_3), .Z(f0_round_4_t_n15) );
  XNOR2_X1 f0_round_4_t_U31 ( .A(f0_round_3_io_state_out_0_2), .B(
        f0_round_4_t_n15), .ZN(f0_round_4_t_n13) );
  XOR2_X1 f0_round_4_t_U30 ( .A(f0_round_3_io_state_out_0_1), .B(
        f0_round_3_io_state_out_0_0), .Z(f0_round_4_t_n14) );
  XNOR2_X1 f0_round_4_t_U29 ( .A(f0_round_4_t_n13), .B(f0_round_4_t_n14), .ZN(
        f0_round_4_t_n2) );
  XOR2_X1 f0_round_4_t_U28 ( .A(f0_round_4_t_n6), .B(f0_round_4_t_n2), .Z(
        f0_round_4_t_n12) );
  XOR2_X1 f0_round_4_t_U27 ( .A(f0_round_3_io_state_out_1_0), .B(
        f0_round_4_t_n12), .Z(f0_round_4_p_io_state_out_0_2) );
  XOR2_X1 f0_round_4_t_U26 ( .A(f0_round_3_io_state_out_1_1), .B(
        f0_round_4_t_n12), .Z(f0_round_4_p_io_state_out_1_0) );
  XOR2_X1 f0_round_4_t_U25 ( .A(f0_round_3_io_state_out_1_2), .B(
        f0_round_4_t_n12), .Z(f0_round_4_p_io_state_out_2_3) );
  XOR2_X1 f0_round_4_t_U24 ( .A(f0_round_3_io_state_out_1_3), .B(
        f0_round_4_t_n12), .Z(f0_round_4_p_io_state_out_3_1) );
  XOR2_X1 f0_round_4_t_U23 ( .A(f0_round_3_io_state_out_1_4), .B(
        f0_round_4_t_n12), .Z(f0_round_4_p_io_state_out_4_4) );
  XOR2_X1 f0_round_4_t_U22 ( .A(f0_round_3_io_state_out_3_4), .B(
        f0_round_3_io_state_out_3_3), .Z(f0_round_4_t_n11) );
  XNOR2_X1 f0_round_4_t_U21 ( .A(f0_round_3_io_state_out_3_2), .B(
        f0_round_4_t_n11), .ZN(f0_round_4_t_n9) );
  XOR2_X1 f0_round_4_t_U20 ( .A(f0_round_3_io_state_out_3_1), .B(
        f0_round_3_io_state_out_3_0), .Z(f0_round_4_t_n10) );
  XNOR2_X1 f0_round_4_t_U19 ( .A(f0_round_4_t_n9), .B(f0_round_4_t_n10), .ZN(
        f0_round_4_t_n3) );
  XNOR2_X1 f0_round_4_t_U18 ( .A(f0_round_4_t_n8), .B(f0_round_4_t_n3), .ZN(
        f0_round_4_t_n7) );
  XOR2_X1 f0_round_4_t_U17 ( .A(f0_round_3_io_state_out_2_0), .B(
        f0_round_4_t_n7), .Z(f0_round_4_p_io_state_out_0_4) );
  XOR2_X1 f0_round_4_t_U16 ( .A(f0_round_3_io_state_out_2_1), .B(
        f0_round_4_t_n7), .Z(f0_round_4_p_io_state_out_1_2) );
  XOR2_X1 f0_round_4_t_U15 ( .A(f0_round_3_io_state_out_2_2), .B(
        f0_round_4_t_n7), .Z(f0_round_4_p_io_state_out_2_0) );
  XOR2_X1 f0_round_4_t_U14 ( .A(f0_round_3_io_state_out_2_3), .B(
        f0_round_4_t_n7), .Z(f0_round_4_p_io_state_out_3_3) );
  XOR2_X1 f0_round_4_t_U13 ( .A(f0_round_3_io_state_out_2_4), .B(
        f0_round_4_t_n7), .Z(f0_round_4_p_io_state_out_4_1) );
  XOR2_X1 f0_round_4_t_U12 ( .A(f0_round_4_t_n5), .B(f0_round_4_t_n6), .Z(
        f0_round_4_t_n4) );
  XOR2_X1 f0_round_4_t_U11 ( .A(f0_round_3_io_state_out_3_0), .B(
        f0_round_4_t_n4), .Z(f0_round_4_p_io_state_out_0_1) );
  XOR2_X1 f0_round_4_t_U10 ( .A(f0_round_3_io_state_out_3_1), .B(
        f0_round_4_t_n4), .Z(f0_round_4_p_io_state_out_1_4) );
  XOR2_X1 f0_round_4_t_U9 ( .A(f0_round_3_io_state_out_3_2), .B(
        f0_round_4_t_n4), .Z(f0_round_4_p_io_state_out_2_2) );
  XOR2_X1 f0_round_4_t_U8 ( .A(f0_round_3_io_state_out_3_3), .B(
        f0_round_4_t_n4), .Z(f0_round_4_p_io_state_out_3_0) );
  XOR2_X1 f0_round_4_t_U7 ( .A(f0_round_3_io_state_out_3_4), .B(
        f0_round_4_t_n4), .Z(f0_round_4_p_io_state_out_4_3) );
  XOR2_X1 f0_round_4_t_U6 ( .A(f0_round_4_t_n2), .B(f0_round_4_t_n3), .Z(
        f0_round_4_t_n1) );
  XOR2_X1 f0_round_4_t_U5 ( .A(f0_round_3_io_state_out_4_0), .B(
        f0_round_4_t_n1), .Z(f0_round_4_p_io_state_out_0_3) );
  XOR2_X1 f0_round_4_t_U4 ( .A(f0_round_3_io_state_out_4_1), .B(
        f0_round_4_t_n1), .Z(f0_round_4_p_io_state_out_1_1) );
  XOR2_X1 f0_round_4_t_U3 ( .A(f0_round_3_io_state_out_4_2), .B(
        f0_round_4_t_n1), .Z(f0_round_4_p_io_state_out_2_4) );
  XOR2_X1 f0_round_4_t_U2 ( .A(f0_round_3_io_state_out_4_3), .B(
        f0_round_4_t_n1), .Z(f0_round_4_p_io_state_out_3_2) );
  XOR2_X1 f0_round_4_t_U1 ( .A(f0_round_3_io_state_out_4_4), .B(
        f0_round_4_t_n1), .Z(f0_round_4_p_io_state_out_4_0) );
  NAND2_X1 f0_round_4_c_U50 ( .A1(f0_round_4_p_io_state_out_2_0), .A2(
        f0_round_4_p_io_state_out_1_0), .ZN(f0_round_4_c_n25) );
  XOR2_X1 f0_round_4_c_U49 ( .A(f0_round_4_c_n25), .B(
        f0_round_4_p_io_state_out_0_0), .Z(f0_round_4_c_io_state_out_0_0) );
  NAND2_X1 f0_round_4_c_U48 ( .A1(f0_round_4_p_io_state_out_2_1), .A2(
        f0_round_4_p_io_state_out_1_1), .ZN(f0_round_4_c_n24) );
  XOR2_X1 f0_round_4_c_U47 ( .A(f0_round_4_c_n24), .B(
        f0_round_4_p_io_state_out_0_1), .Z(f0_round_4_io_state_out_0_1) );
  NAND2_X1 f0_round_4_c_U46 ( .A1(f0_round_4_p_io_state_out_2_2), .A2(
        f0_round_4_p_io_state_out_1_2), .ZN(f0_round_4_c_n23) );
  XOR2_X1 f0_round_4_c_U45 ( .A(f0_round_4_c_n23), .B(
        f0_round_4_p_io_state_out_0_2), .Z(f0_round_4_io_state_out_0_2) );
  NAND2_X1 f0_round_4_c_U44 ( .A1(f0_round_4_p_io_state_out_2_3), .A2(
        f0_round_4_p_io_state_out_1_3), .ZN(f0_round_4_c_n22) );
  XOR2_X1 f0_round_4_c_U43 ( .A(f0_round_4_c_n22), .B(
        f0_round_4_p_io_state_out_0_3), .Z(f0_round_4_io_state_out_0_3) );
  NAND2_X1 f0_round_4_c_U42 ( .A1(f0_round_4_p_io_state_out_2_4), .A2(
        f0_round_4_p_io_state_out_1_4), .ZN(f0_round_4_c_n21) );
  XOR2_X1 f0_round_4_c_U41 ( .A(f0_round_4_c_n21), .B(
        f0_round_4_p_io_state_out_0_4), .Z(f0_round_4_io_state_out_0_4) );
  NAND2_X1 f0_round_4_c_U40 ( .A1(f0_round_4_p_io_state_out_2_0), .A2(
        f0_round_4_p_io_state_out_3_0), .ZN(f0_round_4_c_n20) );
  XOR2_X1 f0_round_4_c_U39 ( .A(f0_round_4_c_n20), .B(
        f0_round_4_p_io_state_out_1_0), .Z(f0_round_4_io_state_out_1_0) );
  NAND2_X1 f0_round_4_c_U38 ( .A1(f0_round_4_p_io_state_out_2_1), .A2(
        f0_round_4_p_io_state_out_3_1), .ZN(f0_round_4_c_n19) );
  XOR2_X1 f0_round_4_c_U37 ( .A(f0_round_4_c_n19), .B(
        f0_round_4_p_io_state_out_1_1), .Z(f0_round_4_io_state_out_1_1) );
  NAND2_X1 f0_round_4_c_U36 ( .A1(f0_round_4_p_io_state_out_2_2), .A2(
        f0_round_4_p_io_state_out_3_2), .ZN(f0_round_4_c_n18) );
  XOR2_X1 f0_round_4_c_U35 ( .A(f0_round_4_c_n18), .B(
        f0_round_4_p_io_state_out_1_2), .Z(f0_round_4_io_state_out_1_2) );
  NAND2_X1 f0_round_4_c_U34 ( .A1(f0_round_4_p_io_state_out_2_3), .A2(
        f0_round_4_p_io_state_out_3_3), .ZN(f0_round_4_c_n17) );
  XOR2_X1 f0_round_4_c_U33 ( .A(f0_round_4_c_n17), .B(
        f0_round_4_p_io_state_out_1_3), .Z(f0_round_4_io_state_out_1_3) );
  NAND2_X1 f0_round_4_c_U32 ( .A1(f0_round_4_p_io_state_out_2_4), .A2(
        f0_round_4_p_io_state_out_3_4), .ZN(f0_round_4_c_n16) );
  XOR2_X1 f0_round_4_c_U31 ( .A(f0_round_4_c_n16), .B(
        f0_round_4_p_io_state_out_1_4), .Z(f0_round_4_io_state_out_1_4) );
  NAND2_X1 f0_round_4_c_U30 ( .A1(f0_round_4_p_io_state_out_3_0), .A2(
        f0_round_4_p_io_state_out_4_0), .ZN(f0_round_4_c_n15) );
  XOR2_X1 f0_round_4_c_U29 ( .A(f0_round_4_c_n15), .B(
        f0_round_4_p_io_state_out_2_0), .Z(f0_round_4_io_state_out_2_0) );
  NAND2_X1 f0_round_4_c_U28 ( .A1(f0_round_4_p_io_state_out_3_1), .A2(
        f0_round_4_p_io_state_out_4_1), .ZN(f0_round_4_c_n14) );
  XOR2_X1 f0_round_4_c_U27 ( .A(f0_round_4_c_n14), .B(
        f0_round_4_p_io_state_out_2_1), .Z(f0_round_4_io_state_out_2_1) );
  NAND2_X1 f0_round_4_c_U26 ( .A1(f0_round_4_p_io_state_out_3_2), .A2(
        f0_round_4_p_io_state_out_4_2), .ZN(f0_round_4_c_n13) );
  XOR2_X1 f0_round_4_c_U25 ( .A(f0_round_4_c_n13), .B(
        f0_round_4_p_io_state_out_2_2), .Z(f0_round_4_io_state_out_2_2) );
  NAND2_X1 f0_round_4_c_U24 ( .A1(f0_round_4_p_io_state_out_3_3), .A2(
        f0_round_4_p_io_state_out_4_3), .ZN(f0_round_4_c_n12) );
  XOR2_X1 f0_round_4_c_U23 ( .A(f0_round_4_c_n12), .B(
        f0_round_4_p_io_state_out_2_3), .Z(f0_round_4_io_state_out_2_3) );
  NAND2_X1 f0_round_4_c_U22 ( .A1(f0_round_4_p_io_state_out_3_4), .A2(
        f0_round_4_p_io_state_out_4_4), .ZN(f0_round_4_c_n11) );
  XOR2_X1 f0_round_4_c_U21 ( .A(f0_round_4_c_n11), .B(
        f0_round_4_p_io_state_out_2_4), .Z(f0_round_4_io_state_out_2_4) );
  NAND2_X1 f0_round_4_c_U20 ( .A1(f0_round_4_p_io_state_out_4_0), .A2(
        f0_round_4_p_io_state_out_0_0), .ZN(f0_round_4_c_n10) );
  XOR2_X1 f0_round_4_c_U19 ( .A(f0_round_4_c_n10), .B(
        f0_round_4_p_io_state_out_3_0), .Z(f0_round_4_io_state_out_3_0) );
  NAND2_X1 f0_round_4_c_U18 ( .A1(f0_round_4_p_io_state_out_4_1), .A2(
        f0_round_4_p_io_state_out_0_1), .ZN(f0_round_4_c_n9) );
  XOR2_X1 f0_round_4_c_U17 ( .A(f0_round_4_c_n9), .B(
        f0_round_4_p_io_state_out_3_1), .Z(f0_round_4_io_state_out_3_1) );
  NAND2_X1 f0_round_4_c_U16 ( .A1(f0_round_4_p_io_state_out_4_2), .A2(
        f0_round_4_p_io_state_out_0_2), .ZN(f0_round_4_c_n8) );
  XOR2_X1 f0_round_4_c_U15 ( .A(f0_round_4_c_n8), .B(
        f0_round_4_p_io_state_out_3_2), .Z(f0_round_4_io_state_out_3_2) );
  NAND2_X1 f0_round_4_c_U14 ( .A1(f0_round_4_p_io_state_out_4_3), .A2(
        f0_round_4_p_io_state_out_0_3), .ZN(f0_round_4_c_n7) );
  XOR2_X1 f0_round_4_c_U13 ( .A(f0_round_4_c_n7), .B(
        f0_round_4_p_io_state_out_3_3), .Z(f0_round_4_io_state_out_3_3) );
  NAND2_X1 f0_round_4_c_U12 ( .A1(f0_round_4_p_io_state_out_4_4), .A2(
        f0_round_4_p_io_state_out_0_4), .ZN(f0_round_4_c_n6) );
  XOR2_X1 f0_round_4_c_U11 ( .A(f0_round_4_c_n6), .B(
        f0_round_4_p_io_state_out_3_4), .Z(f0_round_4_io_state_out_3_4) );
  NAND2_X1 f0_round_4_c_U10 ( .A1(f0_round_4_p_io_state_out_1_0), .A2(
        f0_round_4_p_io_state_out_0_0), .ZN(f0_round_4_c_n5) );
  XOR2_X1 f0_round_4_c_U9 ( .A(f0_round_4_c_n5), .B(
        f0_round_4_p_io_state_out_4_0), .Z(f0_round_4_io_state_out_4_0) );
  NAND2_X1 f0_round_4_c_U8 ( .A1(f0_round_4_p_io_state_out_1_1), .A2(
        f0_round_4_p_io_state_out_0_1), .ZN(f0_round_4_c_n4) );
  XOR2_X1 f0_round_4_c_U7 ( .A(f0_round_4_c_n4), .B(
        f0_round_4_p_io_state_out_4_1), .Z(f0_round_4_io_state_out_4_1) );
  NAND2_X1 f0_round_4_c_U6 ( .A1(f0_round_4_p_io_state_out_1_2), .A2(
        f0_round_4_p_io_state_out_0_2), .ZN(f0_round_4_c_n3) );
  XOR2_X1 f0_round_4_c_U5 ( .A(f0_round_4_c_n3), .B(
        f0_round_4_p_io_state_out_4_2), .Z(f0_round_4_io_state_out_4_2) );
  NAND2_X1 f0_round_4_c_U4 ( .A1(f0_round_4_p_io_state_out_1_3), .A2(
        f0_round_4_p_io_state_out_0_3), .ZN(f0_round_4_c_n2) );
  XOR2_X1 f0_round_4_c_U3 ( .A(f0_round_4_c_n2), .B(
        f0_round_4_p_io_state_out_4_3), .Z(f0_round_4_io_state_out_4_3) );
  NAND2_X1 f0_round_4_c_U2 ( .A1(f0_round_4_p_io_state_out_1_4), .A2(
        f0_round_4_p_io_state_out_0_4), .ZN(f0_round_4_c_n1) );
  XOR2_X1 f0_round_4_c_U1 ( .A(f0_round_4_c_n1), .B(
        f0_round_4_p_io_state_out_4_4), .Z(f0_round_4_io_state_out_4_4) );
  INV_X1 f0_round_4_i_U1 ( .A(f0_round_4_c_io_state_out_0_0), .ZN(
        f0_round_4_io_state_out_0_0) );
  XOR2_X1 f0_round_5_t_U50 ( .A(f0_round_4_io_state_out_1_4), .B(
        f0_round_4_io_state_out_1_3), .Z(f0_round_5_t_n25) );
  XNOR2_X1 f0_round_5_t_U49 ( .A(f0_round_4_io_state_out_1_2), .B(
        f0_round_5_t_n25), .ZN(f0_round_5_t_n23) );
  XOR2_X1 f0_round_5_t_U48 ( .A(f0_round_4_io_state_out_1_1), .B(
        f0_round_4_io_state_out_1_0), .Z(f0_round_5_t_n24) );
  XOR2_X1 f0_round_5_t_U47 ( .A(f0_round_5_t_n23), .B(f0_round_5_t_n24), .Z(
        f0_round_5_t_n8) );
  XOR2_X1 f0_round_5_t_U46 ( .A(f0_round_4_io_state_out_4_4), .B(
        f0_round_4_io_state_out_4_3), .Z(f0_round_5_t_n22) );
  XNOR2_X1 f0_round_5_t_U45 ( .A(f0_round_4_io_state_out_4_2), .B(
        f0_round_5_t_n22), .ZN(f0_round_5_t_n20) );
  XOR2_X1 f0_round_5_t_U44 ( .A(f0_round_4_io_state_out_4_1), .B(
        f0_round_4_io_state_out_4_0), .Z(f0_round_5_t_n21) );
  XNOR2_X1 f0_round_5_t_U43 ( .A(f0_round_5_t_n20), .B(f0_round_5_t_n21), .ZN(
        f0_round_5_t_n5) );
  XNOR2_X1 f0_round_5_t_U42 ( .A(f0_round_5_t_n8), .B(f0_round_5_t_n5), .ZN(
        f0_round_5_t_n19) );
  XOR2_X1 f0_round_5_t_U41 ( .A(f0_round_4_io_state_out_0_0), .B(
        f0_round_5_t_n19), .Z(f0_round_5_p_io_state_out_0_0) );
  XOR2_X1 f0_round_5_t_U40 ( .A(f0_round_4_io_state_out_0_1), .B(
        f0_round_5_t_n19), .Z(f0_round_5_p_io_state_out_1_3) );
  XOR2_X1 f0_round_5_t_U39 ( .A(f0_round_4_io_state_out_0_2), .B(
        f0_round_5_t_n19), .Z(f0_round_5_p_io_state_out_2_1) );
  XOR2_X1 f0_round_5_t_U38 ( .A(f0_round_4_io_state_out_0_3), .B(
        f0_round_5_t_n19), .Z(f0_round_5_p_io_state_out_3_4) );
  XOR2_X1 f0_round_5_t_U37 ( .A(f0_round_4_io_state_out_0_4), .B(
        f0_round_5_t_n19), .Z(f0_round_5_p_io_state_out_4_2) );
  XOR2_X1 f0_round_5_t_U36 ( .A(f0_round_4_io_state_out_2_4), .B(
        f0_round_4_io_state_out_2_3), .Z(f0_round_5_t_n18) );
  XNOR2_X1 f0_round_5_t_U35 ( .A(f0_round_4_io_state_out_2_2), .B(
        f0_round_5_t_n18), .ZN(f0_round_5_t_n16) );
  XOR2_X1 f0_round_5_t_U34 ( .A(f0_round_4_io_state_out_2_1), .B(
        f0_round_4_io_state_out_2_0), .Z(f0_round_5_t_n17) );
  XNOR2_X1 f0_round_5_t_U33 ( .A(f0_round_5_t_n16), .B(f0_round_5_t_n17), .ZN(
        f0_round_5_t_n6) );
  XOR2_X1 f0_round_5_t_U32 ( .A(f0_round_4_io_state_out_0_4), .B(
        f0_round_4_io_state_out_0_3), .Z(f0_round_5_t_n15) );
  XNOR2_X1 f0_round_5_t_U31 ( .A(f0_round_4_io_state_out_0_2), .B(
        f0_round_5_t_n15), .ZN(f0_round_5_t_n13) );
  XOR2_X1 f0_round_5_t_U30 ( .A(f0_round_4_io_state_out_0_1), .B(
        f0_round_4_io_state_out_0_0), .Z(f0_round_5_t_n14) );
  XNOR2_X1 f0_round_5_t_U29 ( .A(f0_round_5_t_n13), .B(f0_round_5_t_n14), .ZN(
        f0_round_5_t_n2) );
  XOR2_X1 f0_round_5_t_U28 ( .A(f0_round_5_t_n6), .B(f0_round_5_t_n2), .Z(
        f0_round_5_t_n12) );
  XOR2_X1 f0_round_5_t_U27 ( .A(f0_round_4_io_state_out_1_0), .B(
        f0_round_5_t_n12), .Z(f0_round_5_p_io_state_out_0_2) );
  XOR2_X1 f0_round_5_t_U26 ( .A(f0_round_4_io_state_out_1_1), .B(
        f0_round_5_t_n12), .Z(f0_round_5_p_io_state_out_1_0) );
  XOR2_X1 f0_round_5_t_U25 ( .A(f0_round_4_io_state_out_1_2), .B(
        f0_round_5_t_n12), .Z(f0_round_5_p_io_state_out_2_3) );
  XOR2_X1 f0_round_5_t_U24 ( .A(f0_round_4_io_state_out_1_3), .B(
        f0_round_5_t_n12), .Z(f0_round_5_p_io_state_out_3_1) );
  XOR2_X1 f0_round_5_t_U23 ( .A(f0_round_4_io_state_out_1_4), .B(
        f0_round_5_t_n12), .Z(f0_round_5_p_io_state_out_4_4) );
  XOR2_X1 f0_round_5_t_U22 ( .A(f0_round_4_io_state_out_3_4), .B(
        f0_round_4_io_state_out_3_3), .Z(f0_round_5_t_n11) );
  XNOR2_X1 f0_round_5_t_U21 ( .A(f0_round_4_io_state_out_3_2), .B(
        f0_round_5_t_n11), .ZN(f0_round_5_t_n9) );
  XOR2_X1 f0_round_5_t_U20 ( .A(f0_round_4_io_state_out_3_1), .B(
        f0_round_4_io_state_out_3_0), .Z(f0_round_5_t_n10) );
  XNOR2_X1 f0_round_5_t_U19 ( .A(f0_round_5_t_n9), .B(f0_round_5_t_n10), .ZN(
        f0_round_5_t_n3) );
  XNOR2_X1 f0_round_5_t_U18 ( .A(f0_round_5_t_n8), .B(f0_round_5_t_n3), .ZN(
        f0_round_5_t_n7) );
  XOR2_X1 f0_round_5_t_U17 ( .A(f0_round_4_io_state_out_2_0), .B(
        f0_round_5_t_n7), .Z(f0_round_5_p_io_state_out_0_4) );
  XOR2_X1 f0_round_5_t_U16 ( .A(f0_round_4_io_state_out_2_1), .B(
        f0_round_5_t_n7), .Z(f0_round_5_p_io_state_out_1_2) );
  XOR2_X1 f0_round_5_t_U15 ( .A(f0_round_4_io_state_out_2_2), .B(
        f0_round_5_t_n7), .Z(f0_round_5_p_io_state_out_2_0) );
  XOR2_X1 f0_round_5_t_U14 ( .A(f0_round_4_io_state_out_2_3), .B(
        f0_round_5_t_n7), .Z(f0_round_5_p_io_state_out_3_3) );
  XOR2_X1 f0_round_5_t_U13 ( .A(f0_round_4_io_state_out_2_4), .B(
        f0_round_5_t_n7), .Z(f0_round_5_p_io_state_out_4_1) );
  XOR2_X1 f0_round_5_t_U12 ( .A(f0_round_5_t_n5), .B(f0_round_5_t_n6), .Z(
        f0_round_5_t_n4) );
  XOR2_X1 f0_round_5_t_U11 ( .A(f0_round_4_io_state_out_3_0), .B(
        f0_round_5_t_n4), .Z(f0_round_5_p_io_state_out_0_1) );
  XOR2_X1 f0_round_5_t_U10 ( .A(f0_round_4_io_state_out_3_1), .B(
        f0_round_5_t_n4), .Z(f0_round_5_p_io_state_out_1_4) );
  XOR2_X1 f0_round_5_t_U9 ( .A(f0_round_4_io_state_out_3_2), .B(
        f0_round_5_t_n4), .Z(f0_round_5_p_io_state_out_2_2) );
  XOR2_X1 f0_round_5_t_U8 ( .A(f0_round_4_io_state_out_3_3), .B(
        f0_round_5_t_n4), .Z(f0_round_5_p_io_state_out_3_0) );
  XOR2_X1 f0_round_5_t_U7 ( .A(f0_round_4_io_state_out_3_4), .B(
        f0_round_5_t_n4), .Z(f0_round_5_p_io_state_out_4_3) );
  XOR2_X1 f0_round_5_t_U6 ( .A(f0_round_5_t_n2), .B(f0_round_5_t_n3), .Z(
        f0_round_5_t_n1) );
  XOR2_X1 f0_round_5_t_U5 ( .A(f0_round_4_io_state_out_4_0), .B(
        f0_round_5_t_n1), .Z(f0_round_5_p_io_state_out_0_3) );
  XOR2_X1 f0_round_5_t_U4 ( .A(f0_round_4_io_state_out_4_1), .B(
        f0_round_5_t_n1), .Z(f0_round_5_p_io_state_out_1_1) );
  XOR2_X1 f0_round_5_t_U3 ( .A(f0_round_4_io_state_out_4_2), .B(
        f0_round_5_t_n1), .Z(f0_round_5_p_io_state_out_2_4) );
  XOR2_X1 f0_round_5_t_U2 ( .A(f0_round_4_io_state_out_4_3), .B(
        f0_round_5_t_n1), .Z(f0_round_5_p_io_state_out_3_2) );
  XOR2_X1 f0_round_5_t_U1 ( .A(f0_round_4_io_state_out_4_4), .B(
        f0_round_5_t_n1), .Z(f0_round_5_p_io_state_out_4_0) );
  NAND2_X1 f0_round_5_c_U50 ( .A1(f0_round_5_p_io_state_out_2_0), .A2(
        f0_round_5_p_io_state_out_1_0), .ZN(f0_round_5_c_n25) );
  XOR2_X1 f0_round_5_c_U49 ( .A(f0_round_5_c_n25), .B(
        f0_round_5_p_io_state_out_0_0), .Z(f0_round_5_c_io_state_out_0_0) );
  NAND2_X1 f0_round_5_c_U48 ( .A1(f0_round_5_p_io_state_out_2_1), .A2(
        f0_round_5_p_io_state_out_1_1), .ZN(f0_round_5_c_n24) );
  XOR2_X1 f0_round_5_c_U47 ( .A(f0_round_5_c_n24), .B(
        f0_round_5_p_io_state_out_0_1), .Z(f0_round_5_io_state_out_0_1) );
  NAND2_X1 f0_round_5_c_U46 ( .A1(f0_round_5_p_io_state_out_2_2), .A2(
        f0_round_5_p_io_state_out_1_2), .ZN(f0_round_5_c_n23) );
  XOR2_X1 f0_round_5_c_U45 ( .A(f0_round_5_c_n23), .B(
        f0_round_5_p_io_state_out_0_2), .Z(f0_round_5_io_state_out_0_2) );
  NAND2_X1 f0_round_5_c_U44 ( .A1(f0_round_5_p_io_state_out_2_3), .A2(
        f0_round_5_p_io_state_out_1_3), .ZN(f0_round_5_c_n22) );
  XOR2_X1 f0_round_5_c_U43 ( .A(f0_round_5_c_n22), .B(
        f0_round_5_p_io_state_out_0_3), .Z(f0_round_5_io_state_out_0_3) );
  NAND2_X1 f0_round_5_c_U42 ( .A1(f0_round_5_p_io_state_out_2_4), .A2(
        f0_round_5_p_io_state_out_1_4), .ZN(f0_round_5_c_n21) );
  XOR2_X1 f0_round_5_c_U41 ( .A(f0_round_5_c_n21), .B(
        f0_round_5_p_io_state_out_0_4), .Z(f0_round_5_io_state_out_0_4) );
  NAND2_X1 f0_round_5_c_U40 ( .A1(f0_round_5_p_io_state_out_2_0), .A2(
        f0_round_5_p_io_state_out_3_0), .ZN(f0_round_5_c_n20) );
  XOR2_X1 f0_round_5_c_U39 ( .A(f0_round_5_c_n20), .B(
        f0_round_5_p_io_state_out_1_0), .Z(f0_round_5_io_state_out_1_0) );
  NAND2_X1 f0_round_5_c_U38 ( .A1(f0_round_5_p_io_state_out_2_1), .A2(
        f0_round_5_p_io_state_out_3_1), .ZN(f0_round_5_c_n19) );
  XOR2_X1 f0_round_5_c_U37 ( .A(f0_round_5_c_n19), .B(
        f0_round_5_p_io_state_out_1_1), .Z(f0_round_5_io_state_out_1_1) );
  NAND2_X1 f0_round_5_c_U36 ( .A1(f0_round_5_p_io_state_out_2_2), .A2(
        f0_round_5_p_io_state_out_3_2), .ZN(f0_round_5_c_n18) );
  XOR2_X1 f0_round_5_c_U35 ( .A(f0_round_5_c_n18), .B(
        f0_round_5_p_io_state_out_1_2), .Z(f0_round_5_io_state_out_1_2) );
  NAND2_X1 f0_round_5_c_U34 ( .A1(f0_round_5_p_io_state_out_2_3), .A2(
        f0_round_5_p_io_state_out_3_3), .ZN(f0_round_5_c_n17) );
  XOR2_X1 f0_round_5_c_U33 ( .A(f0_round_5_c_n17), .B(
        f0_round_5_p_io_state_out_1_3), .Z(f0_round_5_io_state_out_1_3) );
  NAND2_X1 f0_round_5_c_U32 ( .A1(f0_round_5_p_io_state_out_2_4), .A2(
        f0_round_5_p_io_state_out_3_4), .ZN(f0_round_5_c_n16) );
  XOR2_X1 f0_round_5_c_U31 ( .A(f0_round_5_c_n16), .B(
        f0_round_5_p_io_state_out_1_4), .Z(f0_round_5_io_state_out_1_4) );
  NAND2_X1 f0_round_5_c_U30 ( .A1(f0_round_5_p_io_state_out_3_0), .A2(
        f0_round_5_p_io_state_out_4_0), .ZN(f0_round_5_c_n15) );
  XOR2_X1 f0_round_5_c_U29 ( .A(f0_round_5_c_n15), .B(
        f0_round_5_p_io_state_out_2_0), .Z(f0_round_5_io_state_out_2_0) );
  NAND2_X1 f0_round_5_c_U28 ( .A1(f0_round_5_p_io_state_out_3_1), .A2(
        f0_round_5_p_io_state_out_4_1), .ZN(f0_round_5_c_n14) );
  XOR2_X1 f0_round_5_c_U27 ( .A(f0_round_5_c_n14), .B(
        f0_round_5_p_io_state_out_2_1), .Z(f0_round_5_io_state_out_2_1) );
  NAND2_X1 f0_round_5_c_U26 ( .A1(f0_round_5_p_io_state_out_3_2), .A2(
        f0_round_5_p_io_state_out_4_2), .ZN(f0_round_5_c_n13) );
  XOR2_X1 f0_round_5_c_U25 ( .A(f0_round_5_c_n13), .B(
        f0_round_5_p_io_state_out_2_2), .Z(f0_round_5_io_state_out_2_2) );
  NAND2_X1 f0_round_5_c_U24 ( .A1(f0_round_5_p_io_state_out_3_3), .A2(
        f0_round_5_p_io_state_out_4_3), .ZN(f0_round_5_c_n12) );
  XOR2_X1 f0_round_5_c_U23 ( .A(f0_round_5_c_n12), .B(
        f0_round_5_p_io_state_out_2_3), .Z(f0_round_5_io_state_out_2_3) );
  NAND2_X1 f0_round_5_c_U22 ( .A1(f0_round_5_p_io_state_out_3_4), .A2(
        f0_round_5_p_io_state_out_4_4), .ZN(f0_round_5_c_n11) );
  XOR2_X1 f0_round_5_c_U21 ( .A(f0_round_5_c_n11), .B(
        f0_round_5_p_io_state_out_2_4), .Z(f0_round_5_io_state_out_2_4) );
  NAND2_X1 f0_round_5_c_U20 ( .A1(f0_round_5_p_io_state_out_4_0), .A2(
        f0_round_5_p_io_state_out_0_0), .ZN(f0_round_5_c_n10) );
  XOR2_X1 f0_round_5_c_U19 ( .A(f0_round_5_c_n10), .B(
        f0_round_5_p_io_state_out_3_0), .Z(f0_round_5_io_state_out_3_0) );
  NAND2_X1 f0_round_5_c_U18 ( .A1(f0_round_5_p_io_state_out_4_1), .A2(
        f0_round_5_p_io_state_out_0_1), .ZN(f0_round_5_c_n9) );
  XOR2_X1 f0_round_5_c_U17 ( .A(f0_round_5_c_n9), .B(
        f0_round_5_p_io_state_out_3_1), .Z(f0_round_5_io_state_out_3_1) );
  NAND2_X1 f0_round_5_c_U16 ( .A1(f0_round_5_p_io_state_out_4_2), .A2(
        f0_round_5_p_io_state_out_0_2), .ZN(f0_round_5_c_n8) );
  XOR2_X1 f0_round_5_c_U15 ( .A(f0_round_5_c_n8), .B(
        f0_round_5_p_io_state_out_3_2), .Z(f0_round_5_io_state_out_3_2) );
  NAND2_X1 f0_round_5_c_U14 ( .A1(f0_round_5_p_io_state_out_4_3), .A2(
        f0_round_5_p_io_state_out_0_3), .ZN(f0_round_5_c_n7) );
  XOR2_X1 f0_round_5_c_U13 ( .A(f0_round_5_c_n7), .B(
        f0_round_5_p_io_state_out_3_3), .Z(f0_round_5_io_state_out_3_3) );
  NAND2_X1 f0_round_5_c_U12 ( .A1(f0_round_5_p_io_state_out_4_4), .A2(
        f0_round_5_p_io_state_out_0_4), .ZN(f0_round_5_c_n6) );
  XOR2_X1 f0_round_5_c_U11 ( .A(f0_round_5_c_n6), .B(
        f0_round_5_p_io_state_out_3_4), .Z(f0_round_5_io_state_out_3_4) );
  NAND2_X1 f0_round_5_c_U10 ( .A1(f0_round_5_p_io_state_out_1_0), .A2(
        f0_round_5_p_io_state_out_0_0), .ZN(f0_round_5_c_n5) );
  XOR2_X1 f0_round_5_c_U9 ( .A(f0_round_5_c_n5), .B(
        f0_round_5_p_io_state_out_4_0), .Z(f0_round_5_io_state_out_4_0) );
  NAND2_X1 f0_round_5_c_U8 ( .A1(f0_round_5_p_io_state_out_1_1), .A2(
        f0_round_5_p_io_state_out_0_1), .ZN(f0_round_5_c_n4) );
  XOR2_X1 f0_round_5_c_U7 ( .A(f0_round_5_c_n4), .B(
        f0_round_5_p_io_state_out_4_1), .Z(f0_round_5_io_state_out_4_1) );
  NAND2_X1 f0_round_5_c_U6 ( .A1(f0_round_5_p_io_state_out_1_2), .A2(
        f0_round_5_p_io_state_out_0_2), .ZN(f0_round_5_c_n3) );
  XOR2_X1 f0_round_5_c_U5 ( .A(f0_round_5_c_n3), .B(
        f0_round_5_p_io_state_out_4_2), .Z(f0_round_5_io_state_out_4_2) );
  NAND2_X1 f0_round_5_c_U4 ( .A1(f0_round_5_p_io_state_out_1_3), .A2(
        f0_round_5_p_io_state_out_0_3), .ZN(f0_round_5_c_n2) );
  XOR2_X1 f0_round_5_c_U3 ( .A(f0_round_5_c_n2), .B(
        f0_round_5_p_io_state_out_4_3), .Z(f0_round_5_io_state_out_4_3) );
  NAND2_X1 f0_round_5_c_U2 ( .A1(f0_round_5_p_io_state_out_1_4), .A2(
        f0_round_5_p_io_state_out_0_4), .ZN(f0_round_5_c_n1) );
  XOR2_X1 f0_round_5_c_U1 ( .A(f0_round_5_c_n1), .B(
        f0_round_5_p_io_state_out_4_4), .Z(f0_round_5_io_state_out_4_4) );
  INV_X1 f0_round_5_i_U1 ( .A(f0_round_5_c_io_state_out_0_0), .ZN(
        f0_round_5_io_state_out_0_0) );
  XOR2_X1 f0_round_6_t_U50 ( .A(f0_round_5_io_state_out_1_4), .B(
        f0_round_5_io_state_out_1_3), .Z(f0_round_6_t_n25) );
  XNOR2_X1 f0_round_6_t_U49 ( .A(f0_round_5_io_state_out_1_2), .B(
        f0_round_6_t_n25), .ZN(f0_round_6_t_n23) );
  XOR2_X1 f0_round_6_t_U48 ( .A(f0_round_5_io_state_out_1_1), .B(
        f0_round_5_io_state_out_1_0), .Z(f0_round_6_t_n24) );
  XOR2_X1 f0_round_6_t_U47 ( .A(f0_round_6_t_n23), .B(f0_round_6_t_n24), .Z(
        f0_round_6_t_n8) );
  XOR2_X1 f0_round_6_t_U46 ( .A(f0_round_5_io_state_out_4_4), .B(
        f0_round_5_io_state_out_4_3), .Z(f0_round_6_t_n22) );
  XNOR2_X1 f0_round_6_t_U45 ( .A(f0_round_5_io_state_out_4_2), .B(
        f0_round_6_t_n22), .ZN(f0_round_6_t_n20) );
  XOR2_X1 f0_round_6_t_U44 ( .A(f0_round_5_io_state_out_4_1), .B(
        f0_round_5_io_state_out_4_0), .Z(f0_round_6_t_n21) );
  XNOR2_X1 f0_round_6_t_U43 ( .A(f0_round_6_t_n20), .B(f0_round_6_t_n21), .ZN(
        f0_round_6_t_n5) );
  XNOR2_X1 f0_round_6_t_U42 ( .A(f0_round_6_t_n8), .B(f0_round_6_t_n5), .ZN(
        f0_round_6_t_n19) );
  XOR2_X1 f0_round_6_t_U41 ( .A(f0_round_5_io_state_out_0_0), .B(
        f0_round_6_t_n19), .Z(f0_round_6_p_io_state_out_0_0) );
  XOR2_X1 f0_round_6_t_U40 ( .A(f0_round_5_io_state_out_0_1), .B(
        f0_round_6_t_n19), .Z(f0_round_6_p_io_state_out_1_3) );
  XOR2_X1 f0_round_6_t_U39 ( .A(f0_round_5_io_state_out_0_2), .B(
        f0_round_6_t_n19), .Z(f0_round_6_p_io_state_out_2_1) );
  XOR2_X1 f0_round_6_t_U38 ( .A(f0_round_5_io_state_out_0_3), .B(
        f0_round_6_t_n19), .Z(f0_round_6_p_io_state_out_3_4) );
  XOR2_X1 f0_round_6_t_U37 ( .A(f0_round_5_io_state_out_0_4), .B(
        f0_round_6_t_n19), .Z(f0_round_6_p_io_state_out_4_2) );
  XOR2_X1 f0_round_6_t_U36 ( .A(f0_round_5_io_state_out_2_4), .B(
        f0_round_5_io_state_out_2_3), .Z(f0_round_6_t_n18) );
  XNOR2_X1 f0_round_6_t_U35 ( .A(f0_round_5_io_state_out_2_2), .B(
        f0_round_6_t_n18), .ZN(f0_round_6_t_n16) );
  XOR2_X1 f0_round_6_t_U34 ( .A(f0_round_5_io_state_out_2_1), .B(
        f0_round_5_io_state_out_2_0), .Z(f0_round_6_t_n17) );
  XNOR2_X1 f0_round_6_t_U33 ( .A(f0_round_6_t_n16), .B(f0_round_6_t_n17), .ZN(
        f0_round_6_t_n6) );
  XOR2_X1 f0_round_6_t_U32 ( .A(f0_round_5_io_state_out_0_4), .B(
        f0_round_5_io_state_out_0_3), .Z(f0_round_6_t_n15) );
  XNOR2_X1 f0_round_6_t_U31 ( .A(f0_round_5_io_state_out_0_2), .B(
        f0_round_6_t_n15), .ZN(f0_round_6_t_n13) );
  XOR2_X1 f0_round_6_t_U30 ( .A(f0_round_5_io_state_out_0_1), .B(
        f0_round_5_io_state_out_0_0), .Z(f0_round_6_t_n14) );
  XNOR2_X1 f0_round_6_t_U29 ( .A(f0_round_6_t_n13), .B(f0_round_6_t_n14), .ZN(
        f0_round_6_t_n2) );
  XOR2_X1 f0_round_6_t_U28 ( .A(f0_round_6_t_n6), .B(f0_round_6_t_n2), .Z(
        f0_round_6_t_n12) );
  XOR2_X1 f0_round_6_t_U27 ( .A(f0_round_5_io_state_out_1_0), .B(
        f0_round_6_t_n12), .Z(f0_round_6_p_io_state_out_0_2) );
  XOR2_X1 f0_round_6_t_U26 ( .A(f0_round_5_io_state_out_1_1), .B(
        f0_round_6_t_n12), .Z(f0_round_6_p_io_state_out_1_0) );
  XOR2_X1 f0_round_6_t_U25 ( .A(f0_round_5_io_state_out_1_2), .B(
        f0_round_6_t_n12), .Z(f0_round_6_p_io_state_out_2_3) );
  XOR2_X1 f0_round_6_t_U24 ( .A(f0_round_5_io_state_out_1_3), .B(
        f0_round_6_t_n12), .Z(f0_round_6_p_io_state_out_3_1) );
  XOR2_X1 f0_round_6_t_U23 ( .A(f0_round_5_io_state_out_1_4), .B(
        f0_round_6_t_n12), .Z(f0_round_6_p_io_state_out_4_4) );
  XOR2_X1 f0_round_6_t_U22 ( .A(f0_round_5_io_state_out_3_4), .B(
        f0_round_5_io_state_out_3_3), .Z(f0_round_6_t_n11) );
  XNOR2_X1 f0_round_6_t_U21 ( .A(f0_round_5_io_state_out_3_2), .B(
        f0_round_6_t_n11), .ZN(f0_round_6_t_n9) );
  XOR2_X1 f0_round_6_t_U20 ( .A(f0_round_5_io_state_out_3_1), .B(
        f0_round_5_io_state_out_3_0), .Z(f0_round_6_t_n10) );
  XNOR2_X1 f0_round_6_t_U19 ( .A(f0_round_6_t_n9), .B(f0_round_6_t_n10), .ZN(
        f0_round_6_t_n3) );
  XNOR2_X1 f0_round_6_t_U18 ( .A(f0_round_6_t_n8), .B(f0_round_6_t_n3), .ZN(
        f0_round_6_t_n7) );
  XOR2_X1 f0_round_6_t_U17 ( .A(f0_round_5_io_state_out_2_0), .B(
        f0_round_6_t_n7), .Z(f0_round_6_p_io_state_out_0_4) );
  XOR2_X1 f0_round_6_t_U16 ( .A(f0_round_5_io_state_out_2_1), .B(
        f0_round_6_t_n7), .Z(f0_round_6_p_io_state_out_1_2) );
  XOR2_X1 f0_round_6_t_U15 ( .A(f0_round_5_io_state_out_2_2), .B(
        f0_round_6_t_n7), .Z(f0_round_6_p_io_state_out_2_0) );
  XOR2_X1 f0_round_6_t_U14 ( .A(f0_round_5_io_state_out_2_3), .B(
        f0_round_6_t_n7), .Z(f0_round_6_p_io_state_out_3_3) );
  XOR2_X1 f0_round_6_t_U13 ( .A(f0_round_5_io_state_out_2_4), .B(
        f0_round_6_t_n7), .Z(f0_round_6_p_io_state_out_4_1) );
  XOR2_X1 f0_round_6_t_U12 ( .A(f0_round_6_t_n5), .B(f0_round_6_t_n6), .Z(
        f0_round_6_t_n4) );
  XOR2_X1 f0_round_6_t_U11 ( .A(f0_round_5_io_state_out_3_0), .B(
        f0_round_6_t_n4), .Z(f0_round_6_p_io_state_out_0_1) );
  XOR2_X1 f0_round_6_t_U10 ( .A(f0_round_5_io_state_out_3_1), .B(
        f0_round_6_t_n4), .Z(f0_round_6_p_io_state_out_1_4) );
  XOR2_X1 f0_round_6_t_U9 ( .A(f0_round_5_io_state_out_3_2), .B(
        f0_round_6_t_n4), .Z(f0_round_6_p_io_state_out_2_2) );
  XOR2_X1 f0_round_6_t_U8 ( .A(f0_round_5_io_state_out_3_3), .B(
        f0_round_6_t_n4), .Z(f0_round_6_p_io_state_out_3_0) );
  XOR2_X1 f0_round_6_t_U7 ( .A(f0_round_5_io_state_out_3_4), .B(
        f0_round_6_t_n4), .Z(f0_round_6_p_io_state_out_4_3) );
  XOR2_X1 f0_round_6_t_U6 ( .A(f0_round_6_t_n2), .B(f0_round_6_t_n3), .Z(
        f0_round_6_t_n1) );
  XOR2_X1 f0_round_6_t_U5 ( .A(f0_round_5_io_state_out_4_0), .B(
        f0_round_6_t_n1), .Z(f0_round_6_p_io_state_out_0_3) );
  XOR2_X1 f0_round_6_t_U4 ( .A(f0_round_5_io_state_out_4_1), .B(
        f0_round_6_t_n1), .Z(f0_round_6_p_io_state_out_1_1) );
  XOR2_X1 f0_round_6_t_U3 ( .A(f0_round_5_io_state_out_4_2), .B(
        f0_round_6_t_n1), .Z(f0_round_6_p_io_state_out_2_4) );
  XOR2_X1 f0_round_6_t_U2 ( .A(f0_round_5_io_state_out_4_3), .B(
        f0_round_6_t_n1), .Z(f0_round_6_p_io_state_out_3_2) );
  XOR2_X1 f0_round_6_t_U1 ( .A(f0_round_5_io_state_out_4_4), .B(
        f0_round_6_t_n1), .Z(f0_round_6_p_io_state_out_4_0) );
  NAND2_X1 f0_round_6_c_U50 ( .A1(f0_round_6_p_io_state_out_2_0), .A2(
        f0_round_6_p_io_state_out_1_0), .ZN(f0_round_6_c_n25) );
  XOR2_X1 f0_round_6_c_U49 ( .A(f0_round_6_c_n25), .B(
        f0_round_6_p_io_state_out_0_0), .Z(f0_round_6_c_io_state_out_0_0) );
  NAND2_X1 f0_round_6_c_U48 ( .A1(f0_round_6_p_io_state_out_2_1), .A2(
        f0_round_6_p_io_state_out_1_1), .ZN(f0_round_6_c_n24) );
  XOR2_X1 f0_round_6_c_U47 ( .A(f0_round_6_c_n24), .B(
        f0_round_6_p_io_state_out_0_1), .Z(f0_round_6_io_state_out_0_1) );
  NAND2_X1 f0_round_6_c_U46 ( .A1(f0_round_6_p_io_state_out_2_2), .A2(
        f0_round_6_p_io_state_out_1_2), .ZN(f0_round_6_c_n23) );
  XOR2_X1 f0_round_6_c_U45 ( .A(f0_round_6_c_n23), .B(
        f0_round_6_p_io_state_out_0_2), .Z(f0_round_6_io_state_out_0_2) );
  NAND2_X1 f0_round_6_c_U44 ( .A1(f0_round_6_p_io_state_out_2_3), .A2(
        f0_round_6_p_io_state_out_1_3), .ZN(f0_round_6_c_n22) );
  XOR2_X1 f0_round_6_c_U43 ( .A(f0_round_6_c_n22), .B(
        f0_round_6_p_io_state_out_0_3), .Z(f0_round_6_io_state_out_0_3) );
  NAND2_X1 f0_round_6_c_U42 ( .A1(f0_round_6_p_io_state_out_2_4), .A2(
        f0_round_6_p_io_state_out_1_4), .ZN(f0_round_6_c_n21) );
  XOR2_X1 f0_round_6_c_U41 ( .A(f0_round_6_c_n21), .B(
        f0_round_6_p_io_state_out_0_4), .Z(f0_round_6_io_state_out_0_4) );
  NAND2_X1 f0_round_6_c_U40 ( .A1(f0_round_6_p_io_state_out_2_0), .A2(
        f0_round_6_p_io_state_out_3_0), .ZN(f0_round_6_c_n20) );
  XOR2_X1 f0_round_6_c_U39 ( .A(f0_round_6_c_n20), .B(
        f0_round_6_p_io_state_out_1_0), .Z(f0_round_6_io_state_out_1_0) );
  NAND2_X1 f0_round_6_c_U38 ( .A1(f0_round_6_p_io_state_out_2_1), .A2(
        f0_round_6_p_io_state_out_3_1), .ZN(f0_round_6_c_n19) );
  XOR2_X1 f0_round_6_c_U37 ( .A(f0_round_6_c_n19), .B(
        f0_round_6_p_io_state_out_1_1), .Z(f0_round_6_io_state_out_1_1) );
  NAND2_X1 f0_round_6_c_U36 ( .A1(f0_round_6_p_io_state_out_2_2), .A2(
        f0_round_6_p_io_state_out_3_2), .ZN(f0_round_6_c_n18) );
  XOR2_X1 f0_round_6_c_U35 ( .A(f0_round_6_c_n18), .B(
        f0_round_6_p_io_state_out_1_2), .Z(f0_round_6_io_state_out_1_2) );
  NAND2_X1 f0_round_6_c_U34 ( .A1(f0_round_6_p_io_state_out_2_3), .A2(
        f0_round_6_p_io_state_out_3_3), .ZN(f0_round_6_c_n17) );
  XOR2_X1 f0_round_6_c_U33 ( .A(f0_round_6_c_n17), .B(
        f0_round_6_p_io_state_out_1_3), .Z(f0_round_6_io_state_out_1_3) );
  NAND2_X1 f0_round_6_c_U32 ( .A1(f0_round_6_p_io_state_out_2_4), .A2(
        f0_round_6_p_io_state_out_3_4), .ZN(f0_round_6_c_n16) );
  XOR2_X1 f0_round_6_c_U31 ( .A(f0_round_6_c_n16), .B(
        f0_round_6_p_io_state_out_1_4), .Z(f0_round_6_io_state_out_1_4) );
  NAND2_X1 f0_round_6_c_U30 ( .A1(f0_round_6_p_io_state_out_3_0), .A2(
        f0_round_6_p_io_state_out_4_0), .ZN(f0_round_6_c_n15) );
  XOR2_X1 f0_round_6_c_U29 ( .A(f0_round_6_c_n15), .B(
        f0_round_6_p_io_state_out_2_0), .Z(f0_round_6_io_state_out_2_0) );
  NAND2_X1 f0_round_6_c_U28 ( .A1(f0_round_6_p_io_state_out_3_1), .A2(
        f0_round_6_p_io_state_out_4_1), .ZN(f0_round_6_c_n14) );
  XOR2_X1 f0_round_6_c_U27 ( .A(f0_round_6_c_n14), .B(
        f0_round_6_p_io_state_out_2_1), .Z(f0_round_6_io_state_out_2_1) );
  NAND2_X1 f0_round_6_c_U26 ( .A1(f0_round_6_p_io_state_out_3_2), .A2(
        f0_round_6_p_io_state_out_4_2), .ZN(f0_round_6_c_n13) );
  XOR2_X1 f0_round_6_c_U25 ( .A(f0_round_6_c_n13), .B(
        f0_round_6_p_io_state_out_2_2), .Z(f0_round_6_io_state_out_2_2) );
  NAND2_X1 f0_round_6_c_U24 ( .A1(f0_round_6_p_io_state_out_3_3), .A2(
        f0_round_6_p_io_state_out_4_3), .ZN(f0_round_6_c_n12) );
  XOR2_X1 f0_round_6_c_U23 ( .A(f0_round_6_c_n12), .B(
        f0_round_6_p_io_state_out_2_3), .Z(f0_round_6_io_state_out_2_3) );
  NAND2_X1 f0_round_6_c_U22 ( .A1(f0_round_6_p_io_state_out_3_4), .A2(
        f0_round_6_p_io_state_out_4_4), .ZN(f0_round_6_c_n11) );
  XOR2_X1 f0_round_6_c_U21 ( .A(f0_round_6_c_n11), .B(
        f0_round_6_p_io_state_out_2_4), .Z(f0_round_6_io_state_out_2_4) );
  NAND2_X1 f0_round_6_c_U20 ( .A1(f0_round_6_p_io_state_out_4_0), .A2(
        f0_round_6_p_io_state_out_0_0), .ZN(f0_round_6_c_n10) );
  XOR2_X1 f0_round_6_c_U19 ( .A(f0_round_6_c_n10), .B(
        f0_round_6_p_io_state_out_3_0), .Z(f0_round_6_io_state_out_3_0) );
  NAND2_X1 f0_round_6_c_U18 ( .A1(f0_round_6_p_io_state_out_4_1), .A2(
        f0_round_6_p_io_state_out_0_1), .ZN(f0_round_6_c_n9) );
  XOR2_X1 f0_round_6_c_U17 ( .A(f0_round_6_c_n9), .B(
        f0_round_6_p_io_state_out_3_1), .Z(f0_round_6_io_state_out_3_1) );
  NAND2_X1 f0_round_6_c_U16 ( .A1(f0_round_6_p_io_state_out_4_2), .A2(
        f0_round_6_p_io_state_out_0_2), .ZN(f0_round_6_c_n8) );
  XOR2_X1 f0_round_6_c_U15 ( .A(f0_round_6_c_n8), .B(
        f0_round_6_p_io_state_out_3_2), .Z(f0_round_6_io_state_out_3_2) );
  NAND2_X1 f0_round_6_c_U14 ( .A1(f0_round_6_p_io_state_out_4_3), .A2(
        f0_round_6_p_io_state_out_0_3), .ZN(f0_round_6_c_n7) );
  XOR2_X1 f0_round_6_c_U13 ( .A(f0_round_6_c_n7), .B(
        f0_round_6_p_io_state_out_3_3), .Z(f0_round_6_io_state_out_3_3) );
  NAND2_X1 f0_round_6_c_U12 ( .A1(f0_round_6_p_io_state_out_4_4), .A2(
        f0_round_6_p_io_state_out_0_4), .ZN(f0_round_6_c_n6) );
  XOR2_X1 f0_round_6_c_U11 ( .A(f0_round_6_c_n6), .B(
        f0_round_6_p_io_state_out_3_4), .Z(f0_round_6_io_state_out_3_4) );
  NAND2_X1 f0_round_6_c_U10 ( .A1(f0_round_6_p_io_state_out_1_0), .A2(
        f0_round_6_p_io_state_out_0_0), .ZN(f0_round_6_c_n5) );
  XOR2_X1 f0_round_6_c_U9 ( .A(f0_round_6_c_n5), .B(
        f0_round_6_p_io_state_out_4_0), .Z(f0_round_6_io_state_out_4_0) );
  NAND2_X1 f0_round_6_c_U8 ( .A1(f0_round_6_p_io_state_out_1_1), .A2(
        f0_round_6_p_io_state_out_0_1), .ZN(f0_round_6_c_n4) );
  XOR2_X1 f0_round_6_c_U7 ( .A(f0_round_6_c_n4), .B(
        f0_round_6_p_io_state_out_4_1), .Z(f0_round_6_io_state_out_4_1) );
  NAND2_X1 f0_round_6_c_U6 ( .A1(f0_round_6_p_io_state_out_1_2), .A2(
        f0_round_6_p_io_state_out_0_2), .ZN(f0_round_6_c_n3) );
  XOR2_X1 f0_round_6_c_U5 ( .A(f0_round_6_c_n3), .B(
        f0_round_6_p_io_state_out_4_2), .Z(f0_round_6_io_state_out_4_2) );
  NAND2_X1 f0_round_6_c_U4 ( .A1(f0_round_6_p_io_state_out_1_3), .A2(
        f0_round_6_p_io_state_out_0_3), .ZN(f0_round_6_c_n2) );
  XOR2_X1 f0_round_6_c_U3 ( .A(f0_round_6_c_n2), .B(
        f0_round_6_p_io_state_out_4_3), .Z(f0_round_6_io_state_out_4_3) );
  NAND2_X1 f0_round_6_c_U2 ( .A1(f0_round_6_p_io_state_out_1_4), .A2(
        f0_round_6_p_io_state_out_0_4), .ZN(f0_round_6_c_n1) );
  XOR2_X1 f0_round_6_c_U1 ( .A(f0_round_6_c_n1), .B(
        f0_round_6_p_io_state_out_4_4), .Z(f0_round_6_io_state_out_4_4) );
  INV_X1 f0_round_6_i_U1 ( .A(f0_round_6_c_io_state_out_0_0), .ZN(
        f0_round_6_io_state_out_0_0) );
  XOR2_X1 f0_round_7_t_U50 ( .A(f0_round_6_io_state_out_1_4), .B(
        f0_round_6_io_state_out_1_3), .Z(f0_round_7_t_n25) );
  XNOR2_X1 f0_round_7_t_U49 ( .A(f0_round_6_io_state_out_1_2), .B(
        f0_round_7_t_n25), .ZN(f0_round_7_t_n23) );
  XOR2_X1 f0_round_7_t_U48 ( .A(f0_round_6_io_state_out_1_1), .B(
        f0_round_6_io_state_out_1_0), .Z(f0_round_7_t_n24) );
  XOR2_X1 f0_round_7_t_U47 ( .A(f0_round_7_t_n23), .B(f0_round_7_t_n24), .Z(
        f0_round_7_t_n8) );
  XOR2_X1 f0_round_7_t_U46 ( .A(f0_round_6_io_state_out_4_4), .B(
        f0_round_6_io_state_out_4_3), .Z(f0_round_7_t_n22) );
  XNOR2_X1 f0_round_7_t_U45 ( .A(f0_round_6_io_state_out_4_2), .B(
        f0_round_7_t_n22), .ZN(f0_round_7_t_n20) );
  XOR2_X1 f0_round_7_t_U44 ( .A(f0_round_6_io_state_out_4_1), .B(
        f0_round_6_io_state_out_4_0), .Z(f0_round_7_t_n21) );
  XNOR2_X1 f0_round_7_t_U43 ( .A(f0_round_7_t_n20), .B(f0_round_7_t_n21), .ZN(
        f0_round_7_t_n5) );
  XNOR2_X1 f0_round_7_t_U42 ( .A(f0_round_7_t_n8), .B(f0_round_7_t_n5), .ZN(
        f0_round_7_t_n19) );
  XOR2_X1 f0_round_7_t_U41 ( .A(f0_round_6_io_state_out_0_0), .B(
        f0_round_7_t_n19), .Z(f0_round_7_p_io_state_out_0_0) );
  XOR2_X1 f0_round_7_t_U40 ( .A(f0_round_6_io_state_out_0_1), .B(
        f0_round_7_t_n19), .Z(f0_round_7_p_io_state_out_1_3) );
  XOR2_X1 f0_round_7_t_U39 ( .A(f0_round_6_io_state_out_0_2), .B(
        f0_round_7_t_n19), .Z(f0_round_7_p_io_state_out_2_1) );
  XOR2_X1 f0_round_7_t_U38 ( .A(f0_round_6_io_state_out_0_3), .B(
        f0_round_7_t_n19), .Z(f0_round_7_p_io_state_out_3_4) );
  XOR2_X1 f0_round_7_t_U37 ( .A(f0_round_6_io_state_out_0_4), .B(
        f0_round_7_t_n19), .Z(f0_round_7_p_io_state_out_4_2) );
  XOR2_X1 f0_round_7_t_U36 ( .A(f0_round_6_io_state_out_2_4), .B(
        f0_round_6_io_state_out_2_3), .Z(f0_round_7_t_n18) );
  XNOR2_X1 f0_round_7_t_U35 ( .A(f0_round_6_io_state_out_2_2), .B(
        f0_round_7_t_n18), .ZN(f0_round_7_t_n16) );
  XOR2_X1 f0_round_7_t_U34 ( .A(f0_round_6_io_state_out_2_1), .B(
        f0_round_6_io_state_out_2_0), .Z(f0_round_7_t_n17) );
  XNOR2_X1 f0_round_7_t_U33 ( .A(f0_round_7_t_n16), .B(f0_round_7_t_n17), .ZN(
        f0_round_7_t_n6) );
  XOR2_X1 f0_round_7_t_U32 ( .A(f0_round_6_io_state_out_0_4), .B(
        f0_round_6_io_state_out_0_3), .Z(f0_round_7_t_n15) );
  XNOR2_X1 f0_round_7_t_U31 ( .A(f0_round_6_io_state_out_0_2), .B(
        f0_round_7_t_n15), .ZN(f0_round_7_t_n13) );
  XOR2_X1 f0_round_7_t_U30 ( .A(f0_round_6_io_state_out_0_1), .B(
        f0_round_6_io_state_out_0_0), .Z(f0_round_7_t_n14) );
  XNOR2_X1 f0_round_7_t_U29 ( .A(f0_round_7_t_n13), .B(f0_round_7_t_n14), .ZN(
        f0_round_7_t_n2) );
  XOR2_X1 f0_round_7_t_U28 ( .A(f0_round_7_t_n6), .B(f0_round_7_t_n2), .Z(
        f0_round_7_t_n12) );
  XOR2_X1 f0_round_7_t_U27 ( .A(f0_round_6_io_state_out_1_0), .B(
        f0_round_7_t_n12), .Z(f0_round_7_p_io_state_out_0_2) );
  XOR2_X1 f0_round_7_t_U26 ( .A(f0_round_6_io_state_out_1_1), .B(
        f0_round_7_t_n12), .Z(f0_round_7_p_io_state_out_1_0) );
  XOR2_X1 f0_round_7_t_U25 ( .A(f0_round_6_io_state_out_1_2), .B(
        f0_round_7_t_n12), .Z(f0_round_7_p_io_state_out_2_3) );
  XOR2_X1 f0_round_7_t_U24 ( .A(f0_round_6_io_state_out_1_3), .B(
        f0_round_7_t_n12), .Z(f0_round_7_p_io_state_out_3_1) );
  XOR2_X1 f0_round_7_t_U23 ( .A(f0_round_6_io_state_out_1_4), .B(
        f0_round_7_t_n12), .Z(f0_round_7_p_io_state_out_4_4) );
  XOR2_X1 f0_round_7_t_U22 ( .A(f0_round_6_io_state_out_3_4), .B(
        f0_round_6_io_state_out_3_3), .Z(f0_round_7_t_n11) );
  XNOR2_X1 f0_round_7_t_U21 ( .A(f0_round_6_io_state_out_3_2), .B(
        f0_round_7_t_n11), .ZN(f0_round_7_t_n9) );
  XOR2_X1 f0_round_7_t_U20 ( .A(f0_round_6_io_state_out_3_1), .B(
        f0_round_6_io_state_out_3_0), .Z(f0_round_7_t_n10) );
  XNOR2_X1 f0_round_7_t_U19 ( .A(f0_round_7_t_n9), .B(f0_round_7_t_n10), .ZN(
        f0_round_7_t_n3) );
  XNOR2_X1 f0_round_7_t_U18 ( .A(f0_round_7_t_n8), .B(f0_round_7_t_n3), .ZN(
        f0_round_7_t_n7) );
  XOR2_X1 f0_round_7_t_U17 ( .A(f0_round_6_io_state_out_2_0), .B(
        f0_round_7_t_n7), .Z(f0_round_7_p_io_state_out_0_4) );
  XOR2_X1 f0_round_7_t_U16 ( .A(f0_round_6_io_state_out_2_1), .B(
        f0_round_7_t_n7), .Z(f0_round_7_p_io_state_out_1_2) );
  XOR2_X1 f0_round_7_t_U15 ( .A(f0_round_6_io_state_out_2_2), .B(
        f0_round_7_t_n7), .Z(f0_round_7_p_io_state_out_2_0) );
  XOR2_X1 f0_round_7_t_U14 ( .A(f0_round_6_io_state_out_2_3), .B(
        f0_round_7_t_n7), .Z(f0_round_7_p_io_state_out_3_3) );
  XOR2_X1 f0_round_7_t_U13 ( .A(f0_round_6_io_state_out_2_4), .B(
        f0_round_7_t_n7), .Z(f0_round_7_p_io_state_out_4_1) );
  XOR2_X1 f0_round_7_t_U12 ( .A(f0_round_7_t_n5), .B(f0_round_7_t_n6), .Z(
        f0_round_7_t_n4) );
  XOR2_X1 f0_round_7_t_U11 ( .A(f0_round_6_io_state_out_3_0), .B(
        f0_round_7_t_n4), .Z(f0_round_7_p_io_state_out_0_1) );
  XOR2_X1 f0_round_7_t_U10 ( .A(f0_round_6_io_state_out_3_1), .B(
        f0_round_7_t_n4), .Z(f0_round_7_p_io_state_out_1_4) );
  XOR2_X1 f0_round_7_t_U9 ( .A(f0_round_6_io_state_out_3_2), .B(
        f0_round_7_t_n4), .Z(f0_round_7_p_io_state_out_2_2) );
  XOR2_X1 f0_round_7_t_U8 ( .A(f0_round_6_io_state_out_3_3), .B(
        f0_round_7_t_n4), .Z(f0_round_7_p_io_state_out_3_0) );
  XOR2_X1 f0_round_7_t_U7 ( .A(f0_round_6_io_state_out_3_4), .B(
        f0_round_7_t_n4), .Z(f0_round_7_p_io_state_out_4_3) );
  XOR2_X1 f0_round_7_t_U6 ( .A(f0_round_7_t_n2), .B(f0_round_7_t_n3), .Z(
        f0_round_7_t_n1) );
  XOR2_X1 f0_round_7_t_U5 ( .A(f0_round_6_io_state_out_4_0), .B(
        f0_round_7_t_n1), .Z(f0_round_7_p_io_state_out_0_3) );
  XOR2_X1 f0_round_7_t_U4 ( .A(f0_round_6_io_state_out_4_1), .B(
        f0_round_7_t_n1), .Z(f0_round_7_p_io_state_out_1_1) );
  XOR2_X1 f0_round_7_t_U3 ( .A(f0_round_6_io_state_out_4_2), .B(
        f0_round_7_t_n1), .Z(f0_round_7_p_io_state_out_2_4) );
  XOR2_X1 f0_round_7_t_U2 ( .A(f0_round_6_io_state_out_4_3), .B(
        f0_round_7_t_n1), .Z(f0_round_7_p_io_state_out_3_2) );
  XOR2_X1 f0_round_7_t_U1 ( .A(f0_round_6_io_state_out_4_4), .B(
        f0_round_7_t_n1), .Z(f0_round_7_p_io_state_out_4_0) );
  NAND2_X1 f0_round_7_c_U50 ( .A1(f0_round_7_p_io_state_out_2_0), .A2(
        f0_round_7_p_io_state_out_1_0), .ZN(f0_round_7_c_n25) );
  XOR2_X1 f0_round_7_c_U49 ( .A(f0_round_7_c_n25), .B(
        f0_round_7_p_io_state_out_0_0), .Z(f0_round_7_io_state_out_0_0) );
  NAND2_X1 f0_round_7_c_U48 ( .A1(f0_round_7_p_io_state_out_2_1), .A2(
        f0_round_7_p_io_state_out_1_1), .ZN(f0_round_7_c_n24) );
  XOR2_X1 f0_round_7_c_U47 ( .A(f0_round_7_c_n24), .B(
        f0_round_7_p_io_state_out_0_1), .Z(f0_round_7_io_state_out_0_1) );
  NAND2_X1 f0_round_7_c_U46 ( .A1(f0_round_7_p_io_state_out_2_2), .A2(
        f0_round_7_p_io_state_out_1_2), .ZN(f0_round_7_c_n23) );
  XOR2_X1 f0_round_7_c_U45 ( .A(f0_round_7_c_n23), .B(
        f0_round_7_p_io_state_out_0_2), .Z(f0_round_7_io_state_out_0_2) );
  NAND2_X1 f0_round_7_c_U44 ( .A1(f0_round_7_p_io_state_out_2_3), .A2(
        f0_round_7_p_io_state_out_1_3), .ZN(f0_round_7_c_n22) );
  XOR2_X1 f0_round_7_c_U43 ( .A(f0_round_7_c_n22), .B(
        f0_round_7_p_io_state_out_0_3), .Z(f0_round_7_io_state_out_0_3) );
  NAND2_X1 f0_round_7_c_U42 ( .A1(f0_round_7_p_io_state_out_2_4), .A2(
        f0_round_7_p_io_state_out_1_4), .ZN(f0_round_7_c_n21) );
  XOR2_X1 f0_round_7_c_U41 ( .A(f0_round_7_c_n21), .B(
        f0_round_7_p_io_state_out_0_4), .Z(f0_round_7_io_state_out_0_4) );
  NAND2_X1 f0_round_7_c_U40 ( .A1(f0_round_7_p_io_state_out_2_0), .A2(
        f0_round_7_p_io_state_out_3_0), .ZN(f0_round_7_c_n20) );
  XOR2_X1 f0_round_7_c_U39 ( .A(f0_round_7_c_n20), .B(
        f0_round_7_p_io_state_out_1_0), .Z(f0_round_7_io_state_out_1_0) );
  NAND2_X1 f0_round_7_c_U38 ( .A1(f0_round_7_p_io_state_out_2_1), .A2(
        f0_round_7_p_io_state_out_3_1), .ZN(f0_round_7_c_n19) );
  XOR2_X1 f0_round_7_c_U37 ( .A(f0_round_7_c_n19), .B(
        f0_round_7_p_io_state_out_1_1), .Z(f0_round_7_io_state_out_1_1) );
  NAND2_X1 f0_round_7_c_U36 ( .A1(f0_round_7_p_io_state_out_2_2), .A2(
        f0_round_7_p_io_state_out_3_2), .ZN(f0_round_7_c_n18) );
  XOR2_X1 f0_round_7_c_U35 ( .A(f0_round_7_c_n18), .B(
        f0_round_7_p_io_state_out_1_2), .Z(f0_round_7_io_state_out_1_2) );
  NAND2_X1 f0_round_7_c_U34 ( .A1(f0_round_7_p_io_state_out_2_3), .A2(
        f0_round_7_p_io_state_out_3_3), .ZN(f0_round_7_c_n17) );
  XOR2_X1 f0_round_7_c_U33 ( .A(f0_round_7_c_n17), .B(
        f0_round_7_p_io_state_out_1_3), .Z(f0_round_7_io_state_out_1_3) );
  NAND2_X1 f0_round_7_c_U32 ( .A1(f0_round_7_p_io_state_out_2_4), .A2(
        f0_round_7_p_io_state_out_3_4), .ZN(f0_round_7_c_n16) );
  XOR2_X1 f0_round_7_c_U31 ( .A(f0_round_7_c_n16), .B(
        f0_round_7_p_io_state_out_1_4), .Z(f0_round_7_io_state_out_1_4) );
  NAND2_X1 f0_round_7_c_U30 ( .A1(f0_round_7_p_io_state_out_3_0), .A2(
        f0_round_7_p_io_state_out_4_0), .ZN(f0_round_7_c_n15) );
  XOR2_X1 f0_round_7_c_U29 ( .A(f0_round_7_c_n15), .B(
        f0_round_7_p_io_state_out_2_0), .Z(f0_round_7_io_state_out_2_0) );
  NAND2_X1 f0_round_7_c_U28 ( .A1(f0_round_7_p_io_state_out_3_1), .A2(
        f0_round_7_p_io_state_out_4_1), .ZN(f0_round_7_c_n14) );
  XOR2_X1 f0_round_7_c_U27 ( .A(f0_round_7_c_n14), .B(
        f0_round_7_p_io_state_out_2_1), .Z(f0_round_7_io_state_out_2_1) );
  NAND2_X1 f0_round_7_c_U26 ( .A1(f0_round_7_p_io_state_out_3_2), .A2(
        f0_round_7_p_io_state_out_4_2), .ZN(f0_round_7_c_n13) );
  XOR2_X1 f0_round_7_c_U25 ( .A(f0_round_7_c_n13), .B(
        f0_round_7_p_io_state_out_2_2), .Z(f0_round_7_io_state_out_2_2) );
  NAND2_X1 f0_round_7_c_U24 ( .A1(f0_round_7_p_io_state_out_3_3), .A2(
        f0_round_7_p_io_state_out_4_3), .ZN(f0_round_7_c_n12) );
  XOR2_X1 f0_round_7_c_U23 ( .A(f0_round_7_c_n12), .B(
        f0_round_7_p_io_state_out_2_3), .Z(f0_round_7_io_state_out_2_3) );
  NAND2_X1 f0_round_7_c_U22 ( .A1(f0_round_7_p_io_state_out_3_4), .A2(
        f0_round_7_p_io_state_out_4_4), .ZN(f0_round_7_c_n11) );
  XOR2_X1 f0_round_7_c_U21 ( .A(f0_round_7_c_n11), .B(
        f0_round_7_p_io_state_out_2_4), .Z(f0_round_7_io_state_out_2_4) );
  NAND2_X1 f0_round_7_c_U20 ( .A1(f0_round_7_p_io_state_out_4_0), .A2(
        f0_round_7_p_io_state_out_0_0), .ZN(f0_round_7_c_n10) );
  XOR2_X1 f0_round_7_c_U19 ( .A(f0_round_7_c_n10), .B(
        f0_round_7_p_io_state_out_3_0), .Z(f0_round_7_io_state_out_3_0) );
  NAND2_X1 f0_round_7_c_U18 ( .A1(f0_round_7_p_io_state_out_4_1), .A2(
        f0_round_7_p_io_state_out_0_1), .ZN(f0_round_7_c_n9) );
  XOR2_X1 f0_round_7_c_U17 ( .A(f0_round_7_c_n9), .B(
        f0_round_7_p_io_state_out_3_1), .Z(f0_round_7_io_state_out_3_1) );
  NAND2_X1 f0_round_7_c_U16 ( .A1(f0_round_7_p_io_state_out_4_2), .A2(
        f0_round_7_p_io_state_out_0_2), .ZN(f0_round_7_c_n8) );
  XOR2_X1 f0_round_7_c_U15 ( .A(f0_round_7_c_n8), .B(
        f0_round_7_p_io_state_out_3_2), .Z(f0_round_7_io_state_out_3_2) );
  NAND2_X1 f0_round_7_c_U14 ( .A1(f0_round_7_p_io_state_out_4_3), .A2(
        f0_round_7_p_io_state_out_0_3), .ZN(f0_round_7_c_n7) );
  XOR2_X1 f0_round_7_c_U13 ( .A(f0_round_7_c_n7), .B(
        f0_round_7_p_io_state_out_3_3), .Z(f0_round_7_io_state_out_3_3) );
  NAND2_X1 f0_round_7_c_U12 ( .A1(f0_round_7_p_io_state_out_4_4), .A2(
        f0_round_7_p_io_state_out_0_4), .ZN(f0_round_7_c_n6) );
  XOR2_X1 f0_round_7_c_U11 ( .A(f0_round_7_c_n6), .B(
        f0_round_7_p_io_state_out_3_4), .Z(f0_round_7_io_state_out_3_4) );
  NAND2_X1 f0_round_7_c_U10 ( .A1(f0_round_7_p_io_state_out_1_0), .A2(
        f0_round_7_p_io_state_out_0_0), .ZN(f0_round_7_c_n5) );
  XOR2_X1 f0_round_7_c_U9 ( .A(f0_round_7_c_n5), .B(
        f0_round_7_p_io_state_out_4_0), .Z(f0_round_7_io_state_out_4_0) );
  NAND2_X1 f0_round_7_c_U8 ( .A1(f0_round_7_p_io_state_out_1_1), .A2(
        f0_round_7_p_io_state_out_0_1), .ZN(f0_round_7_c_n4) );
  XOR2_X1 f0_round_7_c_U7 ( .A(f0_round_7_c_n4), .B(
        f0_round_7_p_io_state_out_4_1), .Z(f0_round_7_io_state_out_4_1) );
  NAND2_X1 f0_round_7_c_U6 ( .A1(f0_round_7_p_io_state_out_1_2), .A2(
        f0_round_7_p_io_state_out_0_2), .ZN(f0_round_7_c_n3) );
  XOR2_X1 f0_round_7_c_U5 ( .A(f0_round_7_c_n3), .B(
        f0_round_7_p_io_state_out_4_2), .Z(f0_round_7_io_state_out_4_2) );
  NAND2_X1 f0_round_7_c_U4 ( .A1(f0_round_7_p_io_state_out_1_3), .A2(
        f0_round_7_p_io_state_out_0_3), .ZN(f0_round_7_c_n2) );
  XOR2_X1 f0_round_7_c_U3 ( .A(f0_round_7_c_n2), .B(
        f0_round_7_p_io_state_out_4_3), .Z(f0_round_7_io_state_out_4_3) );
  NAND2_X1 f0_round_7_c_U2 ( .A1(f0_round_7_p_io_state_out_1_4), .A2(
        f0_round_7_p_io_state_out_0_4), .ZN(f0_round_7_c_n1) );
  XOR2_X1 f0_round_7_c_U1 ( .A(f0_round_7_c_n1), .B(
        f0_round_7_p_io_state_out_4_4), .Z(f0_round_7_io_state_out_4_4) );
  XOR2_X1 f0_round_8_t_U50 ( .A(f0_round_7_io_state_out_1_4), .B(
        f0_round_7_io_state_out_1_3), .Z(f0_round_8_t_n25) );
  XNOR2_X1 f0_round_8_t_U49 ( .A(f0_round_7_io_state_out_1_2), .B(
        f0_round_8_t_n25), .ZN(f0_round_8_t_n23) );
  XOR2_X1 f0_round_8_t_U48 ( .A(f0_round_7_io_state_out_1_1), .B(
        f0_round_7_io_state_out_1_0), .Z(f0_round_8_t_n24) );
  XOR2_X1 f0_round_8_t_U47 ( .A(f0_round_8_t_n23), .B(f0_round_8_t_n24), .Z(
        f0_round_8_t_n8) );
  XOR2_X1 f0_round_8_t_U46 ( .A(f0_round_7_io_state_out_4_4), .B(
        f0_round_7_io_state_out_4_3), .Z(f0_round_8_t_n22) );
  XNOR2_X1 f0_round_8_t_U45 ( .A(f0_round_7_io_state_out_4_2), .B(
        f0_round_8_t_n22), .ZN(f0_round_8_t_n20) );
  XOR2_X1 f0_round_8_t_U44 ( .A(f0_round_7_io_state_out_4_1), .B(
        f0_round_7_io_state_out_4_0), .Z(f0_round_8_t_n21) );
  XNOR2_X1 f0_round_8_t_U43 ( .A(f0_round_8_t_n20), .B(f0_round_8_t_n21), .ZN(
        f0_round_8_t_n5) );
  XNOR2_X1 f0_round_8_t_U42 ( .A(f0_round_8_t_n8), .B(f0_round_8_t_n5), .ZN(
        f0_round_8_t_n19) );
  XOR2_X1 f0_round_8_t_U41 ( .A(f0_round_7_io_state_out_0_0), .B(
        f0_round_8_t_n19), .Z(f0_round_8_p_io_state_out_0_0) );
  XOR2_X1 f0_round_8_t_U40 ( .A(f0_round_7_io_state_out_0_1), .B(
        f0_round_8_t_n19), .Z(f0_round_8_p_io_state_out_1_3) );
  XOR2_X1 f0_round_8_t_U39 ( .A(f0_round_7_io_state_out_0_2), .B(
        f0_round_8_t_n19), .Z(f0_round_8_p_io_state_out_2_1) );
  XOR2_X1 f0_round_8_t_U38 ( .A(f0_round_7_io_state_out_0_3), .B(
        f0_round_8_t_n19), .Z(f0_round_8_p_io_state_out_3_4) );
  XOR2_X1 f0_round_8_t_U37 ( .A(f0_round_7_io_state_out_0_4), .B(
        f0_round_8_t_n19), .Z(f0_round_8_p_io_state_out_4_2) );
  XOR2_X1 f0_round_8_t_U36 ( .A(f0_round_7_io_state_out_2_4), .B(
        f0_round_7_io_state_out_2_3), .Z(f0_round_8_t_n18) );
  XNOR2_X1 f0_round_8_t_U35 ( .A(f0_round_7_io_state_out_2_2), .B(
        f0_round_8_t_n18), .ZN(f0_round_8_t_n16) );
  XOR2_X1 f0_round_8_t_U34 ( .A(f0_round_7_io_state_out_2_1), .B(
        f0_round_7_io_state_out_2_0), .Z(f0_round_8_t_n17) );
  XNOR2_X1 f0_round_8_t_U33 ( .A(f0_round_8_t_n16), .B(f0_round_8_t_n17), .ZN(
        f0_round_8_t_n6) );
  XOR2_X1 f0_round_8_t_U32 ( .A(f0_round_7_io_state_out_0_4), .B(
        f0_round_7_io_state_out_0_3), .Z(f0_round_8_t_n15) );
  XNOR2_X1 f0_round_8_t_U31 ( .A(f0_round_7_io_state_out_0_2), .B(
        f0_round_8_t_n15), .ZN(f0_round_8_t_n13) );
  XOR2_X1 f0_round_8_t_U30 ( .A(f0_round_7_io_state_out_0_1), .B(
        f0_round_7_io_state_out_0_0), .Z(f0_round_8_t_n14) );
  XNOR2_X1 f0_round_8_t_U29 ( .A(f0_round_8_t_n13), .B(f0_round_8_t_n14), .ZN(
        f0_round_8_t_n2) );
  XOR2_X1 f0_round_8_t_U28 ( .A(f0_round_8_t_n6), .B(f0_round_8_t_n2), .Z(
        f0_round_8_t_n12) );
  XOR2_X1 f0_round_8_t_U27 ( .A(f0_round_7_io_state_out_1_0), .B(
        f0_round_8_t_n12), .Z(f0_round_8_p_io_state_out_0_2) );
  XOR2_X1 f0_round_8_t_U26 ( .A(f0_round_7_io_state_out_1_1), .B(
        f0_round_8_t_n12), .Z(f0_round_8_p_io_state_out_1_0) );
  XOR2_X1 f0_round_8_t_U25 ( .A(f0_round_7_io_state_out_1_2), .B(
        f0_round_8_t_n12), .Z(f0_round_8_p_io_state_out_2_3) );
  XOR2_X1 f0_round_8_t_U24 ( .A(f0_round_7_io_state_out_1_3), .B(
        f0_round_8_t_n12), .Z(f0_round_8_p_io_state_out_3_1) );
  XOR2_X1 f0_round_8_t_U23 ( .A(f0_round_7_io_state_out_1_4), .B(
        f0_round_8_t_n12), .Z(f0_round_8_p_io_state_out_4_4) );
  XOR2_X1 f0_round_8_t_U22 ( .A(f0_round_7_io_state_out_3_4), .B(
        f0_round_7_io_state_out_3_3), .Z(f0_round_8_t_n11) );
  XNOR2_X1 f0_round_8_t_U21 ( .A(f0_round_7_io_state_out_3_2), .B(
        f0_round_8_t_n11), .ZN(f0_round_8_t_n9) );
  XOR2_X1 f0_round_8_t_U20 ( .A(f0_round_7_io_state_out_3_1), .B(
        f0_round_7_io_state_out_3_0), .Z(f0_round_8_t_n10) );
  XNOR2_X1 f0_round_8_t_U19 ( .A(f0_round_8_t_n9), .B(f0_round_8_t_n10), .ZN(
        f0_round_8_t_n3) );
  XNOR2_X1 f0_round_8_t_U18 ( .A(f0_round_8_t_n8), .B(f0_round_8_t_n3), .ZN(
        f0_round_8_t_n7) );
  XOR2_X1 f0_round_8_t_U17 ( .A(f0_round_7_io_state_out_2_0), .B(
        f0_round_8_t_n7), .Z(f0_round_8_p_io_state_out_0_4) );
  XOR2_X1 f0_round_8_t_U16 ( .A(f0_round_7_io_state_out_2_1), .B(
        f0_round_8_t_n7), .Z(f0_round_8_p_io_state_out_1_2) );
  XOR2_X1 f0_round_8_t_U15 ( .A(f0_round_7_io_state_out_2_2), .B(
        f0_round_8_t_n7), .Z(f0_round_8_p_io_state_out_2_0) );
  XOR2_X1 f0_round_8_t_U14 ( .A(f0_round_7_io_state_out_2_3), .B(
        f0_round_8_t_n7), .Z(f0_round_8_p_io_state_out_3_3) );
  XOR2_X1 f0_round_8_t_U13 ( .A(f0_round_7_io_state_out_2_4), .B(
        f0_round_8_t_n7), .Z(f0_round_8_p_io_state_out_4_1) );
  XOR2_X1 f0_round_8_t_U12 ( .A(f0_round_8_t_n5), .B(f0_round_8_t_n6), .Z(
        f0_round_8_t_n4) );
  XOR2_X1 f0_round_8_t_U11 ( .A(f0_round_7_io_state_out_3_0), .B(
        f0_round_8_t_n4), .Z(f0_round_8_p_io_state_out_0_1) );
  XOR2_X1 f0_round_8_t_U10 ( .A(f0_round_7_io_state_out_3_1), .B(
        f0_round_8_t_n4), .Z(f0_round_8_p_io_state_out_1_4) );
  XOR2_X1 f0_round_8_t_U9 ( .A(f0_round_7_io_state_out_3_2), .B(
        f0_round_8_t_n4), .Z(f0_round_8_p_io_state_out_2_2) );
  XOR2_X1 f0_round_8_t_U8 ( .A(f0_round_7_io_state_out_3_3), .B(
        f0_round_8_t_n4), .Z(f0_round_8_p_io_state_out_3_0) );
  XOR2_X1 f0_round_8_t_U7 ( .A(f0_round_7_io_state_out_3_4), .B(
        f0_round_8_t_n4), .Z(f0_round_8_p_io_state_out_4_3) );
  XOR2_X1 f0_round_8_t_U6 ( .A(f0_round_8_t_n2), .B(f0_round_8_t_n3), .Z(
        f0_round_8_t_n1) );
  XOR2_X1 f0_round_8_t_U5 ( .A(f0_round_7_io_state_out_4_0), .B(
        f0_round_8_t_n1), .Z(f0_round_8_p_io_state_out_0_3) );
  XOR2_X1 f0_round_8_t_U4 ( .A(f0_round_7_io_state_out_4_1), .B(
        f0_round_8_t_n1), .Z(f0_round_8_p_io_state_out_1_1) );
  XOR2_X1 f0_round_8_t_U3 ( .A(f0_round_7_io_state_out_4_2), .B(
        f0_round_8_t_n1), .Z(f0_round_8_p_io_state_out_2_4) );
  XOR2_X1 f0_round_8_t_U2 ( .A(f0_round_7_io_state_out_4_3), .B(
        f0_round_8_t_n1), .Z(f0_round_8_p_io_state_out_3_2) );
  XOR2_X1 f0_round_8_t_U1 ( .A(f0_round_7_io_state_out_4_4), .B(
        f0_round_8_t_n1), .Z(f0_round_8_p_io_state_out_4_0) );
  NAND2_X1 f0_round_8_c_U50 ( .A1(f0_round_8_p_io_state_out_2_0), .A2(
        f0_round_8_p_io_state_out_1_0), .ZN(f0_round_8_c_n25) );
  XOR2_X1 f0_round_8_c_U49 ( .A(f0_round_8_c_n25), .B(
        f0_round_8_p_io_state_out_0_0), .Z(f0_round_8_io_state_out_0_0) );
  NAND2_X1 f0_round_8_c_U48 ( .A1(f0_round_8_p_io_state_out_2_1), .A2(
        f0_round_8_p_io_state_out_1_1), .ZN(f0_round_8_c_n24) );
  XOR2_X1 f0_round_8_c_U47 ( .A(f0_round_8_c_n24), .B(
        f0_round_8_p_io_state_out_0_1), .Z(f0_round_8_io_state_out_0_1) );
  NAND2_X1 f0_round_8_c_U46 ( .A1(f0_round_8_p_io_state_out_2_2), .A2(
        f0_round_8_p_io_state_out_1_2), .ZN(f0_round_8_c_n23) );
  XOR2_X1 f0_round_8_c_U45 ( .A(f0_round_8_c_n23), .B(
        f0_round_8_p_io_state_out_0_2), .Z(f0_round_8_io_state_out_0_2) );
  NAND2_X1 f0_round_8_c_U44 ( .A1(f0_round_8_p_io_state_out_2_3), .A2(
        f0_round_8_p_io_state_out_1_3), .ZN(f0_round_8_c_n22) );
  XOR2_X1 f0_round_8_c_U43 ( .A(f0_round_8_c_n22), .B(
        f0_round_8_p_io_state_out_0_3), .Z(f0_round_8_io_state_out_0_3) );
  NAND2_X1 f0_round_8_c_U42 ( .A1(f0_round_8_p_io_state_out_2_4), .A2(
        f0_round_8_p_io_state_out_1_4), .ZN(f0_round_8_c_n21) );
  XOR2_X1 f0_round_8_c_U41 ( .A(f0_round_8_c_n21), .B(
        f0_round_8_p_io_state_out_0_4), .Z(f0_round_8_io_state_out_0_4) );
  NAND2_X1 f0_round_8_c_U40 ( .A1(f0_round_8_p_io_state_out_2_0), .A2(
        f0_round_8_p_io_state_out_3_0), .ZN(f0_round_8_c_n20) );
  XOR2_X1 f0_round_8_c_U39 ( .A(f0_round_8_c_n20), .B(
        f0_round_8_p_io_state_out_1_0), .Z(f0_round_8_io_state_out_1_0) );
  NAND2_X1 f0_round_8_c_U38 ( .A1(f0_round_8_p_io_state_out_2_1), .A2(
        f0_round_8_p_io_state_out_3_1), .ZN(f0_round_8_c_n19) );
  XOR2_X1 f0_round_8_c_U37 ( .A(f0_round_8_c_n19), .B(
        f0_round_8_p_io_state_out_1_1), .Z(f0_round_8_io_state_out_1_1) );
  NAND2_X1 f0_round_8_c_U36 ( .A1(f0_round_8_p_io_state_out_2_2), .A2(
        f0_round_8_p_io_state_out_3_2), .ZN(f0_round_8_c_n18) );
  XOR2_X1 f0_round_8_c_U35 ( .A(f0_round_8_c_n18), .B(
        f0_round_8_p_io_state_out_1_2), .Z(f0_round_8_io_state_out_1_2) );
  NAND2_X1 f0_round_8_c_U34 ( .A1(f0_round_8_p_io_state_out_2_3), .A2(
        f0_round_8_p_io_state_out_3_3), .ZN(f0_round_8_c_n17) );
  XOR2_X1 f0_round_8_c_U33 ( .A(f0_round_8_c_n17), .B(
        f0_round_8_p_io_state_out_1_3), .Z(f0_round_8_io_state_out_1_3) );
  NAND2_X1 f0_round_8_c_U32 ( .A1(f0_round_8_p_io_state_out_2_4), .A2(
        f0_round_8_p_io_state_out_3_4), .ZN(f0_round_8_c_n16) );
  XOR2_X1 f0_round_8_c_U31 ( .A(f0_round_8_c_n16), .B(
        f0_round_8_p_io_state_out_1_4), .Z(f0_round_8_io_state_out_1_4) );
  NAND2_X1 f0_round_8_c_U30 ( .A1(f0_round_8_p_io_state_out_3_0), .A2(
        f0_round_8_p_io_state_out_4_0), .ZN(f0_round_8_c_n15) );
  XOR2_X1 f0_round_8_c_U29 ( .A(f0_round_8_c_n15), .B(
        f0_round_8_p_io_state_out_2_0), .Z(f0_round_8_io_state_out_2_0) );
  NAND2_X1 f0_round_8_c_U28 ( .A1(f0_round_8_p_io_state_out_3_1), .A2(
        f0_round_8_p_io_state_out_4_1), .ZN(f0_round_8_c_n14) );
  XOR2_X1 f0_round_8_c_U27 ( .A(f0_round_8_c_n14), .B(
        f0_round_8_p_io_state_out_2_1), .Z(f0_round_8_io_state_out_2_1) );
  NAND2_X1 f0_round_8_c_U26 ( .A1(f0_round_8_p_io_state_out_3_2), .A2(
        f0_round_8_p_io_state_out_4_2), .ZN(f0_round_8_c_n13) );
  XOR2_X1 f0_round_8_c_U25 ( .A(f0_round_8_c_n13), .B(
        f0_round_8_p_io_state_out_2_2), .Z(f0_round_8_io_state_out_2_2) );
  NAND2_X1 f0_round_8_c_U24 ( .A1(f0_round_8_p_io_state_out_3_3), .A2(
        f0_round_8_p_io_state_out_4_3), .ZN(f0_round_8_c_n12) );
  XOR2_X1 f0_round_8_c_U23 ( .A(f0_round_8_c_n12), .B(
        f0_round_8_p_io_state_out_2_3), .Z(f0_round_8_io_state_out_2_3) );
  NAND2_X1 f0_round_8_c_U22 ( .A1(f0_round_8_p_io_state_out_3_4), .A2(
        f0_round_8_p_io_state_out_4_4), .ZN(f0_round_8_c_n11) );
  XOR2_X1 f0_round_8_c_U21 ( .A(f0_round_8_c_n11), .B(
        f0_round_8_p_io_state_out_2_4), .Z(f0_round_8_io_state_out_2_4) );
  NAND2_X1 f0_round_8_c_U20 ( .A1(f0_round_8_p_io_state_out_4_0), .A2(
        f0_round_8_p_io_state_out_0_0), .ZN(f0_round_8_c_n10) );
  XOR2_X1 f0_round_8_c_U19 ( .A(f0_round_8_c_n10), .B(
        f0_round_8_p_io_state_out_3_0), .Z(f0_round_8_io_state_out_3_0) );
  NAND2_X1 f0_round_8_c_U18 ( .A1(f0_round_8_p_io_state_out_4_1), .A2(
        f0_round_8_p_io_state_out_0_1), .ZN(f0_round_8_c_n9) );
  XOR2_X1 f0_round_8_c_U17 ( .A(f0_round_8_c_n9), .B(
        f0_round_8_p_io_state_out_3_1), .Z(f0_round_8_io_state_out_3_1) );
  NAND2_X1 f0_round_8_c_U16 ( .A1(f0_round_8_p_io_state_out_4_2), .A2(
        f0_round_8_p_io_state_out_0_2), .ZN(f0_round_8_c_n8) );
  XOR2_X1 f0_round_8_c_U15 ( .A(f0_round_8_c_n8), .B(
        f0_round_8_p_io_state_out_3_2), .Z(f0_round_8_io_state_out_3_2) );
  NAND2_X1 f0_round_8_c_U14 ( .A1(f0_round_8_p_io_state_out_4_3), .A2(
        f0_round_8_p_io_state_out_0_3), .ZN(f0_round_8_c_n7) );
  XOR2_X1 f0_round_8_c_U13 ( .A(f0_round_8_c_n7), .B(
        f0_round_8_p_io_state_out_3_3), .Z(f0_round_8_io_state_out_3_3) );
  NAND2_X1 f0_round_8_c_U12 ( .A1(f0_round_8_p_io_state_out_4_4), .A2(
        f0_round_8_p_io_state_out_0_4), .ZN(f0_round_8_c_n6) );
  XOR2_X1 f0_round_8_c_U11 ( .A(f0_round_8_c_n6), .B(
        f0_round_8_p_io_state_out_3_4), .Z(f0_round_8_io_state_out_3_4) );
  NAND2_X1 f0_round_8_c_U10 ( .A1(f0_round_8_p_io_state_out_1_0), .A2(
        f0_round_8_p_io_state_out_0_0), .ZN(f0_round_8_c_n5) );
  XOR2_X1 f0_round_8_c_U9 ( .A(f0_round_8_c_n5), .B(
        f0_round_8_p_io_state_out_4_0), .Z(f0_round_8_io_state_out_4_0) );
  NAND2_X1 f0_round_8_c_U8 ( .A1(f0_round_8_p_io_state_out_1_1), .A2(
        f0_round_8_p_io_state_out_0_1), .ZN(f0_round_8_c_n4) );
  XOR2_X1 f0_round_8_c_U7 ( .A(f0_round_8_c_n4), .B(
        f0_round_8_p_io_state_out_4_1), .Z(f0_round_8_io_state_out_4_1) );
  NAND2_X1 f0_round_8_c_U6 ( .A1(f0_round_8_p_io_state_out_1_2), .A2(
        f0_round_8_p_io_state_out_0_2), .ZN(f0_round_8_c_n3) );
  XOR2_X1 f0_round_8_c_U5 ( .A(f0_round_8_c_n3), .B(
        f0_round_8_p_io_state_out_4_2), .Z(f0_round_8_io_state_out_4_2) );
  NAND2_X1 f0_round_8_c_U4 ( .A1(f0_round_8_p_io_state_out_1_3), .A2(
        f0_round_8_p_io_state_out_0_3), .ZN(f0_round_8_c_n2) );
  XOR2_X1 f0_round_8_c_U3 ( .A(f0_round_8_c_n2), .B(
        f0_round_8_p_io_state_out_4_3), .Z(f0_round_8_io_state_out_4_3) );
  NAND2_X1 f0_round_8_c_U2 ( .A1(f0_round_8_p_io_state_out_1_4), .A2(
        f0_round_8_p_io_state_out_0_4), .ZN(f0_round_8_c_n1) );
  XOR2_X1 f0_round_8_c_U1 ( .A(f0_round_8_c_n1), .B(
        f0_round_8_p_io_state_out_4_4), .Z(f0_round_8_io_state_out_4_4) );
  XOR2_X1 f0_round_9_t_U50 ( .A(f0_round_8_io_state_out_1_4), .B(
        f0_round_8_io_state_out_1_3), .Z(f0_round_9_t_n25) );
  XNOR2_X1 f0_round_9_t_U49 ( .A(f0_round_8_io_state_out_1_2), .B(
        f0_round_9_t_n25), .ZN(f0_round_9_t_n23) );
  XOR2_X1 f0_round_9_t_U48 ( .A(f0_round_8_io_state_out_1_1), .B(
        f0_round_8_io_state_out_1_0), .Z(f0_round_9_t_n24) );
  XOR2_X1 f0_round_9_t_U47 ( .A(f0_round_9_t_n23), .B(f0_round_9_t_n24), .Z(
        f0_round_9_t_n8) );
  XOR2_X1 f0_round_9_t_U46 ( .A(f0_round_8_io_state_out_4_4), .B(
        f0_round_8_io_state_out_4_3), .Z(f0_round_9_t_n22) );
  XNOR2_X1 f0_round_9_t_U45 ( .A(f0_round_8_io_state_out_4_2), .B(
        f0_round_9_t_n22), .ZN(f0_round_9_t_n20) );
  XOR2_X1 f0_round_9_t_U44 ( .A(f0_round_8_io_state_out_4_1), .B(
        f0_round_8_io_state_out_4_0), .Z(f0_round_9_t_n21) );
  XNOR2_X1 f0_round_9_t_U43 ( .A(f0_round_9_t_n20), .B(f0_round_9_t_n21), .ZN(
        f0_round_9_t_n5) );
  XNOR2_X1 f0_round_9_t_U42 ( .A(f0_round_9_t_n8), .B(f0_round_9_t_n5), .ZN(
        f0_round_9_t_n19) );
  XOR2_X1 f0_round_9_t_U41 ( .A(f0_round_8_io_state_out_0_0), .B(
        f0_round_9_t_n19), .Z(f0_round_9_p_io_state_out_0_0) );
  XOR2_X1 f0_round_9_t_U40 ( .A(f0_round_8_io_state_out_0_1), .B(
        f0_round_9_t_n19), .Z(f0_round_9_p_io_state_out_1_3) );
  XOR2_X1 f0_round_9_t_U39 ( .A(f0_round_8_io_state_out_0_2), .B(
        f0_round_9_t_n19), .Z(f0_round_9_p_io_state_out_2_1) );
  XOR2_X1 f0_round_9_t_U38 ( .A(f0_round_8_io_state_out_0_3), .B(
        f0_round_9_t_n19), .Z(f0_round_9_p_io_state_out_3_4) );
  XOR2_X1 f0_round_9_t_U37 ( .A(f0_round_8_io_state_out_0_4), .B(
        f0_round_9_t_n19), .Z(f0_round_9_p_io_state_out_4_2) );
  XOR2_X1 f0_round_9_t_U36 ( .A(f0_round_8_io_state_out_2_4), .B(
        f0_round_8_io_state_out_2_3), .Z(f0_round_9_t_n18) );
  XNOR2_X1 f0_round_9_t_U35 ( .A(f0_round_8_io_state_out_2_2), .B(
        f0_round_9_t_n18), .ZN(f0_round_9_t_n16) );
  XOR2_X1 f0_round_9_t_U34 ( .A(f0_round_8_io_state_out_2_1), .B(
        f0_round_8_io_state_out_2_0), .Z(f0_round_9_t_n17) );
  XNOR2_X1 f0_round_9_t_U33 ( .A(f0_round_9_t_n16), .B(f0_round_9_t_n17), .ZN(
        f0_round_9_t_n6) );
  XOR2_X1 f0_round_9_t_U32 ( .A(f0_round_8_io_state_out_0_4), .B(
        f0_round_8_io_state_out_0_3), .Z(f0_round_9_t_n15) );
  XNOR2_X1 f0_round_9_t_U31 ( .A(f0_round_8_io_state_out_0_2), .B(
        f0_round_9_t_n15), .ZN(f0_round_9_t_n13) );
  XOR2_X1 f0_round_9_t_U30 ( .A(f0_round_8_io_state_out_0_1), .B(
        f0_round_8_io_state_out_0_0), .Z(f0_round_9_t_n14) );
  XNOR2_X1 f0_round_9_t_U29 ( .A(f0_round_9_t_n13), .B(f0_round_9_t_n14), .ZN(
        f0_round_9_t_n2) );
  XOR2_X1 f0_round_9_t_U28 ( .A(f0_round_9_t_n6), .B(f0_round_9_t_n2), .Z(
        f0_round_9_t_n12) );
  XOR2_X1 f0_round_9_t_U27 ( .A(f0_round_8_io_state_out_1_0), .B(
        f0_round_9_t_n12), .Z(f0_round_9_p_io_state_out_0_2) );
  XOR2_X1 f0_round_9_t_U26 ( .A(f0_round_8_io_state_out_1_1), .B(
        f0_round_9_t_n12), .Z(f0_round_9_p_io_state_out_1_0) );
  XOR2_X1 f0_round_9_t_U25 ( .A(f0_round_8_io_state_out_1_2), .B(
        f0_round_9_t_n12), .Z(f0_round_9_p_io_state_out_2_3) );
  XOR2_X1 f0_round_9_t_U24 ( .A(f0_round_8_io_state_out_1_3), .B(
        f0_round_9_t_n12), .Z(f0_round_9_p_io_state_out_3_1) );
  XOR2_X1 f0_round_9_t_U23 ( .A(f0_round_8_io_state_out_1_4), .B(
        f0_round_9_t_n12), .Z(f0_round_9_p_io_state_out_4_4) );
  XOR2_X1 f0_round_9_t_U22 ( .A(f0_round_8_io_state_out_3_4), .B(
        f0_round_8_io_state_out_3_3), .Z(f0_round_9_t_n11) );
  XNOR2_X1 f0_round_9_t_U21 ( .A(f0_round_8_io_state_out_3_2), .B(
        f0_round_9_t_n11), .ZN(f0_round_9_t_n9) );
  XOR2_X1 f0_round_9_t_U20 ( .A(f0_round_8_io_state_out_3_1), .B(
        f0_round_8_io_state_out_3_0), .Z(f0_round_9_t_n10) );
  XNOR2_X1 f0_round_9_t_U19 ( .A(f0_round_9_t_n9), .B(f0_round_9_t_n10), .ZN(
        f0_round_9_t_n3) );
  XNOR2_X1 f0_round_9_t_U18 ( .A(f0_round_9_t_n8), .B(f0_round_9_t_n3), .ZN(
        f0_round_9_t_n7) );
  XOR2_X1 f0_round_9_t_U17 ( .A(f0_round_8_io_state_out_2_0), .B(
        f0_round_9_t_n7), .Z(f0_round_9_p_io_state_out_0_4) );
  XOR2_X1 f0_round_9_t_U16 ( .A(f0_round_8_io_state_out_2_1), .B(
        f0_round_9_t_n7), .Z(f0_round_9_p_io_state_out_1_2) );
  XOR2_X1 f0_round_9_t_U15 ( .A(f0_round_8_io_state_out_2_2), .B(
        f0_round_9_t_n7), .Z(f0_round_9_p_io_state_out_2_0) );
  XOR2_X1 f0_round_9_t_U14 ( .A(f0_round_8_io_state_out_2_3), .B(
        f0_round_9_t_n7), .Z(f0_round_9_p_io_state_out_3_3) );
  XOR2_X1 f0_round_9_t_U13 ( .A(f0_round_8_io_state_out_2_4), .B(
        f0_round_9_t_n7), .Z(f0_round_9_p_io_state_out_4_1) );
  XOR2_X1 f0_round_9_t_U12 ( .A(f0_round_9_t_n5), .B(f0_round_9_t_n6), .Z(
        f0_round_9_t_n4) );
  XOR2_X1 f0_round_9_t_U11 ( .A(f0_round_8_io_state_out_3_0), .B(
        f0_round_9_t_n4), .Z(f0_round_9_p_io_state_out_0_1) );
  XOR2_X1 f0_round_9_t_U10 ( .A(f0_round_8_io_state_out_3_1), .B(
        f0_round_9_t_n4), .Z(f0_round_9_p_io_state_out_1_4) );
  XOR2_X1 f0_round_9_t_U9 ( .A(f0_round_8_io_state_out_3_2), .B(
        f0_round_9_t_n4), .Z(f0_round_9_p_io_state_out_2_2) );
  XOR2_X1 f0_round_9_t_U8 ( .A(f0_round_8_io_state_out_3_3), .B(
        f0_round_9_t_n4), .Z(f0_round_9_p_io_state_out_3_0) );
  XOR2_X1 f0_round_9_t_U7 ( .A(f0_round_8_io_state_out_3_4), .B(
        f0_round_9_t_n4), .Z(f0_round_9_p_io_state_out_4_3) );
  XOR2_X1 f0_round_9_t_U6 ( .A(f0_round_9_t_n2), .B(f0_round_9_t_n3), .Z(
        f0_round_9_t_n1) );
  XOR2_X1 f0_round_9_t_U5 ( .A(f0_round_8_io_state_out_4_0), .B(
        f0_round_9_t_n1), .Z(f0_round_9_p_io_state_out_0_3) );
  XOR2_X1 f0_round_9_t_U4 ( .A(f0_round_8_io_state_out_4_1), .B(
        f0_round_9_t_n1), .Z(f0_round_9_p_io_state_out_1_1) );
  XOR2_X1 f0_round_9_t_U3 ( .A(f0_round_8_io_state_out_4_2), .B(
        f0_round_9_t_n1), .Z(f0_round_9_p_io_state_out_2_4) );
  XOR2_X1 f0_round_9_t_U2 ( .A(f0_round_8_io_state_out_4_3), .B(
        f0_round_9_t_n1), .Z(f0_round_9_p_io_state_out_3_2) );
  XOR2_X1 f0_round_9_t_U1 ( .A(f0_round_8_io_state_out_4_4), .B(
        f0_round_9_t_n1), .Z(f0_round_9_p_io_state_out_4_0) );
  NAND2_X1 f0_round_9_c_U50 ( .A1(f0_round_9_p_io_state_out_2_0), .A2(
        f0_round_9_p_io_state_out_1_0), .ZN(f0_round_9_c_n25) );
  XOR2_X1 f0_round_9_c_U49 ( .A(f0_round_9_c_n25), .B(
        f0_round_9_p_io_state_out_0_0), .Z(f0_round_9_c_io_state_out_0_0) );
  NAND2_X1 f0_round_9_c_U48 ( .A1(f0_round_9_p_io_state_out_2_1), .A2(
        f0_round_9_p_io_state_out_1_1), .ZN(f0_round_9_c_n24) );
  XOR2_X1 f0_round_9_c_U47 ( .A(f0_round_9_c_n24), .B(
        f0_round_9_p_io_state_out_0_1), .Z(f0_round_9_io_state_out_0_1) );
  NAND2_X1 f0_round_9_c_U46 ( .A1(f0_round_9_p_io_state_out_2_2), .A2(
        f0_round_9_p_io_state_out_1_2), .ZN(f0_round_9_c_n23) );
  XOR2_X1 f0_round_9_c_U45 ( .A(f0_round_9_c_n23), .B(
        f0_round_9_p_io_state_out_0_2), .Z(f0_round_9_io_state_out_0_2) );
  NAND2_X1 f0_round_9_c_U44 ( .A1(f0_round_9_p_io_state_out_2_3), .A2(
        f0_round_9_p_io_state_out_1_3), .ZN(f0_round_9_c_n22) );
  XOR2_X1 f0_round_9_c_U43 ( .A(f0_round_9_c_n22), .B(
        f0_round_9_p_io_state_out_0_3), .Z(f0_round_9_io_state_out_0_3) );
  NAND2_X1 f0_round_9_c_U42 ( .A1(f0_round_9_p_io_state_out_2_4), .A2(
        f0_round_9_p_io_state_out_1_4), .ZN(f0_round_9_c_n21) );
  XOR2_X1 f0_round_9_c_U41 ( .A(f0_round_9_c_n21), .B(
        f0_round_9_p_io_state_out_0_4), .Z(f0_round_9_io_state_out_0_4) );
  NAND2_X1 f0_round_9_c_U40 ( .A1(f0_round_9_p_io_state_out_2_0), .A2(
        f0_round_9_p_io_state_out_3_0), .ZN(f0_round_9_c_n20) );
  XOR2_X1 f0_round_9_c_U39 ( .A(f0_round_9_c_n20), .B(
        f0_round_9_p_io_state_out_1_0), .Z(f0_round_9_io_state_out_1_0) );
  NAND2_X1 f0_round_9_c_U38 ( .A1(f0_round_9_p_io_state_out_2_1), .A2(
        f0_round_9_p_io_state_out_3_1), .ZN(f0_round_9_c_n19) );
  XOR2_X1 f0_round_9_c_U37 ( .A(f0_round_9_c_n19), .B(
        f0_round_9_p_io_state_out_1_1), .Z(f0_round_9_io_state_out_1_1) );
  NAND2_X1 f0_round_9_c_U36 ( .A1(f0_round_9_p_io_state_out_2_2), .A2(
        f0_round_9_p_io_state_out_3_2), .ZN(f0_round_9_c_n18) );
  XOR2_X1 f0_round_9_c_U35 ( .A(f0_round_9_c_n18), .B(
        f0_round_9_p_io_state_out_1_2), .Z(f0_round_9_io_state_out_1_2) );
  NAND2_X1 f0_round_9_c_U34 ( .A1(f0_round_9_p_io_state_out_2_3), .A2(
        f0_round_9_p_io_state_out_3_3), .ZN(f0_round_9_c_n17) );
  XOR2_X1 f0_round_9_c_U33 ( .A(f0_round_9_c_n17), .B(
        f0_round_9_p_io_state_out_1_3), .Z(f0_round_9_io_state_out_1_3) );
  NAND2_X1 f0_round_9_c_U32 ( .A1(f0_round_9_p_io_state_out_2_4), .A2(
        f0_round_9_p_io_state_out_3_4), .ZN(f0_round_9_c_n16) );
  XOR2_X1 f0_round_9_c_U31 ( .A(f0_round_9_c_n16), .B(
        f0_round_9_p_io_state_out_1_4), .Z(f0_round_9_io_state_out_1_4) );
  NAND2_X1 f0_round_9_c_U30 ( .A1(f0_round_9_p_io_state_out_3_0), .A2(
        f0_round_9_p_io_state_out_4_0), .ZN(f0_round_9_c_n15) );
  XOR2_X1 f0_round_9_c_U29 ( .A(f0_round_9_c_n15), .B(
        f0_round_9_p_io_state_out_2_0), .Z(f0_round_9_io_state_out_2_0) );
  NAND2_X1 f0_round_9_c_U28 ( .A1(f0_round_9_p_io_state_out_3_1), .A2(
        f0_round_9_p_io_state_out_4_1), .ZN(f0_round_9_c_n14) );
  XOR2_X1 f0_round_9_c_U27 ( .A(f0_round_9_c_n14), .B(
        f0_round_9_p_io_state_out_2_1), .Z(f0_round_9_io_state_out_2_1) );
  NAND2_X1 f0_round_9_c_U26 ( .A1(f0_round_9_p_io_state_out_3_2), .A2(
        f0_round_9_p_io_state_out_4_2), .ZN(f0_round_9_c_n13) );
  XOR2_X1 f0_round_9_c_U25 ( .A(f0_round_9_c_n13), .B(
        f0_round_9_p_io_state_out_2_2), .Z(f0_round_9_io_state_out_2_2) );
  NAND2_X1 f0_round_9_c_U24 ( .A1(f0_round_9_p_io_state_out_3_3), .A2(
        f0_round_9_p_io_state_out_4_3), .ZN(f0_round_9_c_n12) );
  XOR2_X1 f0_round_9_c_U23 ( .A(f0_round_9_c_n12), .B(
        f0_round_9_p_io_state_out_2_3), .Z(f0_round_9_io_state_out_2_3) );
  NAND2_X1 f0_round_9_c_U22 ( .A1(f0_round_9_p_io_state_out_3_4), .A2(
        f0_round_9_p_io_state_out_4_4), .ZN(f0_round_9_c_n11) );
  XOR2_X1 f0_round_9_c_U21 ( .A(f0_round_9_c_n11), .B(
        f0_round_9_p_io_state_out_2_4), .Z(f0_round_9_io_state_out_2_4) );
  NAND2_X1 f0_round_9_c_U20 ( .A1(f0_round_9_p_io_state_out_4_0), .A2(
        f0_round_9_p_io_state_out_0_0), .ZN(f0_round_9_c_n10) );
  XOR2_X1 f0_round_9_c_U19 ( .A(f0_round_9_c_n10), .B(
        f0_round_9_p_io_state_out_3_0), .Z(f0_round_9_io_state_out_3_0) );
  NAND2_X1 f0_round_9_c_U18 ( .A1(f0_round_9_p_io_state_out_4_1), .A2(
        f0_round_9_p_io_state_out_0_1), .ZN(f0_round_9_c_n9) );
  XOR2_X1 f0_round_9_c_U17 ( .A(f0_round_9_c_n9), .B(
        f0_round_9_p_io_state_out_3_1), .Z(f0_round_9_io_state_out_3_1) );
  NAND2_X1 f0_round_9_c_U16 ( .A1(f0_round_9_p_io_state_out_4_2), .A2(
        f0_round_9_p_io_state_out_0_2), .ZN(f0_round_9_c_n8) );
  XOR2_X1 f0_round_9_c_U15 ( .A(f0_round_9_c_n8), .B(
        f0_round_9_p_io_state_out_3_2), .Z(f0_round_9_io_state_out_3_2) );
  NAND2_X1 f0_round_9_c_U14 ( .A1(f0_round_9_p_io_state_out_4_3), .A2(
        f0_round_9_p_io_state_out_0_3), .ZN(f0_round_9_c_n7) );
  XOR2_X1 f0_round_9_c_U13 ( .A(f0_round_9_c_n7), .B(
        f0_round_9_p_io_state_out_3_3), .Z(f0_round_9_io_state_out_3_3) );
  NAND2_X1 f0_round_9_c_U12 ( .A1(f0_round_9_p_io_state_out_4_4), .A2(
        f0_round_9_p_io_state_out_0_4), .ZN(f0_round_9_c_n6) );
  XOR2_X1 f0_round_9_c_U11 ( .A(f0_round_9_c_n6), .B(
        f0_round_9_p_io_state_out_3_4), .Z(f0_round_9_io_state_out_3_4) );
  NAND2_X1 f0_round_9_c_U10 ( .A1(f0_round_9_p_io_state_out_1_0), .A2(
        f0_round_9_p_io_state_out_0_0), .ZN(f0_round_9_c_n5) );
  XOR2_X1 f0_round_9_c_U9 ( .A(f0_round_9_c_n5), .B(
        f0_round_9_p_io_state_out_4_0), .Z(f0_round_9_io_state_out_4_0) );
  NAND2_X1 f0_round_9_c_U8 ( .A1(f0_round_9_p_io_state_out_1_1), .A2(
        f0_round_9_p_io_state_out_0_1), .ZN(f0_round_9_c_n4) );
  XOR2_X1 f0_round_9_c_U7 ( .A(f0_round_9_c_n4), .B(
        f0_round_9_p_io_state_out_4_1), .Z(f0_round_9_io_state_out_4_1) );
  NAND2_X1 f0_round_9_c_U6 ( .A1(f0_round_9_p_io_state_out_1_2), .A2(
        f0_round_9_p_io_state_out_0_2), .ZN(f0_round_9_c_n3) );
  XOR2_X1 f0_round_9_c_U5 ( .A(f0_round_9_c_n3), .B(
        f0_round_9_p_io_state_out_4_2), .Z(f0_round_9_io_state_out_4_2) );
  NAND2_X1 f0_round_9_c_U4 ( .A1(f0_round_9_p_io_state_out_1_3), .A2(
        f0_round_9_p_io_state_out_0_3), .ZN(f0_round_9_c_n2) );
  XOR2_X1 f0_round_9_c_U3 ( .A(f0_round_9_c_n2), .B(
        f0_round_9_p_io_state_out_4_3), .Z(f0_round_9_io_state_out_4_3) );
  NAND2_X1 f0_round_9_c_U2 ( .A1(f0_round_9_p_io_state_out_1_4), .A2(
        f0_round_9_p_io_state_out_0_4), .ZN(f0_round_9_c_n1) );
  XOR2_X1 f0_round_9_c_U1 ( .A(f0_round_9_c_n1), .B(
        f0_round_9_p_io_state_out_4_4), .Z(f0_round_9_io_state_out_4_4) );
  INV_X1 f0_round_9_i_U1 ( .A(f0_round_9_c_io_state_out_0_0), .ZN(
        f0_round_9_io_state_out_0_0) );
  XOR2_X1 f0_round_10_t_U50 ( .A(f0_round_9_io_state_out_1_4), .B(
        f0_round_9_io_state_out_1_3), .Z(f0_round_10_t_n25) );
  XNOR2_X1 f0_round_10_t_U49 ( .A(f0_round_9_io_state_out_1_2), .B(
        f0_round_10_t_n25), .ZN(f0_round_10_t_n23) );
  XOR2_X1 f0_round_10_t_U48 ( .A(f0_round_9_io_state_out_1_1), .B(
        f0_round_9_io_state_out_1_0), .Z(f0_round_10_t_n24) );
  XOR2_X1 f0_round_10_t_U47 ( .A(f0_round_10_t_n23), .B(f0_round_10_t_n24), 
        .Z(f0_round_10_t_n8) );
  XOR2_X1 f0_round_10_t_U46 ( .A(f0_round_9_io_state_out_4_4), .B(
        f0_round_9_io_state_out_4_3), .Z(f0_round_10_t_n22) );
  XNOR2_X1 f0_round_10_t_U45 ( .A(f0_round_9_io_state_out_4_2), .B(
        f0_round_10_t_n22), .ZN(f0_round_10_t_n20) );
  XOR2_X1 f0_round_10_t_U44 ( .A(f0_round_9_io_state_out_4_1), .B(
        f0_round_9_io_state_out_4_0), .Z(f0_round_10_t_n21) );
  XNOR2_X1 f0_round_10_t_U43 ( .A(f0_round_10_t_n20), .B(f0_round_10_t_n21), 
        .ZN(f0_round_10_t_n5) );
  XNOR2_X1 f0_round_10_t_U42 ( .A(f0_round_10_t_n8), .B(f0_round_10_t_n5), 
        .ZN(f0_round_10_t_n19) );
  XOR2_X1 f0_round_10_t_U41 ( .A(f0_round_9_io_state_out_0_0), .B(
        f0_round_10_t_n19), .Z(f0_round_10_p_io_state_out_0_0) );
  XOR2_X1 f0_round_10_t_U40 ( .A(f0_round_9_io_state_out_0_1), .B(
        f0_round_10_t_n19), .Z(f0_round_10_p_io_state_out_1_3) );
  XOR2_X1 f0_round_10_t_U39 ( .A(f0_round_9_io_state_out_0_2), .B(
        f0_round_10_t_n19), .Z(f0_round_10_p_io_state_out_2_1) );
  XOR2_X1 f0_round_10_t_U38 ( .A(f0_round_9_io_state_out_0_3), .B(
        f0_round_10_t_n19), .Z(f0_round_10_p_io_state_out_3_4) );
  XOR2_X1 f0_round_10_t_U37 ( .A(f0_round_9_io_state_out_0_4), .B(
        f0_round_10_t_n19), .Z(f0_round_10_p_io_state_out_4_2) );
  XOR2_X1 f0_round_10_t_U36 ( .A(f0_round_9_io_state_out_2_4), .B(
        f0_round_9_io_state_out_2_3), .Z(f0_round_10_t_n18) );
  XNOR2_X1 f0_round_10_t_U35 ( .A(f0_round_9_io_state_out_2_2), .B(
        f0_round_10_t_n18), .ZN(f0_round_10_t_n16) );
  XOR2_X1 f0_round_10_t_U34 ( .A(f0_round_9_io_state_out_2_1), .B(
        f0_round_9_io_state_out_2_0), .Z(f0_round_10_t_n17) );
  XNOR2_X1 f0_round_10_t_U33 ( .A(f0_round_10_t_n16), .B(f0_round_10_t_n17), 
        .ZN(f0_round_10_t_n6) );
  XOR2_X1 f0_round_10_t_U32 ( .A(f0_round_9_io_state_out_0_4), .B(
        f0_round_9_io_state_out_0_3), .Z(f0_round_10_t_n15) );
  XNOR2_X1 f0_round_10_t_U31 ( .A(f0_round_9_io_state_out_0_2), .B(
        f0_round_10_t_n15), .ZN(f0_round_10_t_n13) );
  XOR2_X1 f0_round_10_t_U30 ( .A(f0_round_9_io_state_out_0_1), .B(
        f0_round_9_io_state_out_0_0), .Z(f0_round_10_t_n14) );
  XNOR2_X1 f0_round_10_t_U29 ( .A(f0_round_10_t_n13), .B(f0_round_10_t_n14), 
        .ZN(f0_round_10_t_n2) );
  XOR2_X1 f0_round_10_t_U28 ( .A(f0_round_10_t_n6), .B(f0_round_10_t_n2), .Z(
        f0_round_10_t_n12) );
  XOR2_X1 f0_round_10_t_U27 ( .A(f0_round_9_io_state_out_1_0), .B(
        f0_round_10_t_n12), .Z(f0_round_10_p_io_state_out_0_2) );
  XOR2_X1 f0_round_10_t_U26 ( .A(f0_round_9_io_state_out_1_1), .B(
        f0_round_10_t_n12), .Z(f0_round_10_p_io_state_out_1_0) );
  XOR2_X1 f0_round_10_t_U25 ( .A(f0_round_9_io_state_out_1_2), .B(
        f0_round_10_t_n12), .Z(f0_round_10_p_io_state_out_2_3) );
  XOR2_X1 f0_round_10_t_U24 ( .A(f0_round_9_io_state_out_1_3), .B(
        f0_round_10_t_n12), .Z(f0_round_10_p_io_state_out_3_1) );
  XOR2_X1 f0_round_10_t_U23 ( .A(f0_round_9_io_state_out_1_4), .B(
        f0_round_10_t_n12), .Z(f0_round_10_p_io_state_out_4_4) );
  XOR2_X1 f0_round_10_t_U22 ( .A(f0_round_9_io_state_out_3_4), .B(
        f0_round_9_io_state_out_3_3), .Z(f0_round_10_t_n11) );
  XNOR2_X1 f0_round_10_t_U21 ( .A(f0_round_9_io_state_out_3_2), .B(
        f0_round_10_t_n11), .ZN(f0_round_10_t_n9) );
  XOR2_X1 f0_round_10_t_U20 ( .A(f0_round_9_io_state_out_3_1), .B(
        f0_round_9_io_state_out_3_0), .Z(f0_round_10_t_n10) );
  XNOR2_X1 f0_round_10_t_U19 ( .A(f0_round_10_t_n9), .B(f0_round_10_t_n10), 
        .ZN(f0_round_10_t_n3) );
  XNOR2_X1 f0_round_10_t_U18 ( .A(f0_round_10_t_n8), .B(f0_round_10_t_n3), 
        .ZN(f0_round_10_t_n7) );
  XOR2_X1 f0_round_10_t_U17 ( .A(f0_round_9_io_state_out_2_0), .B(
        f0_round_10_t_n7), .Z(f0_round_10_p_io_state_out_0_4) );
  XOR2_X1 f0_round_10_t_U16 ( .A(f0_round_9_io_state_out_2_1), .B(
        f0_round_10_t_n7), .Z(f0_round_10_p_io_state_out_1_2) );
  XOR2_X1 f0_round_10_t_U15 ( .A(f0_round_9_io_state_out_2_2), .B(
        f0_round_10_t_n7), .Z(f0_round_10_p_io_state_out_2_0) );
  XOR2_X1 f0_round_10_t_U14 ( .A(f0_round_9_io_state_out_2_3), .B(
        f0_round_10_t_n7), .Z(f0_round_10_p_io_state_out_3_3) );
  XOR2_X1 f0_round_10_t_U13 ( .A(f0_round_9_io_state_out_2_4), .B(
        f0_round_10_t_n7), .Z(f0_round_10_p_io_state_out_4_1) );
  XOR2_X1 f0_round_10_t_U12 ( .A(f0_round_10_t_n5), .B(f0_round_10_t_n6), .Z(
        f0_round_10_t_n4) );
  XOR2_X1 f0_round_10_t_U11 ( .A(f0_round_9_io_state_out_3_0), .B(
        f0_round_10_t_n4), .Z(f0_round_10_p_io_state_out_0_1) );
  XOR2_X1 f0_round_10_t_U10 ( .A(f0_round_9_io_state_out_3_1), .B(
        f0_round_10_t_n4), .Z(f0_round_10_p_io_state_out_1_4) );
  XOR2_X1 f0_round_10_t_U9 ( .A(f0_round_9_io_state_out_3_2), .B(
        f0_round_10_t_n4), .Z(f0_round_10_p_io_state_out_2_2) );
  XOR2_X1 f0_round_10_t_U8 ( .A(f0_round_9_io_state_out_3_3), .B(
        f0_round_10_t_n4), .Z(f0_round_10_p_io_state_out_3_0) );
  XOR2_X1 f0_round_10_t_U7 ( .A(f0_round_9_io_state_out_3_4), .B(
        f0_round_10_t_n4), .Z(f0_round_10_p_io_state_out_4_3) );
  XOR2_X1 f0_round_10_t_U6 ( .A(f0_round_10_t_n2), .B(f0_round_10_t_n3), .Z(
        f0_round_10_t_n1) );
  XOR2_X1 f0_round_10_t_U5 ( .A(f0_round_9_io_state_out_4_0), .B(
        f0_round_10_t_n1), .Z(f0_round_10_p_io_state_out_0_3) );
  XOR2_X1 f0_round_10_t_U4 ( .A(f0_round_9_io_state_out_4_1), .B(
        f0_round_10_t_n1), .Z(f0_round_10_p_io_state_out_1_1) );
  XOR2_X1 f0_round_10_t_U3 ( .A(f0_round_9_io_state_out_4_2), .B(
        f0_round_10_t_n1), .Z(f0_round_10_p_io_state_out_2_4) );
  XOR2_X1 f0_round_10_t_U2 ( .A(f0_round_9_io_state_out_4_3), .B(
        f0_round_10_t_n1), .Z(f0_round_10_p_io_state_out_3_2) );
  XOR2_X1 f0_round_10_t_U1 ( .A(f0_round_9_io_state_out_4_4), .B(
        f0_round_10_t_n1), .Z(f0_round_10_p_io_state_out_4_0) );
  NAND2_X1 f0_round_10_c_U50 ( .A1(f0_round_10_p_io_state_out_2_0), .A2(
        f0_round_10_p_io_state_out_1_0), .ZN(f0_round_10_c_n25) );
  XOR2_X1 f0_round_10_c_U49 ( .A(f0_round_10_c_n25), .B(
        f0_round_10_p_io_state_out_0_0), .Z(f0_io_state_out_0_0) );
  NAND2_X1 f0_round_10_c_U48 ( .A1(f0_round_10_p_io_state_out_2_1), .A2(
        f0_round_10_p_io_state_out_1_1), .ZN(f0_round_10_c_n24) );
  XOR2_X1 f0_round_10_c_U47 ( .A(f0_round_10_c_n24), .B(
        f0_round_10_p_io_state_out_0_1), .Z(f0_io_state_out_0_1) );
  NAND2_X1 f0_round_10_c_U46 ( .A1(f0_round_10_p_io_state_out_2_2), .A2(
        f0_round_10_p_io_state_out_1_2), .ZN(f0_round_10_c_n23) );
  XOR2_X1 f0_round_10_c_U45 ( .A(f0_round_10_c_n23), .B(
        f0_round_10_p_io_state_out_0_2), .Z(abs1_io_state_out_0_2) );
  NAND2_X1 f0_round_10_c_U44 ( .A1(f0_round_10_p_io_state_out_2_3), .A2(
        f0_round_10_p_io_state_out_1_3), .ZN(f0_round_10_c_n22) );
  XOR2_X1 f0_round_10_c_U43 ( .A(f0_round_10_c_n22), .B(
        f0_round_10_p_io_state_out_0_3), .Z(abs1_io_state_out_0_3) );
  NAND2_X1 f0_round_10_c_U42 ( .A1(f0_round_10_p_io_state_out_2_4), .A2(
        f0_round_10_p_io_state_out_1_4), .ZN(f0_round_10_c_n21) );
  XOR2_X1 f0_round_10_c_U41 ( .A(f0_round_10_c_n21), .B(
        f0_round_10_p_io_state_out_0_4), .Z(abs1_io_state_out_0_4) );
  NAND2_X1 f0_round_10_c_U40 ( .A1(f0_round_10_p_io_state_out_2_0), .A2(
        f0_round_10_p_io_state_out_3_0), .ZN(f0_round_10_c_n20) );
  XOR2_X1 f0_round_10_c_U39 ( .A(f0_round_10_c_n20), .B(
        f0_round_10_p_io_state_out_1_0), .Z(f0_io_state_out_1_0) );
  NAND2_X1 f0_round_10_c_U38 ( .A1(f0_round_10_p_io_state_out_2_1), .A2(
        f0_round_10_p_io_state_out_3_1), .ZN(f0_round_10_c_n19) );
  XOR2_X1 f0_round_10_c_U37 ( .A(f0_round_10_c_n19), .B(
        f0_round_10_p_io_state_out_1_1), .Z(f0_io_state_out_1_1) );
  NAND2_X1 f0_round_10_c_U36 ( .A1(f0_round_10_p_io_state_out_2_2), .A2(
        f0_round_10_p_io_state_out_3_2), .ZN(f0_round_10_c_n18) );
  XOR2_X1 f0_round_10_c_U35 ( .A(f0_round_10_c_n18), .B(
        f0_round_10_p_io_state_out_1_2), .Z(abs1_io_state_out_1_2) );
  NAND2_X1 f0_round_10_c_U34 ( .A1(f0_round_10_p_io_state_out_2_3), .A2(
        f0_round_10_p_io_state_out_3_3), .ZN(f0_round_10_c_n17) );
  XOR2_X1 f0_round_10_c_U33 ( .A(f0_round_10_c_n17), .B(
        f0_round_10_p_io_state_out_1_3), .Z(abs1_io_state_out_1_3) );
  NAND2_X1 f0_round_10_c_U32 ( .A1(f0_round_10_p_io_state_out_2_4), .A2(
        f0_round_10_p_io_state_out_3_4), .ZN(f0_round_10_c_n16) );
  XOR2_X1 f0_round_10_c_U31 ( .A(f0_round_10_c_n16), .B(
        f0_round_10_p_io_state_out_1_4), .Z(abs1_io_state_out_1_4) );
  NAND2_X1 f0_round_10_c_U30 ( .A1(f0_round_10_p_io_state_out_3_0), .A2(
        f0_round_10_p_io_state_out_4_0), .ZN(f0_round_10_c_n15) );
  XOR2_X1 f0_round_10_c_U29 ( .A(f0_round_10_c_n15), .B(
        f0_round_10_p_io_state_out_2_0), .Z(f0_io_state_out_2_0) );
  NAND2_X1 f0_round_10_c_U28 ( .A1(f0_round_10_p_io_state_out_3_1), .A2(
        f0_round_10_p_io_state_out_4_1), .ZN(f0_round_10_c_n14) );
  XOR2_X1 f0_round_10_c_U27 ( .A(f0_round_10_c_n14), .B(
        f0_round_10_p_io_state_out_2_1), .Z(f0_io_state_out_2_1) );
  NAND2_X1 f0_round_10_c_U26 ( .A1(f0_round_10_p_io_state_out_3_2), .A2(
        f0_round_10_p_io_state_out_4_2), .ZN(f0_round_10_c_n13) );
  XOR2_X1 f0_round_10_c_U25 ( .A(f0_round_10_c_n13), .B(
        f0_round_10_p_io_state_out_2_2), .Z(abs1_io_state_out_2_2) );
  NAND2_X1 f0_round_10_c_U24 ( .A1(f0_round_10_p_io_state_out_3_3), .A2(
        f0_round_10_p_io_state_out_4_3), .ZN(f0_round_10_c_n12) );
  XOR2_X1 f0_round_10_c_U23 ( .A(f0_round_10_c_n12), .B(
        f0_round_10_p_io_state_out_2_3), .Z(abs1_io_state_out_2_3) );
  NAND2_X1 f0_round_10_c_U22 ( .A1(f0_round_10_p_io_state_out_3_4), .A2(
        f0_round_10_p_io_state_out_4_4), .ZN(f0_round_10_c_n11) );
  XOR2_X1 f0_round_10_c_U21 ( .A(f0_round_10_c_n11), .B(
        f0_round_10_p_io_state_out_2_4), .Z(abs1_io_state_out_2_4) );
  NAND2_X1 f0_round_10_c_U20 ( .A1(f0_round_10_p_io_state_out_4_0), .A2(
        f0_round_10_p_io_state_out_0_0), .ZN(f0_round_10_c_n10) );
  XOR2_X1 f0_round_10_c_U19 ( .A(f0_round_10_c_n10), .B(
        f0_round_10_p_io_state_out_3_0), .Z(f0_io_state_out_3_0) );
  NAND2_X1 f0_round_10_c_U18 ( .A1(f0_round_10_p_io_state_out_4_1), .A2(
        f0_round_10_p_io_state_out_0_1), .ZN(f0_round_10_c_n9) );
  XOR2_X1 f0_round_10_c_U17 ( .A(f0_round_10_c_n9), .B(
        f0_round_10_p_io_state_out_3_1), .Z(f0_io_state_out_3_1) );
  NAND2_X1 f0_round_10_c_U16 ( .A1(f0_round_10_p_io_state_out_4_2), .A2(
        f0_round_10_p_io_state_out_0_2), .ZN(f0_round_10_c_n8) );
  XOR2_X1 f0_round_10_c_U15 ( .A(f0_round_10_c_n8), .B(
        f0_round_10_p_io_state_out_3_2), .Z(abs1_io_state_out_3_2) );
  NAND2_X1 f0_round_10_c_U14 ( .A1(f0_round_10_p_io_state_out_4_3), .A2(
        f0_round_10_p_io_state_out_0_3), .ZN(f0_round_10_c_n7) );
  XOR2_X1 f0_round_10_c_U13 ( .A(f0_round_10_c_n7), .B(
        f0_round_10_p_io_state_out_3_3), .Z(abs1_io_state_out_3_3) );
  NAND2_X1 f0_round_10_c_U12 ( .A1(f0_round_10_p_io_state_out_4_4), .A2(
        f0_round_10_p_io_state_out_0_4), .ZN(f0_round_10_c_n6) );
  XOR2_X1 f0_round_10_c_U11 ( .A(f0_round_10_c_n6), .B(
        f0_round_10_p_io_state_out_3_4), .Z(abs1_io_state_out_3_4) );
  NAND2_X1 f0_round_10_c_U10 ( .A1(f0_round_10_p_io_state_out_1_0), .A2(
        f0_round_10_p_io_state_out_0_0), .ZN(f0_round_10_c_n5) );
  XOR2_X1 f0_round_10_c_U9 ( .A(f0_round_10_c_n5), .B(
        f0_round_10_p_io_state_out_4_0), .Z(f0_io_state_out_4_0) );
  NAND2_X1 f0_round_10_c_U8 ( .A1(f0_round_10_p_io_state_out_1_1), .A2(
        f0_round_10_p_io_state_out_0_1), .ZN(f0_round_10_c_n4) );
  XOR2_X1 f0_round_10_c_U7 ( .A(f0_round_10_c_n4), .B(
        f0_round_10_p_io_state_out_4_1), .Z(f0_io_state_out_4_1) );
  NAND2_X1 f0_round_10_c_U6 ( .A1(f0_round_10_p_io_state_out_1_2), .A2(
        f0_round_10_p_io_state_out_0_2), .ZN(f0_round_10_c_n3) );
  XOR2_X1 f0_round_10_c_U5 ( .A(f0_round_10_c_n3), .B(
        f0_round_10_p_io_state_out_4_2), .Z(abs1_io_state_out_4_2) );
  NAND2_X1 f0_round_10_c_U4 ( .A1(f0_round_10_p_io_state_out_1_3), .A2(
        f0_round_10_p_io_state_out_0_3), .ZN(f0_round_10_c_n2) );
  XOR2_X1 f0_round_10_c_U3 ( .A(f0_round_10_c_n2), .B(
        f0_round_10_p_io_state_out_4_3), .Z(abs1_io_state_out_4_3) );
  NAND2_X1 f0_round_10_c_U2 ( .A1(f0_round_10_p_io_state_out_1_4), .A2(
        f0_round_10_p_io_state_out_0_4), .ZN(f0_round_10_c_n1) );
  XOR2_X1 f0_round_10_c_U1 ( .A(f0_round_10_c_n1), .B(
        f0_round_10_p_io_state_out_4_4), .Z(abs1_io_state_out_4_4) );
  XOR2_X1 abs1_U10 ( .A(f0_io_state_out_0_0), .B(io_block_i1[0]), .Z(
        abs1_io_state_out_0_0) );
  XOR2_X1 abs1_U9 ( .A(f0_io_state_out_0_1), .B(io_block_i1[5]), .Z(
        abs1_io_state_out_0_1) );
  XOR2_X1 abs1_U8 ( .A(f0_io_state_out_1_0), .B(io_block_i1[1]), .Z(
        abs1_io_state_out_1_0) );
  XOR2_X1 abs1_U7 ( .A(f0_io_state_out_1_1), .B(io_block_i1[6]), .Z(
        abs1_io_state_out_1_1) );
  XOR2_X1 abs1_U6 ( .A(f0_io_state_out_2_0), .B(io_block_i1[2]), .Z(
        abs1_io_state_out_2_0) );
  XOR2_X1 abs1_U5 ( .A(f0_io_state_out_2_1), .B(io_block_i1[7]), .Z(
        abs1_io_state_out_2_1) );
  XOR2_X1 abs1_U4 ( .A(f0_io_state_out_3_0), .B(io_block_i1[3]), .Z(
        abs1_io_state_out_3_0) );
  XOR2_X1 abs1_U3 ( .A(f0_io_state_out_3_1), .B(io_block_i1[8]), .Z(
        abs1_io_state_out_3_1) );
  XOR2_X1 abs1_U2 ( .A(f0_io_state_out_4_0), .B(io_block_i1[4]), .Z(
        abs1_io_state_out_4_0) );
  XOR2_X1 abs1_U1 ( .A(f0_io_state_out_4_1), .B(io_block_i1[9]), .Z(
        abs1_io_state_out_4_1) );
  XOR2_X1 f1_round_t_U50 ( .A(abs1_io_state_out_1_4), .B(abs1_io_state_out_1_3), .Z(f1_round_t_n25) );
  XNOR2_X1 f1_round_t_U49 ( .A(abs1_io_state_out_1_2), .B(f1_round_t_n25), 
        .ZN(f1_round_t_n23) );
  XOR2_X1 f1_round_t_U48 ( .A(abs1_io_state_out_1_1), .B(abs1_io_state_out_1_0), .Z(f1_round_t_n24) );
  XOR2_X1 f1_round_t_U47 ( .A(f1_round_t_n23), .B(f1_round_t_n24), .Z(
        f1_round_t_n8) );
  XOR2_X1 f1_round_t_U46 ( .A(abs1_io_state_out_4_4), .B(abs1_io_state_out_4_3), .Z(f1_round_t_n22) );
  XNOR2_X1 f1_round_t_U45 ( .A(abs1_io_state_out_4_2), .B(f1_round_t_n22), 
        .ZN(f1_round_t_n20) );
  XOR2_X1 f1_round_t_U44 ( .A(abs1_io_state_out_4_1), .B(abs1_io_state_out_4_0), .Z(f1_round_t_n21) );
  XNOR2_X1 f1_round_t_U43 ( .A(f1_round_t_n20), .B(f1_round_t_n21), .ZN(
        f1_round_t_n5) );
  XNOR2_X1 f1_round_t_U42 ( .A(f1_round_t_n8), .B(f1_round_t_n5), .ZN(
        f1_round_t_n19) );
  XOR2_X1 f1_round_t_U41 ( .A(abs1_io_state_out_0_0), .B(f1_round_t_n19), .Z(
        f1_round_p_io_state_out_0_0) );
  XOR2_X1 f1_round_t_U40 ( .A(abs1_io_state_out_0_1), .B(f1_round_t_n19), .Z(
        f1_round_p_io_state_out_1_3) );
  XOR2_X1 f1_round_t_U39 ( .A(abs1_io_state_out_0_2), .B(f1_round_t_n19), .Z(
        f1_round_p_io_state_out_2_1) );
  XOR2_X1 f1_round_t_U38 ( .A(abs1_io_state_out_0_3), .B(f1_round_t_n19), .Z(
        f1_round_p_io_state_out_3_4) );
  XOR2_X1 f1_round_t_U37 ( .A(abs1_io_state_out_0_4), .B(f1_round_t_n19), .Z(
        f1_round_p_io_state_out_4_2) );
  XOR2_X1 f1_round_t_U36 ( .A(abs1_io_state_out_2_4), .B(abs1_io_state_out_2_3), .Z(f1_round_t_n18) );
  XNOR2_X1 f1_round_t_U35 ( .A(abs1_io_state_out_2_2), .B(f1_round_t_n18), 
        .ZN(f1_round_t_n16) );
  XOR2_X1 f1_round_t_U34 ( .A(abs1_io_state_out_2_1), .B(abs1_io_state_out_2_0), .Z(f1_round_t_n17) );
  XNOR2_X1 f1_round_t_U33 ( .A(f1_round_t_n16), .B(f1_round_t_n17), .ZN(
        f1_round_t_n6) );
  XOR2_X1 f1_round_t_U32 ( .A(abs1_io_state_out_0_4), .B(abs1_io_state_out_0_3), .Z(f1_round_t_n15) );
  XNOR2_X1 f1_round_t_U31 ( .A(abs1_io_state_out_0_2), .B(f1_round_t_n15), 
        .ZN(f1_round_t_n13) );
  XOR2_X1 f1_round_t_U30 ( .A(abs1_io_state_out_0_1), .B(abs1_io_state_out_0_0), .Z(f1_round_t_n14) );
  XNOR2_X1 f1_round_t_U29 ( .A(f1_round_t_n13), .B(f1_round_t_n14), .ZN(
        f1_round_t_n2) );
  XOR2_X1 f1_round_t_U28 ( .A(f1_round_t_n6), .B(f1_round_t_n2), .Z(
        f1_round_t_n12) );
  XOR2_X1 f1_round_t_U27 ( .A(abs1_io_state_out_1_0), .B(f1_round_t_n12), .Z(
        f1_round_p_io_state_out_0_2) );
  XOR2_X1 f1_round_t_U26 ( .A(abs1_io_state_out_1_1), .B(f1_round_t_n12), .Z(
        f1_round_p_io_state_out_1_0) );
  XOR2_X1 f1_round_t_U25 ( .A(abs1_io_state_out_1_2), .B(f1_round_t_n12), .Z(
        f1_round_p_io_state_out_2_3) );
  XOR2_X1 f1_round_t_U24 ( .A(abs1_io_state_out_1_3), .B(f1_round_t_n12), .Z(
        f1_round_p_io_state_out_3_1) );
  XOR2_X1 f1_round_t_U23 ( .A(abs1_io_state_out_1_4), .B(f1_round_t_n12), .Z(
        f1_round_p_io_state_out_4_4) );
  XOR2_X1 f1_round_t_U22 ( .A(abs1_io_state_out_3_4), .B(abs1_io_state_out_3_3), .Z(f1_round_t_n11) );
  XNOR2_X1 f1_round_t_U21 ( .A(abs1_io_state_out_3_2), .B(f1_round_t_n11), 
        .ZN(f1_round_t_n9) );
  XOR2_X1 f1_round_t_U20 ( .A(abs1_io_state_out_3_1), .B(abs1_io_state_out_3_0), .Z(f1_round_t_n10) );
  XNOR2_X1 f1_round_t_U19 ( .A(f1_round_t_n9), .B(f1_round_t_n10), .ZN(
        f1_round_t_n3) );
  XNOR2_X1 f1_round_t_U18 ( .A(f1_round_t_n8), .B(f1_round_t_n3), .ZN(
        f1_round_t_n7) );
  XOR2_X1 f1_round_t_U17 ( .A(abs1_io_state_out_2_0), .B(f1_round_t_n7), .Z(
        f1_round_p_io_state_out_0_4) );
  XOR2_X1 f1_round_t_U16 ( .A(abs1_io_state_out_2_1), .B(f1_round_t_n7), .Z(
        f1_round_p_io_state_out_1_2) );
  XOR2_X1 f1_round_t_U15 ( .A(abs1_io_state_out_2_2), .B(f1_round_t_n7), .Z(
        f1_round_p_io_state_out_2_0) );
  XOR2_X1 f1_round_t_U14 ( .A(abs1_io_state_out_2_3), .B(f1_round_t_n7), .Z(
        f1_round_p_io_state_out_3_3) );
  XOR2_X1 f1_round_t_U13 ( .A(abs1_io_state_out_2_4), .B(f1_round_t_n7), .Z(
        f1_round_p_io_state_out_4_1) );
  XOR2_X1 f1_round_t_U12 ( .A(f1_round_t_n5), .B(f1_round_t_n6), .Z(
        f1_round_t_n4) );
  XOR2_X1 f1_round_t_U11 ( .A(abs1_io_state_out_3_0), .B(f1_round_t_n4), .Z(
        f1_round_p_io_state_out_0_1) );
  XOR2_X1 f1_round_t_U10 ( .A(abs1_io_state_out_3_1), .B(f1_round_t_n4), .Z(
        f1_round_p_io_state_out_1_4) );
  XOR2_X1 f1_round_t_U9 ( .A(abs1_io_state_out_3_2), .B(f1_round_t_n4), .Z(
        f1_round_p_io_state_out_2_2) );
  XOR2_X1 f1_round_t_U8 ( .A(abs1_io_state_out_3_3), .B(f1_round_t_n4), .Z(
        f1_round_p_io_state_out_3_0) );
  XOR2_X1 f1_round_t_U7 ( .A(abs1_io_state_out_3_4), .B(f1_round_t_n4), .Z(
        f1_round_p_io_state_out_4_3) );
  XOR2_X1 f1_round_t_U6 ( .A(f1_round_t_n2), .B(f1_round_t_n3), .Z(
        f1_round_t_n1) );
  XOR2_X1 f1_round_t_U5 ( .A(abs1_io_state_out_4_0), .B(f1_round_t_n1), .Z(
        f1_round_p_io_state_out_0_3) );
  XOR2_X1 f1_round_t_U4 ( .A(abs1_io_state_out_4_1), .B(f1_round_t_n1), .Z(
        f1_round_p_io_state_out_1_1) );
  XOR2_X1 f1_round_t_U3 ( .A(abs1_io_state_out_4_2), .B(f1_round_t_n1), .Z(
        f1_round_p_io_state_out_2_4) );
  XOR2_X1 f1_round_t_U2 ( .A(abs1_io_state_out_4_3), .B(f1_round_t_n1), .Z(
        f1_round_p_io_state_out_3_2) );
  XOR2_X1 f1_round_t_U1 ( .A(abs1_io_state_out_4_4), .B(f1_round_t_n1), .Z(
        f1_round_p_io_state_out_4_0) );
  NAND2_X1 f1_round_c_U50 ( .A1(f1_round_p_io_state_out_2_0), .A2(
        f1_round_p_io_state_out_1_0), .ZN(f1_round_c_n25) );
  XOR2_X1 f1_round_c_U49 ( .A(f1_round_c_n25), .B(f1_round_p_io_state_out_0_0), 
        .Z(f1_round_c_io_state_out_0_0) );
  NAND2_X1 f1_round_c_U48 ( .A1(f1_round_p_io_state_out_2_1), .A2(
        f1_round_p_io_state_out_1_1), .ZN(f1_round_c_n24) );
  XOR2_X1 f1_round_c_U47 ( .A(f1_round_c_n24), .B(f1_round_p_io_state_out_0_1), 
        .Z(f1_round_io_state_out_0_1) );
  NAND2_X1 f1_round_c_U46 ( .A1(f1_round_p_io_state_out_2_2), .A2(
        f1_round_p_io_state_out_1_2), .ZN(f1_round_c_n23) );
  XOR2_X1 f1_round_c_U45 ( .A(f1_round_c_n23), .B(f1_round_p_io_state_out_0_2), 
        .Z(f1_round_io_state_out_0_2) );
  NAND2_X1 f1_round_c_U44 ( .A1(f1_round_p_io_state_out_2_3), .A2(
        f1_round_p_io_state_out_1_3), .ZN(f1_round_c_n22) );
  XOR2_X1 f1_round_c_U43 ( .A(f1_round_c_n22), .B(f1_round_p_io_state_out_0_3), 
        .Z(f1_round_io_state_out_0_3) );
  NAND2_X1 f1_round_c_U42 ( .A1(f1_round_p_io_state_out_2_4), .A2(
        f1_round_p_io_state_out_1_4), .ZN(f1_round_c_n21) );
  XOR2_X1 f1_round_c_U41 ( .A(f1_round_c_n21), .B(f1_round_p_io_state_out_0_4), 
        .Z(f1_round_io_state_out_0_4) );
  NAND2_X1 f1_round_c_U40 ( .A1(f1_round_p_io_state_out_2_0), .A2(
        f1_round_p_io_state_out_3_0), .ZN(f1_round_c_n20) );
  XOR2_X1 f1_round_c_U39 ( .A(f1_round_c_n20), .B(f1_round_p_io_state_out_1_0), 
        .Z(f1_round_io_state_out_1_0) );
  NAND2_X1 f1_round_c_U38 ( .A1(f1_round_p_io_state_out_2_1), .A2(
        f1_round_p_io_state_out_3_1), .ZN(f1_round_c_n19) );
  XOR2_X1 f1_round_c_U37 ( .A(f1_round_c_n19), .B(f1_round_p_io_state_out_1_1), 
        .Z(f1_round_io_state_out_1_1) );
  NAND2_X1 f1_round_c_U36 ( .A1(f1_round_p_io_state_out_2_2), .A2(
        f1_round_p_io_state_out_3_2), .ZN(f1_round_c_n18) );
  XOR2_X1 f1_round_c_U35 ( .A(f1_round_c_n18), .B(f1_round_p_io_state_out_1_2), 
        .Z(f1_round_io_state_out_1_2) );
  NAND2_X1 f1_round_c_U34 ( .A1(f1_round_p_io_state_out_2_3), .A2(
        f1_round_p_io_state_out_3_3), .ZN(f1_round_c_n17) );
  XOR2_X1 f1_round_c_U33 ( .A(f1_round_c_n17), .B(f1_round_p_io_state_out_1_3), 
        .Z(f1_round_io_state_out_1_3) );
  NAND2_X1 f1_round_c_U32 ( .A1(f1_round_p_io_state_out_2_4), .A2(
        f1_round_p_io_state_out_3_4), .ZN(f1_round_c_n16) );
  XOR2_X1 f1_round_c_U31 ( .A(f1_round_c_n16), .B(f1_round_p_io_state_out_1_4), 
        .Z(f1_round_io_state_out_1_4) );
  NAND2_X1 f1_round_c_U30 ( .A1(f1_round_p_io_state_out_3_0), .A2(
        f1_round_p_io_state_out_4_0), .ZN(f1_round_c_n15) );
  XOR2_X1 f1_round_c_U29 ( .A(f1_round_c_n15), .B(f1_round_p_io_state_out_2_0), 
        .Z(f1_round_io_state_out_2_0) );
  NAND2_X1 f1_round_c_U28 ( .A1(f1_round_p_io_state_out_3_1), .A2(
        f1_round_p_io_state_out_4_1), .ZN(f1_round_c_n14) );
  XOR2_X1 f1_round_c_U27 ( .A(f1_round_c_n14), .B(f1_round_p_io_state_out_2_1), 
        .Z(f1_round_io_state_out_2_1) );
  NAND2_X1 f1_round_c_U26 ( .A1(f1_round_p_io_state_out_3_2), .A2(
        f1_round_p_io_state_out_4_2), .ZN(f1_round_c_n13) );
  XOR2_X1 f1_round_c_U25 ( .A(f1_round_c_n13), .B(f1_round_p_io_state_out_2_2), 
        .Z(f1_round_io_state_out_2_2) );
  NAND2_X1 f1_round_c_U24 ( .A1(f1_round_p_io_state_out_3_3), .A2(
        f1_round_p_io_state_out_4_3), .ZN(f1_round_c_n12) );
  XOR2_X1 f1_round_c_U23 ( .A(f1_round_c_n12), .B(f1_round_p_io_state_out_2_3), 
        .Z(f1_round_io_state_out_2_3) );
  NAND2_X1 f1_round_c_U22 ( .A1(f1_round_p_io_state_out_3_4), .A2(
        f1_round_p_io_state_out_4_4), .ZN(f1_round_c_n11) );
  XOR2_X1 f1_round_c_U21 ( .A(f1_round_c_n11), .B(f1_round_p_io_state_out_2_4), 
        .Z(f1_round_io_state_out_2_4) );
  NAND2_X1 f1_round_c_U20 ( .A1(f1_round_p_io_state_out_4_0), .A2(
        f1_round_p_io_state_out_0_0), .ZN(f1_round_c_n10) );
  XOR2_X1 f1_round_c_U19 ( .A(f1_round_c_n10), .B(f1_round_p_io_state_out_3_0), 
        .Z(f1_round_io_state_out_3_0) );
  NAND2_X1 f1_round_c_U18 ( .A1(f1_round_p_io_state_out_4_1), .A2(
        f1_round_p_io_state_out_0_1), .ZN(f1_round_c_n9) );
  XOR2_X1 f1_round_c_U17 ( .A(f1_round_c_n9), .B(f1_round_p_io_state_out_3_1), 
        .Z(f1_round_io_state_out_3_1) );
  NAND2_X1 f1_round_c_U16 ( .A1(f1_round_p_io_state_out_4_2), .A2(
        f1_round_p_io_state_out_0_2), .ZN(f1_round_c_n8) );
  XOR2_X1 f1_round_c_U15 ( .A(f1_round_c_n8), .B(f1_round_p_io_state_out_3_2), 
        .Z(f1_round_io_state_out_3_2) );
  NAND2_X1 f1_round_c_U14 ( .A1(f1_round_p_io_state_out_4_3), .A2(
        f1_round_p_io_state_out_0_3), .ZN(f1_round_c_n7) );
  XOR2_X1 f1_round_c_U13 ( .A(f1_round_c_n7), .B(f1_round_p_io_state_out_3_3), 
        .Z(f1_round_io_state_out_3_3) );
  NAND2_X1 f1_round_c_U12 ( .A1(f1_round_p_io_state_out_4_4), .A2(
        f1_round_p_io_state_out_0_4), .ZN(f1_round_c_n6) );
  XOR2_X1 f1_round_c_U11 ( .A(f1_round_c_n6), .B(f1_round_p_io_state_out_3_4), 
        .Z(f1_round_io_state_out_3_4) );
  NAND2_X1 f1_round_c_U10 ( .A1(f1_round_p_io_state_out_1_0), .A2(
        f1_round_p_io_state_out_0_0), .ZN(f1_round_c_n5) );
  XOR2_X1 f1_round_c_U9 ( .A(f1_round_c_n5), .B(f1_round_p_io_state_out_4_0), 
        .Z(f1_round_io_state_out_4_0) );
  NAND2_X1 f1_round_c_U8 ( .A1(f1_round_p_io_state_out_1_1), .A2(
        f1_round_p_io_state_out_0_1), .ZN(f1_round_c_n4) );
  XOR2_X1 f1_round_c_U7 ( .A(f1_round_c_n4), .B(f1_round_p_io_state_out_4_1), 
        .Z(f1_round_io_state_out_4_1) );
  NAND2_X1 f1_round_c_U6 ( .A1(f1_round_p_io_state_out_1_2), .A2(
        f1_round_p_io_state_out_0_2), .ZN(f1_round_c_n3) );
  XOR2_X1 f1_round_c_U5 ( .A(f1_round_c_n3), .B(f1_round_p_io_state_out_4_2), 
        .Z(f1_round_io_state_out_4_2) );
  NAND2_X1 f1_round_c_U4 ( .A1(f1_round_p_io_state_out_1_3), .A2(
        f1_round_p_io_state_out_0_3), .ZN(f1_round_c_n2) );
  XOR2_X1 f1_round_c_U3 ( .A(f1_round_c_n2), .B(f1_round_p_io_state_out_4_3), 
        .Z(f1_round_io_state_out_4_3) );
  NAND2_X1 f1_round_c_U2 ( .A1(f1_round_p_io_state_out_1_4), .A2(
        f1_round_p_io_state_out_0_4), .ZN(f1_round_c_n1) );
  XOR2_X1 f1_round_c_U1 ( .A(f1_round_c_n1), .B(f1_round_p_io_state_out_4_4), 
        .Z(f1_round_io_state_out_4_4) );
  INV_X1 f1_round_i_U1 ( .A(f1_round_c_io_state_out_0_0), .ZN(
        f1_round_io_state_out_0_0) );
  XOR2_X1 f1_round_1_t_U50 ( .A(f1_round_io_state_out_1_4), .B(
        f1_round_io_state_out_1_3), .Z(f1_round_1_t_n25) );
  XNOR2_X1 f1_round_1_t_U49 ( .A(f1_round_io_state_out_1_2), .B(
        f1_round_1_t_n25), .ZN(f1_round_1_t_n23) );
  XOR2_X1 f1_round_1_t_U48 ( .A(f1_round_io_state_out_1_1), .B(
        f1_round_io_state_out_1_0), .Z(f1_round_1_t_n24) );
  XOR2_X1 f1_round_1_t_U47 ( .A(f1_round_1_t_n23), .B(f1_round_1_t_n24), .Z(
        f1_round_1_t_n8) );
  XOR2_X1 f1_round_1_t_U46 ( .A(f1_round_io_state_out_4_4), .B(
        f1_round_io_state_out_4_3), .Z(f1_round_1_t_n22) );
  XNOR2_X1 f1_round_1_t_U45 ( .A(f1_round_io_state_out_4_2), .B(
        f1_round_1_t_n22), .ZN(f1_round_1_t_n20) );
  XOR2_X1 f1_round_1_t_U44 ( .A(f1_round_io_state_out_4_1), .B(
        f1_round_io_state_out_4_0), .Z(f1_round_1_t_n21) );
  XNOR2_X1 f1_round_1_t_U43 ( .A(f1_round_1_t_n20), .B(f1_round_1_t_n21), .ZN(
        f1_round_1_t_n5) );
  XNOR2_X1 f1_round_1_t_U42 ( .A(f1_round_1_t_n8), .B(f1_round_1_t_n5), .ZN(
        f1_round_1_t_n19) );
  XOR2_X1 f1_round_1_t_U41 ( .A(f1_round_io_state_out_0_0), .B(
        f1_round_1_t_n19), .Z(f1_round_1_p_io_state_out_0_0) );
  XOR2_X1 f1_round_1_t_U40 ( .A(f1_round_io_state_out_0_1), .B(
        f1_round_1_t_n19), .Z(f1_round_1_p_io_state_out_1_3) );
  XOR2_X1 f1_round_1_t_U39 ( .A(f1_round_io_state_out_0_2), .B(
        f1_round_1_t_n19), .Z(f1_round_1_p_io_state_out_2_1) );
  XOR2_X1 f1_round_1_t_U38 ( .A(f1_round_io_state_out_0_3), .B(
        f1_round_1_t_n19), .Z(f1_round_1_p_io_state_out_3_4) );
  XOR2_X1 f1_round_1_t_U37 ( .A(f1_round_io_state_out_0_4), .B(
        f1_round_1_t_n19), .Z(f1_round_1_p_io_state_out_4_2) );
  XOR2_X1 f1_round_1_t_U36 ( .A(f1_round_io_state_out_2_4), .B(
        f1_round_io_state_out_2_3), .Z(f1_round_1_t_n18) );
  XNOR2_X1 f1_round_1_t_U35 ( .A(f1_round_io_state_out_2_2), .B(
        f1_round_1_t_n18), .ZN(f1_round_1_t_n16) );
  XOR2_X1 f1_round_1_t_U34 ( .A(f1_round_io_state_out_2_1), .B(
        f1_round_io_state_out_2_0), .Z(f1_round_1_t_n17) );
  XNOR2_X1 f1_round_1_t_U33 ( .A(f1_round_1_t_n16), .B(f1_round_1_t_n17), .ZN(
        f1_round_1_t_n6) );
  XOR2_X1 f1_round_1_t_U32 ( .A(f1_round_io_state_out_0_4), .B(
        f1_round_io_state_out_0_3), .Z(f1_round_1_t_n15) );
  XNOR2_X1 f1_round_1_t_U31 ( .A(f1_round_io_state_out_0_2), .B(
        f1_round_1_t_n15), .ZN(f1_round_1_t_n13) );
  XOR2_X1 f1_round_1_t_U30 ( .A(f1_round_io_state_out_0_1), .B(
        f1_round_io_state_out_0_0), .Z(f1_round_1_t_n14) );
  XNOR2_X1 f1_round_1_t_U29 ( .A(f1_round_1_t_n13), .B(f1_round_1_t_n14), .ZN(
        f1_round_1_t_n2) );
  XOR2_X1 f1_round_1_t_U28 ( .A(f1_round_1_t_n6), .B(f1_round_1_t_n2), .Z(
        f1_round_1_t_n12) );
  XOR2_X1 f1_round_1_t_U27 ( .A(f1_round_io_state_out_1_0), .B(
        f1_round_1_t_n12), .Z(f1_round_1_p_io_state_out_0_2) );
  XOR2_X1 f1_round_1_t_U26 ( .A(f1_round_io_state_out_1_1), .B(
        f1_round_1_t_n12), .Z(f1_round_1_p_io_state_out_1_0) );
  XOR2_X1 f1_round_1_t_U25 ( .A(f1_round_io_state_out_1_2), .B(
        f1_round_1_t_n12), .Z(f1_round_1_p_io_state_out_2_3) );
  XOR2_X1 f1_round_1_t_U24 ( .A(f1_round_io_state_out_1_3), .B(
        f1_round_1_t_n12), .Z(f1_round_1_p_io_state_out_3_1) );
  XOR2_X1 f1_round_1_t_U23 ( .A(f1_round_io_state_out_1_4), .B(
        f1_round_1_t_n12), .Z(f1_round_1_p_io_state_out_4_4) );
  XOR2_X1 f1_round_1_t_U22 ( .A(f1_round_io_state_out_3_4), .B(
        f1_round_io_state_out_3_3), .Z(f1_round_1_t_n11) );
  XNOR2_X1 f1_round_1_t_U21 ( .A(f1_round_io_state_out_3_2), .B(
        f1_round_1_t_n11), .ZN(f1_round_1_t_n9) );
  XOR2_X1 f1_round_1_t_U20 ( .A(f1_round_io_state_out_3_1), .B(
        f1_round_io_state_out_3_0), .Z(f1_round_1_t_n10) );
  XNOR2_X1 f1_round_1_t_U19 ( .A(f1_round_1_t_n9), .B(f1_round_1_t_n10), .ZN(
        f1_round_1_t_n3) );
  XNOR2_X1 f1_round_1_t_U18 ( .A(f1_round_1_t_n8), .B(f1_round_1_t_n3), .ZN(
        f1_round_1_t_n7) );
  XOR2_X1 f1_round_1_t_U17 ( .A(f1_round_io_state_out_2_0), .B(f1_round_1_t_n7), .Z(f1_round_1_p_io_state_out_0_4) );
  XOR2_X1 f1_round_1_t_U16 ( .A(f1_round_io_state_out_2_1), .B(f1_round_1_t_n7), .Z(f1_round_1_p_io_state_out_1_2) );
  XOR2_X1 f1_round_1_t_U15 ( .A(f1_round_io_state_out_2_2), .B(f1_round_1_t_n7), .Z(f1_round_1_p_io_state_out_2_0) );
  XOR2_X1 f1_round_1_t_U14 ( .A(f1_round_io_state_out_2_3), .B(f1_round_1_t_n7), .Z(f1_round_1_p_io_state_out_3_3) );
  XOR2_X1 f1_round_1_t_U13 ( .A(f1_round_io_state_out_2_4), .B(f1_round_1_t_n7), .Z(f1_round_1_p_io_state_out_4_1) );
  XOR2_X1 f1_round_1_t_U12 ( .A(f1_round_1_t_n5), .B(f1_round_1_t_n6), .Z(
        f1_round_1_t_n4) );
  XOR2_X1 f1_round_1_t_U11 ( .A(f1_round_io_state_out_3_0), .B(f1_round_1_t_n4), .Z(f1_round_1_p_io_state_out_0_1) );
  XOR2_X1 f1_round_1_t_U10 ( .A(f1_round_io_state_out_3_1), .B(f1_round_1_t_n4), .Z(f1_round_1_p_io_state_out_1_4) );
  XOR2_X1 f1_round_1_t_U9 ( .A(f1_round_io_state_out_3_2), .B(f1_round_1_t_n4), 
        .Z(f1_round_1_p_io_state_out_2_2) );
  XOR2_X1 f1_round_1_t_U8 ( .A(f1_round_io_state_out_3_3), .B(f1_round_1_t_n4), 
        .Z(f1_round_1_p_io_state_out_3_0) );
  XOR2_X1 f1_round_1_t_U7 ( .A(f1_round_io_state_out_3_4), .B(f1_round_1_t_n4), 
        .Z(f1_round_1_p_io_state_out_4_3) );
  XOR2_X1 f1_round_1_t_U6 ( .A(f1_round_1_t_n2), .B(f1_round_1_t_n3), .Z(
        f1_round_1_t_n1) );
  XOR2_X1 f1_round_1_t_U5 ( .A(f1_round_io_state_out_4_0), .B(f1_round_1_t_n1), 
        .Z(f1_round_1_p_io_state_out_0_3) );
  XOR2_X1 f1_round_1_t_U4 ( .A(f1_round_io_state_out_4_1), .B(f1_round_1_t_n1), 
        .Z(f1_round_1_p_io_state_out_1_1) );
  XOR2_X1 f1_round_1_t_U3 ( .A(f1_round_io_state_out_4_2), .B(f1_round_1_t_n1), 
        .Z(f1_round_1_p_io_state_out_2_4) );
  XOR2_X1 f1_round_1_t_U2 ( .A(f1_round_io_state_out_4_3), .B(f1_round_1_t_n1), 
        .Z(f1_round_1_p_io_state_out_3_2) );
  XOR2_X1 f1_round_1_t_U1 ( .A(f1_round_io_state_out_4_4), .B(f1_round_1_t_n1), 
        .Z(f1_round_1_p_io_state_out_4_0) );
  NAND2_X1 f1_round_1_c_U50 ( .A1(f1_round_1_p_io_state_out_2_0), .A2(
        f1_round_1_p_io_state_out_1_0), .ZN(f1_round_1_c_n25) );
  XOR2_X1 f1_round_1_c_U49 ( .A(f1_round_1_c_n25), .B(
        f1_round_1_p_io_state_out_0_0), .Z(f1_round_1_io_state_out_0_0) );
  NAND2_X1 f1_round_1_c_U48 ( .A1(f1_round_1_p_io_state_out_2_1), .A2(
        f1_round_1_p_io_state_out_1_1), .ZN(f1_round_1_c_n24) );
  XOR2_X1 f1_round_1_c_U47 ( .A(f1_round_1_c_n24), .B(
        f1_round_1_p_io_state_out_0_1), .Z(f1_round_1_io_state_out_0_1) );
  NAND2_X1 f1_round_1_c_U46 ( .A1(f1_round_1_p_io_state_out_2_2), .A2(
        f1_round_1_p_io_state_out_1_2), .ZN(f1_round_1_c_n23) );
  XOR2_X1 f1_round_1_c_U45 ( .A(f1_round_1_c_n23), .B(
        f1_round_1_p_io_state_out_0_2), .Z(f1_round_1_io_state_out_0_2) );
  NAND2_X1 f1_round_1_c_U44 ( .A1(f1_round_1_p_io_state_out_2_3), .A2(
        f1_round_1_p_io_state_out_1_3), .ZN(f1_round_1_c_n22) );
  XOR2_X1 f1_round_1_c_U43 ( .A(f1_round_1_c_n22), .B(
        f1_round_1_p_io_state_out_0_3), .Z(f1_round_1_io_state_out_0_3) );
  NAND2_X1 f1_round_1_c_U42 ( .A1(f1_round_1_p_io_state_out_2_4), .A2(
        f1_round_1_p_io_state_out_1_4), .ZN(f1_round_1_c_n21) );
  XOR2_X1 f1_round_1_c_U41 ( .A(f1_round_1_c_n21), .B(
        f1_round_1_p_io_state_out_0_4), .Z(f1_round_1_io_state_out_0_4) );
  NAND2_X1 f1_round_1_c_U40 ( .A1(f1_round_1_p_io_state_out_2_0), .A2(
        f1_round_1_p_io_state_out_3_0), .ZN(f1_round_1_c_n20) );
  XOR2_X1 f1_round_1_c_U39 ( .A(f1_round_1_c_n20), .B(
        f1_round_1_p_io_state_out_1_0), .Z(f1_round_1_io_state_out_1_0) );
  NAND2_X1 f1_round_1_c_U38 ( .A1(f1_round_1_p_io_state_out_2_1), .A2(
        f1_round_1_p_io_state_out_3_1), .ZN(f1_round_1_c_n19) );
  XOR2_X1 f1_round_1_c_U37 ( .A(f1_round_1_c_n19), .B(
        f1_round_1_p_io_state_out_1_1), .Z(f1_round_1_io_state_out_1_1) );
  NAND2_X1 f1_round_1_c_U36 ( .A1(f1_round_1_p_io_state_out_2_2), .A2(
        f1_round_1_p_io_state_out_3_2), .ZN(f1_round_1_c_n18) );
  XOR2_X1 f1_round_1_c_U35 ( .A(f1_round_1_c_n18), .B(
        f1_round_1_p_io_state_out_1_2), .Z(f1_round_1_io_state_out_1_2) );
  NAND2_X1 f1_round_1_c_U34 ( .A1(f1_round_1_p_io_state_out_2_3), .A2(
        f1_round_1_p_io_state_out_3_3), .ZN(f1_round_1_c_n17) );
  XOR2_X1 f1_round_1_c_U33 ( .A(f1_round_1_c_n17), .B(
        f1_round_1_p_io_state_out_1_3), .Z(f1_round_1_io_state_out_1_3) );
  NAND2_X1 f1_round_1_c_U32 ( .A1(f1_round_1_p_io_state_out_2_4), .A2(
        f1_round_1_p_io_state_out_3_4), .ZN(f1_round_1_c_n16) );
  XOR2_X1 f1_round_1_c_U31 ( .A(f1_round_1_c_n16), .B(
        f1_round_1_p_io_state_out_1_4), .Z(f1_round_1_io_state_out_1_4) );
  NAND2_X1 f1_round_1_c_U30 ( .A1(f1_round_1_p_io_state_out_3_0), .A2(
        f1_round_1_p_io_state_out_4_0), .ZN(f1_round_1_c_n15) );
  XOR2_X1 f1_round_1_c_U29 ( .A(f1_round_1_c_n15), .B(
        f1_round_1_p_io_state_out_2_0), .Z(f1_round_1_io_state_out_2_0) );
  NAND2_X1 f1_round_1_c_U28 ( .A1(f1_round_1_p_io_state_out_3_1), .A2(
        f1_round_1_p_io_state_out_4_1), .ZN(f1_round_1_c_n14) );
  XOR2_X1 f1_round_1_c_U27 ( .A(f1_round_1_c_n14), .B(
        f1_round_1_p_io_state_out_2_1), .Z(f1_round_1_io_state_out_2_1) );
  NAND2_X1 f1_round_1_c_U26 ( .A1(f1_round_1_p_io_state_out_3_2), .A2(
        f1_round_1_p_io_state_out_4_2), .ZN(f1_round_1_c_n13) );
  XOR2_X1 f1_round_1_c_U25 ( .A(f1_round_1_c_n13), .B(
        f1_round_1_p_io_state_out_2_2), .Z(f1_round_1_io_state_out_2_2) );
  NAND2_X1 f1_round_1_c_U24 ( .A1(f1_round_1_p_io_state_out_3_3), .A2(
        f1_round_1_p_io_state_out_4_3), .ZN(f1_round_1_c_n12) );
  XOR2_X1 f1_round_1_c_U23 ( .A(f1_round_1_c_n12), .B(
        f1_round_1_p_io_state_out_2_3), .Z(f1_round_1_io_state_out_2_3) );
  NAND2_X1 f1_round_1_c_U22 ( .A1(f1_round_1_p_io_state_out_3_4), .A2(
        f1_round_1_p_io_state_out_4_4), .ZN(f1_round_1_c_n11) );
  XOR2_X1 f1_round_1_c_U21 ( .A(f1_round_1_c_n11), .B(
        f1_round_1_p_io_state_out_2_4), .Z(f1_round_1_io_state_out_2_4) );
  NAND2_X1 f1_round_1_c_U20 ( .A1(f1_round_1_p_io_state_out_4_0), .A2(
        f1_round_1_p_io_state_out_0_0), .ZN(f1_round_1_c_n10) );
  XOR2_X1 f1_round_1_c_U19 ( .A(f1_round_1_c_n10), .B(
        f1_round_1_p_io_state_out_3_0), .Z(f1_round_1_io_state_out_3_0) );
  NAND2_X1 f1_round_1_c_U18 ( .A1(f1_round_1_p_io_state_out_4_1), .A2(
        f1_round_1_p_io_state_out_0_1), .ZN(f1_round_1_c_n9) );
  XOR2_X1 f1_round_1_c_U17 ( .A(f1_round_1_c_n9), .B(
        f1_round_1_p_io_state_out_3_1), .Z(f1_round_1_io_state_out_3_1) );
  NAND2_X1 f1_round_1_c_U16 ( .A1(f1_round_1_p_io_state_out_4_2), .A2(
        f1_round_1_p_io_state_out_0_2), .ZN(f1_round_1_c_n8) );
  XOR2_X1 f1_round_1_c_U15 ( .A(f1_round_1_c_n8), .B(
        f1_round_1_p_io_state_out_3_2), .Z(f1_round_1_io_state_out_3_2) );
  NAND2_X1 f1_round_1_c_U14 ( .A1(f1_round_1_p_io_state_out_4_3), .A2(
        f1_round_1_p_io_state_out_0_3), .ZN(f1_round_1_c_n7) );
  XOR2_X1 f1_round_1_c_U13 ( .A(f1_round_1_c_n7), .B(
        f1_round_1_p_io_state_out_3_3), .Z(f1_round_1_io_state_out_3_3) );
  NAND2_X1 f1_round_1_c_U12 ( .A1(f1_round_1_p_io_state_out_4_4), .A2(
        f1_round_1_p_io_state_out_0_4), .ZN(f1_round_1_c_n6) );
  XOR2_X1 f1_round_1_c_U11 ( .A(f1_round_1_c_n6), .B(
        f1_round_1_p_io_state_out_3_4), .Z(f1_round_1_io_state_out_3_4) );
  NAND2_X1 f1_round_1_c_U10 ( .A1(f1_round_1_p_io_state_out_1_0), .A2(
        f1_round_1_p_io_state_out_0_0), .ZN(f1_round_1_c_n5) );
  XOR2_X1 f1_round_1_c_U9 ( .A(f1_round_1_c_n5), .B(
        f1_round_1_p_io_state_out_4_0), .Z(f1_round_1_io_state_out_4_0) );
  NAND2_X1 f1_round_1_c_U8 ( .A1(f1_round_1_p_io_state_out_1_1), .A2(
        f1_round_1_p_io_state_out_0_1), .ZN(f1_round_1_c_n4) );
  XOR2_X1 f1_round_1_c_U7 ( .A(f1_round_1_c_n4), .B(
        f1_round_1_p_io_state_out_4_1), .Z(f1_round_1_io_state_out_4_1) );
  NAND2_X1 f1_round_1_c_U6 ( .A1(f1_round_1_p_io_state_out_1_2), .A2(
        f1_round_1_p_io_state_out_0_2), .ZN(f1_round_1_c_n3) );
  XOR2_X1 f1_round_1_c_U5 ( .A(f1_round_1_c_n3), .B(
        f1_round_1_p_io_state_out_4_2), .Z(f1_round_1_io_state_out_4_2) );
  NAND2_X1 f1_round_1_c_U4 ( .A1(f1_round_1_p_io_state_out_1_3), .A2(
        f1_round_1_p_io_state_out_0_3), .ZN(f1_round_1_c_n2) );
  XOR2_X1 f1_round_1_c_U3 ( .A(f1_round_1_c_n2), .B(
        f1_round_1_p_io_state_out_4_3), .Z(f1_round_1_io_state_out_4_3) );
  NAND2_X1 f1_round_1_c_U2 ( .A1(f1_round_1_p_io_state_out_1_4), .A2(
        f1_round_1_p_io_state_out_0_4), .ZN(f1_round_1_c_n1) );
  XOR2_X1 f1_round_1_c_U1 ( .A(f1_round_1_c_n1), .B(
        f1_round_1_p_io_state_out_4_4), .Z(f1_round_1_io_state_out_4_4) );
  XOR2_X1 f1_round_2_t_U50 ( .A(f1_round_1_io_state_out_1_4), .B(
        f1_round_1_io_state_out_1_3), .Z(f1_round_2_t_n25) );
  XNOR2_X1 f1_round_2_t_U49 ( .A(f1_round_1_io_state_out_1_2), .B(
        f1_round_2_t_n25), .ZN(f1_round_2_t_n23) );
  XOR2_X1 f1_round_2_t_U48 ( .A(f1_round_1_io_state_out_1_1), .B(
        f1_round_1_io_state_out_1_0), .Z(f1_round_2_t_n24) );
  XOR2_X1 f1_round_2_t_U47 ( .A(f1_round_2_t_n23), .B(f1_round_2_t_n24), .Z(
        f1_round_2_t_n8) );
  XOR2_X1 f1_round_2_t_U46 ( .A(f1_round_1_io_state_out_4_4), .B(
        f1_round_1_io_state_out_4_3), .Z(f1_round_2_t_n22) );
  XNOR2_X1 f1_round_2_t_U45 ( .A(f1_round_1_io_state_out_4_2), .B(
        f1_round_2_t_n22), .ZN(f1_round_2_t_n20) );
  XOR2_X1 f1_round_2_t_U44 ( .A(f1_round_1_io_state_out_4_1), .B(
        f1_round_1_io_state_out_4_0), .Z(f1_round_2_t_n21) );
  XNOR2_X1 f1_round_2_t_U43 ( .A(f1_round_2_t_n20), .B(f1_round_2_t_n21), .ZN(
        f1_round_2_t_n5) );
  XNOR2_X1 f1_round_2_t_U42 ( .A(f1_round_2_t_n8), .B(f1_round_2_t_n5), .ZN(
        f1_round_2_t_n19) );
  XOR2_X1 f1_round_2_t_U41 ( .A(f1_round_1_io_state_out_0_0), .B(
        f1_round_2_t_n19), .Z(f1_round_2_p_io_state_out_0_0) );
  XOR2_X1 f1_round_2_t_U40 ( .A(f1_round_1_io_state_out_0_1), .B(
        f1_round_2_t_n19), .Z(f1_round_2_p_io_state_out_1_3) );
  XOR2_X1 f1_round_2_t_U39 ( .A(f1_round_1_io_state_out_0_2), .B(
        f1_round_2_t_n19), .Z(f1_round_2_p_io_state_out_2_1) );
  XOR2_X1 f1_round_2_t_U38 ( .A(f1_round_1_io_state_out_0_3), .B(
        f1_round_2_t_n19), .Z(f1_round_2_p_io_state_out_3_4) );
  XOR2_X1 f1_round_2_t_U37 ( .A(f1_round_1_io_state_out_0_4), .B(
        f1_round_2_t_n19), .Z(f1_round_2_p_io_state_out_4_2) );
  XOR2_X1 f1_round_2_t_U36 ( .A(f1_round_1_io_state_out_2_4), .B(
        f1_round_1_io_state_out_2_3), .Z(f1_round_2_t_n18) );
  XNOR2_X1 f1_round_2_t_U35 ( .A(f1_round_1_io_state_out_2_2), .B(
        f1_round_2_t_n18), .ZN(f1_round_2_t_n16) );
  XOR2_X1 f1_round_2_t_U34 ( .A(f1_round_1_io_state_out_2_1), .B(
        f1_round_1_io_state_out_2_0), .Z(f1_round_2_t_n17) );
  XNOR2_X1 f1_round_2_t_U33 ( .A(f1_round_2_t_n16), .B(f1_round_2_t_n17), .ZN(
        f1_round_2_t_n6) );
  XOR2_X1 f1_round_2_t_U32 ( .A(f1_round_1_io_state_out_0_4), .B(
        f1_round_1_io_state_out_0_3), .Z(f1_round_2_t_n15) );
  XNOR2_X1 f1_round_2_t_U31 ( .A(f1_round_1_io_state_out_0_2), .B(
        f1_round_2_t_n15), .ZN(f1_round_2_t_n13) );
  XOR2_X1 f1_round_2_t_U30 ( .A(f1_round_1_io_state_out_0_1), .B(
        f1_round_1_io_state_out_0_0), .Z(f1_round_2_t_n14) );
  XNOR2_X1 f1_round_2_t_U29 ( .A(f1_round_2_t_n13), .B(f1_round_2_t_n14), .ZN(
        f1_round_2_t_n2) );
  XOR2_X1 f1_round_2_t_U28 ( .A(f1_round_2_t_n6), .B(f1_round_2_t_n2), .Z(
        f1_round_2_t_n12) );
  XOR2_X1 f1_round_2_t_U27 ( .A(f1_round_1_io_state_out_1_0), .B(
        f1_round_2_t_n12), .Z(f1_round_2_p_io_state_out_0_2) );
  XOR2_X1 f1_round_2_t_U26 ( .A(f1_round_1_io_state_out_1_1), .B(
        f1_round_2_t_n12), .Z(f1_round_2_p_io_state_out_1_0) );
  XOR2_X1 f1_round_2_t_U25 ( .A(f1_round_1_io_state_out_1_2), .B(
        f1_round_2_t_n12), .Z(f1_round_2_p_io_state_out_2_3) );
  XOR2_X1 f1_round_2_t_U24 ( .A(f1_round_1_io_state_out_1_3), .B(
        f1_round_2_t_n12), .Z(f1_round_2_p_io_state_out_3_1) );
  XOR2_X1 f1_round_2_t_U23 ( .A(f1_round_1_io_state_out_1_4), .B(
        f1_round_2_t_n12), .Z(f1_round_2_p_io_state_out_4_4) );
  XOR2_X1 f1_round_2_t_U22 ( .A(f1_round_1_io_state_out_3_4), .B(
        f1_round_1_io_state_out_3_3), .Z(f1_round_2_t_n11) );
  XNOR2_X1 f1_round_2_t_U21 ( .A(f1_round_1_io_state_out_3_2), .B(
        f1_round_2_t_n11), .ZN(f1_round_2_t_n9) );
  XOR2_X1 f1_round_2_t_U20 ( .A(f1_round_1_io_state_out_3_1), .B(
        f1_round_1_io_state_out_3_0), .Z(f1_round_2_t_n10) );
  XNOR2_X1 f1_round_2_t_U19 ( .A(f1_round_2_t_n9), .B(f1_round_2_t_n10), .ZN(
        f1_round_2_t_n3) );
  XNOR2_X1 f1_round_2_t_U18 ( .A(f1_round_2_t_n8), .B(f1_round_2_t_n3), .ZN(
        f1_round_2_t_n7) );
  XOR2_X1 f1_round_2_t_U17 ( .A(f1_round_1_io_state_out_2_0), .B(
        f1_round_2_t_n7), .Z(f1_round_2_p_io_state_out_0_4) );
  XOR2_X1 f1_round_2_t_U16 ( .A(f1_round_1_io_state_out_2_1), .B(
        f1_round_2_t_n7), .Z(f1_round_2_p_io_state_out_1_2) );
  XOR2_X1 f1_round_2_t_U15 ( .A(f1_round_1_io_state_out_2_2), .B(
        f1_round_2_t_n7), .Z(f1_round_2_p_io_state_out_2_0) );
  XOR2_X1 f1_round_2_t_U14 ( .A(f1_round_1_io_state_out_2_3), .B(
        f1_round_2_t_n7), .Z(f1_round_2_p_io_state_out_3_3) );
  XOR2_X1 f1_round_2_t_U13 ( .A(f1_round_1_io_state_out_2_4), .B(
        f1_round_2_t_n7), .Z(f1_round_2_p_io_state_out_4_1) );
  XOR2_X1 f1_round_2_t_U12 ( .A(f1_round_2_t_n5), .B(f1_round_2_t_n6), .Z(
        f1_round_2_t_n4) );
  XOR2_X1 f1_round_2_t_U11 ( .A(f1_round_1_io_state_out_3_0), .B(
        f1_round_2_t_n4), .Z(f1_round_2_p_io_state_out_0_1) );
  XOR2_X1 f1_round_2_t_U10 ( .A(f1_round_1_io_state_out_3_1), .B(
        f1_round_2_t_n4), .Z(f1_round_2_p_io_state_out_1_4) );
  XOR2_X1 f1_round_2_t_U9 ( .A(f1_round_1_io_state_out_3_2), .B(
        f1_round_2_t_n4), .Z(f1_round_2_p_io_state_out_2_2) );
  XOR2_X1 f1_round_2_t_U8 ( .A(f1_round_1_io_state_out_3_3), .B(
        f1_round_2_t_n4), .Z(f1_round_2_p_io_state_out_3_0) );
  XOR2_X1 f1_round_2_t_U7 ( .A(f1_round_1_io_state_out_3_4), .B(
        f1_round_2_t_n4), .Z(f1_round_2_p_io_state_out_4_3) );
  XOR2_X1 f1_round_2_t_U6 ( .A(f1_round_2_t_n2), .B(f1_round_2_t_n3), .Z(
        f1_round_2_t_n1) );
  XOR2_X1 f1_round_2_t_U5 ( .A(f1_round_1_io_state_out_4_0), .B(
        f1_round_2_t_n1), .Z(f1_round_2_p_io_state_out_0_3) );
  XOR2_X1 f1_round_2_t_U4 ( .A(f1_round_1_io_state_out_4_1), .B(
        f1_round_2_t_n1), .Z(f1_round_2_p_io_state_out_1_1) );
  XOR2_X1 f1_round_2_t_U3 ( .A(f1_round_1_io_state_out_4_2), .B(
        f1_round_2_t_n1), .Z(f1_round_2_p_io_state_out_2_4) );
  XOR2_X1 f1_round_2_t_U2 ( .A(f1_round_1_io_state_out_4_3), .B(
        f1_round_2_t_n1), .Z(f1_round_2_p_io_state_out_3_2) );
  XOR2_X1 f1_round_2_t_U1 ( .A(f1_round_1_io_state_out_4_4), .B(
        f1_round_2_t_n1), .Z(f1_round_2_p_io_state_out_4_0) );
  NAND2_X1 f1_round_2_c_U50 ( .A1(f1_round_2_p_io_state_out_2_0), .A2(
        f1_round_2_p_io_state_out_1_0), .ZN(f1_round_2_c_n25) );
  XOR2_X1 f1_round_2_c_U49 ( .A(f1_round_2_c_n25), .B(
        f1_round_2_p_io_state_out_0_0), .Z(f1_round_2_io_state_out_0_0) );
  NAND2_X1 f1_round_2_c_U48 ( .A1(f1_round_2_p_io_state_out_2_1), .A2(
        f1_round_2_p_io_state_out_1_1), .ZN(f1_round_2_c_n24) );
  XOR2_X1 f1_round_2_c_U47 ( .A(f1_round_2_c_n24), .B(
        f1_round_2_p_io_state_out_0_1), .Z(f1_round_2_io_state_out_0_1) );
  NAND2_X1 f1_round_2_c_U46 ( .A1(f1_round_2_p_io_state_out_2_2), .A2(
        f1_round_2_p_io_state_out_1_2), .ZN(f1_round_2_c_n23) );
  XOR2_X1 f1_round_2_c_U45 ( .A(f1_round_2_c_n23), .B(
        f1_round_2_p_io_state_out_0_2), .Z(f1_round_2_io_state_out_0_2) );
  NAND2_X1 f1_round_2_c_U44 ( .A1(f1_round_2_p_io_state_out_2_3), .A2(
        f1_round_2_p_io_state_out_1_3), .ZN(f1_round_2_c_n22) );
  XOR2_X1 f1_round_2_c_U43 ( .A(f1_round_2_c_n22), .B(
        f1_round_2_p_io_state_out_0_3), .Z(f1_round_2_io_state_out_0_3) );
  NAND2_X1 f1_round_2_c_U42 ( .A1(f1_round_2_p_io_state_out_2_4), .A2(
        f1_round_2_p_io_state_out_1_4), .ZN(f1_round_2_c_n21) );
  XOR2_X1 f1_round_2_c_U41 ( .A(f1_round_2_c_n21), .B(
        f1_round_2_p_io_state_out_0_4), .Z(f1_round_2_io_state_out_0_4) );
  NAND2_X1 f1_round_2_c_U40 ( .A1(f1_round_2_p_io_state_out_2_0), .A2(
        f1_round_2_p_io_state_out_3_0), .ZN(f1_round_2_c_n20) );
  XOR2_X1 f1_round_2_c_U39 ( .A(f1_round_2_c_n20), .B(
        f1_round_2_p_io_state_out_1_0), .Z(f1_round_2_io_state_out_1_0) );
  NAND2_X1 f1_round_2_c_U38 ( .A1(f1_round_2_p_io_state_out_2_1), .A2(
        f1_round_2_p_io_state_out_3_1), .ZN(f1_round_2_c_n19) );
  XOR2_X1 f1_round_2_c_U37 ( .A(f1_round_2_c_n19), .B(
        f1_round_2_p_io_state_out_1_1), .Z(f1_round_2_io_state_out_1_1) );
  NAND2_X1 f1_round_2_c_U36 ( .A1(f1_round_2_p_io_state_out_2_2), .A2(
        f1_round_2_p_io_state_out_3_2), .ZN(f1_round_2_c_n18) );
  XOR2_X1 f1_round_2_c_U35 ( .A(f1_round_2_c_n18), .B(
        f1_round_2_p_io_state_out_1_2), .Z(f1_round_2_io_state_out_1_2) );
  NAND2_X1 f1_round_2_c_U34 ( .A1(f1_round_2_p_io_state_out_2_3), .A2(
        f1_round_2_p_io_state_out_3_3), .ZN(f1_round_2_c_n17) );
  XOR2_X1 f1_round_2_c_U33 ( .A(f1_round_2_c_n17), .B(
        f1_round_2_p_io_state_out_1_3), .Z(f1_round_2_io_state_out_1_3) );
  NAND2_X1 f1_round_2_c_U32 ( .A1(f1_round_2_p_io_state_out_2_4), .A2(
        f1_round_2_p_io_state_out_3_4), .ZN(f1_round_2_c_n16) );
  XOR2_X1 f1_round_2_c_U31 ( .A(f1_round_2_c_n16), .B(
        f1_round_2_p_io_state_out_1_4), .Z(f1_round_2_io_state_out_1_4) );
  NAND2_X1 f1_round_2_c_U30 ( .A1(f1_round_2_p_io_state_out_3_0), .A2(
        f1_round_2_p_io_state_out_4_0), .ZN(f1_round_2_c_n15) );
  XOR2_X1 f1_round_2_c_U29 ( .A(f1_round_2_c_n15), .B(
        f1_round_2_p_io_state_out_2_0), .Z(f1_round_2_io_state_out_2_0) );
  NAND2_X1 f1_round_2_c_U28 ( .A1(f1_round_2_p_io_state_out_3_1), .A2(
        f1_round_2_p_io_state_out_4_1), .ZN(f1_round_2_c_n14) );
  XOR2_X1 f1_round_2_c_U27 ( .A(f1_round_2_c_n14), .B(
        f1_round_2_p_io_state_out_2_1), .Z(f1_round_2_io_state_out_2_1) );
  NAND2_X1 f1_round_2_c_U26 ( .A1(f1_round_2_p_io_state_out_3_2), .A2(
        f1_round_2_p_io_state_out_4_2), .ZN(f1_round_2_c_n13) );
  XOR2_X1 f1_round_2_c_U25 ( .A(f1_round_2_c_n13), .B(
        f1_round_2_p_io_state_out_2_2), .Z(f1_round_2_io_state_out_2_2) );
  NAND2_X1 f1_round_2_c_U24 ( .A1(f1_round_2_p_io_state_out_3_3), .A2(
        f1_round_2_p_io_state_out_4_3), .ZN(f1_round_2_c_n12) );
  XOR2_X1 f1_round_2_c_U23 ( .A(f1_round_2_c_n12), .B(
        f1_round_2_p_io_state_out_2_3), .Z(f1_round_2_io_state_out_2_3) );
  NAND2_X1 f1_round_2_c_U22 ( .A1(f1_round_2_p_io_state_out_3_4), .A2(
        f1_round_2_p_io_state_out_4_4), .ZN(f1_round_2_c_n11) );
  XOR2_X1 f1_round_2_c_U21 ( .A(f1_round_2_c_n11), .B(
        f1_round_2_p_io_state_out_2_4), .Z(f1_round_2_io_state_out_2_4) );
  NAND2_X1 f1_round_2_c_U20 ( .A1(f1_round_2_p_io_state_out_4_0), .A2(
        f1_round_2_p_io_state_out_0_0), .ZN(f1_round_2_c_n10) );
  XOR2_X1 f1_round_2_c_U19 ( .A(f1_round_2_c_n10), .B(
        f1_round_2_p_io_state_out_3_0), .Z(f1_round_2_io_state_out_3_0) );
  NAND2_X1 f1_round_2_c_U18 ( .A1(f1_round_2_p_io_state_out_4_1), .A2(
        f1_round_2_p_io_state_out_0_1), .ZN(f1_round_2_c_n9) );
  XOR2_X1 f1_round_2_c_U17 ( .A(f1_round_2_c_n9), .B(
        f1_round_2_p_io_state_out_3_1), .Z(f1_round_2_io_state_out_3_1) );
  NAND2_X1 f1_round_2_c_U16 ( .A1(f1_round_2_p_io_state_out_4_2), .A2(
        f1_round_2_p_io_state_out_0_2), .ZN(f1_round_2_c_n8) );
  XOR2_X1 f1_round_2_c_U15 ( .A(f1_round_2_c_n8), .B(
        f1_round_2_p_io_state_out_3_2), .Z(f1_round_2_io_state_out_3_2) );
  NAND2_X1 f1_round_2_c_U14 ( .A1(f1_round_2_p_io_state_out_4_3), .A2(
        f1_round_2_p_io_state_out_0_3), .ZN(f1_round_2_c_n7) );
  XOR2_X1 f1_round_2_c_U13 ( .A(f1_round_2_c_n7), .B(
        f1_round_2_p_io_state_out_3_3), .Z(f1_round_2_io_state_out_3_3) );
  NAND2_X1 f1_round_2_c_U12 ( .A1(f1_round_2_p_io_state_out_4_4), .A2(
        f1_round_2_p_io_state_out_0_4), .ZN(f1_round_2_c_n6) );
  XOR2_X1 f1_round_2_c_U11 ( .A(f1_round_2_c_n6), .B(
        f1_round_2_p_io_state_out_3_4), .Z(f1_round_2_io_state_out_3_4) );
  NAND2_X1 f1_round_2_c_U10 ( .A1(f1_round_2_p_io_state_out_1_0), .A2(
        f1_round_2_p_io_state_out_0_0), .ZN(f1_round_2_c_n5) );
  XOR2_X1 f1_round_2_c_U9 ( .A(f1_round_2_c_n5), .B(
        f1_round_2_p_io_state_out_4_0), .Z(f1_round_2_io_state_out_4_0) );
  NAND2_X1 f1_round_2_c_U8 ( .A1(f1_round_2_p_io_state_out_1_1), .A2(
        f1_round_2_p_io_state_out_0_1), .ZN(f1_round_2_c_n4) );
  XOR2_X1 f1_round_2_c_U7 ( .A(f1_round_2_c_n4), .B(
        f1_round_2_p_io_state_out_4_1), .Z(f1_round_2_io_state_out_4_1) );
  NAND2_X1 f1_round_2_c_U6 ( .A1(f1_round_2_p_io_state_out_1_2), .A2(
        f1_round_2_p_io_state_out_0_2), .ZN(f1_round_2_c_n3) );
  XOR2_X1 f1_round_2_c_U5 ( .A(f1_round_2_c_n3), .B(
        f1_round_2_p_io_state_out_4_2), .Z(f1_round_2_io_state_out_4_2) );
  NAND2_X1 f1_round_2_c_U4 ( .A1(f1_round_2_p_io_state_out_1_3), .A2(
        f1_round_2_p_io_state_out_0_3), .ZN(f1_round_2_c_n2) );
  XOR2_X1 f1_round_2_c_U3 ( .A(f1_round_2_c_n2), .B(
        f1_round_2_p_io_state_out_4_3), .Z(f1_round_2_io_state_out_4_3) );
  NAND2_X1 f1_round_2_c_U2 ( .A1(f1_round_2_p_io_state_out_1_4), .A2(
        f1_round_2_p_io_state_out_0_4), .ZN(f1_round_2_c_n1) );
  XOR2_X1 f1_round_2_c_U1 ( .A(f1_round_2_c_n1), .B(
        f1_round_2_p_io_state_out_4_4), .Z(f1_round_2_io_state_out_4_4) );
  XOR2_X1 f1_round_3_t_U50 ( .A(f1_round_2_io_state_out_1_4), .B(
        f1_round_2_io_state_out_1_3), .Z(f1_round_3_t_n25) );
  XNOR2_X1 f1_round_3_t_U49 ( .A(f1_round_2_io_state_out_1_2), .B(
        f1_round_3_t_n25), .ZN(f1_round_3_t_n23) );
  XOR2_X1 f1_round_3_t_U48 ( .A(f1_round_2_io_state_out_1_1), .B(
        f1_round_2_io_state_out_1_0), .Z(f1_round_3_t_n24) );
  XOR2_X1 f1_round_3_t_U47 ( .A(f1_round_3_t_n23), .B(f1_round_3_t_n24), .Z(
        f1_round_3_t_n8) );
  XOR2_X1 f1_round_3_t_U46 ( .A(f1_round_2_io_state_out_4_4), .B(
        f1_round_2_io_state_out_4_3), .Z(f1_round_3_t_n22) );
  XNOR2_X1 f1_round_3_t_U45 ( .A(f1_round_2_io_state_out_4_2), .B(
        f1_round_3_t_n22), .ZN(f1_round_3_t_n20) );
  XOR2_X1 f1_round_3_t_U44 ( .A(f1_round_2_io_state_out_4_1), .B(
        f1_round_2_io_state_out_4_0), .Z(f1_round_3_t_n21) );
  XNOR2_X1 f1_round_3_t_U43 ( .A(f1_round_3_t_n20), .B(f1_round_3_t_n21), .ZN(
        f1_round_3_t_n5) );
  XNOR2_X1 f1_round_3_t_U42 ( .A(f1_round_3_t_n8), .B(f1_round_3_t_n5), .ZN(
        f1_round_3_t_n19) );
  XOR2_X1 f1_round_3_t_U41 ( .A(f1_round_2_io_state_out_0_0), .B(
        f1_round_3_t_n19), .Z(f1_round_3_p_io_state_out_0_0) );
  XOR2_X1 f1_round_3_t_U40 ( .A(f1_round_2_io_state_out_0_1), .B(
        f1_round_3_t_n19), .Z(f1_round_3_p_io_state_out_1_3) );
  XOR2_X1 f1_round_3_t_U39 ( .A(f1_round_2_io_state_out_0_2), .B(
        f1_round_3_t_n19), .Z(f1_round_3_p_io_state_out_2_1) );
  XOR2_X1 f1_round_3_t_U38 ( .A(f1_round_2_io_state_out_0_3), .B(
        f1_round_3_t_n19), .Z(f1_round_3_p_io_state_out_3_4) );
  XOR2_X1 f1_round_3_t_U37 ( .A(f1_round_2_io_state_out_0_4), .B(
        f1_round_3_t_n19), .Z(f1_round_3_p_io_state_out_4_2) );
  XOR2_X1 f1_round_3_t_U36 ( .A(f1_round_2_io_state_out_2_4), .B(
        f1_round_2_io_state_out_2_3), .Z(f1_round_3_t_n18) );
  XNOR2_X1 f1_round_3_t_U35 ( .A(f1_round_2_io_state_out_2_2), .B(
        f1_round_3_t_n18), .ZN(f1_round_3_t_n16) );
  XOR2_X1 f1_round_3_t_U34 ( .A(f1_round_2_io_state_out_2_1), .B(
        f1_round_2_io_state_out_2_0), .Z(f1_round_3_t_n17) );
  XNOR2_X1 f1_round_3_t_U33 ( .A(f1_round_3_t_n16), .B(f1_round_3_t_n17), .ZN(
        f1_round_3_t_n6) );
  XOR2_X1 f1_round_3_t_U32 ( .A(f1_round_2_io_state_out_0_4), .B(
        f1_round_2_io_state_out_0_3), .Z(f1_round_3_t_n15) );
  XNOR2_X1 f1_round_3_t_U31 ( .A(f1_round_2_io_state_out_0_2), .B(
        f1_round_3_t_n15), .ZN(f1_round_3_t_n13) );
  XOR2_X1 f1_round_3_t_U30 ( .A(f1_round_2_io_state_out_0_1), .B(
        f1_round_2_io_state_out_0_0), .Z(f1_round_3_t_n14) );
  XNOR2_X1 f1_round_3_t_U29 ( .A(f1_round_3_t_n13), .B(f1_round_3_t_n14), .ZN(
        f1_round_3_t_n2) );
  XOR2_X1 f1_round_3_t_U28 ( .A(f1_round_3_t_n6), .B(f1_round_3_t_n2), .Z(
        f1_round_3_t_n12) );
  XOR2_X1 f1_round_3_t_U27 ( .A(f1_round_2_io_state_out_1_0), .B(
        f1_round_3_t_n12), .Z(f1_round_3_p_io_state_out_0_2) );
  XOR2_X1 f1_round_3_t_U26 ( .A(f1_round_2_io_state_out_1_1), .B(
        f1_round_3_t_n12), .Z(f1_round_3_p_io_state_out_1_0) );
  XOR2_X1 f1_round_3_t_U25 ( .A(f1_round_2_io_state_out_1_2), .B(
        f1_round_3_t_n12), .Z(f1_round_3_p_io_state_out_2_3) );
  XOR2_X1 f1_round_3_t_U24 ( .A(f1_round_2_io_state_out_1_3), .B(
        f1_round_3_t_n12), .Z(f1_round_3_p_io_state_out_3_1) );
  XOR2_X1 f1_round_3_t_U23 ( .A(f1_round_2_io_state_out_1_4), .B(
        f1_round_3_t_n12), .Z(f1_round_3_p_io_state_out_4_4) );
  XOR2_X1 f1_round_3_t_U22 ( .A(f1_round_2_io_state_out_3_4), .B(
        f1_round_2_io_state_out_3_3), .Z(f1_round_3_t_n11) );
  XNOR2_X1 f1_round_3_t_U21 ( .A(f1_round_2_io_state_out_3_2), .B(
        f1_round_3_t_n11), .ZN(f1_round_3_t_n9) );
  XOR2_X1 f1_round_3_t_U20 ( .A(f1_round_2_io_state_out_3_1), .B(
        f1_round_2_io_state_out_3_0), .Z(f1_round_3_t_n10) );
  XNOR2_X1 f1_round_3_t_U19 ( .A(f1_round_3_t_n9), .B(f1_round_3_t_n10), .ZN(
        f1_round_3_t_n3) );
  XNOR2_X1 f1_round_3_t_U18 ( .A(f1_round_3_t_n8), .B(f1_round_3_t_n3), .ZN(
        f1_round_3_t_n7) );
  XOR2_X1 f1_round_3_t_U17 ( .A(f1_round_2_io_state_out_2_0), .B(
        f1_round_3_t_n7), .Z(f1_round_3_p_io_state_out_0_4) );
  XOR2_X1 f1_round_3_t_U16 ( .A(f1_round_2_io_state_out_2_1), .B(
        f1_round_3_t_n7), .Z(f1_round_3_p_io_state_out_1_2) );
  XOR2_X1 f1_round_3_t_U15 ( .A(f1_round_2_io_state_out_2_2), .B(
        f1_round_3_t_n7), .Z(f1_round_3_p_io_state_out_2_0) );
  XOR2_X1 f1_round_3_t_U14 ( .A(f1_round_2_io_state_out_2_3), .B(
        f1_round_3_t_n7), .Z(f1_round_3_p_io_state_out_3_3) );
  XOR2_X1 f1_round_3_t_U13 ( .A(f1_round_2_io_state_out_2_4), .B(
        f1_round_3_t_n7), .Z(f1_round_3_p_io_state_out_4_1) );
  XOR2_X1 f1_round_3_t_U12 ( .A(f1_round_3_t_n5), .B(f1_round_3_t_n6), .Z(
        f1_round_3_t_n4) );
  XOR2_X1 f1_round_3_t_U11 ( .A(f1_round_2_io_state_out_3_0), .B(
        f1_round_3_t_n4), .Z(f1_round_3_p_io_state_out_0_1) );
  XOR2_X1 f1_round_3_t_U10 ( .A(f1_round_2_io_state_out_3_1), .B(
        f1_round_3_t_n4), .Z(f1_round_3_p_io_state_out_1_4) );
  XOR2_X1 f1_round_3_t_U9 ( .A(f1_round_2_io_state_out_3_2), .B(
        f1_round_3_t_n4), .Z(f1_round_3_p_io_state_out_2_2) );
  XOR2_X1 f1_round_3_t_U8 ( .A(f1_round_2_io_state_out_3_3), .B(
        f1_round_3_t_n4), .Z(f1_round_3_p_io_state_out_3_0) );
  XOR2_X1 f1_round_3_t_U7 ( .A(f1_round_2_io_state_out_3_4), .B(
        f1_round_3_t_n4), .Z(f1_round_3_p_io_state_out_4_3) );
  XOR2_X1 f1_round_3_t_U6 ( .A(f1_round_3_t_n2), .B(f1_round_3_t_n3), .Z(
        f1_round_3_t_n1) );
  XOR2_X1 f1_round_3_t_U5 ( .A(f1_round_2_io_state_out_4_0), .B(
        f1_round_3_t_n1), .Z(f1_round_3_p_io_state_out_0_3) );
  XOR2_X1 f1_round_3_t_U4 ( .A(f1_round_2_io_state_out_4_1), .B(
        f1_round_3_t_n1), .Z(f1_round_3_p_io_state_out_1_1) );
  XOR2_X1 f1_round_3_t_U3 ( .A(f1_round_2_io_state_out_4_2), .B(
        f1_round_3_t_n1), .Z(f1_round_3_p_io_state_out_2_4) );
  XOR2_X1 f1_round_3_t_U2 ( .A(f1_round_2_io_state_out_4_3), .B(
        f1_round_3_t_n1), .Z(f1_round_3_p_io_state_out_3_2) );
  XOR2_X1 f1_round_3_t_U1 ( .A(f1_round_2_io_state_out_4_4), .B(
        f1_round_3_t_n1), .Z(f1_round_3_p_io_state_out_4_0) );
  NAND2_X1 f1_round_3_c_U50 ( .A1(f1_round_3_p_io_state_out_2_0), .A2(
        f1_round_3_p_io_state_out_1_0), .ZN(f1_round_3_c_n25) );
  XOR2_X1 f1_round_3_c_U49 ( .A(f1_round_3_c_n25), .B(
        f1_round_3_p_io_state_out_0_0), .Z(f1_round_3_io_state_out_0_0) );
  NAND2_X1 f1_round_3_c_U48 ( .A1(f1_round_3_p_io_state_out_2_1), .A2(
        f1_round_3_p_io_state_out_1_1), .ZN(f1_round_3_c_n24) );
  XOR2_X1 f1_round_3_c_U47 ( .A(f1_round_3_c_n24), .B(
        f1_round_3_p_io_state_out_0_1), .Z(f1_round_3_io_state_out_0_1) );
  NAND2_X1 f1_round_3_c_U46 ( .A1(f1_round_3_p_io_state_out_2_2), .A2(
        f1_round_3_p_io_state_out_1_2), .ZN(f1_round_3_c_n23) );
  XOR2_X1 f1_round_3_c_U45 ( .A(f1_round_3_c_n23), .B(
        f1_round_3_p_io_state_out_0_2), .Z(f1_round_3_io_state_out_0_2) );
  NAND2_X1 f1_round_3_c_U44 ( .A1(f1_round_3_p_io_state_out_2_3), .A2(
        f1_round_3_p_io_state_out_1_3), .ZN(f1_round_3_c_n22) );
  XOR2_X1 f1_round_3_c_U43 ( .A(f1_round_3_c_n22), .B(
        f1_round_3_p_io_state_out_0_3), .Z(f1_round_3_io_state_out_0_3) );
  NAND2_X1 f1_round_3_c_U42 ( .A1(f1_round_3_p_io_state_out_2_4), .A2(
        f1_round_3_p_io_state_out_1_4), .ZN(f1_round_3_c_n21) );
  XOR2_X1 f1_round_3_c_U41 ( .A(f1_round_3_c_n21), .B(
        f1_round_3_p_io_state_out_0_4), .Z(f1_round_3_io_state_out_0_4) );
  NAND2_X1 f1_round_3_c_U40 ( .A1(f1_round_3_p_io_state_out_2_0), .A2(
        f1_round_3_p_io_state_out_3_0), .ZN(f1_round_3_c_n20) );
  XOR2_X1 f1_round_3_c_U39 ( .A(f1_round_3_c_n20), .B(
        f1_round_3_p_io_state_out_1_0), .Z(f1_round_3_io_state_out_1_0) );
  NAND2_X1 f1_round_3_c_U38 ( .A1(f1_round_3_p_io_state_out_2_1), .A2(
        f1_round_3_p_io_state_out_3_1), .ZN(f1_round_3_c_n19) );
  XOR2_X1 f1_round_3_c_U37 ( .A(f1_round_3_c_n19), .B(
        f1_round_3_p_io_state_out_1_1), .Z(f1_round_3_io_state_out_1_1) );
  NAND2_X1 f1_round_3_c_U36 ( .A1(f1_round_3_p_io_state_out_2_2), .A2(
        f1_round_3_p_io_state_out_3_2), .ZN(f1_round_3_c_n18) );
  XOR2_X1 f1_round_3_c_U35 ( .A(f1_round_3_c_n18), .B(
        f1_round_3_p_io_state_out_1_2), .Z(f1_round_3_io_state_out_1_2) );
  NAND2_X1 f1_round_3_c_U34 ( .A1(f1_round_3_p_io_state_out_2_3), .A2(
        f1_round_3_p_io_state_out_3_3), .ZN(f1_round_3_c_n17) );
  XOR2_X1 f1_round_3_c_U33 ( .A(f1_round_3_c_n17), .B(
        f1_round_3_p_io_state_out_1_3), .Z(f1_round_3_io_state_out_1_3) );
  NAND2_X1 f1_round_3_c_U32 ( .A1(f1_round_3_p_io_state_out_2_4), .A2(
        f1_round_3_p_io_state_out_3_4), .ZN(f1_round_3_c_n16) );
  XOR2_X1 f1_round_3_c_U31 ( .A(f1_round_3_c_n16), .B(
        f1_round_3_p_io_state_out_1_4), .Z(f1_round_3_io_state_out_1_4) );
  NAND2_X1 f1_round_3_c_U30 ( .A1(f1_round_3_p_io_state_out_3_0), .A2(
        f1_round_3_p_io_state_out_4_0), .ZN(f1_round_3_c_n15) );
  XOR2_X1 f1_round_3_c_U29 ( .A(f1_round_3_c_n15), .B(
        f1_round_3_p_io_state_out_2_0), .Z(f1_round_3_io_state_out_2_0) );
  NAND2_X1 f1_round_3_c_U28 ( .A1(f1_round_3_p_io_state_out_3_1), .A2(
        f1_round_3_p_io_state_out_4_1), .ZN(f1_round_3_c_n14) );
  XOR2_X1 f1_round_3_c_U27 ( .A(f1_round_3_c_n14), .B(
        f1_round_3_p_io_state_out_2_1), .Z(f1_round_3_io_state_out_2_1) );
  NAND2_X1 f1_round_3_c_U26 ( .A1(f1_round_3_p_io_state_out_3_2), .A2(
        f1_round_3_p_io_state_out_4_2), .ZN(f1_round_3_c_n13) );
  XOR2_X1 f1_round_3_c_U25 ( .A(f1_round_3_c_n13), .B(
        f1_round_3_p_io_state_out_2_2), .Z(f1_round_3_io_state_out_2_2) );
  NAND2_X1 f1_round_3_c_U24 ( .A1(f1_round_3_p_io_state_out_3_3), .A2(
        f1_round_3_p_io_state_out_4_3), .ZN(f1_round_3_c_n12) );
  XOR2_X1 f1_round_3_c_U23 ( .A(f1_round_3_c_n12), .B(
        f1_round_3_p_io_state_out_2_3), .Z(f1_round_3_io_state_out_2_3) );
  NAND2_X1 f1_round_3_c_U22 ( .A1(f1_round_3_p_io_state_out_3_4), .A2(
        f1_round_3_p_io_state_out_4_4), .ZN(f1_round_3_c_n11) );
  XOR2_X1 f1_round_3_c_U21 ( .A(f1_round_3_c_n11), .B(
        f1_round_3_p_io_state_out_2_4), .Z(f1_round_3_io_state_out_2_4) );
  NAND2_X1 f1_round_3_c_U20 ( .A1(f1_round_3_p_io_state_out_4_0), .A2(
        f1_round_3_p_io_state_out_0_0), .ZN(f1_round_3_c_n10) );
  XOR2_X1 f1_round_3_c_U19 ( .A(f1_round_3_c_n10), .B(
        f1_round_3_p_io_state_out_3_0), .Z(f1_round_3_io_state_out_3_0) );
  NAND2_X1 f1_round_3_c_U18 ( .A1(f1_round_3_p_io_state_out_4_1), .A2(
        f1_round_3_p_io_state_out_0_1), .ZN(f1_round_3_c_n9) );
  XOR2_X1 f1_round_3_c_U17 ( .A(f1_round_3_c_n9), .B(
        f1_round_3_p_io_state_out_3_1), .Z(f1_round_3_io_state_out_3_1) );
  NAND2_X1 f1_round_3_c_U16 ( .A1(f1_round_3_p_io_state_out_4_2), .A2(
        f1_round_3_p_io_state_out_0_2), .ZN(f1_round_3_c_n8) );
  XOR2_X1 f1_round_3_c_U15 ( .A(f1_round_3_c_n8), .B(
        f1_round_3_p_io_state_out_3_2), .Z(f1_round_3_io_state_out_3_2) );
  NAND2_X1 f1_round_3_c_U14 ( .A1(f1_round_3_p_io_state_out_4_3), .A2(
        f1_round_3_p_io_state_out_0_3), .ZN(f1_round_3_c_n7) );
  XOR2_X1 f1_round_3_c_U13 ( .A(f1_round_3_c_n7), .B(
        f1_round_3_p_io_state_out_3_3), .Z(f1_round_3_io_state_out_3_3) );
  NAND2_X1 f1_round_3_c_U12 ( .A1(f1_round_3_p_io_state_out_4_4), .A2(
        f1_round_3_p_io_state_out_0_4), .ZN(f1_round_3_c_n6) );
  XOR2_X1 f1_round_3_c_U11 ( .A(f1_round_3_c_n6), .B(
        f1_round_3_p_io_state_out_3_4), .Z(f1_round_3_io_state_out_3_4) );
  NAND2_X1 f1_round_3_c_U10 ( .A1(f1_round_3_p_io_state_out_1_0), .A2(
        f1_round_3_p_io_state_out_0_0), .ZN(f1_round_3_c_n5) );
  XOR2_X1 f1_round_3_c_U9 ( .A(f1_round_3_c_n5), .B(
        f1_round_3_p_io_state_out_4_0), .Z(f1_round_3_io_state_out_4_0) );
  NAND2_X1 f1_round_3_c_U8 ( .A1(f1_round_3_p_io_state_out_1_1), .A2(
        f1_round_3_p_io_state_out_0_1), .ZN(f1_round_3_c_n4) );
  XOR2_X1 f1_round_3_c_U7 ( .A(f1_round_3_c_n4), .B(
        f1_round_3_p_io_state_out_4_1), .Z(f1_round_3_io_state_out_4_1) );
  NAND2_X1 f1_round_3_c_U6 ( .A1(f1_round_3_p_io_state_out_1_2), .A2(
        f1_round_3_p_io_state_out_0_2), .ZN(f1_round_3_c_n3) );
  XOR2_X1 f1_round_3_c_U5 ( .A(f1_round_3_c_n3), .B(
        f1_round_3_p_io_state_out_4_2), .Z(f1_round_3_io_state_out_4_2) );
  NAND2_X1 f1_round_3_c_U4 ( .A1(f1_round_3_p_io_state_out_1_3), .A2(
        f1_round_3_p_io_state_out_0_3), .ZN(f1_round_3_c_n2) );
  XOR2_X1 f1_round_3_c_U3 ( .A(f1_round_3_c_n2), .B(
        f1_round_3_p_io_state_out_4_3), .Z(f1_round_3_io_state_out_4_3) );
  NAND2_X1 f1_round_3_c_U2 ( .A1(f1_round_3_p_io_state_out_1_4), .A2(
        f1_round_3_p_io_state_out_0_4), .ZN(f1_round_3_c_n1) );
  XOR2_X1 f1_round_3_c_U1 ( .A(f1_round_3_c_n1), .B(
        f1_round_3_p_io_state_out_4_4), .Z(f1_round_3_io_state_out_4_4) );
  XOR2_X1 f1_round_4_t_U50 ( .A(f1_round_3_io_state_out_1_4), .B(
        f1_round_3_io_state_out_1_3), .Z(f1_round_4_t_n25) );
  XNOR2_X1 f1_round_4_t_U49 ( .A(f1_round_3_io_state_out_1_2), .B(
        f1_round_4_t_n25), .ZN(f1_round_4_t_n23) );
  XOR2_X1 f1_round_4_t_U48 ( .A(f1_round_3_io_state_out_1_1), .B(
        f1_round_3_io_state_out_1_0), .Z(f1_round_4_t_n24) );
  XOR2_X1 f1_round_4_t_U47 ( .A(f1_round_4_t_n23), .B(f1_round_4_t_n24), .Z(
        f1_round_4_t_n8) );
  XOR2_X1 f1_round_4_t_U46 ( .A(f1_round_3_io_state_out_4_4), .B(
        f1_round_3_io_state_out_4_3), .Z(f1_round_4_t_n22) );
  XNOR2_X1 f1_round_4_t_U45 ( .A(f1_round_3_io_state_out_4_2), .B(
        f1_round_4_t_n22), .ZN(f1_round_4_t_n20) );
  XOR2_X1 f1_round_4_t_U44 ( .A(f1_round_3_io_state_out_4_1), .B(
        f1_round_3_io_state_out_4_0), .Z(f1_round_4_t_n21) );
  XNOR2_X1 f1_round_4_t_U43 ( .A(f1_round_4_t_n20), .B(f1_round_4_t_n21), .ZN(
        f1_round_4_t_n5) );
  XNOR2_X1 f1_round_4_t_U42 ( .A(f1_round_4_t_n8), .B(f1_round_4_t_n5), .ZN(
        f1_round_4_t_n19) );
  XOR2_X1 f1_round_4_t_U41 ( .A(f1_round_3_io_state_out_0_0), .B(
        f1_round_4_t_n19), .Z(f1_round_4_p_io_state_out_0_0) );
  XOR2_X1 f1_round_4_t_U40 ( .A(f1_round_3_io_state_out_0_1), .B(
        f1_round_4_t_n19), .Z(f1_round_4_p_io_state_out_1_3) );
  XOR2_X1 f1_round_4_t_U39 ( .A(f1_round_3_io_state_out_0_2), .B(
        f1_round_4_t_n19), .Z(f1_round_4_p_io_state_out_2_1) );
  XOR2_X1 f1_round_4_t_U38 ( .A(f1_round_3_io_state_out_0_3), .B(
        f1_round_4_t_n19), .Z(f1_round_4_p_io_state_out_3_4) );
  XOR2_X1 f1_round_4_t_U37 ( .A(f1_round_3_io_state_out_0_4), .B(
        f1_round_4_t_n19), .Z(f1_round_4_p_io_state_out_4_2) );
  XOR2_X1 f1_round_4_t_U36 ( .A(f1_round_3_io_state_out_2_4), .B(
        f1_round_3_io_state_out_2_3), .Z(f1_round_4_t_n18) );
  XNOR2_X1 f1_round_4_t_U35 ( .A(f1_round_3_io_state_out_2_2), .B(
        f1_round_4_t_n18), .ZN(f1_round_4_t_n16) );
  XOR2_X1 f1_round_4_t_U34 ( .A(f1_round_3_io_state_out_2_1), .B(
        f1_round_3_io_state_out_2_0), .Z(f1_round_4_t_n17) );
  XNOR2_X1 f1_round_4_t_U33 ( .A(f1_round_4_t_n16), .B(f1_round_4_t_n17), .ZN(
        f1_round_4_t_n6) );
  XOR2_X1 f1_round_4_t_U32 ( .A(f1_round_3_io_state_out_0_4), .B(
        f1_round_3_io_state_out_0_3), .Z(f1_round_4_t_n15) );
  XNOR2_X1 f1_round_4_t_U31 ( .A(f1_round_3_io_state_out_0_2), .B(
        f1_round_4_t_n15), .ZN(f1_round_4_t_n13) );
  XOR2_X1 f1_round_4_t_U30 ( .A(f1_round_3_io_state_out_0_1), .B(
        f1_round_3_io_state_out_0_0), .Z(f1_round_4_t_n14) );
  XNOR2_X1 f1_round_4_t_U29 ( .A(f1_round_4_t_n13), .B(f1_round_4_t_n14), .ZN(
        f1_round_4_t_n2) );
  XOR2_X1 f1_round_4_t_U28 ( .A(f1_round_4_t_n6), .B(f1_round_4_t_n2), .Z(
        f1_round_4_t_n12) );
  XOR2_X1 f1_round_4_t_U27 ( .A(f1_round_3_io_state_out_1_0), .B(
        f1_round_4_t_n12), .Z(f1_round_4_p_io_state_out_0_2) );
  XOR2_X1 f1_round_4_t_U26 ( .A(f1_round_3_io_state_out_1_1), .B(
        f1_round_4_t_n12), .Z(f1_round_4_p_io_state_out_1_0) );
  XOR2_X1 f1_round_4_t_U25 ( .A(f1_round_3_io_state_out_1_2), .B(
        f1_round_4_t_n12), .Z(f1_round_4_p_io_state_out_2_3) );
  XOR2_X1 f1_round_4_t_U24 ( .A(f1_round_3_io_state_out_1_3), .B(
        f1_round_4_t_n12), .Z(f1_round_4_p_io_state_out_3_1) );
  XOR2_X1 f1_round_4_t_U23 ( .A(f1_round_3_io_state_out_1_4), .B(
        f1_round_4_t_n12), .Z(f1_round_4_p_io_state_out_4_4) );
  XOR2_X1 f1_round_4_t_U22 ( .A(f1_round_3_io_state_out_3_4), .B(
        f1_round_3_io_state_out_3_3), .Z(f1_round_4_t_n11) );
  XNOR2_X1 f1_round_4_t_U21 ( .A(f1_round_3_io_state_out_3_2), .B(
        f1_round_4_t_n11), .ZN(f1_round_4_t_n9) );
  XOR2_X1 f1_round_4_t_U20 ( .A(f1_round_3_io_state_out_3_1), .B(
        f1_round_3_io_state_out_3_0), .Z(f1_round_4_t_n10) );
  XNOR2_X1 f1_round_4_t_U19 ( .A(f1_round_4_t_n9), .B(f1_round_4_t_n10), .ZN(
        f1_round_4_t_n3) );
  XNOR2_X1 f1_round_4_t_U18 ( .A(f1_round_4_t_n8), .B(f1_round_4_t_n3), .ZN(
        f1_round_4_t_n7) );
  XOR2_X1 f1_round_4_t_U17 ( .A(f1_round_3_io_state_out_2_0), .B(
        f1_round_4_t_n7), .Z(f1_round_4_p_io_state_out_0_4) );
  XOR2_X1 f1_round_4_t_U16 ( .A(f1_round_3_io_state_out_2_1), .B(
        f1_round_4_t_n7), .Z(f1_round_4_p_io_state_out_1_2) );
  XOR2_X1 f1_round_4_t_U15 ( .A(f1_round_3_io_state_out_2_2), .B(
        f1_round_4_t_n7), .Z(f1_round_4_p_io_state_out_2_0) );
  XOR2_X1 f1_round_4_t_U14 ( .A(f1_round_3_io_state_out_2_3), .B(
        f1_round_4_t_n7), .Z(f1_round_4_p_io_state_out_3_3) );
  XOR2_X1 f1_round_4_t_U13 ( .A(f1_round_3_io_state_out_2_4), .B(
        f1_round_4_t_n7), .Z(f1_round_4_p_io_state_out_4_1) );
  XOR2_X1 f1_round_4_t_U12 ( .A(f1_round_4_t_n5), .B(f1_round_4_t_n6), .Z(
        f1_round_4_t_n4) );
  XOR2_X1 f1_round_4_t_U11 ( .A(f1_round_3_io_state_out_3_0), .B(
        f1_round_4_t_n4), .Z(f1_round_4_p_io_state_out_0_1) );
  XOR2_X1 f1_round_4_t_U10 ( .A(f1_round_3_io_state_out_3_1), .B(
        f1_round_4_t_n4), .Z(f1_round_4_p_io_state_out_1_4) );
  XOR2_X1 f1_round_4_t_U9 ( .A(f1_round_3_io_state_out_3_2), .B(
        f1_round_4_t_n4), .Z(f1_round_4_p_io_state_out_2_2) );
  XOR2_X1 f1_round_4_t_U8 ( .A(f1_round_3_io_state_out_3_3), .B(
        f1_round_4_t_n4), .Z(f1_round_4_p_io_state_out_3_0) );
  XOR2_X1 f1_round_4_t_U7 ( .A(f1_round_3_io_state_out_3_4), .B(
        f1_round_4_t_n4), .Z(f1_round_4_p_io_state_out_4_3) );
  XOR2_X1 f1_round_4_t_U6 ( .A(f1_round_4_t_n2), .B(f1_round_4_t_n3), .Z(
        f1_round_4_t_n1) );
  XOR2_X1 f1_round_4_t_U5 ( .A(f1_round_3_io_state_out_4_0), .B(
        f1_round_4_t_n1), .Z(f1_round_4_p_io_state_out_0_3) );
  XOR2_X1 f1_round_4_t_U4 ( .A(f1_round_3_io_state_out_4_1), .B(
        f1_round_4_t_n1), .Z(f1_round_4_p_io_state_out_1_1) );
  XOR2_X1 f1_round_4_t_U3 ( .A(f1_round_3_io_state_out_4_2), .B(
        f1_round_4_t_n1), .Z(f1_round_4_p_io_state_out_2_4) );
  XOR2_X1 f1_round_4_t_U2 ( .A(f1_round_3_io_state_out_4_3), .B(
        f1_round_4_t_n1), .Z(f1_round_4_p_io_state_out_3_2) );
  XOR2_X1 f1_round_4_t_U1 ( .A(f1_round_3_io_state_out_4_4), .B(
        f1_round_4_t_n1), .Z(f1_round_4_p_io_state_out_4_0) );
  NAND2_X1 f1_round_4_c_U50 ( .A1(f1_round_4_p_io_state_out_2_0), .A2(
        f1_round_4_p_io_state_out_1_0), .ZN(f1_round_4_c_n25) );
  XOR2_X1 f1_round_4_c_U49 ( .A(f1_round_4_c_n25), .B(
        f1_round_4_p_io_state_out_0_0), .Z(f1_round_4_c_io_state_out_0_0) );
  NAND2_X1 f1_round_4_c_U48 ( .A1(f1_round_4_p_io_state_out_2_1), .A2(
        f1_round_4_p_io_state_out_1_1), .ZN(f1_round_4_c_n24) );
  XOR2_X1 f1_round_4_c_U47 ( .A(f1_round_4_c_n24), .B(
        f1_round_4_p_io_state_out_0_1), .Z(f1_round_4_io_state_out_0_1) );
  NAND2_X1 f1_round_4_c_U46 ( .A1(f1_round_4_p_io_state_out_2_2), .A2(
        f1_round_4_p_io_state_out_1_2), .ZN(f1_round_4_c_n23) );
  XOR2_X1 f1_round_4_c_U45 ( .A(f1_round_4_c_n23), .B(
        f1_round_4_p_io_state_out_0_2), .Z(f1_round_4_io_state_out_0_2) );
  NAND2_X1 f1_round_4_c_U44 ( .A1(f1_round_4_p_io_state_out_2_3), .A2(
        f1_round_4_p_io_state_out_1_3), .ZN(f1_round_4_c_n22) );
  XOR2_X1 f1_round_4_c_U43 ( .A(f1_round_4_c_n22), .B(
        f1_round_4_p_io_state_out_0_3), .Z(f1_round_4_io_state_out_0_3) );
  NAND2_X1 f1_round_4_c_U42 ( .A1(f1_round_4_p_io_state_out_2_4), .A2(
        f1_round_4_p_io_state_out_1_4), .ZN(f1_round_4_c_n21) );
  XOR2_X1 f1_round_4_c_U41 ( .A(f1_round_4_c_n21), .B(
        f1_round_4_p_io_state_out_0_4), .Z(f1_round_4_io_state_out_0_4) );
  NAND2_X1 f1_round_4_c_U40 ( .A1(f1_round_4_p_io_state_out_2_0), .A2(
        f1_round_4_p_io_state_out_3_0), .ZN(f1_round_4_c_n20) );
  XOR2_X1 f1_round_4_c_U39 ( .A(f1_round_4_c_n20), .B(
        f1_round_4_p_io_state_out_1_0), .Z(f1_round_4_io_state_out_1_0) );
  NAND2_X1 f1_round_4_c_U38 ( .A1(f1_round_4_p_io_state_out_2_1), .A2(
        f1_round_4_p_io_state_out_3_1), .ZN(f1_round_4_c_n19) );
  XOR2_X1 f1_round_4_c_U37 ( .A(f1_round_4_c_n19), .B(
        f1_round_4_p_io_state_out_1_1), .Z(f1_round_4_io_state_out_1_1) );
  NAND2_X1 f1_round_4_c_U36 ( .A1(f1_round_4_p_io_state_out_2_2), .A2(
        f1_round_4_p_io_state_out_3_2), .ZN(f1_round_4_c_n18) );
  XOR2_X1 f1_round_4_c_U35 ( .A(f1_round_4_c_n18), .B(
        f1_round_4_p_io_state_out_1_2), .Z(f1_round_4_io_state_out_1_2) );
  NAND2_X1 f1_round_4_c_U34 ( .A1(f1_round_4_p_io_state_out_2_3), .A2(
        f1_round_4_p_io_state_out_3_3), .ZN(f1_round_4_c_n17) );
  XOR2_X1 f1_round_4_c_U33 ( .A(f1_round_4_c_n17), .B(
        f1_round_4_p_io_state_out_1_3), .Z(f1_round_4_io_state_out_1_3) );
  NAND2_X1 f1_round_4_c_U32 ( .A1(f1_round_4_p_io_state_out_2_4), .A2(
        f1_round_4_p_io_state_out_3_4), .ZN(f1_round_4_c_n16) );
  XOR2_X1 f1_round_4_c_U31 ( .A(f1_round_4_c_n16), .B(
        f1_round_4_p_io_state_out_1_4), .Z(f1_round_4_io_state_out_1_4) );
  NAND2_X1 f1_round_4_c_U30 ( .A1(f1_round_4_p_io_state_out_3_0), .A2(
        f1_round_4_p_io_state_out_4_0), .ZN(f1_round_4_c_n15) );
  XOR2_X1 f1_round_4_c_U29 ( .A(f1_round_4_c_n15), .B(
        f1_round_4_p_io_state_out_2_0), .Z(f1_round_4_io_state_out_2_0) );
  NAND2_X1 f1_round_4_c_U28 ( .A1(f1_round_4_p_io_state_out_3_1), .A2(
        f1_round_4_p_io_state_out_4_1), .ZN(f1_round_4_c_n14) );
  XOR2_X1 f1_round_4_c_U27 ( .A(f1_round_4_c_n14), .B(
        f1_round_4_p_io_state_out_2_1), .Z(f1_round_4_io_state_out_2_1) );
  NAND2_X1 f1_round_4_c_U26 ( .A1(f1_round_4_p_io_state_out_3_2), .A2(
        f1_round_4_p_io_state_out_4_2), .ZN(f1_round_4_c_n13) );
  XOR2_X1 f1_round_4_c_U25 ( .A(f1_round_4_c_n13), .B(
        f1_round_4_p_io_state_out_2_2), .Z(f1_round_4_io_state_out_2_2) );
  NAND2_X1 f1_round_4_c_U24 ( .A1(f1_round_4_p_io_state_out_3_3), .A2(
        f1_round_4_p_io_state_out_4_3), .ZN(f1_round_4_c_n12) );
  XOR2_X1 f1_round_4_c_U23 ( .A(f1_round_4_c_n12), .B(
        f1_round_4_p_io_state_out_2_3), .Z(f1_round_4_io_state_out_2_3) );
  NAND2_X1 f1_round_4_c_U22 ( .A1(f1_round_4_p_io_state_out_3_4), .A2(
        f1_round_4_p_io_state_out_4_4), .ZN(f1_round_4_c_n11) );
  XOR2_X1 f1_round_4_c_U21 ( .A(f1_round_4_c_n11), .B(
        f1_round_4_p_io_state_out_2_4), .Z(f1_round_4_io_state_out_2_4) );
  NAND2_X1 f1_round_4_c_U20 ( .A1(f1_round_4_p_io_state_out_4_0), .A2(
        f1_round_4_p_io_state_out_0_0), .ZN(f1_round_4_c_n10) );
  XOR2_X1 f1_round_4_c_U19 ( .A(f1_round_4_c_n10), .B(
        f1_round_4_p_io_state_out_3_0), .Z(f1_round_4_io_state_out_3_0) );
  NAND2_X1 f1_round_4_c_U18 ( .A1(f1_round_4_p_io_state_out_4_1), .A2(
        f1_round_4_p_io_state_out_0_1), .ZN(f1_round_4_c_n9) );
  XOR2_X1 f1_round_4_c_U17 ( .A(f1_round_4_c_n9), .B(
        f1_round_4_p_io_state_out_3_1), .Z(f1_round_4_io_state_out_3_1) );
  NAND2_X1 f1_round_4_c_U16 ( .A1(f1_round_4_p_io_state_out_4_2), .A2(
        f1_round_4_p_io_state_out_0_2), .ZN(f1_round_4_c_n8) );
  XOR2_X1 f1_round_4_c_U15 ( .A(f1_round_4_c_n8), .B(
        f1_round_4_p_io_state_out_3_2), .Z(f1_round_4_io_state_out_3_2) );
  NAND2_X1 f1_round_4_c_U14 ( .A1(f1_round_4_p_io_state_out_4_3), .A2(
        f1_round_4_p_io_state_out_0_3), .ZN(f1_round_4_c_n7) );
  XOR2_X1 f1_round_4_c_U13 ( .A(f1_round_4_c_n7), .B(
        f1_round_4_p_io_state_out_3_3), .Z(f1_round_4_io_state_out_3_3) );
  NAND2_X1 f1_round_4_c_U12 ( .A1(f1_round_4_p_io_state_out_4_4), .A2(
        f1_round_4_p_io_state_out_0_4), .ZN(f1_round_4_c_n6) );
  XOR2_X1 f1_round_4_c_U11 ( .A(f1_round_4_c_n6), .B(
        f1_round_4_p_io_state_out_3_4), .Z(f1_round_4_io_state_out_3_4) );
  NAND2_X1 f1_round_4_c_U10 ( .A1(f1_round_4_p_io_state_out_1_0), .A2(
        f1_round_4_p_io_state_out_0_0), .ZN(f1_round_4_c_n5) );
  XOR2_X1 f1_round_4_c_U9 ( .A(f1_round_4_c_n5), .B(
        f1_round_4_p_io_state_out_4_0), .Z(f1_round_4_io_state_out_4_0) );
  NAND2_X1 f1_round_4_c_U8 ( .A1(f1_round_4_p_io_state_out_1_1), .A2(
        f1_round_4_p_io_state_out_0_1), .ZN(f1_round_4_c_n4) );
  XOR2_X1 f1_round_4_c_U7 ( .A(f1_round_4_c_n4), .B(
        f1_round_4_p_io_state_out_4_1), .Z(f1_round_4_io_state_out_4_1) );
  NAND2_X1 f1_round_4_c_U6 ( .A1(f1_round_4_p_io_state_out_1_2), .A2(
        f1_round_4_p_io_state_out_0_2), .ZN(f1_round_4_c_n3) );
  XOR2_X1 f1_round_4_c_U5 ( .A(f1_round_4_c_n3), .B(
        f1_round_4_p_io_state_out_4_2), .Z(f1_round_4_io_state_out_4_2) );
  NAND2_X1 f1_round_4_c_U4 ( .A1(f1_round_4_p_io_state_out_1_3), .A2(
        f1_round_4_p_io_state_out_0_3), .ZN(f1_round_4_c_n2) );
  XOR2_X1 f1_round_4_c_U3 ( .A(f1_round_4_c_n2), .B(
        f1_round_4_p_io_state_out_4_3), .Z(f1_round_4_io_state_out_4_3) );
  NAND2_X1 f1_round_4_c_U2 ( .A1(f1_round_4_p_io_state_out_1_4), .A2(
        f1_round_4_p_io_state_out_0_4), .ZN(f1_round_4_c_n1) );
  XOR2_X1 f1_round_4_c_U1 ( .A(f1_round_4_c_n1), .B(
        f1_round_4_p_io_state_out_4_4), .Z(f1_round_4_io_state_out_4_4) );
  INV_X1 f1_round_4_i_U1 ( .A(f1_round_4_c_io_state_out_0_0), .ZN(
        f1_round_4_io_state_out_0_0) );
  XOR2_X1 f1_round_5_t_U50 ( .A(f1_round_4_io_state_out_1_4), .B(
        f1_round_4_io_state_out_1_3), .Z(f1_round_5_t_n25) );
  XNOR2_X1 f1_round_5_t_U49 ( .A(f1_round_4_io_state_out_1_2), .B(
        f1_round_5_t_n25), .ZN(f1_round_5_t_n23) );
  XOR2_X1 f1_round_5_t_U48 ( .A(f1_round_4_io_state_out_1_1), .B(
        f1_round_4_io_state_out_1_0), .Z(f1_round_5_t_n24) );
  XOR2_X1 f1_round_5_t_U47 ( .A(f1_round_5_t_n23), .B(f1_round_5_t_n24), .Z(
        f1_round_5_t_n8) );
  XOR2_X1 f1_round_5_t_U46 ( .A(f1_round_4_io_state_out_4_4), .B(
        f1_round_4_io_state_out_4_3), .Z(f1_round_5_t_n22) );
  XNOR2_X1 f1_round_5_t_U45 ( .A(f1_round_4_io_state_out_4_2), .B(
        f1_round_5_t_n22), .ZN(f1_round_5_t_n20) );
  XOR2_X1 f1_round_5_t_U44 ( .A(f1_round_4_io_state_out_4_1), .B(
        f1_round_4_io_state_out_4_0), .Z(f1_round_5_t_n21) );
  XNOR2_X1 f1_round_5_t_U43 ( .A(f1_round_5_t_n20), .B(f1_round_5_t_n21), .ZN(
        f1_round_5_t_n5) );
  XNOR2_X1 f1_round_5_t_U42 ( .A(f1_round_5_t_n8), .B(f1_round_5_t_n5), .ZN(
        f1_round_5_t_n19) );
  XOR2_X1 f1_round_5_t_U41 ( .A(f1_round_4_io_state_out_0_0), .B(
        f1_round_5_t_n19), .Z(f1_round_5_p_io_state_out_0_0) );
  XOR2_X1 f1_round_5_t_U40 ( .A(f1_round_4_io_state_out_0_1), .B(
        f1_round_5_t_n19), .Z(f1_round_5_p_io_state_out_1_3) );
  XOR2_X1 f1_round_5_t_U39 ( .A(f1_round_4_io_state_out_0_2), .B(
        f1_round_5_t_n19), .Z(f1_round_5_p_io_state_out_2_1) );
  XOR2_X1 f1_round_5_t_U38 ( .A(f1_round_4_io_state_out_0_3), .B(
        f1_round_5_t_n19), .Z(f1_round_5_p_io_state_out_3_4) );
  XOR2_X1 f1_round_5_t_U37 ( .A(f1_round_4_io_state_out_0_4), .B(
        f1_round_5_t_n19), .Z(f1_round_5_p_io_state_out_4_2) );
  XOR2_X1 f1_round_5_t_U36 ( .A(f1_round_4_io_state_out_2_4), .B(
        f1_round_4_io_state_out_2_3), .Z(f1_round_5_t_n18) );
  XNOR2_X1 f1_round_5_t_U35 ( .A(f1_round_4_io_state_out_2_2), .B(
        f1_round_5_t_n18), .ZN(f1_round_5_t_n16) );
  XOR2_X1 f1_round_5_t_U34 ( .A(f1_round_4_io_state_out_2_1), .B(
        f1_round_4_io_state_out_2_0), .Z(f1_round_5_t_n17) );
  XNOR2_X1 f1_round_5_t_U33 ( .A(f1_round_5_t_n16), .B(f1_round_5_t_n17), .ZN(
        f1_round_5_t_n6) );
  XOR2_X1 f1_round_5_t_U32 ( .A(f1_round_4_io_state_out_0_4), .B(
        f1_round_4_io_state_out_0_3), .Z(f1_round_5_t_n15) );
  XNOR2_X1 f1_round_5_t_U31 ( .A(f1_round_4_io_state_out_0_2), .B(
        f1_round_5_t_n15), .ZN(f1_round_5_t_n13) );
  XOR2_X1 f1_round_5_t_U30 ( .A(f1_round_4_io_state_out_0_1), .B(
        f1_round_4_io_state_out_0_0), .Z(f1_round_5_t_n14) );
  XNOR2_X1 f1_round_5_t_U29 ( .A(f1_round_5_t_n13), .B(f1_round_5_t_n14), .ZN(
        f1_round_5_t_n2) );
  XOR2_X1 f1_round_5_t_U28 ( .A(f1_round_5_t_n6), .B(f1_round_5_t_n2), .Z(
        f1_round_5_t_n12) );
  XOR2_X1 f1_round_5_t_U27 ( .A(f1_round_4_io_state_out_1_0), .B(
        f1_round_5_t_n12), .Z(f1_round_5_p_io_state_out_0_2) );
  XOR2_X1 f1_round_5_t_U26 ( .A(f1_round_4_io_state_out_1_1), .B(
        f1_round_5_t_n12), .Z(f1_round_5_p_io_state_out_1_0) );
  XOR2_X1 f1_round_5_t_U25 ( .A(f1_round_4_io_state_out_1_2), .B(
        f1_round_5_t_n12), .Z(f1_round_5_p_io_state_out_2_3) );
  XOR2_X1 f1_round_5_t_U24 ( .A(f1_round_4_io_state_out_1_3), .B(
        f1_round_5_t_n12), .Z(f1_round_5_p_io_state_out_3_1) );
  XOR2_X1 f1_round_5_t_U23 ( .A(f1_round_4_io_state_out_1_4), .B(
        f1_round_5_t_n12), .Z(f1_round_5_p_io_state_out_4_4) );
  XOR2_X1 f1_round_5_t_U22 ( .A(f1_round_4_io_state_out_3_4), .B(
        f1_round_4_io_state_out_3_3), .Z(f1_round_5_t_n11) );
  XNOR2_X1 f1_round_5_t_U21 ( .A(f1_round_4_io_state_out_3_2), .B(
        f1_round_5_t_n11), .ZN(f1_round_5_t_n9) );
  XOR2_X1 f1_round_5_t_U20 ( .A(f1_round_4_io_state_out_3_1), .B(
        f1_round_4_io_state_out_3_0), .Z(f1_round_5_t_n10) );
  XNOR2_X1 f1_round_5_t_U19 ( .A(f1_round_5_t_n9), .B(f1_round_5_t_n10), .ZN(
        f1_round_5_t_n3) );
  XNOR2_X1 f1_round_5_t_U18 ( .A(f1_round_5_t_n8), .B(f1_round_5_t_n3), .ZN(
        f1_round_5_t_n7) );
  XOR2_X1 f1_round_5_t_U17 ( .A(f1_round_4_io_state_out_2_0), .B(
        f1_round_5_t_n7), .Z(f1_round_5_p_io_state_out_0_4) );
  XOR2_X1 f1_round_5_t_U16 ( .A(f1_round_4_io_state_out_2_1), .B(
        f1_round_5_t_n7), .Z(f1_round_5_p_io_state_out_1_2) );
  XOR2_X1 f1_round_5_t_U15 ( .A(f1_round_4_io_state_out_2_2), .B(
        f1_round_5_t_n7), .Z(f1_round_5_p_io_state_out_2_0) );
  XOR2_X1 f1_round_5_t_U14 ( .A(f1_round_4_io_state_out_2_3), .B(
        f1_round_5_t_n7), .Z(f1_round_5_p_io_state_out_3_3) );
  XOR2_X1 f1_round_5_t_U13 ( .A(f1_round_4_io_state_out_2_4), .B(
        f1_round_5_t_n7), .Z(f1_round_5_p_io_state_out_4_1) );
  XOR2_X1 f1_round_5_t_U12 ( .A(f1_round_5_t_n5), .B(f1_round_5_t_n6), .Z(
        f1_round_5_t_n4) );
  XOR2_X1 f1_round_5_t_U11 ( .A(f1_round_4_io_state_out_3_0), .B(
        f1_round_5_t_n4), .Z(f1_round_5_p_io_state_out_0_1) );
  XOR2_X1 f1_round_5_t_U10 ( .A(f1_round_4_io_state_out_3_1), .B(
        f1_round_5_t_n4), .Z(f1_round_5_p_io_state_out_1_4) );
  XOR2_X1 f1_round_5_t_U9 ( .A(f1_round_4_io_state_out_3_2), .B(
        f1_round_5_t_n4), .Z(f1_round_5_p_io_state_out_2_2) );
  XOR2_X1 f1_round_5_t_U8 ( .A(f1_round_4_io_state_out_3_3), .B(
        f1_round_5_t_n4), .Z(f1_round_5_p_io_state_out_3_0) );
  XOR2_X1 f1_round_5_t_U7 ( .A(f1_round_4_io_state_out_3_4), .B(
        f1_round_5_t_n4), .Z(f1_round_5_p_io_state_out_4_3) );
  XOR2_X1 f1_round_5_t_U6 ( .A(f1_round_5_t_n2), .B(f1_round_5_t_n3), .Z(
        f1_round_5_t_n1) );
  XOR2_X1 f1_round_5_t_U5 ( .A(f1_round_4_io_state_out_4_0), .B(
        f1_round_5_t_n1), .Z(f1_round_5_p_io_state_out_0_3) );
  XOR2_X1 f1_round_5_t_U4 ( .A(f1_round_4_io_state_out_4_1), .B(
        f1_round_5_t_n1), .Z(f1_round_5_p_io_state_out_1_1) );
  XOR2_X1 f1_round_5_t_U3 ( .A(f1_round_4_io_state_out_4_2), .B(
        f1_round_5_t_n1), .Z(f1_round_5_p_io_state_out_2_4) );
  XOR2_X1 f1_round_5_t_U2 ( .A(f1_round_4_io_state_out_4_3), .B(
        f1_round_5_t_n1), .Z(f1_round_5_p_io_state_out_3_2) );
  XOR2_X1 f1_round_5_t_U1 ( .A(f1_round_4_io_state_out_4_4), .B(
        f1_round_5_t_n1), .Z(f1_round_5_p_io_state_out_4_0) );
  NAND2_X1 f1_round_5_c_U50 ( .A1(f1_round_5_p_io_state_out_2_0), .A2(
        f1_round_5_p_io_state_out_1_0), .ZN(f1_round_5_c_n25) );
  XOR2_X1 f1_round_5_c_U49 ( .A(f1_round_5_c_n25), .B(
        f1_round_5_p_io_state_out_0_0), .Z(f1_round_5_c_io_state_out_0_0) );
  NAND2_X1 f1_round_5_c_U48 ( .A1(f1_round_5_p_io_state_out_2_1), .A2(
        f1_round_5_p_io_state_out_1_1), .ZN(f1_round_5_c_n24) );
  XOR2_X1 f1_round_5_c_U47 ( .A(f1_round_5_c_n24), .B(
        f1_round_5_p_io_state_out_0_1), .Z(f1_round_5_io_state_out_0_1) );
  NAND2_X1 f1_round_5_c_U46 ( .A1(f1_round_5_p_io_state_out_2_2), .A2(
        f1_round_5_p_io_state_out_1_2), .ZN(f1_round_5_c_n23) );
  XOR2_X1 f1_round_5_c_U45 ( .A(f1_round_5_c_n23), .B(
        f1_round_5_p_io_state_out_0_2), .Z(f1_round_5_io_state_out_0_2) );
  NAND2_X1 f1_round_5_c_U44 ( .A1(f1_round_5_p_io_state_out_2_3), .A2(
        f1_round_5_p_io_state_out_1_3), .ZN(f1_round_5_c_n22) );
  XOR2_X1 f1_round_5_c_U43 ( .A(f1_round_5_c_n22), .B(
        f1_round_5_p_io_state_out_0_3), .Z(f1_round_5_io_state_out_0_3) );
  NAND2_X1 f1_round_5_c_U42 ( .A1(f1_round_5_p_io_state_out_2_4), .A2(
        f1_round_5_p_io_state_out_1_4), .ZN(f1_round_5_c_n21) );
  XOR2_X1 f1_round_5_c_U41 ( .A(f1_round_5_c_n21), .B(
        f1_round_5_p_io_state_out_0_4), .Z(f1_round_5_io_state_out_0_4) );
  NAND2_X1 f1_round_5_c_U40 ( .A1(f1_round_5_p_io_state_out_2_0), .A2(
        f1_round_5_p_io_state_out_3_0), .ZN(f1_round_5_c_n20) );
  XOR2_X1 f1_round_5_c_U39 ( .A(f1_round_5_c_n20), .B(
        f1_round_5_p_io_state_out_1_0), .Z(f1_round_5_io_state_out_1_0) );
  NAND2_X1 f1_round_5_c_U38 ( .A1(f1_round_5_p_io_state_out_2_1), .A2(
        f1_round_5_p_io_state_out_3_1), .ZN(f1_round_5_c_n19) );
  XOR2_X1 f1_round_5_c_U37 ( .A(f1_round_5_c_n19), .B(
        f1_round_5_p_io_state_out_1_1), .Z(f1_round_5_io_state_out_1_1) );
  NAND2_X1 f1_round_5_c_U36 ( .A1(f1_round_5_p_io_state_out_2_2), .A2(
        f1_round_5_p_io_state_out_3_2), .ZN(f1_round_5_c_n18) );
  XOR2_X1 f1_round_5_c_U35 ( .A(f1_round_5_c_n18), .B(
        f1_round_5_p_io_state_out_1_2), .Z(f1_round_5_io_state_out_1_2) );
  NAND2_X1 f1_round_5_c_U34 ( .A1(f1_round_5_p_io_state_out_2_3), .A2(
        f1_round_5_p_io_state_out_3_3), .ZN(f1_round_5_c_n17) );
  XOR2_X1 f1_round_5_c_U33 ( .A(f1_round_5_c_n17), .B(
        f1_round_5_p_io_state_out_1_3), .Z(f1_round_5_io_state_out_1_3) );
  NAND2_X1 f1_round_5_c_U32 ( .A1(f1_round_5_p_io_state_out_2_4), .A2(
        f1_round_5_p_io_state_out_3_4), .ZN(f1_round_5_c_n16) );
  XOR2_X1 f1_round_5_c_U31 ( .A(f1_round_5_c_n16), .B(
        f1_round_5_p_io_state_out_1_4), .Z(f1_round_5_io_state_out_1_4) );
  NAND2_X1 f1_round_5_c_U30 ( .A1(f1_round_5_p_io_state_out_3_0), .A2(
        f1_round_5_p_io_state_out_4_0), .ZN(f1_round_5_c_n15) );
  XOR2_X1 f1_round_5_c_U29 ( .A(f1_round_5_c_n15), .B(
        f1_round_5_p_io_state_out_2_0), .Z(f1_round_5_io_state_out_2_0) );
  NAND2_X1 f1_round_5_c_U28 ( .A1(f1_round_5_p_io_state_out_3_1), .A2(
        f1_round_5_p_io_state_out_4_1), .ZN(f1_round_5_c_n14) );
  XOR2_X1 f1_round_5_c_U27 ( .A(f1_round_5_c_n14), .B(
        f1_round_5_p_io_state_out_2_1), .Z(f1_round_5_io_state_out_2_1) );
  NAND2_X1 f1_round_5_c_U26 ( .A1(f1_round_5_p_io_state_out_3_2), .A2(
        f1_round_5_p_io_state_out_4_2), .ZN(f1_round_5_c_n13) );
  XOR2_X1 f1_round_5_c_U25 ( .A(f1_round_5_c_n13), .B(
        f1_round_5_p_io_state_out_2_2), .Z(f1_round_5_io_state_out_2_2) );
  NAND2_X1 f1_round_5_c_U24 ( .A1(f1_round_5_p_io_state_out_3_3), .A2(
        f1_round_5_p_io_state_out_4_3), .ZN(f1_round_5_c_n12) );
  XOR2_X1 f1_round_5_c_U23 ( .A(f1_round_5_c_n12), .B(
        f1_round_5_p_io_state_out_2_3), .Z(f1_round_5_io_state_out_2_3) );
  NAND2_X1 f1_round_5_c_U22 ( .A1(f1_round_5_p_io_state_out_3_4), .A2(
        f1_round_5_p_io_state_out_4_4), .ZN(f1_round_5_c_n11) );
  XOR2_X1 f1_round_5_c_U21 ( .A(f1_round_5_c_n11), .B(
        f1_round_5_p_io_state_out_2_4), .Z(f1_round_5_io_state_out_2_4) );
  NAND2_X1 f1_round_5_c_U20 ( .A1(f1_round_5_p_io_state_out_4_0), .A2(
        f1_round_5_p_io_state_out_0_0), .ZN(f1_round_5_c_n10) );
  XOR2_X1 f1_round_5_c_U19 ( .A(f1_round_5_c_n10), .B(
        f1_round_5_p_io_state_out_3_0), .Z(f1_round_5_io_state_out_3_0) );
  NAND2_X1 f1_round_5_c_U18 ( .A1(f1_round_5_p_io_state_out_4_1), .A2(
        f1_round_5_p_io_state_out_0_1), .ZN(f1_round_5_c_n9) );
  XOR2_X1 f1_round_5_c_U17 ( .A(f1_round_5_c_n9), .B(
        f1_round_5_p_io_state_out_3_1), .Z(f1_round_5_io_state_out_3_1) );
  NAND2_X1 f1_round_5_c_U16 ( .A1(f1_round_5_p_io_state_out_4_2), .A2(
        f1_round_5_p_io_state_out_0_2), .ZN(f1_round_5_c_n8) );
  XOR2_X1 f1_round_5_c_U15 ( .A(f1_round_5_c_n8), .B(
        f1_round_5_p_io_state_out_3_2), .Z(f1_round_5_io_state_out_3_2) );
  NAND2_X1 f1_round_5_c_U14 ( .A1(f1_round_5_p_io_state_out_4_3), .A2(
        f1_round_5_p_io_state_out_0_3), .ZN(f1_round_5_c_n7) );
  XOR2_X1 f1_round_5_c_U13 ( .A(f1_round_5_c_n7), .B(
        f1_round_5_p_io_state_out_3_3), .Z(f1_round_5_io_state_out_3_3) );
  NAND2_X1 f1_round_5_c_U12 ( .A1(f1_round_5_p_io_state_out_4_4), .A2(
        f1_round_5_p_io_state_out_0_4), .ZN(f1_round_5_c_n6) );
  XOR2_X1 f1_round_5_c_U11 ( .A(f1_round_5_c_n6), .B(
        f1_round_5_p_io_state_out_3_4), .Z(f1_round_5_io_state_out_3_4) );
  NAND2_X1 f1_round_5_c_U10 ( .A1(f1_round_5_p_io_state_out_1_0), .A2(
        f1_round_5_p_io_state_out_0_0), .ZN(f1_round_5_c_n5) );
  XOR2_X1 f1_round_5_c_U9 ( .A(f1_round_5_c_n5), .B(
        f1_round_5_p_io_state_out_4_0), .Z(f1_round_5_io_state_out_4_0) );
  NAND2_X1 f1_round_5_c_U8 ( .A1(f1_round_5_p_io_state_out_1_1), .A2(
        f1_round_5_p_io_state_out_0_1), .ZN(f1_round_5_c_n4) );
  XOR2_X1 f1_round_5_c_U7 ( .A(f1_round_5_c_n4), .B(
        f1_round_5_p_io_state_out_4_1), .Z(f1_round_5_io_state_out_4_1) );
  NAND2_X1 f1_round_5_c_U6 ( .A1(f1_round_5_p_io_state_out_1_2), .A2(
        f1_round_5_p_io_state_out_0_2), .ZN(f1_round_5_c_n3) );
  XOR2_X1 f1_round_5_c_U5 ( .A(f1_round_5_c_n3), .B(
        f1_round_5_p_io_state_out_4_2), .Z(f1_round_5_io_state_out_4_2) );
  NAND2_X1 f1_round_5_c_U4 ( .A1(f1_round_5_p_io_state_out_1_3), .A2(
        f1_round_5_p_io_state_out_0_3), .ZN(f1_round_5_c_n2) );
  XOR2_X1 f1_round_5_c_U3 ( .A(f1_round_5_c_n2), .B(
        f1_round_5_p_io_state_out_4_3), .Z(f1_round_5_io_state_out_4_3) );
  NAND2_X1 f1_round_5_c_U2 ( .A1(f1_round_5_p_io_state_out_1_4), .A2(
        f1_round_5_p_io_state_out_0_4), .ZN(f1_round_5_c_n1) );
  XOR2_X1 f1_round_5_c_U1 ( .A(f1_round_5_c_n1), .B(
        f1_round_5_p_io_state_out_4_4), .Z(f1_round_5_io_state_out_4_4) );
  INV_X1 f1_round_5_i_U1 ( .A(f1_round_5_c_io_state_out_0_0), .ZN(
        f1_round_5_io_state_out_0_0) );
  XOR2_X1 f1_round_6_t_U50 ( .A(f1_round_5_io_state_out_1_4), .B(
        f1_round_5_io_state_out_1_3), .Z(f1_round_6_t_n25) );
  XNOR2_X1 f1_round_6_t_U49 ( .A(f1_round_5_io_state_out_1_2), .B(
        f1_round_6_t_n25), .ZN(f1_round_6_t_n23) );
  XOR2_X1 f1_round_6_t_U48 ( .A(f1_round_5_io_state_out_1_1), .B(
        f1_round_5_io_state_out_1_0), .Z(f1_round_6_t_n24) );
  XOR2_X1 f1_round_6_t_U47 ( .A(f1_round_6_t_n23), .B(f1_round_6_t_n24), .Z(
        f1_round_6_t_n8) );
  XOR2_X1 f1_round_6_t_U46 ( .A(f1_round_5_io_state_out_4_4), .B(
        f1_round_5_io_state_out_4_3), .Z(f1_round_6_t_n22) );
  XNOR2_X1 f1_round_6_t_U45 ( .A(f1_round_5_io_state_out_4_2), .B(
        f1_round_6_t_n22), .ZN(f1_round_6_t_n20) );
  XOR2_X1 f1_round_6_t_U44 ( .A(f1_round_5_io_state_out_4_1), .B(
        f1_round_5_io_state_out_4_0), .Z(f1_round_6_t_n21) );
  XNOR2_X1 f1_round_6_t_U43 ( .A(f1_round_6_t_n20), .B(f1_round_6_t_n21), .ZN(
        f1_round_6_t_n5) );
  XNOR2_X1 f1_round_6_t_U42 ( .A(f1_round_6_t_n8), .B(f1_round_6_t_n5), .ZN(
        f1_round_6_t_n19) );
  XOR2_X1 f1_round_6_t_U41 ( .A(f1_round_5_io_state_out_0_0), .B(
        f1_round_6_t_n19), .Z(f1_round_6_p_io_state_out_0_0) );
  XOR2_X1 f1_round_6_t_U40 ( .A(f1_round_5_io_state_out_0_1), .B(
        f1_round_6_t_n19), .Z(f1_round_6_p_io_state_out_1_3) );
  XOR2_X1 f1_round_6_t_U39 ( .A(f1_round_5_io_state_out_0_2), .B(
        f1_round_6_t_n19), .Z(f1_round_6_p_io_state_out_2_1) );
  XOR2_X1 f1_round_6_t_U38 ( .A(f1_round_5_io_state_out_0_3), .B(
        f1_round_6_t_n19), .Z(f1_round_6_p_io_state_out_3_4) );
  XOR2_X1 f1_round_6_t_U37 ( .A(f1_round_5_io_state_out_0_4), .B(
        f1_round_6_t_n19), .Z(f1_round_6_p_io_state_out_4_2) );
  XOR2_X1 f1_round_6_t_U36 ( .A(f1_round_5_io_state_out_2_4), .B(
        f1_round_5_io_state_out_2_3), .Z(f1_round_6_t_n18) );
  XNOR2_X1 f1_round_6_t_U35 ( .A(f1_round_5_io_state_out_2_2), .B(
        f1_round_6_t_n18), .ZN(f1_round_6_t_n16) );
  XOR2_X1 f1_round_6_t_U34 ( .A(f1_round_5_io_state_out_2_1), .B(
        f1_round_5_io_state_out_2_0), .Z(f1_round_6_t_n17) );
  XNOR2_X1 f1_round_6_t_U33 ( .A(f1_round_6_t_n16), .B(f1_round_6_t_n17), .ZN(
        f1_round_6_t_n6) );
  XOR2_X1 f1_round_6_t_U32 ( .A(f1_round_5_io_state_out_0_4), .B(
        f1_round_5_io_state_out_0_3), .Z(f1_round_6_t_n15) );
  XNOR2_X1 f1_round_6_t_U31 ( .A(f1_round_5_io_state_out_0_2), .B(
        f1_round_6_t_n15), .ZN(f1_round_6_t_n13) );
  XOR2_X1 f1_round_6_t_U30 ( .A(f1_round_5_io_state_out_0_1), .B(
        f1_round_5_io_state_out_0_0), .Z(f1_round_6_t_n14) );
  XNOR2_X1 f1_round_6_t_U29 ( .A(f1_round_6_t_n13), .B(f1_round_6_t_n14), .ZN(
        f1_round_6_t_n2) );
  XOR2_X1 f1_round_6_t_U28 ( .A(f1_round_6_t_n6), .B(f1_round_6_t_n2), .Z(
        f1_round_6_t_n12) );
  XOR2_X1 f1_round_6_t_U27 ( .A(f1_round_5_io_state_out_1_0), .B(
        f1_round_6_t_n12), .Z(f1_round_6_p_io_state_out_0_2) );
  XOR2_X1 f1_round_6_t_U26 ( .A(f1_round_5_io_state_out_1_1), .B(
        f1_round_6_t_n12), .Z(f1_round_6_p_io_state_out_1_0) );
  XOR2_X1 f1_round_6_t_U25 ( .A(f1_round_5_io_state_out_1_2), .B(
        f1_round_6_t_n12), .Z(f1_round_6_p_io_state_out_2_3) );
  XOR2_X1 f1_round_6_t_U24 ( .A(f1_round_5_io_state_out_1_3), .B(
        f1_round_6_t_n12), .Z(f1_round_6_p_io_state_out_3_1) );
  XOR2_X1 f1_round_6_t_U23 ( .A(f1_round_5_io_state_out_1_4), .B(
        f1_round_6_t_n12), .Z(f1_round_6_p_io_state_out_4_4) );
  XOR2_X1 f1_round_6_t_U22 ( .A(f1_round_5_io_state_out_3_4), .B(
        f1_round_5_io_state_out_3_3), .Z(f1_round_6_t_n11) );
  XNOR2_X1 f1_round_6_t_U21 ( .A(f1_round_5_io_state_out_3_2), .B(
        f1_round_6_t_n11), .ZN(f1_round_6_t_n9) );
  XOR2_X1 f1_round_6_t_U20 ( .A(f1_round_5_io_state_out_3_1), .B(
        f1_round_5_io_state_out_3_0), .Z(f1_round_6_t_n10) );
  XNOR2_X1 f1_round_6_t_U19 ( .A(f1_round_6_t_n9), .B(f1_round_6_t_n10), .ZN(
        f1_round_6_t_n3) );
  XNOR2_X1 f1_round_6_t_U18 ( .A(f1_round_6_t_n8), .B(f1_round_6_t_n3), .ZN(
        f1_round_6_t_n7) );
  XOR2_X1 f1_round_6_t_U17 ( .A(f1_round_5_io_state_out_2_0), .B(
        f1_round_6_t_n7), .Z(f1_round_6_p_io_state_out_0_4) );
  XOR2_X1 f1_round_6_t_U16 ( .A(f1_round_5_io_state_out_2_1), .B(
        f1_round_6_t_n7), .Z(f1_round_6_p_io_state_out_1_2) );
  XOR2_X1 f1_round_6_t_U15 ( .A(f1_round_5_io_state_out_2_2), .B(
        f1_round_6_t_n7), .Z(f1_round_6_p_io_state_out_2_0) );
  XOR2_X1 f1_round_6_t_U14 ( .A(f1_round_5_io_state_out_2_3), .B(
        f1_round_6_t_n7), .Z(f1_round_6_p_io_state_out_3_3) );
  XOR2_X1 f1_round_6_t_U13 ( .A(f1_round_5_io_state_out_2_4), .B(
        f1_round_6_t_n7), .Z(f1_round_6_p_io_state_out_4_1) );
  XOR2_X1 f1_round_6_t_U12 ( .A(f1_round_6_t_n5), .B(f1_round_6_t_n6), .Z(
        f1_round_6_t_n4) );
  XOR2_X1 f1_round_6_t_U11 ( .A(f1_round_5_io_state_out_3_0), .B(
        f1_round_6_t_n4), .Z(f1_round_6_p_io_state_out_0_1) );
  XOR2_X1 f1_round_6_t_U10 ( .A(f1_round_5_io_state_out_3_1), .B(
        f1_round_6_t_n4), .Z(f1_round_6_p_io_state_out_1_4) );
  XOR2_X1 f1_round_6_t_U9 ( .A(f1_round_5_io_state_out_3_2), .B(
        f1_round_6_t_n4), .Z(f1_round_6_p_io_state_out_2_2) );
  XOR2_X1 f1_round_6_t_U8 ( .A(f1_round_5_io_state_out_3_3), .B(
        f1_round_6_t_n4), .Z(f1_round_6_p_io_state_out_3_0) );
  XOR2_X1 f1_round_6_t_U7 ( .A(f1_round_5_io_state_out_3_4), .B(
        f1_round_6_t_n4), .Z(f1_round_6_p_io_state_out_4_3) );
  XOR2_X1 f1_round_6_t_U6 ( .A(f1_round_6_t_n2), .B(f1_round_6_t_n3), .Z(
        f1_round_6_t_n1) );
  XOR2_X1 f1_round_6_t_U5 ( .A(f1_round_5_io_state_out_4_0), .B(
        f1_round_6_t_n1), .Z(f1_round_6_p_io_state_out_0_3) );
  XOR2_X1 f1_round_6_t_U4 ( .A(f1_round_5_io_state_out_4_1), .B(
        f1_round_6_t_n1), .Z(f1_round_6_p_io_state_out_1_1) );
  XOR2_X1 f1_round_6_t_U3 ( .A(f1_round_5_io_state_out_4_2), .B(
        f1_round_6_t_n1), .Z(f1_round_6_p_io_state_out_2_4) );
  XOR2_X1 f1_round_6_t_U2 ( .A(f1_round_5_io_state_out_4_3), .B(
        f1_round_6_t_n1), .Z(f1_round_6_p_io_state_out_3_2) );
  XOR2_X1 f1_round_6_t_U1 ( .A(f1_round_5_io_state_out_4_4), .B(
        f1_round_6_t_n1), .Z(f1_round_6_p_io_state_out_4_0) );
  NAND2_X1 f1_round_6_c_U50 ( .A1(f1_round_6_p_io_state_out_2_0), .A2(
        f1_round_6_p_io_state_out_1_0), .ZN(f1_round_6_c_n25) );
  XOR2_X1 f1_round_6_c_U49 ( .A(f1_round_6_c_n25), .B(
        f1_round_6_p_io_state_out_0_0), .Z(f1_round_6_c_io_state_out_0_0) );
  NAND2_X1 f1_round_6_c_U48 ( .A1(f1_round_6_p_io_state_out_2_1), .A2(
        f1_round_6_p_io_state_out_1_1), .ZN(f1_round_6_c_n24) );
  XOR2_X1 f1_round_6_c_U47 ( .A(f1_round_6_c_n24), .B(
        f1_round_6_p_io_state_out_0_1), .Z(f1_round_6_io_state_out_0_1) );
  NAND2_X1 f1_round_6_c_U46 ( .A1(f1_round_6_p_io_state_out_2_2), .A2(
        f1_round_6_p_io_state_out_1_2), .ZN(f1_round_6_c_n23) );
  XOR2_X1 f1_round_6_c_U45 ( .A(f1_round_6_c_n23), .B(
        f1_round_6_p_io_state_out_0_2), .Z(f1_round_6_io_state_out_0_2) );
  NAND2_X1 f1_round_6_c_U44 ( .A1(f1_round_6_p_io_state_out_2_3), .A2(
        f1_round_6_p_io_state_out_1_3), .ZN(f1_round_6_c_n22) );
  XOR2_X1 f1_round_6_c_U43 ( .A(f1_round_6_c_n22), .B(
        f1_round_6_p_io_state_out_0_3), .Z(f1_round_6_io_state_out_0_3) );
  NAND2_X1 f1_round_6_c_U42 ( .A1(f1_round_6_p_io_state_out_2_4), .A2(
        f1_round_6_p_io_state_out_1_4), .ZN(f1_round_6_c_n21) );
  XOR2_X1 f1_round_6_c_U41 ( .A(f1_round_6_c_n21), .B(
        f1_round_6_p_io_state_out_0_4), .Z(f1_round_6_io_state_out_0_4) );
  NAND2_X1 f1_round_6_c_U40 ( .A1(f1_round_6_p_io_state_out_2_0), .A2(
        f1_round_6_p_io_state_out_3_0), .ZN(f1_round_6_c_n20) );
  XOR2_X1 f1_round_6_c_U39 ( .A(f1_round_6_c_n20), .B(
        f1_round_6_p_io_state_out_1_0), .Z(f1_round_6_io_state_out_1_0) );
  NAND2_X1 f1_round_6_c_U38 ( .A1(f1_round_6_p_io_state_out_2_1), .A2(
        f1_round_6_p_io_state_out_3_1), .ZN(f1_round_6_c_n19) );
  XOR2_X1 f1_round_6_c_U37 ( .A(f1_round_6_c_n19), .B(
        f1_round_6_p_io_state_out_1_1), .Z(f1_round_6_io_state_out_1_1) );
  NAND2_X1 f1_round_6_c_U36 ( .A1(f1_round_6_p_io_state_out_2_2), .A2(
        f1_round_6_p_io_state_out_3_2), .ZN(f1_round_6_c_n18) );
  XOR2_X1 f1_round_6_c_U35 ( .A(f1_round_6_c_n18), .B(
        f1_round_6_p_io_state_out_1_2), .Z(f1_round_6_io_state_out_1_2) );
  NAND2_X1 f1_round_6_c_U34 ( .A1(f1_round_6_p_io_state_out_2_3), .A2(
        f1_round_6_p_io_state_out_3_3), .ZN(f1_round_6_c_n17) );
  XOR2_X1 f1_round_6_c_U33 ( .A(f1_round_6_c_n17), .B(
        f1_round_6_p_io_state_out_1_3), .Z(f1_round_6_io_state_out_1_3) );
  NAND2_X1 f1_round_6_c_U32 ( .A1(f1_round_6_p_io_state_out_2_4), .A2(
        f1_round_6_p_io_state_out_3_4), .ZN(f1_round_6_c_n16) );
  XOR2_X1 f1_round_6_c_U31 ( .A(f1_round_6_c_n16), .B(
        f1_round_6_p_io_state_out_1_4), .Z(f1_round_6_io_state_out_1_4) );
  NAND2_X1 f1_round_6_c_U30 ( .A1(f1_round_6_p_io_state_out_3_0), .A2(
        f1_round_6_p_io_state_out_4_0), .ZN(f1_round_6_c_n15) );
  XOR2_X1 f1_round_6_c_U29 ( .A(f1_round_6_c_n15), .B(
        f1_round_6_p_io_state_out_2_0), .Z(f1_round_6_io_state_out_2_0) );
  NAND2_X1 f1_round_6_c_U28 ( .A1(f1_round_6_p_io_state_out_3_1), .A2(
        f1_round_6_p_io_state_out_4_1), .ZN(f1_round_6_c_n14) );
  XOR2_X1 f1_round_6_c_U27 ( .A(f1_round_6_c_n14), .B(
        f1_round_6_p_io_state_out_2_1), .Z(f1_round_6_io_state_out_2_1) );
  NAND2_X1 f1_round_6_c_U26 ( .A1(f1_round_6_p_io_state_out_3_2), .A2(
        f1_round_6_p_io_state_out_4_2), .ZN(f1_round_6_c_n13) );
  XOR2_X1 f1_round_6_c_U25 ( .A(f1_round_6_c_n13), .B(
        f1_round_6_p_io_state_out_2_2), .Z(f1_round_6_io_state_out_2_2) );
  NAND2_X1 f1_round_6_c_U24 ( .A1(f1_round_6_p_io_state_out_3_3), .A2(
        f1_round_6_p_io_state_out_4_3), .ZN(f1_round_6_c_n12) );
  XOR2_X1 f1_round_6_c_U23 ( .A(f1_round_6_c_n12), .B(
        f1_round_6_p_io_state_out_2_3), .Z(f1_round_6_io_state_out_2_3) );
  NAND2_X1 f1_round_6_c_U22 ( .A1(f1_round_6_p_io_state_out_3_4), .A2(
        f1_round_6_p_io_state_out_4_4), .ZN(f1_round_6_c_n11) );
  XOR2_X1 f1_round_6_c_U21 ( .A(f1_round_6_c_n11), .B(
        f1_round_6_p_io_state_out_2_4), .Z(f1_round_6_io_state_out_2_4) );
  NAND2_X1 f1_round_6_c_U20 ( .A1(f1_round_6_p_io_state_out_4_0), .A2(
        f1_round_6_p_io_state_out_0_0), .ZN(f1_round_6_c_n10) );
  XOR2_X1 f1_round_6_c_U19 ( .A(f1_round_6_c_n10), .B(
        f1_round_6_p_io_state_out_3_0), .Z(f1_round_6_io_state_out_3_0) );
  NAND2_X1 f1_round_6_c_U18 ( .A1(f1_round_6_p_io_state_out_4_1), .A2(
        f1_round_6_p_io_state_out_0_1), .ZN(f1_round_6_c_n9) );
  XOR2_X1 f1_round_6_c_U17 ( .A(f1_round_6_c_n9), .B(
        f1_round_6_p_io_state_out_3_1), .Z(f1_round_6_io_state_out_3_1) );
  NAND2_X1 f1_round_6_c_U16 ( .A1(f1_round_6_p_io_state_out_4_2), .A2(
        f1_round_6_p_io_state_out_0_2), .ZN(f1_round_6_c_n8) );
  XOR2_X1 f1_round_6_c_U15 ( .A(f1_round_6_c_n8), .B(
        f1_round_6_p_io_state_out_3_2), .Z(f1_round_6_io_state_out_3_2) );
  NAND2_X1 f1_round_6_c_U14 ( .A1(f1_round_6_p_io_state_out_4_3), .A2(
        f1_round_6_p_io_state_out_0_3), .ZN(f1_round_6_c_n7) );
  XOR2_X1 f1_round_6_c_U13 ( .A(f1_round_6_c_n7), .B(
        f1_round_6_p_io_state_out_3_3), .Z(f1_round_6_io_state_out_3_3) );
  NAND2_X1 f1_round_6_c_U12 ( .A1(f1_round_6_p_io_state_out_4_4), .A2(
        f1_round_6_p_io_state_out_0_4), .ZN(f1_round_6_c_n6) );
  XOR2_X1 f1_round_6_c_U11 ( .A(f1_round_6_c_n6), .B(
        f1_round_6_p_io_state_out_3_4), .Z(f1_round_6_io_state_out_3_4) );
  NAND2_X1 f1_round_6_c_U10 ( .A1(f1_round_6_p_io_state_out_1_0), .A2(
        f1_round_6_p_io_state_out_0_0), .ZN(f1_round_6_c_n5) );
  XOR2_X1 f1_round_6_c_U9 ( .A(f1_round_6_c_n5), .B(
        f1_round_6_p_io_state_out_4_0), .Z(f1_round_6_io_state_out_4_0) );
  NAND2_X1 f1_round_6_c_U8 ( .A1(f1_round_6_p_io_state_out_1_1), .A2(
        f1_round_6_p_io_state_out_0_1), .ZN(f1_round_6_c_n4) );
  XOR2_X1 f1_round_6_c_U7 ( .A(f1_round_6_c_n4), .B(
        f1_round_6_p_io_state_out_4_1), .Z(f1_round_6_io_state_out_4_1) );
  NAND2_X1 f1_round_6_c_U6 ( .A1(f1_round_6_p_io_state_out_1_2), .A2(
        f1_round_6_p_io_state_out_0_2), .ZN(f1_round_6_c_n3) );
  XOR2_X1 f1_round_6_c_U5 ( .A(f1_round_6_c_n3), .B(
        f1_round_6_p_io_state_out_4_2), .Z(f1_round_6_io_state_out_4_2) );
  NAND2_X1 f1_round_6_c_U4 ( .A1(f1_round_6_p_io_state_out_1_3), .A2(
        f1_round_6_p_io_state_out_0_3), .ZN(f1_round_6_c_n2) );
  XOR2_X1 f1_round_6_c_U3 ( .A(f1_round_6_c_n2), .B(
        f1_round_6_p_io_state_out_4_3), .Z(f1_round_6_io_state_out_4_3) );
  NAND2_X1 f1_round_6_c_U2 ( .A1(f1_round_6_p_io_state_out_1_4), .A2(
        f1_round_6_p_io_state_out_0_4), .ZN(f1_round_6_c_n1) );
  XOR2_X1 f1_round_6_c_U1 ( .A(f1_round_6_c_n1), .B(
        f1_round_6_p_io_state_out_4_4), .Z(f1_round_6_io_state_out_4_4) );
  INV_X1 f1_round_6_i_U1 ( .A(f1_round_6_c_io_state_out_0_0), .ZN(
        f1_round_6_io_state_out_0_0) );
  XOR2_X1 f1_round_7_t_U50 ( .A(f1_round_6_io_state_out_1_4), .B(
        f1_round_6_io_state_out_1_3), .Z(f1_round_7_t_n25) );
  XNOR2_X1 f1_round_7_t_U49 ( .A(f1_round_6_io_state_out_1_2), .B(
        f1_round_7_t_n25), .ZN(f1_round_7_t_n23) );
  XOR2_X1 f1_round_7_t_U48 ( .A(f1_round_6_io_state_out_1_1), .B(
        f1_round_6_io_state_out_1_0), .Z(f1_round_7_t_n24) );
  XOR2_X1 f1_round_7_t_U47 ( .A(f1_round_7_t_n23), .B(f1_round_7_t_n24), .Z(
        f1_round_7_t_n8) );
  XOR2_X1 f1_round_7_t_U46 ( .A(f1_round_6_io_state_out_4_4), .B(
        f1_round_6_io_state_out_4_3), .Z(f1_round_7_t_n22) );
  XNOR2_X1 f1_round_7_t_U45 ( .A(f1_round_6_io_state_out_4_2), .B(
        f1_round_7_t_n22), .ZN(f1_round_7_t_n20) );
  XOR2_X1 f1_round_7_t_U44 ( .A(f1_round_6_io_state_out_4_1), .B(
        f1_round_6_io_state_out_4_0), .Z(f1_round_7_t_n21) );
  XNOR2_X1 f1_round_7_t_U43 ( .A(f1_round_7_t_n20), .B(f1_round_7_t_n21), .ZN(
        f1_round_7_t_n5) );
  XNOR2_X1 f1_round_7_t_U42 ( .A(f1_round_7_t_n8), .B(f1_round_7_t_n5), .ZN(
        f1_round_7_t_n19) );
  XOR2_X1 f1_round_7_t_U41 ( .A(f1_round_6_io_state_out_0_0), .B(
        f1_round_7_t_n19), .Z(f1_round_7_p_io_state_out_0_0) );
  XOR2_X1 f1_round_7_t_U40 ( .A(f1_round_6_io_state_out_0_1), .B(
        f1_round_7_t_n19), .Z(f1_round_7_p_io_state_out_1_3) );
  XOR2_X1 f1_round_7_t_U39 ( .A(f1_round_6_io_state_out_0_2), .B(
        f1_round_7_t_n19), .Z(f1_round_7_p_io_state_out_2_1) );
  XOR2_X1 f1_round_7_t_U38 ( .A(f1_round_6_io_state_out_0_3), .B(
        f1_round_7_t_n19), .Z(f1_round_7_p_io_state_out_3_4) );
  XOR2_X1 f1_round_7_t_U37 ( .A(f1_round_6_io_state_out_0_4), .B(
        f1_round_7_t_n19), .Z(f1_round_7_p_io_state_out_4_2) );
  XOR2_X1 f1_round_7_t_U36 ( .A(f1_round_6_io_state_out_2_4), .B(
        f1_round_6_io_state_out_2_3), .Z(f1_round_7_t_n18) );
  XNOR2_X1 f1_round_7_t_U35 ( .A(f1_round_6_io_state_out_2_2), .B(
        f1_round_7_t_n18), .ZN(f1_round_7_t_n16) );
  XOR2_X1 f1_round_7_t_U34 ( .A(f1_round_6_io_state_out_2_1), .B(
        f1_round_6_io_state_out_2_0), .Z(f1_round_7_t_n17) );
  XNOR2_X1 f1_round_7_t_U33 ( .A(f1_round_7_t_n16), .B(f1_round_7_t_n17), .ZN(
        f1_round_7_t_n6) );
  XOR2_X1 f1_round_7_t_U32 ( .A(f1_round_6_io_state_out_0_4), .B(
        f1_round_6_io_state_out_0_3), .Z(f1_round_7_t_n15) );
  XNOR2_X1 f1_round_7_t_U31 ( .A(f1_round_6_io_state_out_0_2), .B(
        f1_round_7_t_n15), .ZN(f1_round_7_t_n13) );
  XOR2_X1 f1_round_7_t_U30 ( .A(f1_round_6_io_state_out_0_1), .B(
        f1_round_6_io_state_out_0_0), .Z(f1_round_7_t_n14) );
  XNOR2_X1 f1_round_7_t_U29 ( .A(f1_round_7_t_n13), .B(f1_round_7_t_n14), .ZN(
        f1_round_7_t_n2) );
  XOR2_X1 f1_round_7_t_U28 ( .A(f1_round_7_t_n6), .B(f1_round_7_t_n2), .Z(
        f1_round_7_t_n12) );
  XOR2_X1 f1_round_7_t_U27 ( .A(f1_round_6_io_state_out_1_0), .B(
        f1_round_7_t_n12), .Z(f1_round_7_p_io_state_out_0_2) );
  XOR2_X1 f1_round_7_t_U26 ( .A(f1_round_6_io_state_out_1_1), .B(
        f1_round_7_t_n12), .Z(f1_round_7_p_io_state_out_1_0) );
  XOR2_X1 f1_round_7_t_U25 ( .A(f1_round_6_io_state_out_1_2), .B(
        f1_round_7_t_n12), .Z(f1_round_7_p_io_state_out_2_3) );
  XOR2_X1 f1_round_7_t_U24 ( .A(f1_round_6_io_state_out_1_3), .B(
        f1_round_7_t_n12), .Z(f1_round_7_p_io_state_out_3_1) );
  XOR2_X1 f1_round_7_t_U23 ( .A(f1_round_6_io_state_out_1_4), .B(
        f1_round_7_t_n12), .Z(f1_round_7_p_io_state_out_4_4) );
  XOR2_X1 f1_round_7_t_U22 ( .A(f1_round_6_io_state_out_3_4), .B(
        f1_round_6_io_state_out_3_3), .Z(f1_round_7_t_n11) );
  XNOR2_X1 f1_round_7_t_U21 ( .A(f1_round_6_io_state_out_3_2), .B(
        f1_round_7_t_n11), .ZN(f1_round_7_t_n9) );
  XOR2_X1 f1_round_7_t_U20 ( .A(f1_round_6_io_state_out_3_1), .B(
        f1_round_6_io_state_out_3_0), .Z(f1_round_7_t_n10) );
  XNOR2_X1 f1_round_7_t_U19 ( .A(f1_round_7_t_n9), .B(f1_round_7_t_n10), .ZN(
        f1_round_7_t_n3) );
  XNOR2_X1 f1_round_7_t_U18 ( .A(f1_round_7_t_n8), .B(f1_round_7_t_n3), .ZN(
        f1_round_7_t_n7) );
  XOR2_X1 f1_round_7_t_U17 ( .A(f1_round_6_io_state_out_2_0), .B(
        f1_round_7_t_n7), .Z(f1_round_7_p_io_state_out_0_4) );
  XOR2_X1 f1_round_7_t_U16 ( .A(f1_round_6_io_state_out_2_1), .B(
        f1_round_7_t_n7), .Z(f1_round_7_p_io_state_out_1_2) );
  XOR2_X1 f1_round_7_t_U15 ( .A(f1_round_6_io_state_out_2_2), .B(
        f1_round_7_t_n7), .Z(f1_round_7_p_io_state_out_2_0) );
  XOR2_X1 f1_round_7_t_U14 ( .A(f1_round_6_io_state_out_2_3), .B(
        f1_round_7_t_n7), .Z(f1_round_7_p_io_state_out_3_3) );
  XOR2_X1 f1_round_7_t_U13 ( .A(f1_round_6_io_state_out_2_4), .B(
        f1_round_7_t_n7), .Z(f1_round_7_p_io_state_out_4_1) );
  XOR2_X1 f1_round_7_t_U12 ( .A(f1_round_7_t_n5), .B(f1_round_7_t_n6), .Z(
        f1_round_7_t_n4) );
  XOR2_X1 f1_round_7_t_U11 ( .A(f1_round_6_io_state_out_3_0), .B(
        f1_round_7_t_n4), .Z(f1_round_7_p_io_state_out_0_1) );
  XOR2_X1 f1_round_7_t_U10 ( .A(f1_round_6_io_state_out_3_1), .B(
        f1_round_7_t_n4), .Z(f1_round_7_p_io_state_out_1_4) );
  XOR2_X1 f1_round_7_t_U9 ( .A(f1_round_6_io_state_out_3_2), .B(
        f1_round_7_t_n4), .Z(f1_round_7_p_io_state_out_2_2) );
  XOR2_X1 f1_round_7_t_U8 ( .A(f1_round_6_io_state_out_3_3), .B(
        f1_round_7_t_n4), .Z(f1_round_7_p_io_state_out_3_0) );
  XOR2_X1 f1_round_7_t_U7 ( .A(f1_round_6_io_state_out_3_4), .B(
        f1_round_7_t_n4), .Z(f1_round_7_p_io_state_out_4_3) );
  XOR2_X1 f1_round_7_t_U6 ( .A(f1_round_7_t_n2), .B(f1_round_7_t_n3), .Z(
        f1_round_7_t_n1) );
  XOR2_X1 f1_round_7_t_U5 ( .A(f1_round_6_io_state_out_4_0), .B(
        f1_round_7_t_n1), .Z(f1_round_7_p_io_state_out_0_3) );
  XOR2_X1 f1_round_7_t_U4 ( .A(f1_round_6_io_state_out_4_1), .B(
        f1_round_7_t_n1), .Z(f1_round_7_p_io_state_out_1_1) );
  XOR2_X1 f1_round_7_t_U3 ( .A(f1_round_6_io_state_out_4_2), .B(
        f1_round_7_t_n1), .Z(f1_round_7_p_io_state_out_2_4) );
  XOR2_X1 f1_round_7_t_U2 ( .A(f1_round_6_io_state_out_4_3), .B(
        f1_round_7_t_n1), .Z(f1_round_7_p_io_state_out_3_2) );
  XOR2_X1 f1_round_7_t_U1 ( .A(f1_round_6_io_state_out_4_4), .B(
        f1_round_7_t_n1), .Z(f1_round_7_p_io_state_out_4_0) );
  NAND2_X1 f1_round_7_c_U50 ( .A1(f1_round_7_p_io_state_out_2_0), .A2(
        f1_round_7_p_io_state_out_1_0), .ZN(f1_round_7_c_n25) );
  XOR2_X1 f1_round_7_c_U49 ( .A(f1_round_7_c_n25), .B(
        f1_round_7_p_io_state_out_0_0), .Z(f1_round_7_c_io_state_out_0_0) );
  NAND2_X1 f1_round_7_c_U48 ( .A1(f1_round_7_p_io_state_out_2_1), .A2(
        f1_round_7_p_io_state_out_1_1), .ZN(f1_round_7_c_n24) );
  XOR2_X1 f1_round_7_c_U47 ( .A(f1_round_7_c_n24), .B(
        f1_round_7_p_io_state_out_0_1), .Z(f1_round_7_io_state_out_0_1) );
  NAND2_X1 f1_round_7_c_U46 ( .A1(f1_round_7_p_io_state_out_2_2), .A2(
        f1_round_7_p_io_state_out_1_2), .ZN(f1_round_7_c_n23) );
  XOR2_X1 f1_round_7_c_U45 ( .A(f1_round_7_c_n23), .B(
        f1_round_7_p_io_state_out_0_2), .Z(f1_round_7_io_state_out_0_2) );
  NAND2_X1 f1_round_7_c_U44 ( .A1(f1_round_7_p_io_state_out_2_3), .A2(
        f1_round_7_p_io_state_out_1_3), .ZN(f1_round_7_c_n22) );
  XOR2_X1 f1_round_7_c_U43 ( .A(f1_round_7_c_n22), .B(
        f1_round_7_p_io_state_out_0_3), .Z(f1_round_7_io_state_out_0_3) );
  NAND2_X1 f1_round_7_c_U42 ( .A1(f1_round_7_p_io_state_out_2_4), .A2(
        f1_round_7_p_io_state_out_1_4), .ZN(f1_round_7_c_n21) );
  XOR2_X1 f1_round_7_c_U41 ( .A(f1_round_7_c_n21), .B(
        f1_round_7_p_io_state_out_0_4), .Z(f1_round_7_io_state_out_0_4) );
  NAND2_X1 f1_round_7_c_U40 ( .A1(f1_round_7_p_io_state_out_2_0), .A2(
        f1_round_7_p_io_state_out_3_0), .ZN(f1_round_7_c_n20) );
  XOR2_X1 f1_round_7_c_U39 ( .A(f1_round_7_c_n20), .B(
        f1_round_7_p_io_state_out_1_0), .Z(f1_round_7_io_state_out_1_0) );
  NAND2_X1 f1_round_7_c_U38 ( .A1(f1_round_7_p_io_state_out_2_1), .A2(
        f1_round_7_p_io_state_out_3_1), .ZN(f1_round_7_c_n19) );
  XOR2_X1 f1_round_7_c_U37 ( .A(f1_round_7_c_n19), .B(
        f1_round_7_p_io_state_out_1_1), .Z(f1_round_7_io_state_out_1_1) );
  NAND2_X1 f1_round_7_c_U36 ( .A1(f1_round_7_p_io_state_out_2_2), .A2(
        f1_round_7_p_io_state_out_3_2), .ZN(f1_round_7_c_n18) );
  XOR2_X1 f1_round_7_c_U35 ( .A(f1_round_7_c_n18), .B(
        f1_round_7_p_io_state_out_1_2), .Z(f1_round_7_io_state_out_1_2) );
  NAND2_X1 f1_round_7_c_U34 ( .A1(f1_round_7_p_io_state_out_2_3), .A2(
        f1_round_7_p_io_state_out_3_3), .ZN(f1_round_7_c_n17) );
  XOR2_X1 f1_round_7_c_U33 ( .A(f1_round_7_c_n17), .B(
        f1_round_7_p_io_state_out_1_3), .Z(f1_round_7_io_state_out_1_3) );
  NAND2_X1 f1_round_7_c_U32 ( .A1(f1_round_7_p_io_state_out_2_4), .A2(
        f1_round_7_p_io_state_out_3_4), .ZN(f1_round_7_c_n16) );
  XOR2_X1 f1_round_7_c_U31 ( .A(f1_round_7_c_n16), .B(
        f1_round_7_p_io_state_out_1_4), .Z(f1_round_7_io_state_out_1_4) );
  NAND2_X1 f1_round_7_c_U30 ( .A1(f1_round_7_p_io_state_out_3_0), .A2(
        f1_round_7_p_io_state_out_4_0), .ZN(f1_round_7_c_n15) );
  XOR2_X1 f1_round_7_c_U29 ( .A(f1_round_7_c_n15), .B(
        f1_round_7_p_io_state_out_2_0), .Z(f1_round_7_io_state_out_2_0) );
  NAND2_X1 f1_round_7_c_U28 ( .A1(f1_round_7_p_io_state_out_3_1), .A2(
        f1_round_7_p_io_state_out_4_1), .ZN(f1_round_7_c_n14) );
  XOR2_X1 f1_round_7_c_U27 ( .A(f1_round_7_c_n14), .B(
        f1_round_7_p_io_state_out_2_1), .Z(f1_round_7_io_state_out_2_1) );
  NAND2_X1 f1_round_7_c_U26 ( .A1(f1_round_7_p_io_state_out_3_2), .A2(
        f1_round_7_p_io_state_out_4_2), .ZN(f1_round_7_c_n13) );
  XOR2_X1 f1_round_7_c_U25 ( .A(f1_round_7_c_n13), .B(
        f1_round_7_p_io_state_out_2_2), .Z(f1_round_7_io_state_out_2_2) );
  NAND2_X1 f1_round_7_c_U24 ( .A1(f1_round_7_p_io_state_out_3_3), .A2(
        f1_round_7_p_io_state_out_4_3), .ZN(f1_round_7_c_n12) );
  XOR2_X1 f1_round_7_c_U23 ( .A(f1_round_7_c_n12), .B(
        f1_round_7_p_io_state_out_2_3), .Z(f1_round_7_io_state_out_2_3) );
  NAND2_X1 f1_round_7_c_U22 ( .A1(f1_round_7_p_io_state_out_3_4), .A2(
        f1_round_7_p_io_state_out_4_4), .ZN(f1_round_7_c_n11) );
  XOR2_X1 f1_round_7_c_U21 ( .A(f1_round_7_c_n11), .B(
        f1_round_7_p_io_state_out_2_4), .Z(f1_round_7_io_state_out_2_4) );
  NAND2_X1 f1_round_7_c_U20 ( .A1(f1_round_7_p_io_state_out_4_0), .A2(
        f1_round_7_p_io_state_out_0_0), .ZN(f1_round_7_c_n10) );
  XOR2_X1 f1_round_7_c_U19 ( .A(f1_round_7_c_n10), .B(
        f1_round_7_p_io_state_out_3_0), .Z(f1_round_7_io_state_out_3_0) );
  NAND2_X1 f1_round_7_c_U18 ( .A1(f1_round_7_p_io_state_out_4_1), .A2(
        f1_round_7_p_io_state_out_0_1), .ZN(f1_round_7_c_n9) );
  XOR2_X1 f1_round_7_c_U17 ( .A(f1_round_7_c_n9), .B(
        f1_round_7_p_io_state_out_3_1), .Z(f1_round_7_io_state_out_3_1) );
  NAND2_X1 f1_round_7_c_U16 ( .A1(f1_round_7_p_io_state_out_4_2), .A2(
        f1_round_7_p_io_state_out_0_2), .ZN(f1_round_7_c_n8) );
  XOR2_X1 f1_round_7_c_U15 ( .A(f1_round_7_c_n8), .B(
        f1_round_7_p_io_state_out_3_2), .Z(f1_round_7_io_state_out_3_2) );
  NAND2_X1 f1_round_7_c_U14 ( .A1(f1_round_7_p_io_state_out_4_3), .A2(
        f1_round_7_p_io_state_out_0_3), .ZN(f1_round_7_c_n7) );
  XOR2_X1 f1_round_7_c_U13 ( .A(f1_round_7_c_n7), .B(
        f1_round_7_p_io_state_out_3_3), .Z(f1_round_7_io_state_out_3_3) );
  NAND2_X1 f1_round_7_c_U12 ( .A1(f1_round_7_p_io_state_out_4_4), .A2(
        f1_round_7_p_io_state_out_0_4), .ZN(f1_round_7_c_n6) );
  XOR2_X1 f1_round_7_c_U11 ( .A(f1_round_7_c_n6), .B(
        f1_round_7_p_io_state_out_3_4), .Z(f1_round_7_io_state_out_3_4) );
  NAND2_X1 f1_round_7_c_U10 ( .A1(f1_round_7_p_io_state_out_1_0), .A2(
        f1_round_7_p_io_state_out_0_0), .ZN(f1_round_7_c_n5) );
  XOR2_X1 f1_round_7_c_U9 ( .A(f1_round_7_c_n5), .B(
        f1_round_7_p_io_state_out_4_0), .Z(f1_round_7_io_state_out_4_0) );
  NAND2_X1 f1_round_7_c_U8 ( .A1(f1_round_7_p_io_state_out_1_1), .A2(
        f1_round_7_p_io_state_out_0_1), .ZN(f1_round_7_c_n4) );
  XOR2_X1 f1_round_7_c_U7 ( .A(f1_round_7_c_n4), .B(
        f1_round_7_p_io_state_out_4_1), .Z(f1_round_7_io_state_out_4_1) );
  NAND2_X1 f1_round_7_c_U6 ( .A1(f1_round_7_p_io_state_out_1_2), .A2(
        f1_round_7_p_io_state_out_0_2), .ZN(f1_round_7_c_n3) );
  XOR2_X1 f1_round_7_c_U5 ( .A(f1_round_7_c_n3), .B(
        f1_round_7_p_io_state_out_4_2), .Z(f1_round_7_io_state_out_4_2) );
  NAND2_X1 f1_round_7_c_U4 ( .A1(f1_round_7_p_io_state_out_1_3), .A2(
        f1_round_7_p_io_state_out_0_3), .ZN(f1_round_7_c_n2) );
  XOR2_X1 f1_round_7_c_U3 ( .A(f1_round_7_c_n2), .B(
        f1_round_7_p_io_state_out_4_3), .Z(f1_round_7_io_state_out_4_3) );
  NAND2_X1 f1_round_7_c_U2 ( .A1(f1_round_7_p_io_state_out_1_4), .A2(
        f1_round_7_p_io_state_out_0_4), .ZN(f1_round_7_c_n1) );
  XOR2_X1 f1_round_7_c_U1 ( .A(f1_round_7_c_n1), .B(
        f1_round_7_p_io_state_out_4_4), .Z(f1_round_7_io_state_out_4_4) );
  INV_X1 f1_round_7_i_U1 ( .A(f1_round_7_c_io_state_out_0_0), .ZN(
        f1_round_7_io_state_out_0_0) );
  XOR2_X1 f1_round_8_t_U50 ( .A(f1_round_7_io_state_out_1_4), .B(
        f1_round_7_io_state_out_1_3), .Z(f1_round_8_t_n25) );
  XNOR2_X1 f1_round_8_t_U49 ( .A(f1_round_7_io_state_out_1_2), .B(
        f1_round_8_t_n25), .ZN(f1_round_8_t_n23) );
  XOR2_X1 f1_round_8_t_U48 ( .A(f1_round_7_io_state_out_1_1), .B(
        f1_round_7_io_state_out_1_0), .Z(f1_round_8_t_n24) );
  XOR2_X1 f1_round_8_t_U47 ( .A(f1_round_8_t_n23), .B(f1_round_8_t_n24), .Z(
        f1_round_8_t_n8) );
  XOR2_X1 f1_round_8_t_U46 ( .A(f1_round_7_io_state_out_4_4), .B(
        f1_round_7_io_state_out_4_3), .Z(f1_round_8_t_n22) );
  XNOR2_X1 f1_round_8_t_U45 ( .A(f1_round_7_io_state_out_4_2), .B(
        f1_round_8_t_n22), .ZN(f1_round_8_t_n20) );
  XOR2_X1 f1_round_8_t_U44 ( .A(f1_round_7_io_state_out_4_1), .B(
        f1_round_7_io_state_out_4_0), .Z(f1_round_8_t_n21) );
  XNOR2_X1 f1_round_8_t_U43 ( .A(f1_round_8_t_n20), .B(f1_round_8_t_n21), .ZN(
        f1_round_8_t_n5) );
  XNOR2_X1 f1_round_8_t_U42 ( .A(f1_round_8_t_n8), .B(f1_round_8_t_n5), .ZN(
        f1_round_8_t_n19) );
  XOR2_X1 f1_round_8_t_U41 ( .A(f1_round_7_io_state_out_0_0), .B(
        f1_round_8_t_n19), .Z(f1_round_8_p_io_state_out_0_0) );
  XOR2_X1 f1_round_8_t_U40 ( .A(f1_round_7_io_state_out_0_1), .B(
        f1_round_8_t_n19), .Z(f1_round_8_p_io_state_out_1_3) );
  XOR2_X1 f1_round_8_t_U39 ( .A(f1_round_7_io_state_out_0_2), .B(
        f1_round_8_t_n19), .Z(f1_round_8_p_io_state_out_2_1) );
  XOR2_X1 f1_round_8_t_U38 ( .A(f1_round_7_io_state_out_0_3), .B(
        f1_round_8_t_n19), .Z(f1_round_8_p_io_state_out_3_4) );
  XOR2_X1 f1_round_8_t_U37 ( .A(f1_round_7_io_state_out_0_4), .B(
        f1_round_8_t_n19), .Z(f1_round_8_p_io_state_out_4_2) );
  XOR2_X1 f1_round_8_t_U36 ( .A(f1_round_7_io_state_out_2_4), .B(
        f1_round_7_io_state_out_2_3), .Z(f1_round_8_t_n18) );
  XNOR2_X1 f1_round_8_t_U35 ( .A(f1_round_7_io_state_out_2_2), .B(
        f1_round_8_t_n18), .ZN(f1_round_8_t_n16) );
  XOR2_X1 f1_round_8_t_U34 ( .A(f1_round_7_io_state_out_2_1), .B(
        f1_round_7_io_state_out_2_0), .Z(f1_round_8_t_n17) );
  XNOR2_X1 f1_round_8_t_U33 ( .A(f1_round_8_t_n16), .B(f1_round_8_t_n17), .ZN(
        f1_round_8_t_n6) );
  XOR2_X1 f1_round_8_t_U32 ( .A(f1_round_7_io_state_out_0_4), .B(
        f1_round_7_io_state_out_0_3), .Z(f1_round_8_t_n15) );
  XNOR2_X1 f1_round_8_t_U31 ( .A(f1_round_7_io_state_out_0_2), .B(
        f1_round_8_t_n15), .ZN(f1_round_8_t_n13) );
  XOR2_X1 f1_round_8_t_U30 ( .A(f1_round_7_io_state_out_0_1), .B(
        f1_round_7_io_state_out_0_0), .Z(f1_round_8_t_n14) );
  XNOR2_X1 f1_round_8_t_U29 ( .A(f1_round_8_t_n13), .B(f1_round_8_t_n14), .ZN(
        f1_round_8_t_n2) );
  XOR2_X1 f1_round_8_t_U28 ( .A(f1_round_8_t_n6), .B(f1_round_8_t_n2), .Z(
        f1_round_8_t_n12) );
  XOR2_X1 f1_round_8_t_U27 ( .A(f1_round_7_io_state_out_1_0), .B(
        f1_round_8_t_n12), .Z(f1_round_8_p_io_state_out_0_2) );
  XOR2_X1 f1_round_8_t_U26 ( .A(f1_round_7_io_state_out_1_1), .B(
        f1_round_8_t_n12), .Z(f1_round_8_p_io_state_out_1_0) );
  XOR2_X1 f1_round_8_t_U25 ( .A(f1_round_7_io_state_out_1_2), .B(
        f1_round_8_t_n12), .Z(f1_round_8_p_io_state_out_2_3) );
  XOR2_X1 f1_round_8_t_U24 ( .A(f1_round_7_io_state_out_1_3), .B(
        f1_round_8_t_n12), .Z(f1_round_8_p_io_state_out_3_1) );
  XOR2_X1 f1_round_8_t_U23 ( .A(f1_round_7_io_state_out_1_4), .B(
        f1_round_8_t_n12), .Z(f1_round_8_p_io_state_out_4_4) );
  XOR2_X1 f1_round_8_t_U22 ( .A(f1_round_7_io_state_out_3_4), .B(
        f1_round_7_io_state_out_3_3), .Z(f1_round_8_t_n11) );
  XNOR2_X1 f1_round_8_t_U21 ( .A(f1_round_7_io_state_out_3_2), .B(
        f1_round_8_t_n11), .ZN(f1_round_8_t_n9) );
  XOR2_X1 f1_round_8_t_U20 ( .A(f1_round_7_io_state_out_3_1), .B(
        f1_round_7_io_state_out_3_0), .Z(f1_round_8_t_n10) );
  XNOR2_X1 f1_round_8_t_U19 ( .A(f1_round_8_t_n9), .B(f1_round_8_t_n10), .ZN(
        f1_round_8_t_n3) );
  XNOR2_X1 f1_round_8_t_U18 ( .A(f1_round_8_t_n8), .B(f1_round_8_t_n3), .ZN(
        f1_round_8_t_n7) );
  XOR2_X1 f1_round_8_t_U17 ( .A(f1_round_7_io_state_out_2_0), .B(
        f1_round_8_t_n7), .Z(f1_round_8_p_io_state_out_0_4) );
  XOR2_X1 f1_round_8_t_U16 ( .A(f1_round_7_io_state_out_2_1), .B(
        f1_round_8_t_n7), .Z(f1_round_8_p_io_state_out_1_2) );
  XOR2_X1 f1_round_8_t_U15 ( .A(f1_round_7_io_state_out_2_2), .B(
        f1_round_8_t_n7), .Z(f1_round_8_p_io_state_out_2_0) );
  XOR2_X1 f1_round_8_t_U14 ( .A(f1_round_7_io_state_out_2_3), .B(
        f1_round_8_t_n7), .Z(f1_round_8_p_io_state_out_3_3) );
  XOR2_X1 f1_round_8_t_U13 ( .A(f1_round_7_io_state_out_2_4), .B(
        f1_round_8_t_n7), .Z(f1_round_8_p_io_state_out_4_1) );
  XOR2_X1 f1_round_8_t_U12 ( .A(f1_round_8_t_n5), .B(f1_round_8_t_n6), .Z(
        f1_round_8_t_n4) );
  XOR2_X1 f1_round_8_t_U11 ( .A(f1_round_7_io_state_out_3_0), .B(
        f1_round_8_t_n4), .Z(f1_round_8_p_io_state_out_0_1) );
  XOR2_X1 f1_round_8_t_U10 ( .A(f1_round_7_io_state_out_3_1), .B(
        f1_round_8_t_n4), .Z(f1_round_8_p_io_state_out_1_4) );
  XOR2_X1 f1_round_8_t_U9 ( .A(f1_round_7_io_state_out_3_2), .B(
        f1_round_8_t_n4), .Z(f1_round_8_p_io_state_out_2_2) );
  XOR2_X1 f1_round_8_t_U8 ( .A(f1_round_7_io_state_out_3_3), .B(
        f1_round_8_t_n4), .Z(f1_round_8_p_io_state_out_3_0) );
  XOR2_X1 f1_round_8_t_U7 ( .A(f1_round_7_io_state_out_3_4), .B(
        f1_round_8_t_n4), .Z(f1_round_8_p_io_state_out_4_3) );
  XOR2_X1 f1_round_8_t_U6 ( .A(f1_round_8_t_n2), .B(f1_round_8_t_n3), .Z(
        f1_round_8_t_n1) );
  XOR2_X1 f1_round_8_t_U5 ( .A(f1_round_7_io_state_out_4_0), .B(
        f1_round_8_t_n1), .Z(f1_round_8_p_io_state_out_0_3) );
  XOR2_X1 f1_round_8_t_U4 ( .A(f1_round_7_io_state_out_4_1), .B(
        f1_round_8_t_n1), .Z(f1_round_8_p_io_state_out_1_1) );
  XOR2_X1 f1_round_8_t_U3 ( .A(f1_round_7_io_state_out_4_2), .B(
        f1_round_8_t_n1), .Z(f1_round_8_p_io_state_out_2_4) );
  XOR2_X1 f1_round_8_t_U2 ( .A(f1_round_7_io_state_out_4_3), .B(
        f1_round_8_t_n1), .Z(f1_round_8_p_io_state_out_3_2) );
  XOR2_X1 f1_round_8_t_U1 ( .A(f1_round_7_io_state_out_4_4), .B(
        f1_round_8_t_n1), .Z(f1_round_8_p_io_state_out_4_0) );
  NAND2_X1 f1_round_8_c_U50 ( .A1(f1_round_8_p_io_state_out_2_0), .A2(
        f1_round_8_p_io_state_out_1_0), .ZN(f1_round_8_c_n25) );
  XOR2_X1 f1_round_8_c_U49 ( .A(f1_round_8_c_n25), .B(
        f1_round_8_p_io_state_out_0_0), .Z(f1_round_8_io_state_out_0_0) );
  NAND2_X1 f1_round_8_c_U48 ( .A1(f1_round_8_p_io_state_out_2_1), .A2(
        f1_round_8_p_io_state_out_1_1), .ZN(f1_round_8_c_n24) );
  XOR2_X1 f1_round_8_c_U47 ( .A(f1_round_8_c_n24), .B(
        f1_round_8_p_io_state_out_0_1), .Z(f1_round_8_io_state_out_0_1) );
  NAND2_X1 f1_round_8_c_U46 ( .A1(f1_round_8_p_io_state_out_2_2), .A2(
        f1_round_8_p_io_state_out_1_2), .ZN(f1_round_8_c_n23) );
  XOR2_X1 f1_round_8_c_U45 ( .A(f1_round_8_c_n23), .B(
        f1_round_8_p_io_state_out_0_2), .Z(f1_round_8_io_state_out_0_2) );
  NAND2_X1 f1_round_8_c_U44 ( .A1(f1_round_8_p_io_state_out_2_3), .A2(
        f1_round_8_p_io_state_out_1_3), .ZN(f1_round_8_c_n22) );
  XOR2_X1 f1_round_8_c_U43 ( .A(f1_round_8_c_n22), .B(
        f1_round_8_p_io_state_out_0_3), .Z(f1_round_8_io_state_out_0_3) );
  NAND2_X1 f1_round_8_c_U42 ( .A1(f1_round_8_p_io_state_out_2_4), .A2(
        f1_round_8_p_io_state_out_1_4), .ZN(f1_round_8_c_n21) );
  XOR2_X1 f1_round_8_c_U41 ( .A(f1_round_8_c_n21), .B(
        f1_round_8_p_io_state_out_0_4), .Z(f1_round_8_io_state_out_0_4) );
  NAND2_X1 f1_round_8_c_U40 ( .A1(f1_round_8_p_io_state_out_2_0), .A2(
        f1_round_8_p_io_state_out_3_0), .ZN(f1_round_8_c_n20) );
  XOR2_X1 f1_round_8_c_U39 ( .A(f1_round_8_c_n20), .B(
        f1_round_8_p_io_state_out_1_0), .Z(f1_round_8_io_state_out_1_0) );
  NAND2_X1 f1_round_8_c_U38 ( .A1(f1_round_8_p_io_state_out_2_1), .A2(
        f1_round_8_p_io_state_out_3_1), .ZN(f1_round_8_c_n19) );
  XOR2_X1 f1_round_8_c_U37 ( .A(f1_round_8_c_n19), .B(
        f1_round_8_p_io_state_out_1_1), .Z(f1_round_8_io_state_out_1_1) );
  NAND2_X1 f1_round_8_c_U36 ( .A1(f1_round_8_p_io_state_out_2_2), .A2(
        f1_round_8_p_io_state_out_3_2), .ZN(f1_round_8_c_n18) );
  XOR2_X1 f1_round_8_c_U35 ( .A(f1_round_8_c_n18), .B(
        f1_round_8_p_io_state_out_1_2), .Z(f1_round_8_io_state_out_1_2) );
  NAND2_X1 f1_round_8_c_U34 ( .A1(f1_round_8_p_io_state_out_2_3), .A2(
        f1_round_8_p_io_state_out_3_3), .ZN(f1_round_8_c_n17) );
  XOR2_X1 f1_round_8_c_U33 ( .A(f1_round_8_c_n17), .B(
        f1_round_8_p_io_state_out_1_3), .Z(f1_round_8_io_state_out_1_3) );
  NAND2_X1 f1_round_8_c_U32 ( .A1(f1_round_8_p_io_state_out_2_4), .A2(
        f1_round_8_p_io_state_out_3_4), .ZN(f1_round_8_c_n16) );
  XOR2_X1 f1_round_8_c_U31 ( .A(f1_round_8_c_n16), .B(
        f1_round_8_p_io_state_out_1_4), .Z(f1_round_8_io_state_out_1_4) );
  NAND2_X1 f1_round_8_c_U30 ( .A1(f1_round_8_p_io_state_out_3_0), .A2(
        f1_round_8_p_io_state_out_4_0), .ZN(f1_round_8_c_n15) );
  XOR2_X1 f1_round_8_c_U29 ( .A(f1_round_8_c_n15), .B(
        f1_round_8_p_io_state_out_2_0), .Z(f1_round_8_io_state_out_2_0) );
  NAND2_X1 f1_round_8_c_U28 ( .A1(f1_round_8_p_io_state_out_3_1), .A2(
        f1_round_8_p_io_state_out_4_1), .ZN(f1_round_8_c_n14) );
  XOR2_X1 f1_round_8_c_U27 ( .A(f1_round_8_c_n14), .B(
        f1_round_8_p_io_state_out_2_1), .Z(f1_round_8_io_state_out_2_1) );
  NAND2_X1 f1_round_8_c_U26 ( .A1(f1_round_8_p_io_state_out_3_2), .A2(
        f1_round_8_p_io_state_out_4_2), .ZN(f1_round_8_c_n13) );
  XOR2_X1 f1_round_8_c_U25 ( .A(f1_round_8_c_n13), .B(
        f1_round_8_p_io_state_out_2_2), .Z(f1_round_8_io_state_out_2_2) );
  NAND2_X1 f1_round_8_c_U24 ( .A1(f1_round_8_p_io_state_out_3_3), .A2(
        f1_round_8_p_io_state_out_4_3), .ZN(f1_round_8_c_n12) );
  XOR2_X1 f1_round_8_c_U23 ( .A(f1_round_8_c_n12), .B(
        f1_round_8_p_io_state_out_2_3), .Z(f1_round_8_io_state_out_2_3) );
  NAND2_X1 f1_round_8_c_U22 ( .A1(f1_round_8_p_io_state_out_3_4), .A2(
        f1_round_8_p_io_state_out_4_4), .ZN(f1_round_8_c_n11) );
  XOR2_X1 f1_round_8_c_U21 ( .A(f1_round_8_c_n11), .B(
        f1_round_8_p_io_state_out_2_4), .Z(f1_round_8_io_state_out_2_4) );
  NAND2_X1 f1_round_8_c_U20 ( .A1(f1_round_8_p_io_state_out_4_0), .A2(
        f1_round_8_p_io_state_out_0_0), .ZN(f1_round_8_c_n10) );
  XOR2_X1 f1_round_8_c_U19 ( .A(f1_round_8_c_n10), .B(
        f1_round_8_p_io_state_out_3_0), .Z(f1_round_8_io_state_out_3_0) );
  NAND2_X1 f1_round_8_c_U18 ( .A1(f1_round_8_p_io_state_out_4_1), .A2(
        f1_round_8_p_io_state_out_0_1), .ZN(f1_round_8_c_n9) );
  XOR2_X1 f1_round_8_c_U17 ( .A(f1_round_8_c_n9), .B(
        f1_round_8_p_io_state_out_3_1), .Z(f1_round_8_io_state_out_3_1) );
  NAND2_X1 f1_round_8_c_U16 ( .A1(f1_round_8_p_io_state_out_4_2), .A2(
        f1_round_8_p_io_state_out_0_2), .ZN(f1_round_8_c_n8) );
  XOR2_X1 f1_round_8_c_U15 ( .A(f1_round_8_c_n8), .B(
        f1_round_8_p_io_state_out_3_2), .Z(f1_round_8_io_state_out_3_2) );
  NAND2_X1 f1_round_8_c_U14 ( .A1(f1_round_8_p_io_state_out_4_3), .A2(
        f1_round_8_p_io_state_out_0_3), .ZN(f1_round_8_c_n7) );
  XOR2_X1 f1_round_8_c_U13 ( .A(f1_round_8_c_n7), .B(
        f1_round_8_p_io_state_out_3_3), .Z(f1_round_8_io_state_out_3_3) );
  NAND2_X1 f1_round_8_c_U12 ( .A1(f1_round_8_p_io_state_out_4_4), .A2(
        f1_round_8_p_io_state_out_0_4), .ZN(f1_round_8_c_n6) );
  XOR2_X1 f1_round_8_c_U11 ( .A(f1_round_8_c_n6), .B(
        f1_round_8_p_io_state_out_3_4), .Z(f1_round_8_io_state_out_3_4) );
  NAND2_X1 f1_round_8_c_U10 ( .A1(f1_round_8_p_io_state_out_1_0), .A2(
        f1_round_8_p_io_state_out_0_0), .ZN(f1_round_8_c_n5) );
  XOR2_X1 f1_round_8_c_U9 ( .A(f1_round_8_c_n5), .B(
        f1_round_8_p_io_state_out_4_0), .Z(f1_round_8_io_state_out_4_0) );
  NAND2_X1 f1_round_8_c_U8 ( .A1(f1_round_8_p_io_state_out_1_1), .A2(
        f1_round_8_p_io_state_out_0_1), .ZN(f1_round_8_c_n4) );
  XOR2_X1 f1_round_8_c_U7 ( .A(f1_round_8_c_n4), .B(
        f1_round_8_p_io_state_out_4_1), .Z(f1_round_8_io_state_out_4_1) );
  NAND2_X1 f1_round_8_c_U6 ( .A1(f1_round_8_p_io_state_out_1_2), .A2(
        f1_round_8_p_io_state_out_0_2), .ZN(f1_round_8_c_n3) );
  XOR2_X1 f1_round_8_c_U5 ( .A(f1_round_8_c_n3), .B(
        f1_round_8_p_io_state_out_4_2), .Z(f1_round_8_io_state_out_4_2) );
  NAND2_X1 f1_round_8_c_U4 ( .A1(f1_round_8_p_io_state_out_1_3), .A2(
        f1_round_8_p_io_state_out_0_3), .ZN(f1_round_8_c_n2) );
  XOR2_X1 f1_round_8_c_U3 ( .A(f1_round_8_c_n2), .B(
        f1_round_8_p_io_state_out_4_3), .Z(f1_round_8_io_state_out_4_3) );
  NAND2_X1 f1_round_8_c_U2 ( .A1(f1_round_8_p_io_state_out_1_4), .A2(
        f1_round_8_p_io_state_out_0_4), .ZN(f1_round_8_c_n1) );
  XOR2_X1 f1_round_8_c_U1 ( .A(f1_round_8_c_n1), .B(
        f1_round_8_p_io_state_out_4_4), .Z(f1_round_8_io_state_out_4_4) );
  XOR2_X1 f1_round_9_t_U50 ( .A(f1_round_8_io_state_out_1_4), .B(
        f1_round_8_io_state_out_1_3), .Z(f1_round_9_t_n25) );
  XNOR2_X1 f1_round_9_t_U49 ( .A(f1_round_8_io_state_out_1_2), .B(
        f1_round_9_t_n25), .ZN(f1_round_9_t_n23) );
  XOR2_X1 f1_round_9_t_U48 ( .A(f1_round_8_io_state_out_1_1), .B(
        f1_round_8_io_state_out_1_0), .Z(f1_round_9_t_n24) );
  XOR2_X1 f1_round_9_t_U47 ( .A(f1_round_9_t_n23), .B(f1_round_9_t_n24), .Z(
        f1_round_9_t_n8) );
  XOR2_X1 f1_round_9_t_U46 ( .A(f1_round_8_io_state_out_4_4), .B(
        f1_round_8_io_state_out_4_3), .Z(f1_round_9_t_n22) );
  XNOR2_X1 f1_round_9_t_U45 ( .A(f1_round_8_io_state_out_4_2), .B(
        f1_round_9_t_n22), .ZN(f1_round_9_t_n20) );
  XOR2_X1 f1_round_9_t_U44 ( .A(f1_round_8_io_state_out_4_1), .B(
        f1_round_8_io_state_out_4_0), .Z(f1_round_9_t_n21) );
  XNOR2_X1 f1_round_9_t_U43 ( .A(f1_round_9_t_n20), .B(f1_round_9_t_n21), .ZN(
        f1_round_9_t_n5) );
  XNOR2_X1 f1_round_9_t_U42 ( .A(f1_round_9_t_n8), .B(f1_round_9_t_n5), .ZN(
        f1_round_9_t_n19) );
  XOR2_X1 f1_round_9_t_U41 ( .A(f1_round_8_io_state_out_0_0), .B(
        f1_round_9_t_n19), .Z(f1_round_9_p_io_state_out_0_0) );
  XOR2_X1 f1_round_9_t_U40 ( .A(f1_round_8_io_state_out_0_1), .B(
        f1_round_9_t_n19), .Z(f1_round_9_p_io_state_out_1_3) );
  XOR2_X1 f1_round_9_t_U39 ( .A(f1_round_8_io_state_out_0_2), .B(
        f1_round_9_t_n19), .Z(f1_round_9_p_io_state_out_2_1) );
  XOR2_X1 f1_round_9_t_U38 ( .A(f1_round_8_io_state_out_0_3), .B(
        f1_round_9_t_n19), .Z(f1_round_9_p_io_state_out_3_4) );
  XOR2_X1 f1_round_9_t_U37 ( .A(f1_round_8_io_state_out_0_4), .B(
        f1_round_9_t_n19), .Z(f1_round_9_p_io_state_out_4_2) );
  XOR2_X1 f1_round_9_t_U36 ( .A(f1_round_8_io_state_out_2_4), .B(
        f1_round_8_io_state_out_2_3), .Z(f1_round_9_t_n18) );
  XNOR2_X1 f1_round_9_t_U35 ( .A(f1_round_8_io_state_out_2_2), .B(
        f1_round_9_t_n18), .ZN(f1_round_9_t_n16) );
  XOR2_X1 f1_round_9_t_U34 ( .A(f1_round_8_io_state_out_2_1), .B(
        f1_round_8_io_state_out_2_0), .Z(f1_round_9_t_n17) );
  XNOR2_X1 f1_round_9_t_U33 ( .A(f1_round_9_t_n16), .B(f1_round_9_t_n17), .ZN(
        f1_round_9_t_n6) );
  XOR2_X1 f1_round_9_t_U32 ( .A(f1_round_8_io_state_out_0_4), .B(
        f1_round_8_io_state_out_0_3), .Z(f1_round_9_t_n15) );
  XNOR2_X1 f1_round_9_t_U31 ( .A(f1_round_8_io_state_out_0_2), .B(
        f1_round_9_t_n15), .ZN(f1_round_9_t_n13) );
  XOR2_X1 f1_round_9_t_U30 ( .A(f1_round_8_io_state_out_0_1), .B(
        f1_round_8_io_state_out_0_0), .Z(f1_round_9_t_n14) );
  XNOR2_X1 f1_round_9_t_U29 ( .A(f1_round_9_t_n13), .B(f1_round_9_t_n14), .ZN(
        f1_round_9_t_n2) );
  XOR2_X1 f1_round_9_t_U28 ( .A(f1_round_9_t_n6), .B(f1_round_9_t_n2), .Z(
        f1_round_9_t_n12) );
  XOR2_X1 f1_round_9_t_U27 ( .A(f1_round_8_io_state_out_1_0), .B(
        f1_round_9_t_n12), .Z(f1_round_9_p_io_state_out_0_2) );
  XOR2_X1 f1_round_9_t_U26 ( .A(f1_round_8_io_state_out_1_1), .B(
        f1_round_9_t_n12), .Z(f1_round_9_p_io_state_out_1_0) );
  XOR2_X1 f1_round_9_t_U25 ( .A(f1_round_8_io_state_out_1_2), .B(
        f1_round_9_t_n12), .Z(f1_round_9_p_io_state_out_2_3) );
  XOR2_X1 f1_round_9_t_U24 ( .A(f1_round_8_io_state_out_1_3), .B(
        f1_round_9_t_n12), .Z(f1_round_9_p_io_state_out_3_1) );
  XOR2_X1 f1_round_9_t_U23 ( .A(f1_round_8_io_state_out_1_4), .B(
        f1_round_9_t_n12), .Z(f1_round_9_p_io_state_out_4_4) );
  XOR2_X1 f1_round_9_t_U22 ( .A(f1_round_8_io_state_out_3_4), .B(
        f1_round_8_io_state_out_3_3), .Z(f1_round_9_t_n11) );
  XNOR2_X1 f1_round_9_t_U21 ( .A(f1_round_8_io_state_out_3_2), .B(
        f1_round_9_t_n11), .ZN(f1_round_9_t_n9) );
  XOR2_X1 f1_round_9_t_U20 ( .A(f1_round_8_io_state_out_3_1), .B(
        f1_round_8_io_state_out_3_0), .Z(f1_round_9_t_n10) );
  XNOR2_X1 f1_round_9_t_U19 ( .A(f1_round_9_t_n9), .B(f1_round_9_t_n10), .ZN(
        f1_round_9_t_n3) );
  XNOR2_X1 f1_round_9_t_U18 ( .A(f1_round_9_t_n8), .B(f1_round_9_t_n3), .ZN(
        f1_round_9_t_n7) );
  XOR2_X1 f1_round_9_t_U17 ( .A(f1_round_8_io_state_out_2_0), .B(
        f1_round_9_t_n7), .Z(f1_round_9_p_io_state_out_0_4) );
  XOR2_X1 f1_round_9_t_U16 ( .A(f1_round_8_io_state_out_2_1), .B(
        f1_round_9_t_n7), .Z(f1_round_9_p_io_state_out_1_2) );
  XOR2_X1 f1_round_9_t_U15 ( .A(f1_round_8_io_state_out_2_2), .B(
        f1_round_9_t_n7), .Z(f1_round_9_p_io_state_out_2_0) );
  XOR2_X1 f1_round_9_t_U14 ( .A(f1_round_8_io_state_out_2_3), .B(
        f1_round_9_t_n7), .Z(f1_round_9_p_io_state_out_3_3) );
  XOR2_X1 f1_round_9_t_U13 ( .A(f1_round_8_io_state_out_2_4), .B(
        f1_round_9_t_n7), .Z(f1_round_9_p_io_state_out_4_1) );
  XOR2_X1 f1_round_9_t_U12 ( .A(f1_round_9_t_n5), .B(f1_round_9_t_n6), .Z(
        f1_round_9_t_n4) );
  XOR2_X1 f1_round_9_t_U11 ( .A(f1_round_8_io_state_out_3_0), .B(
        f1_round_9_t_n4), .Z(f1_round_9_p_io_state_out_0_1) );
  XOR2_X1 f1_round_9_t_U10 ( .A(f1_round_8_io_state_out_3_1), .B(
        f1_round_9_t_n4), .Z(f1_round_9_p_io_state_out_1_4) );
  XOR2_X1 f1_round_9_t_U9 ( .A(f1_round_8_io_state_out_3_2), .B(
        f1_round_9_t_n4), .Z(f1_round_9_p_io_state_out_2_2) );
  XOR2_X1 f1_round_9_t_U8 ( .A(f1_round_8_io_state_out_3_3), .B(
        f1_round_9_t_n4), .Z(f1_round_9_p_io_state_out_3_0) );
  XOR2_X1 f1_round_9_t_U7 ( .A(f1_round_8_io_state_out_3_4), .B(
        f1_round_9_t_n4), .Z(f1_round_9_p_io_state_out_4_3) );
  XOR2_X1 f1_round_9_t_U6 ( .A(f1_round_9_t_n2), .B(f1_round_9_t_n3), .Z(
        f1_round_9_t_n1) );
  XOR2_X1 f1_round_9_t_U5 ( .A(f1_round_8_io_state_out_4_0), .B(
        f1_round_9_t_n1), .Z(f1_round_9_p_io_state_out_0_3) );
  XOR2_X1 f1_round_9_t_U4 ( .A(f1_round_8_io_state_out_4_1), .B(
        f1_round_9_t_n1), .Z(f1_round_9_p_io_state_out_1_1) );
  XOR2_X1 f1_round_9_t_U3 ( .A(f1_round_8_io_state_out_4_2), .B(
        f1_round_9_t_n1), .Z(f1_round_9_p_io_state_out_2_4) );
  XOR2_X1 f1_round_9_t_U2 ( .A(f1_round_8_io_state_out_4_3), .B(
        f1_round_9_t_n1), .Z(f1_round_9_p_io_state_out_3_2) );
  XOR2_X1 f1_round_9_t_U1 ( .A(f1_round_8_io_state_out_4_4), .B(
        f1_round_9_t_n1), .Z(f1_round_9_p_io_state_out_4_0) );
  NAND2_X1 f1_round_9_c_U50 ( .A1(f1_round_9_p_io_state_out_2_0), .A2(
        f1_round_9_p_io_state_out_1_0), .ZN(f1_round_9_c_n25) );
  XOR2_X1 f1_round_9_c_U49 ( .A(f1_round_9_c_n25), .B(
        f1_round_9_p_io_state_out_0_0), .Z(f1_round_9_io_state_out_0_0) );
  NAND2_X1 f1_round_9_c_U48 ( .A1(f1_round_9_p_io_state_out_2_1), .A2(
        f1_round_9_p_io_state_out_1_1), .ZN(f1_round_9_c_n24) );
  XOR2_X1 f1_round_9_c_U47 ( .A(f1_round_9_c_n24), .B(
        f1_round_9_p_io_state_out_0_1), .Z(f1_round_9_io_state_out_0_1) );
  NAND2_X1 f1_round_9_c_U46 ( .A1(f1_round_9_p_io_state_out_2_2), .A2(
        f1_round_9_p_io_state_out_1_2), .ZN(f1_round_9_c_n23) );
  XOR2_X1 f1_round_9_c_U45 ( .A(f1_round_9_c_n23), .B(
        f1_round_9_p_io_state_out_0_2), .Z(f1_round_9_io_state_out_0_2) );
  NAND2_X1 f1_round_9_c_U44 ( .A1(f1_round_9_p_io_state_out_2_3), .A2(
        f1_round_9_p_io_state_out_1_3), .ZN(f1_round_9_c_n22) );
  XOR2_X1 f1_round_9_c_U43 ( .A(f1_round_9_c_n22), .B(
        f1_round_9_p_io_state_out_0_3), .Z(f1_round_9_io_state_out_0_3) );
  NAND2_X1 f1_round_9_c_U42 ( .A1(f1_round_9_p_io_state_out_2_4), .A2(
        f1_round_9_p_io_state_out_1_4), .ZN(f1_round_9_c_n21) );
  XOR2_X1 f1_round_9_c_U41 ( .A(f1_round_9_c_n21), .B(
        f1_round_9_p_io_state_out_0_4), .Z(f1_round_9_io_state_out_0_4) );
  NAND2_X1 f1_round_9_c_U40 ( .A1(f1_round_9_p_io_state_out_2_0), .A2(
        f1_round_9_p_io_state_out_3_0), .ZN(f1_round_9_c_n20) );
  XOR2_X1 f1_round_9_c_U39 ( .A(f1_round_9_c_n20), .B(
        f1_round_9_p_io_state_out_1_0), .Z(f1_round_9_io_state_out_1_0) );
  NAND2_X1 f1_round_9_c_U38 ( .A1(f1_round_9_p_io_state_out_2_1), .A2(
        f1_round_9_p_io_state_out_3_1), .ZN(f1_round_9_c_n19) );
  XOR2_X1 f1_round_9_c_U37 ( .A(f1_round_9_c_n19), .B(
        f1_round_9_p_io_state_out_1_1), .Z(f1_round_9_io_state_out_1_1) );
  NAND2_X1 f1_round_9_c_U36 ( .A1(f1_round_9_p_io_state_out_2_2), .A2(
        f1_round_9_p_io_state_out_3_2), .ZN(f1_round_9_c_n18) );
  XOR2_X1 f1_round_9_c_U35 ( .A(f1_round_9_c_n18), .B(
        f1_round_9_p_io_state_out_1_2), .Z(f1_round_9_io_state_out_1_2) );
  NAND2_X1 f1_round_9_c_U34 ( .A1(f1_round_9_p_io_state_out_2_3), .A2(
        f1_round_9_p_io_state_out_3_3), .ZN(f1_round_9_c_n17) );
  XOR2_X1 f1_round_9_c_U33 ( .A(f1_round_9_c_n17), .B(
        f1_round_9_p_io_state_out_1_3), .Z(f1_round_9_io_state_out_1_3) );
  NAND2_X1 f1_round_9_c_U32 ( .A1(f1_round_9_p_io_state_out_2_4), .A2(
        f1_round_9_p_io_state_out_3_4), .ZN(f1_round_9_c_n16) );
  XOR2_X1 f1_round_9_c_U31 ( .A(f1_round_9_c_n16), .B(
        f1_round_9_p_io_state_out_1_4), .Z(f1_round_9_io_state_out_1_4) );
  NAND2_X1 f1_round_9_c_U30 ( .A1(f1_round_9_p_io_state_out_3_0), .A2(
        f1_round_9_p_io_state_out_4_0), .ZN(f1_round_9_c_n15) );
  XOR2_X1 f1_round_9_c_U29 ( .A(f1_round_9_c_n15), .B(
        f1_round_9_p_io_state_out_2_0), .Z(f1_round_9_io_state_out_2_0) );
  NAND2_X1 f1_round_9_c_U28 ( .A1(f1_round_9_p_io_state_out_3_1), .A2(
        f1_round_9_p_io_state_out_4_1), .ZN(f1_round_9_c_n14) );
  XOR2_X1 f1_round_9_c_U27 ( .A(f1_round_9_c_n14), .B(
        f1_round_9_p_io_state_out_2_1), .Z(f1_round_9_io_state_out_2_1) );
  NAND2_X1 f1_round_9_c_U26 ( .A1(f1_round_9_p_io_state_out_3_2), .A2(
        f1_round_9_p_io_state_out_4_2), .ZN(f1_round_9_c_n13) );
  XOR2_X1 f1_round_9_c_U25 ( .A(f1_round_9_c_n13), .B(
        f1_round_9_p_io_state_out_2_2), .Z(f1_round_9_io_state_out_2_2) );
  NAND2_X1 f1_round_9_c_U24 ( .A1(f1_round_9_p_io_state_out_3_3), .A2(
        f1_round_9_p_io_state_out_4_3), .ZN(f1_round_9_c_n12) );
  XOR2_X1 f1_round_9_c_U23 ( .A(f1_round_9_c_n12), .B(
        f1_round_9_p_io_state_out_2_3), .Z(f1_round_9_io_state_out_2_3) );
  NAND2_X1 f1_round_9_c_U22 ( .A1(f1_round_9_p_io_state_out_3_4), .A2(
        f1_round_9_p_io_state_out_4_4), .ZN(f1_round_9_c_n11) );
  XOR2_X1 f1_round_9_c_U21 ( .A(f1_round_9_c_n11), .B(
        f1_round_9_p_io_state_out_2_4), .Z(f1_round_9_io_state_out_2_4) );
  NAND2_X1 f1_round_9_c_U20 ( .A1(f1_round_9_p_io_state_out_4_0), .A2(
        f1_round_9_p_io_state_out_0_0), .ZN(f1_round_9_c_n10) );
  XOR2_X1 f1_round_9_c_U19 ( .A(f1_round_9_c_n10), .B(
        f1_round_9_p_io_state_out_3_0), .Z(f1_round_9_io_state_out_3_0) );
  NAND2_X1 f1_round_9_c_U18 ( .A1(f1_round_9_p_io_state_out_4_1), .A2(
        f1_round_9_p_io_state_out_0_1), .ZN(f1_round_9_c_n9) );
  XOR2_X1 f1_round_9_c_U17 ( .A(f1_round_9_c_n9), .B(
        f1_round_9_p_io_state_out_3_1), .Z(f1_round_9_io_state_out_3_1) );
  NAND2_X1 f1_round_9_c_U16 ( .A1(f1_round_9_p_io_state_out_4_2), .A2(
        f1_round_9_p_io_state_out_0_2), .ZN(f1_round_9_c_n8) );
  XOR2_X1 f1_round_9_c_U15 ( .A(f1_round_9_c_n8), .B(
        f1_round_9_p_io_state_out_3_2), .Z(f1_round_9_io_state_out_3_2) );
  NAND2_X1 f1_round_9_c_U14 ( .A1(f1_round_9_p_io_state_out_4_3), .A2(
        f1_round_9_p_io_state_out_0_3), .ZN(f1_round_9_c_n7) );
  XOR2_X1 f1_round_9_c_U13 ( .A(f1_round_9_c_n7), .B(
        f1_round_9_p_io_state_out_3_3), .Z(f1_round_9_io_state_out_3_3) );
  NAND2_X1 f1_round_9_c_U12 ( .A1(f1_round_9_p_io_state_out_4_4), .A2(
        f1_round_9_p_io_state_out_0_4), .ZN(f1_round_9_c_n6) );
  XOR2_X1 f1_round_9_c_U11 ( .A(f1_round_9_c_n6), .B(
        f1_round_9_p_io_state_out_3_4), .Z(f1_round_9_io_state_out_3_4) );
  NAND2_X1 f1_round_9_c_U10 ( .A1(f1_round_9_p_io_state_out_1_0), .A2(
        f1_round_9_p_io_state_out_0_0), .ZN(f1_round_9_c_n5) );
  XOR2_X1 f1_round_9_c_U9 ( .A(f1_round_9_c_n5), .B(
        f1_round_9_p_io_state_out_4_0), .Z(f1_round_9_io_state_out_4_0) );
  NAND2_X1 f1_round_9_c_U8 ( .A1(f1_round_9_p_io_state_out_1_1), .A2(
        f1_round_9_p_io_state_out_0_1), .ZN(f1_round_9_c_n4) );
  XOR2_X1 f1_round_9_c_U7 ( .A(f1_round_9_c_n4), .B(
        f1_round_9_p_io_state_out_4_1), .Z(f1_round_9_io_state_out_4_1) );
  NAND2_X1 f1_round_9_c_U6 ( .A1(f1_round_9_p_io_state_out_1_2), .A2(
        f1_round_9_p_io_state_out_0_2), .ZN(f1_round_9_c_n3) );
  XOR2_X1 f1_round_9_c_U5 ( .A(f1_round_9_c_n3), .B(
        f1_round_9_p_io_state_out_4_2), .Z(f1_round_9_io_state_out_4_2) );
  NAND2_X1 f1_round_9_c_U4 ( .A1(f1_round_9_p_io_state_out_1_3), .A2(
        f1_round_9_p_io_state_out_0_3), .ZN(f1_round_9_c_n2) );
  XOR2_X1 f1_round_9_c_U3 ( .A(f1_round_9_c_n2), .B(
        f1_round_9_p_io_state_out_4_3), .Z(f1_round_9_io_state_out_4_3) );
  NAND2_X1 f1_round_9_c_U2 ( .A1(f1_round_9_p_io_state_out_1_4), .A2(
        f1_round_9_p_io_state_out_0_4), .ZN(f1_round_9_c_n1) );
  XOR2_X1 f1_round_9_c_U1 ( .A(f1_round_9_c_n1), .B(
        f1_round_9_p_io_state_out_4_4), .Z(f1_round_9_io_state_out_4_4) );
  XOR2_X1 f1_round_10_t_U50 ( .A(f1_round_9_io_state_out_1_4), .B(
        f1_round_9_io_state_out_1_3), .Z(f1_round_10_t_n25) );
  XNOR2_X1 f1_round_10_t_U49 ( .A(f1_round_9_io_state_out_1_2), .B(
        f1_round_10_t_n25), .ZN(f1_round_10_t_n23) );
  XOR2_X1 f1_round_10_t_U48 ( .A(f1_round_9_io_state_out_1_1), .B(
        f1_round_9_io_state_out_1_0), .Z(f1_round_10_t_n24) );
  XOR2_X1 f1_round_10_t_U47 ( .A(f1_round_10_t_n23), .B(f1_round_10_t_n24), 
        .Z(f1_round_10_t_n8) );
  XOR2_X1 f1_round_10_t_U46 ( .A(f1_round_9_io_state_out_4_4), .B(
        f1_round_9_io_state_out_4_3), .Z(f1_round_10_t_n22) );
  XNOR2_X1 f1_round_10_t_U45 ( .A(f1_round_9_io_state_out_4_2), .B(
        f1_round_10_t_n22), .ZN(f1_round_10_t_n20) );
  XOR2_X1 f1_round_10_t_U44 ( .A(f1_round_9_io_state_out_4_1), .B(
        f1_round_9_io_state_out_4_0), .Z(f1_round_10_t_n21) );
  XNOR2_X1 f1_round_10_t_U43 ( .A(f1_round_10_t_n20), .B(f1_round_10_t_n21), 
        .ZN(f1_round_10_t_n5) );
  XNOR2_X1 f1_round_10_t_U42 ( .A(f1_round_10_t_n8), .B(f1_round_10_t_n5), 
        .ZN(f1_round_10_t_n19) );
  XOR2_X1 f1_round_10_t_U41 ( .A(f1_round_9_io_state_out_0_0), .B(
        f1_round_10_t_n19), .Z(f1_round_10_p_io_state_out_0_0) );
  XOR2_X1 f1_round_10_t_U40 ( .A(f1_round_9_io_state_out_0_1), .B(
        f1_round_10_t_n19), .Z(f1_round_10_p_io_state_out_1_3) );
  XOR2_X1 f1_round_10_t_U39 ( .A(f1_round_9_io_state_out_0_2), .B(
        f1_round_10_t_n19), .Z(f1_round_10_p_io_state_out_2_1) );
  XOR2_X1 f1_round_10_t_U38 ( .A(f1_round_9_io_state_out_0_3), .B(
        f1_round_10_t_n19), .Z(f1_round_10_p_io_state_out_3_4) );
  XOR2_X1 f1_round_10_t_U37 ( .A(f1_round_9_io_state_out_0_4), .B(
        f1_round_10_t_n19), .Z(f1_round_10_p_io_state_out_4_2) );
  XOR2_X1 f1_round_10_t_U36 ( .A(f1_round_9_io_state_out_2_4), .B(
        f1_round_9_io_state_out_2_3), .Z(f1_round_10_t_n18) );
  XNOR2_X1 f1_round_10_t_U35 ( .A(f1_round_9_io_state_out_2_2), .B(
        f1_round_10_t_n18), .ZN(f1_round_10_t_n16) );
  XOR2_X1 f1_round_10_t_U34 ( .A(f1_round_9_io_state_out_2_1), .B(
        f1_round_9_io_state_out_2_0), .Z(f1_round_10_t_n17) );
  XNOR2_X1 f1_round_10_t_U33 ( .A(f1_round_10_t_n16), .B(f1_round_10_t_n17), 
        .ZN(f1_round_10_t_n6) );
  XOR2_X1 f1_round_10_t_U32 ( .A(f1_round_9_io_state_out_0_4), .B(
        f1_round_9_io_state_out_0_3), .Z(f1_round_10_t_n15) );
  XNOR2_X1 f1_round_10_t_U31 ( .A(f1_round_9_io_state_out_0_2), .B(
        f1_round_10_t_n15), .ZN(f1_round_10_t_n13) );
  XOR2_X1 f1_round_10_t_U30 ( .A(f1_round_9_io_state_out_0_1), .B(
        f1_round_9_io_state_out_0_0), .Z(f1_round_10_t_n14) );
  XNOR2_X1 f1_round_10_t_U29 ( .A(f1_round_10_t_n13), .B(f1_round_10_t_n14), 
        .ZN(f1_round_10_t_n2) );
  XOR2_X1 f1_round_10_t_U28 ( .A(f1_round_10_t_n6), .B(f1_round_10_t_n2), .Z(
        f1_round_10_t_n12) );
  XOR2_X1 f1_round_10_t_U27 ( .A(f1_round_9_io_state_out_1_0), .B(
        f1_round_10_t_n12), .Z(f1_round_10_p_io_state_out_0_2) );
  XOR2_X1 f1_round_10_t_U26 ( .A(f1_round_9_io_state_out_1_1), .B(
        f1_round_10_t_n12), .Z(f1_round_10_p_io_state_out_1_0) );
  XOR2_X1 f1_round_10_t_U25 ( .A(f1_round_9_io_state_out_1_2), .B(
        f1_round_10_t_n12), .Z(f1_round_10_p_io_state_out_2_3) );
  XOR2_X1 f1_round_10_t_U24 ( .A(f1_round_9_io_state_out_1_3), .B(
        f1_round_10_t_n12), .Z(f1_round_10_p_io_state_out_3_1) );
  XOR2_X1 f1_round_10_t_U23 ( .A(f1_round_9_io_state_out_1_4), .B(
        f1_round_10_t_n12), .Z(f1_round_10_p_io_state_out_4_4) );
  XOR2_X1 f1_round_10_t_U22 ( .A(f1_round_9_io_state_out_3_4), .B(
        f1_round_9_io_state_out_3_3), .Z(f1_round_10_t_n11) );
  XNOR2_X1 f1_round_10_t_U21 ( .A(f1_round_9_io_state_out_3_2), .B(
        f1_round_10_t_n11), .ZN(f1_round_10_t_n9) );
  XOR2_X1 f1_round_10_t_U20 ( .A(f1_round_9_io_state_out_3_1), .B(
        f1_round_9_io_state_out_3_0), .Z(f1_round_10_t_n10) );
  XNOR2_X1 f1_round_10_t_U19 ( .A(f1_round_10_t_n9), .B(f1_round_10_t_n10), 
        .ZN(f1_round_10_t_n3) );
  XNOR2_X1 f1_round_10_t_U18 ( .A(f1_round_10_t_n8), .B(f1_round_10_t_n3), 
        .ZN(f1_round_10_t_n7) );
  XOR2_X1 f1_round_10_t_U17 ( .A(f1_round_9_io_state_out_2_0), .B(
        f1_round_10_t_n7), .Z(f1_round_10_p_io_state_out_0_4) );
  XOR2_X1 f1_round_10_t_U16 ( .A(f1_round_9_io_state_out_2_1), .B(
        f1_round_10_t_n7), .Z(f1_round_10_p_io_state_out_1_2) );
  XOR2_X1 f1_round_10_t_U15 ( .A(f1_round_9_io_state_out_2_2), .B(
        f1_round_10_t_n7), .Z(f1_round_10_p_io_state_out_2_0) );
  XOR2_X1 f1_round_10_t_U14 ( .A(f1_round_9_io_state_out_2_3), .B(
        f1_round_10_t_n7), .Z(f1_round_10_p_io_state_out_3_3) );
  XOR2_X1 f1_round_10_t_U13 ( .A(f1_round_9_io_state_out_2_4), .B(
        f1_round_10_t_n7), .Z(f1_round_10_p_io_state_out_4_1) );
  XOR2_X1 f1_round_10_t_U12 ( .A(f1_round_10_t_n5), .B(f1_round_10_t_n6), .Z(
        f1_round_10_t_n4) );
  XOR2_X1 f1_round_10_t_U11 ( .A(f1_round_9_io_state_out_3_0), .B(
        f1_round_10_t_n4), .Z(f1_round_10_p_io_state_out_0_1) );
  XOR2_X1 f1_round_10_t_U10 ( .A(f1_round_9_io_state_out_3_1), .B(
        f1_round_10_t_n4), .Z(f1_round_10_p_io_state_out_1_4) );
  XOR2_X1 f1_round_10_t_U9 ( .A(f1_round_9_io_state_out_3_2), .B(
        f1_round_10_t_n4), .Z(f1_round_10_p_io_state_out_2_2) );
  XOR2_X1 f1_round_10_t_U8 ( .A(f1_round_9_io_state_out_3_3), .B(
        f1_round_10_t_n4), .Z(f1_round_10_p_io_state_out_3_0) );
  XOR2_X1 f1_round_10_t_U7 ( .A(f1_round_9_io_state_out_3_4), .B(
        f1_round_10_t_n4), .Z(f1_round_10_p_io_state_out_4_3) );
  XOR2_X1 f1_round_10_t_U6 ( .A(f1_round_10_t_n2), .B(f1_round_10_t_n3), .Z(
        f1_round_10_t_n1) );
  XOR2_X1 f1_round_10_t_U5 ( .A(f1_round_9_io_state_out_4_0), .B(
        f1_round_10_t_n1), .Z(f1_round_10_p_io_state_out_0_3) );
  XOR2_X1 f1_round_10_t_U4 ( .A(f1_round_9_io_state_out_4_1), .B(
        f1_round_10_t_n1), .Z(f1_round_10_p_io_state_out_1_1) );
  XOR2_X1 f1_round_10_t_U3 ( .A(f1_round_9_io_state_out_4_2), .B(
        f1_round_10_t_n1), .Z(f1_round_10_p_io_state_out_2_4) );
  XOR2_X1 f1_round_10_t_U2 ( .A(f1_round_9_io_state_out_4_3), .B(
        f1_round_10_t_n1), .Z(f1_round_10_p_io_state_out_3_2) );
  XOR2_X1 f1_round_10_t_U1 ( .A(f1_round_9_io_state_out_4_4), .B(
        f1_round_10_t_n1), .Z(f1_round_10_p_io_state_out_4_0) );
  NAND2_X1 f1_round_10_c_U50 ( .A1(f1_round_10_p_io_state_out_2_0), .A2(
        f1_round_10_p_io_state_out_1_0), .ZN(f1_round_10_c_n25) );
  XOR2_X1 f1_round_10_c_U49 ( .A(f1_round_10_c_n25), .B(
        f1_round_10_p_io_state_out_0_0), .Z(f1_round_10_c_io_state_out_0_0) );
  NAND2_X1 f1_round_10_c_U48 ( .A1(f1_round_10_p_io_state_out_2_1), .A2(
        f1_round_10_p_io_state_out_1_1), .ZN(f1_round_10_c_n24) );
  XOR2_X1 f1_round_10_c_U47 ( .A(f1_round_10_c_n24), .B(
        f1_round_10_p_io_state_out_0_1), .Z(f1_round_10_io_state_out_0_1) );
  NAND2_X1 f1_round_10_c_U46 ( .A1(f1_round_10_p_io_state_out_2_2), .A2(
        f1_round_10_p_io_state_out_1_2), .ZN(f1_round_10_c_n23) );
  XOR2_X1 f1_round_10_c_U45 ( .A(f1_round_10_c_n23), .B(
        f1_round_10_p_io_state_out_0_2), .Z(f1_round_10_io_state_out_0_2) );
  NAND2_X1 f1_round_10_c_U44 ( .A1(f1_round_10_p_io_state_out_2_3), .A2(
        f1_round_10_p_io_state_out_1_3), .ZN(f1_round_10_c_n22) );
  XOR2_X1 f1_round_10_c_U43 ( .A(f1_round_10_c_n22), .B(
        f1_round_10_p_io_state_out_0_3), .Z(f1_round_10_io_state_out_0_3) );
  NAND2_X1 f1_round_10_c_U42 ( .A1(f1_round_10_p_io_state_out_2_4), .A2(
        f1_round_10_p_io_state_out_1_4), .ZN(f1_round_10_c_n21) );
  XOR2_X1 f1_round_10_c_U41 ( .A(f1_round_10_c_n21), .B(
        f1_round_10_p_io_state_out_0_4), .Z(f1_round_10_io_state_out_0_4) );
  NAND2_X1 f1_round_10_c_U40 ( .A1(f1_round_10_p_io_state_out_2_0), .A2(
        f1_round_10_p_io_state_out_3_0), .ZN(f1_round_10_c_n20) );
  XOR2_X1 f1_round_10_c_U39 ( .A(f1_round_10_c_n20), .B(
        f1_round_10_p_io_state_out_1_0), .Z(f1_round_10_io_state_out_1_0) );
  NAND2_X1 f1_round_10_c_U38 ( .A1(f1_round_10_p_io_state_out_2_1), .A2(
        f1_round_10_p_io_state_out_3_1), .ZN(f1_round_10_c_n19) );
  XOR2_X1 f1_round_10_c_U37 ( .A(f1_round_10_c_n19), .B(
        f1_round_10_p_io_state_out_1_1), .Z(f1_round_10_io_state_out_1_1) );
  NAND2_X1 f1_round_10_c_U36 ( .A1(f1_round_10_p_io_state_out_2_2), .A2(
        f1_round_10_p_io_state_out_3_2), .ZN(f1_round_10_c_n18) );
  XOR2_X1 f1_round_10_c_U35 ( .A(f1_round_10_c_n18), .B(
        f1_round_10_p_io_state_out_1_2), .Z(f1_round_10_io_state_out_1_2) );
  NAND2_X1 f1_round_10_c_U34 ( .A1(f1_round_10_p_io_state_out_2_3), .A2(
        f1_round_10_p_io_state_out_3_3), .ZN(f1_round_10_c_n17) );
  XOR2_X1 f1_round_10_c_U33 ( .A(f1_round_10_c_n17), .B(
        f1_round_10_p_io_state_out_1_3), .Z(f1_round_10_io_state_out_1_3) );
  NAND2_X1 f1_round_10_c_U32 ( .A1(f1_round_10_p_io_state_out_2_4), .A2(
        f1_round_10_p_io_state_out_3_4), .ZN(f1_round_10_c_n16) );
  XOR2_X1 f1_round_10_c_U31 ( .A(f1_round_10_c_n16), .B(
        f1_round_10_p_io_state_out_1_4), .Z(f1_round_10_io_state_out_1_4) );
  NAND2_X1 f1_round_10_c_U30 ( .A1(f1_round_10_p_io_state_out_3_0), .A2(
        f1_round_10_p_io_state_out_4_0), .ZN(f1_round_10_c_n15) );
  XOR2_X1 f1_round_10_c_U29 ( .A(f1_round_10_c_n15), .B(
        f1_round_10_p_io_state_out_2_0), .Z(f1_round_10_io_state_out_2_0) );
  NAND2_X1 f1_round_10_c_U28 ( .A1(f1_round_10_p_io_state_out_3_1), .A2(
        f1_round_10_p_io_state_out_4_1), .ZN(f1_round_10_c_n14) );
  XOR2_X1 f1_round_10_c_U27 ( .A(f1_round_10_c_n14), .B(
        f1_round_10_p_io_state_out_2_1), .Z(f1_round_10_io_state_out_2_1) );
  NAND2_X1 f1_round_10_c_U26 ( .A1(f1_round_10_p_io_state_out_3_2), .A2(
        f1_round_10_p_io_state_out_4_2), .ZN(f1_round_10_c_n13) );
  XOR2_X1 f1_round_10_c_U25 ( .A(f1_round_10_c_n13), .B(
        f1_round_10_p_io_state_out_2_2), .Z(f1_round_10_io_state_out_2_2) );
  NAND2_X1 f1_round_10_c_U24 ( .A1(f1_round_10_p_io_state_out_3_3), .A2(
        f1_round_10_p_io_state_out_4_3), .ZN(f1_round_10_c_n12) );
  XOR2_X1 f1_round_10_c_U23 ( .A(f1_round_10_c_n12), .B(
        f1_round_10_p_io_state_out_2_3), .Z(f1_round_10_io_state_out_2_3) );
  NAND2_X1 f1_round_10_c_U22 ( .A1(f1_round_10_p_io_state_out_3_4), .A2(
        f1_round_10_p_io_state_out_4_4), .ZN(f1_round_10_c_n11) );
  XOR2_X1 f1_round_10_c_U21 ( .A(f1_round_10_c_n11), .B(
        f1_round_10_p_io_state_out_2_4), .Z(f1_round_10_io_state_out_2_4) );
  NAND2_X1 f1_round_10_c_U20 ( .A1(f1_round_10_p_io_state_out_4_0), .A2(
        f1_round_10_p_io_state_out_0_0), .ZN(f1_round_10_c_n10) );
  XOR2_X1 f1_round_10_c_U19 ( .A(f1_round_10_c_n10), .B(
        f1_round_10_p_io_state_out_3_0), .Z(f1_round_10_io_state_out_3_0) );
  NAND2_X1 f1_round_10_c_U18 ( .A1(f1_round_10_p_io_state_out_4_1), .A2(
        f1_round_10_p_io_state_out_0_1), .ZN(f1_round_10_c_n9) );
  XOR2_X1 f1_round_10_c_U17 ( .A(f1_round_10_c_n9), .B(
        f1_round_10_p_io_state_out_3_1), .Z(f1_round_10_io_state_out_3_1) );
  NAND2_X1 f1_round_10_c_U16 ( .A1(f1_round_10_p_io_state_out_4_2), .A2(
        f1_round_10_p_io_state_out_0_2), .ZN(f1_round_10_c_n8) );
  XOR2_X1 f1_round_10_c_U15 ( .A(f1_round_10_c_n8), .B(
        f1_round_10_p_io_state_out_3_2), .Z(f1_round_10_io_state_out_3_2) );
  NAND2_X1 f1_round_10_c_U14 ( .A1(f1_round_10_p_io_state_out_4_3), .A2(
        f1_round_10_p_io_state_out_0_3), .ZN(f1_round_10_c_n7) );
  XOR2_X1 f1_round_10_c_U13 ( .A(f1_round_10_c_n7), .B(
        f1_round_10_p_io_state_out_3_3), .Z(f1_round_10_io_state_out_3_3) );
  NAND2_X1 f1_round_10_c_U12 ( .A1(f1_round_10_p_io_state_out_4_4), .A2(
        f1_round_10_p_io_state_out_0_4), .ZN(f1_round_10_c_n6) );
  XOR2_X1 f1_round_10_c_U11 ( .A(f1_round_10_c_n6), .B(
        f1_round_10_p_io_state_out_3_4), .Z(f1_round_10_io_state_out_3_4) );
  NAND2_X1 f1_round_10_c_U10 ( .A1(f1_round_10_p_io_state_out_1_0), .A2(
        f1_round_10_p_io_state_out_0_0), .ZN(f1_round_10_c_n5) );
  XOR2_X1 f1_round_10_c_U9 ( .A(f1_round_10_c_n5), .B(
        f1_round_10_p_io_state_out_4_0), .Z(f1_round_10_io_state_out_4_0) );
  NAND2_X1 f1_round_10_c_U8 ( .A1(f1_round_10_p_io_state_out_1_1), .A2(
        f1_round_10_p_io_state_out_0_1), .ZN(f1_round_10_c_n4) );
  XOR2_X1 f1_round_10_c_U7 ( .A(f1_round_10_c_n4), .B(
        f1_round_10_p_io_state_out_4_1), .Z(f1_round_10_io_state_out_4_1) );
  NAND2_X1 f1_round_10_c_U6 ( .A1(f1_round_10_p_io_state_out_1_2), .A2(
        f1_round_10_p_io_state_out_0_2), .ZN(f1_round_10_c_n3) );
  XOR2_X1 f1_round_10_c_U5 ( .A(f1_round_10_c_n3), .B(
        f1_round_10_p_io_state_out_4_2), .Z(f1_round_10_io_state_out_4_2) );
  NAND2_X1 f1_round_10_c_U4 ( .A1(f1_round_10_p_io_state_out_1_3), .A2(
        f1_round_10_p_io_state_out_0_3), .ZN(f1_round_10_c_n2) );
  XOR2_X1 f1_round_10_c_U3 ( .A(f1_round_10_c_n2), .B(
        f1_round_10_p_io_state_out_4_3), .Z(f1_round_10_io_state_out_4_3) );
  NAND2_X1 f1_round_10_c_U2 ( .A1(f1_round_10_p_io_state_out_1_4), .A2(
        f1_round_10_p_io_state_out_0_4), .ZN(f1_round_10_c_n1) );
  XOR2_X1 f1_round_10_c_U1 ( .A(f1_round_10_c_n1), .B(
        f1_round_10_p_io_state_out_4_4), .Z(f1_round_10_io_state_out_4_4) );
  INV_X1 f1_round_10_i_U1 ( .A(f1_round_10_c_io_state_out_0_0), .ZN(
        f1_round_10_io_state_out_0_0) );
  XOR2_X1 f1_round_11_t_U50 ( .A(f1_round_10_io_state_out_1_4), .B(
        f1_round_10_io_state_out_1_3), .Z(f1_round_11_t_n25) );
  XNOR2_X1 f1_round_11_t_U49 ( .A(f1_round_10_io_state_out_1_2), .B(
        f1_round_11_t_n25), .ZN(f1_round_11_t_n23) );
  XOR2_X1 f1_round_11_t_U48 ( .A(f1_round_10_io_state_out_1_1), .B(
        f1_round_10_io_state_out_1_0), .Z(f1_round_11_t_n24) );
  XOR2_X1 f1_round_11_t_U47 ( .A(f1_round_11_t_n23), .B(f1_round_11_t_n24), 
        .Z(f1_round_11_t_n8) );
  XOR2_X1 f1_round_11_t_U46 ( .A(f1_round_10_io_state_out_4_4), .B(
        f1_round_10_io_state_out_4_3), .Z(f1_round_11_t_n22) );
  XNOR2_X1 f1_round_11_t_U45 ( .A(f1_round_10_io_state_out_4_2), .B(
        f1_round_11_t_n22), .ZN(f1_round_11_t_n20) );
  XOR2_X1 f1_round_11_t_U44 ( .A(f1_round_10_io_state_out_4_1), .B(
        f1_round_10_io_state_out_4_0), .Z(f1_round_11_t_n21) );
  XNOR2_X1 f1_round_11_t_U43 ( .A(f1_round_11_t_n20), .B(f1_round_11_t_n21), 
        .ZN(f1_round_11_t_n5) );
  XNOR2_X1 f1_round_11_t_U42 ( .A(f1_round_11_t_n8), .B(f1_round_11_t_n5), 
        .ZN(f1_round_11_t_n19) );
  XOR2_X1 f1_round_11_t_U41 ( .A(f1_round_10_io_state_out_0_0), .B(
        f1_round_11_t_n19), .Z(f1_round_11_p_io_state_out_0_0) );
  XOR2_X1 f1_round_11_t_U40 ( .A(f1_round_10_io_state_out_0_1), .B(
        f1_round_11_t_n19), .Z(f1_round_11_p_io_state_out_1_3) );
  XOR2_X1 f1_round_11_t_U39 ( .A(f1_round_10_io_state_out_0_2), .B(
        f1_round_11_t_n19), .Z(f1_round_11_p_io_state_out_2_1) );
  XOR2_X1 f1_round_11_t_U38 ( .A(f1_round_10_io_state_out_0_3), .B(
        f1_round_11_t_n19), .Z(f1_round_11_p_io_state_out_3_4) );
  XOR2_X1 f1_round_11_t_U37 ( .A(f1_round_10_io_state_out_0_4), .B(
        f1_round_11_t_n19), .Z(f1_round_11_p_io_state_out_4_2) );
  XOR2_X1 f1_round_11_t_U36 ( .A(f1_round_10_io_state_out_2_4), .B(
        f1_round_10_io_state_out_2_3), .Z(f1_round_11_t_n18) );
  XNOR2_X1 f1_round_11_t_U35 ( .A(f1_round_10_io_state_out_2_2), .B(
        f1_round_11_t_n18), .ZN(f1_round_11_t_n16) );
  XOR2_X1 f1_round_11_t_U34 ( .A(f1_round_10_io_state_out_2_1), .B(
        f1_round_10_io_state_out_2_0), .Z(f1_round_11_t_n17) );
  XNOR2_X1 f1_round_11_t_U33 ( .A(f1_round_11_t_n16), .B(f1_round_11_t_n17), 
        .ZN(f1_round_11_t_n6) );
  XOR2_X1 f1_round_11_t_U32 ( .A(f1_round_10_io_state_out_0_4), .B(
        f1_round_10_io_state_out_0_3), .Z(f1_round_11_t_n15) );
  XNOR2_X1 f1_round_11_t_U31 ( .A(f1_round_10_io_state_out_0_2), .B(
        f1_round_11_t_n15), .ZN(f1_round_11_t_n13) );
  XOR2_X1 f1_round_11_t_U30 ( .A(f1_round_10_io_state_out_0_1), .B(
        f1_round_10_io_state_out_0_0), .Z(f1_round_11_t_n14) );
  XNOR2_X1 f1_round_11_t_U29 ( .A(f1_round_11_t_n13), .B(f1_round_11_t_n14), 
        .ZN(f1_round_11_t_n2) );
  XOR2_X1 f1_round_11_t_U28 ( .A(f1_round_11_t_n6), .B(f1_round_11_t_n2), .Z(
        f1_round_11_t_n12) );
  XOR2_X1 f1_round_11_t_U27 ( .A(f1_round_10_io_state_out_1_0), .B(
        f1_round_11_t_n12), .Z(f1_round_11_p_io_state_out_0_2) );
  XOR2_X1 f1_round_11_t_U26 ( .A(f1_round_10_io_state_out_1_1), .B(
        f1_round_11_t_n12), .Z(f1_round_11_p_io_state_out_1_0) );
  XOR2_X1 f1_round_11_t_U25 ( .A(f1_round_10_io_state_out_1_2), .B(
        f1_round_11_t_n12), .Z(f1_round_11_p_io_state_out_2_3) );
  XOR2_X1 f1_round_11_t_U24 ( .A(f1_round_10_io_state_out_1_3), .B(
        f1_round_11_t_n12), .Z(f1_round_11_p_io_state_out_3_1) );
  XOR2_X1 f1_round_11_t_U23 ( .A(f1_round_10_io_state_out_1_4), .B(
        f1_round_11_t_n12), .Z(f1_round_11_p_io_state_out_4_4) );
  XOR2_X1 f1_round_11_t_U22 ( .A(f1_round_10_io_state_out_3_4), .B(
        f1_round_10_io_state_out_3_3), .Z(f1_round_11_t_n11) );
  XNOR2_X1 f1_round_11_t_U21 ( .A(f1_round_10_io_state_out_3_2), .B(
        f1_round_11_t_n11), .ZN(f1_round_11_t_n9) );
  XOR2_X1 f1_round_11_t_U20 ( .A(f1_round_10_io_state_out_3_1), .B(
        f1_round_10_io_state_out_3_0), .Z(f1_round_11_t_n10) );
  XNOR2_X1 f1_round_11_t_U19 ( .A(f1_round_11_t_n9), .B(f1_round_11_t_n10), 
        .ZN(f1_round_11_t_n3) );
  XNOR2_X1 f1_round_11_t_U18 ( .A(f1_round_11_t_n8), .B(f1_round_11_t_n3), 
        .ZN(f1_round_11_t_n7) );
  XOR2_X1 f1_round_11_t_U17 ( .A(f1_round_10_io_state_out_2_0), .B(
        f1_round_11_t_n7), .Z(f1_round_11_p_io_state_out_0_4) );
  XOR2_X1 f1_round_11_t_U16 ( .A(f1_round_10_io_state_out_2_1), .B(
        f1_round_11_t_n7), .Z(f1_round_11_p_io_state_out_1_2) );
  XOR2_X1 f1_round_11_t_U15 ( .A(f1_round_10_io_state_out_2_2), .B(
        f1_round_11_t_n7), .Z(f1_round_11_p_io_state_out_2_0) );
  XOR2_X1 f1_round_11_t_U14 ( .A(f1_round_10_io_state_out_2_3), .B(
        f1_round_11_t_n7), .Z(f1_round_11_p_io_state_out_3_3) );
  XOR2_X1 f1_round_11_t_U13 ( .A(f1_round_10_io_state_out_2_4), .B(
        f1_round_11_t_n7), .Z(f1_round_11_p_io_state_out_4_1) );
  XOR2_X1 f1_round_11_t_U12 ( .A(f1_round_11_t_n5), .B(f1_round_11_t_n6), .Z(
        f1_round_11_t_n4) );
  XOR2_X1 f1_round_11_t_U11 ( .A(f1_round_10_io_state_out_3_0), .B(
        f1_round_11_t_n4), .Z(f1_round_11_p_io_state_out_0_1) );
  XOR2_X1 f1_round_11_t_U10 ( .A(f1_round_10_io_state_out_3_1), .B(
        f1_round_11_t_n4), .Z(f1_round_11_p_io_state_out_1_4) );
  XOR2_X1 f1_round_11_t_U9 ( .A(f1_round_10_io_state_out_3_2), .B(
        f1_round_11_t_n4), .Z(f1_round_11_p_io_state_out_2_2) );
  XOR2_X1 f1_round_11_t_U8 ( .A(f1_round_10_io_state_out_3_3), .B(
        f1_round_11_t_n4), .Z(f1_round_11_p_io_state_out_3_0) );
  XOR2_X1 f1_round_11_t_U7 ( .A(f1_round_10_io_state_out_3_4), .B(
        f1_round_11_t_n4), .Z(f1_round_11_p_io_state_out_4_3) );
  XOR2_X1 f1_round_11_t_U6 ( .A(f1_round_11_t_n2), .B(f1_round_11_t_n3), .Z(
        f1_round_11_t_n1) );
  XOR2_X1 f1_round_11_t_U5 ( .A(f1_round_10_io_state_out_4_0), .B(
        f1_round_11_t_n1), .Z(f1_round_11_p_io_state_out_0_3) );
  XOR2_X1 f1_round_11_t_U4 ( .A(f1_round_10_io_state_out_4_1), .B(
        f1_round_11_t_n1), .Z(f1_round_11_p_io_state_out_1_1) );
  XOR2_X1 f1_round_11_t_U3 ( .A(f1_round_10_io_state_out_4_2), .B(
        f1_round_11_t_n1), .Z(f1_round_11_p_io_state_out_2_4) );
  XOR2_X1 f1_round_11_t_U2 ( .A(f1_round_10_io_state_out_4_3), .B(
        f1_round_11_t_n1), .Z(f1_round_11_p_io_state_out_3_2) );
  XOR2_X1 f1_round_11_t_U1 ( .A(f1_round_10_io_state_out_4_4), .B(
        f1_round_11_t_n1), .Z(f1_round_11_p_io_state_out_4_0) );
  NAND2_X1 f1_round_11_c_U50 ( .A1(f1_round_11_p_io_state_out_2_0), .A2(
        f1_round_11_p_io_state_out_1_0), .ZN(f1_round_11_c_n25) );
  XOR2_X1 f1_round_11_c_U49 ( .A(f1_round_11_c_n25), .B(
        f1_round_11_p_io_state_out_0_0), .Z(io_block_o0[0]) );
  NAND2_X1 f1_round_11_c_U48 ( .A1(f1_round_11_p_io_state_out_2_1), .A2(
        f1_round_11_p_io_state_out_1_1), .ZN(f1_round_11_c_n24) );
  XOR2_X1 f1_round_11_c_U47 ( .A(f1_round_11_c_n24), .B(
        f1_round_11_p_io_state_out_0_1), .Z(io_block_o0[5]) );
  NAND2_X1 f1_round_11_c_U46 ( .A1(f1_round_11_p_io_state_out_2_2), .A2(
        f1_round_11_p_io_state_out_1_2), .ZN(f1_round_11_c_n23) );
  XOR2_X1 f1_round_11_c_U45 ( .A(f1_round_11_c_n23), .B(
        f1_round_11_p_io_state_out_0_2), .Z(f1_round_11_c_io_state_out_0_2) );
  NAND2_X1 f1_round_11_c_U44 ( .A1(f1_round_11_p_io_state_out_2_3), .A2(
        f1_round_11_p_io_state_out_1_3), .ZN(f1_round_11_c_n22) );
  XOR2_X1 f1_round_11_c_U43 ( .A(f1_round_11_c_n22), .B(
        f1_round_11_p_io_state_out_0_3), .Z(f1_round_11_c_io_state_out_0_3) );
  NAND2_X1 f1_round_11_c_U42 ( .A1(f1_round_11_p_io_state_out_2_4), .A2(
        f1_round_11_p_io_state_out_1_4), .ZN(f1_round_11_c_n21) );
  XOR2_X1 f1_round_11_c_U41 ( .A(f1_round_11_c_n21), .B(
        f1_round_11_p_io_state_out_0_4), .Z(f1_round_11_c_io_state_out_0_4) );
  NAND2_X1 f1_round_11_c_U40 ( .A1(f1_round_11_p_io_state_out_2_0), .A2(
        f1_round_11_p_io_state_out_3_0), .ZN(f1_round_11_c_n20) );
  XOR2_X1 f1_round_11_c_U39 ( .A(f1_round_11_c_n20), .B(
        f1_round_11_p_io_state_out_1_0), .Z(io_block_o0[1]) );
  NAND2_X1 f1_round_11_c_U38 ( .A1(f1_round_11_p_io_state_out_2_1), .A2(
        f1_round_11_p_io_state_out_3_1), .ZN(f1_round_11_c_n19) );
  XOR2_X1 f1_round_11_c_U37 ( .A(f1_round_11_c_n19), .B(
        f1_round_11_p_io_state_out_1_1), .Z(io_block_o0[6]) );
  NAND2_X1 f1_round_11_c_U36 ( .A1(f1_round_11_p_io_state_out_2_2), .A2(
        f1_round_11_p_io_state_out_3_2), .ZN(f1_round_11_c_n18) );
  XOR2_X1 f1_round_11_c_U35 ( .A(f1_round_11_c_n18), .B(
        f1_round_11_p_io_state_out_1_2), .Z(f1_round_11_c_io_state_out_1_2) );
  NAND2_X1 f1_round_11_c_U34 ( .A1(f1_round_11_p_io_state_out_2_3), .A2(
        f1_round_11_p_io_state_out_3_3), .ZN(f1_round_11_c_n17) );
  XOR2_X1 f1_round_11_c_U33 ( .A(f1_round_11_c_n17), .B(
        f1_round_11_p_io_state_out_1_3), .Z(f1_round_11_c_io_state_out_1_3) );
  NAND2_X1 f1_round_11_c_U32 ( .A1(f1_round_11_p_io_state_out_2_4), .A2(
        f1_round_11_p_io_state_out_3_4), .ZN(f1_round_11_c_n16) );
  XOR2_X1 f1_round_11_c_U31 ( .A(f1_round_11_c_n16), .B(
        f1_round_11_p_io_state_out_1_4), .Z(f1_round_11_c_io_state_out_1_4) );
  NAND2_X1 f1_round_11_c_U30 ( .A1(f1_round_11_p_io_state_out_3_0), .A2(
        f1_round_11_p_io_state_out_4_0), .ZN(f1_round_11_c_n15) );
  XOR2_X1 f1_round_11_c_U29 ( .A(f1_round_11_c_n15), .B(
        f1_round_11_p_io_state_out_2_0), .Z(io_block_o0[2]) );
  NAND2_X1 f1_round_11_c_U28 ( .A1(f1_round_11_p_io_state_out_3_1), .A2(
        f1_round_11_p_io_state_out_4_1), .ZN(f1_round_11_c_n14) );
  XOR2_X1 f1_round_11_c_U27 ( .A(f1_round_11_c_n14), .B(
        f1_round_11_p_io_state_out_2_1), .Z(io_block_o0[7]) );
  NAND2_X1 f1_round_11_c_U26 ( .A1(f1_round_11_p_io_state_out_3_2), .A2(
        f1_round_11_p_io_state_out_4_2), .ZN(f1_round_11_c_n13) );
  XOR2_X1 f1_round_11_c_U25 ( .A(f1_round_11_c_n13), .B(
        f1_round_11_p_io_state_out_2_2), .Z(f1_round_11_c_io_state_out_2_2) );
  NAND2_X1 f1_round_11_c_U24 ( .A1(f1_round_11_p_io_state_out_3_3), .A2(
        f1_round_11_p_io_state_out_4_3), .ZN(f1_round_11_c_n12) );
  XOR2_X1 f1_round_11_c_U23 ( .A(f1_round_11_c_n12), .B(
        f1_round_11_p_io_state_out_2_3), .Z(f1_round_11_c_io_state_out_2_3) );
  NAND2_X1 f1_round_11_c_U22 ( .A1(f1_round_11_p_io_state_out_3_4), .A2(
        f1_round_11_p_io_state_out_4_4), .ZN(f1_round_11_c_n11) );
  XOR2_X1 f1_round_11_c_U21 ( .A(f1_round_11_c_n11), .B(
        f1_round_11_p_io_state_out_2_4), .Z(f1_round_11_c_io_state_out_2_4) );
  NAND2_X1 f1_round_11_c_U20 ( .A1(f1_round_11_p_io_state_out_4_0), .A2(
        f1_round_11_p_io_state_out_0_0), .ZN(f1_round_11_c_n10) );
  XOR2_X1 f1_round_11_c_U19 ( .A(f1_round_11_c_n10), .B(
        f1_round_11_p_io_state_out_3_0), .Z(io_block_o0[3]) );
  NAND2_X1 f1_round_11_c_U18 ( .A1(f1_round_11_p_io_state_out_4_1), .A2(
        f1_round_11_p_io_state_out_0_1), .ZN(f1_round_11_c_n9) );
  XOR2_X1 f1_round_11_c_U17 ( .A(f1_round_11_c_n9), .B(
        f1_round_11_p_io_state_out_3_1), .Z(io_block_o0[8]) );
  NAND2_X1 f1_round_11_c_U16 ( .A1(f1_round_11_p_io_state_out_4_2), .A2(
        f1_round_11_p_io_state_out_0_2), .ZN(f1_round_11_c_n8) );
  XOR2_X1 f1_round_11_c_U15 ( .A(f1_round_11_c_n8), .B(
        f1_round_11_p_io_state_out_3_2), .Z(f1_round_11_c_io_state_out_3_2) );
  NAND2_X1 f1_round_11_c_U14 ( .A1(f1_round_11_p_io_state_out_4_3), .A2(
        f1_round_11_p_io_state_out_0_3), .ZN(f1_round_11_c_n7) );
  XOR2_X1 f1_round_11_c_U13 ( .A(f1_round_11_c_n7), .B(
        f1_round_11_p_io_state_out_3_3), .Z(f1_round_11_c_io_state_out_3_3) );
  NAND2_X1 f1_round_11_c_U12 ( .A1(f1_round_11_p_io_state_out_4_4), .A2(
        f1_round_11_p_io_state_out_0_4), .ZN(f1_round_11_c_n6) );
  XOR2_X1 f1_round_11_c_U11 ( .A(f1_round_11_c_n6), .B(
        f1_round_11_p_io_state_out_3_4), .Z(f1_round_11_c_io_state_out_3_4) );
  NAND2_X1 f1_round_11_c_U10 ( .A1(f1_round_11_p_io_state_out_1_0), .A2(
        f1_round_11_p_io_state_out_0_0), .ZN(f1_round_11_c_n5) );
  XOR2_X1 f1_round_11_c_U9 ( .A(f1_round_11_c_n5), .B(
        f1_round_11_p_io_state_out_4_0), .Z(io_block_o0[4]) );
  NAND2_X1 f1_round_11_c_U8 ( .A1(f1_round_11_p_io_state_out_1_1), .A2(
        f1_round_11_p_io_state_out_0_1), .ZN(f1_round_11_c_n4) );
  XOR2_X1 f1_round_11_c_U7 ( .A(f1_round_11_c_n4), .B(
        f1_round_11_p_io_state_out_4_1), .Z(io_block_o0[9]) );
  NAND2_X1 f1_round_11_c_U6 ( .A1(f1_round_11_p_io_state_out_1_2), .A2(
        f1_round_11_p_io_state_out_0_2), .ZN(f1_round_11_c_n3) );
  XOR2_X1 f1_round_11_c_U5 ( .A(f1_round_11_c_n3), .B(
        f1_round_11_p_io_state_out_4_2), .Z(f1_round_11_c_io_state_out_4_2) );
  NAND2_X1 f1_round_11_c_U4 ( .A1(f1_round_11_p_io_state_out_1_3), .A2(
        f1_round_11_p_io_state_out_0_3), .ZN(f1_round_11_c_n2) );
  XOR2_X1 f1_round_11_c_U3 ( .A(f1_round_11_c_n2), .B(
        f1_round_11_p_io_state_out_4_3), .Z(f1_round_11_c_io_state_out_4_3) );
  NAND2_X1 f1_round_11_c_U2 ( .A1(f1_round_11_p_io_state_out_1_4), .A2(
        f1_round_11_p_io_state_out_0_4), .ZN(f1_round_11_c_n1) );
  XOR2_X1 f1_round_11_c_U1 ( .A(f1_round_11_c_n1), .B(
        f1_round_11_p_io_state_out_4_4), .Z(f1_round_11_c_io_state_out_4_4) );
endmodule

