
module Sbox_opt ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i1_s0, io_i1_s1, 
        io_i2_s0, io_i2_s1, io_i3_s0, io_i3_s1, io_i4_s0, io_i4_s1, io_i5_s0, 
        io_i5_s1, io_i6_s0, io_i6_s1, io_i7_s0, io_i7_s1, io_k0_s0, io_k0_s1, 
        io_k1_s0, io_k1_s1, io_k2_s0, io_k2_s1, io_k3_s0, io_k3_s1, io_k4_s0, 
        io_k4_s1, io_k5_s0, io_k5_s1, io_k6_s0, io_k6_s1, io_k7_s0, io_k7_s1, 
        p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, 
        p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12, 
        p_rand_13, p_rand_14, p_rand_15, p_rand_16, p_rand_17, p_rand_18, 
        p_rand_19, p_rand_20, p_rand_21, p_rand_22, p_rand_23, p_rand_24, 
        p_rand_25, p_rand_26, p_rand_27, p_rand_28, p_rand_29, p_rand_30, 
        p_rand_31, p_rand_32, p_rand_33, io_o0_s0, io_o0_s1, io_o1_s0, 
        io_o1_s1, io_o2_s0, io_o2_s1, io_o3_s0, io_o3_s1, io_o4_s0, io_o4_s1, 
        io_o5_s0, io_o5_s1, io_o6_s0, io_o6_s1, io_o7_s0, io_o7_s1 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i1_s0, io_i1_s1, io_i2_s0,
         io_i2_s1, io_i3_s0, io_i3_s1, io_i4_s0, io_i4_s1, io_i5_s0, io_i5_s1,
         io_i6_s0, io_i6_s1, io_i7_s0, io_i7_s1, io_k0_s0, io_k0_s1, io_k1_s0,
         io_k1_s1, io_k2_s0, io_k2_s1, io_k3_s0, io_k3_s1, io_k4_s0, io_k4_s1,
         io_k5_s0, io_k5_s1, io_k6_s0, io_k6_s1, io_k7_s0, io_k7_s1, p_rand_0,
         p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6, p_rand_7,
         p_rand_8, p_rand_9, p_rand_10, p_rand_11, p_rand_12, p_rand_13,
         p_rand_14, p_rand_15, p_rand_16, p_rand_17, p_rand_18, p_rand_19,
         p_rand_20, p_rand_21, p_rand_22, p_rand_23, p_rand_24, p_rand_25,
         p_rand_26, p_rand_27, p_rand_28, p_rand_29, p_rand_30, p_rand_31,
         p_rand_32, p_rand_33;
  output io_o0_s0, io_o0_s1, io_o1_s0, io_o1_s1, io_o2_s0, io_o2_s1, io_o3_s0,
         io_o3_s1, io_o4_s0, io_o4_s1, io_o5_s0, io_o5_s1, io_o6_s0, io_o6_s1,
         io_o7_s0, io_o7_s1;
  wire   n_xor_module_1_res, n_xor_module_2_res, n_xor_module_3_res,
         n_xor_module_4_res, n_xor_module_5_res, n_xor_module_6_res,
         n_xor_module_7_res, n_xor_module_8_res, n_xor_module_9_res,
         n_xor_module_10_res, n_xor_module_11_res, n_xor_module_12_res,
         n_xor_module_13_res, n_xor_module_14_res, n_xor_module_15_res,
         n_xor_module_16_res, n_xor_module_17_res, n_xor_module_18_res,
         n_xor_module_19_res, n_xor_module_20_res, n_xor_module_21_res,
         n_xor_module_22_res, n_xor_module_23_res, n_xor_module_24_res,
         n_xor_module_25_res, n_xor_module_26_res, n_xor_module_27_res,
         n_xor_module_28_res, n_xor_module_29_res, n_xor_module_30_res,
         n_xor_module_31_res, n_xor_module_32_res, n_xor_module_33_res,
         n_xor_module_34_res, n_xor_module_35_res, n_xor_module_36_res,
         n_xor_module_37_res, n_xor_module_38_res, n_xor_module_39_res,
         n_xor_module_40_res, n_xor_module_41_res, n_xor_module_42_res,
         n_xor_module_43_res, n_xor_module_44_res, n_xor_module_45_res,
         n_xor_module_46_res, n_xor_module_47_res, n_xor_module_48_res,
         n_xor_module_49_res, n_xor_module_50_res, n_xor_module_51_res,
         n_xor_module_52_res, n_xor_module_53_res, n_xor_module_54_res,
         n_reg_module_1_res, n_not_module_1_res, n_and_module_1_res,
         n_xor_module_55_res, n_not_module_2_res, n_and_module_2_res,
         n_xor_module_56_res, n_reg_module_2_res, n_and_module_3_res,
         n_reg_module_3_res, n_reg_module_4_res, n_and_module_4_res,
         n_reg_module_5_res, n_reg_module_6_res, n_xor_module_57_res,
         n_xor_module_58_res, n_reg_module_7_res, n_and_module_5_res,
         n_reg_module_8_res, n_reg_module_9_res, n_and_module_6_res,
         n_reg_module_10_res, n_reg_module_11_res, n_xor_module_59_res,
         n_xor_module_60_res, n_reg_module_12_res, n_not_module_3_res,
         n_and_module_7_res, n_xor_module_61_res, n_not_module_4_res,
         n_and_module_8_res, n_xor_module_62_res, n_reg_module_13_res,
         n_and_module_9_res, n_reg_module_14_res, n_reg_module_15_res,
         n_and_module_10_res, n_reg_module_16_res, n_reg_module_17_res,
         n_xor_module_63_res, n_xor_module_64_res, n_reg_module_18_res,
         n_and_module_11_res, n_reg_module_19_res, n_reg_module_20_res,
         n_and_module_12_res, n_reg_module_21_res, n_reg_module_22_res,
         n_xor_module_65_res, n_xor_module_66_res, n_xor_module_67_res,
         n_xor_module_68_res, n_reg_module_23_res, n_not_module_5_res,
         n_and_module_13_res, n_xor_module_69_res, n_not_module_6_res,
         n_and_module_14_res, n_xor_module_70_res, n_reg_module_24_res,
         n_and_module_15_res, n_reg_module_25_res, n_reg_module_26_res,
         n_and_module_16_res, n_reg_module_27_res, n_reg_module_28_res,
         n_xor_module_71_res, n_xor_module_72_res, n_reg_module_29_res,
         n_and_module_17_res, n_reg_module_30_res, n_reg_module_31_res,
         n_and_module_18_res, n_reg_module_32_res, n_reg_module_33_res,
         n_xor_module_73_res, n_xor_module_74_res, n_xor_module_75_res,
         n_xor_module_76_res, n_reg_module_34_res, n_not_module_7_res,
         n_and_module_19_res, n_xor_module_77_res, n_not_module_8_res,
         n_and_module_20_res, n_xor_module_78_res, n_reg_module_35_res,
         n_and_module_21_res, n_reg_module_36_res, n_reg_module_37_res,
         n_and_module_22_res, n_reg_module_38_res, n_reg_module_39_res,
         n_xor_module_79_res, n_xor_module_80_res, n_reg_module_40_res,
         n_and_module_23_res, n_reg_module_41_res, n_reg_module_42_res,
         n_and_module_24_res, n_reg_module_43_res, n_reg_module_44_res,
         n_xor_module_81_res, n_xor_module_82_res, n_reg_module_45_res,
         n_not_module_9_res, n_and_module_25_res, n_xor_module_83_res,
         n_not_module_10_res, n_and_module_26_res, n_xor_module_84_res,
         n_reg_module_46_res, n_and_module_27_res, n_reg_module_47_res,
         n_reg_module_48_res, n_and_module_28_res, n_reg_module_49_res,
         n_reg_module_50_res, n_xor_module_85_res, n_xor_module_86_res,
         n_reg_module_51_res, n_and_module_29_res, n_reg_module_52_res,
         n_reg_module_53_res, n_and_module_30_res, n_reg_module_54_res,
         n_reg_module_55_res, n_xor_module_87_res, n_xor_module_88_res,
         n_xor_module_89_res, n_xor_module_90_res, n_reg_module_56_res,
         n_not_module_11_res, n_and_module_31_res, n_xor_module_91_res,
         n_not_module_12_res, n_and_module_32_res, n_xor_module_92_res,
         n_reg_module_57_res, n_and_module_33_res, n_reg_module_58_res,
         n_reg_module_59_res, n_and_module_34_res, n_reg_module_60_res,
         n_reg_module_61_res, n_xor_module_93_res, n_xor_module_94_res,
         n_reg_module_62_res, n_and_module_35_res, n_reg_module_63_res,
         n_reg_module_64_res, n_and_module_36_res, n_reg_module_65_res,
         n_reg_module_66_res, n_xor_module_95_res, n_xor_module_96_res,
         n_xor_module_97_res, n_xor_module_98_res, n_reg_module_67_res,
         n_not_module_13_res, n_and_module_37_res, n_xor_module_99_res,
         n_not_module_14_res, n_and_module_38_res, n_xor_module_100_res,
         n_reg_module_68_res, n_and_module_39_res, n_reg_module_69_res,
         n_reg_module_70_res, n_and_module_40_res, n_reg_module_71_res,
         n_reg_module_72_res, n_xor_module_101_res, n_xor_module_102_res,
         n_reg_module_73_res, n_and_module_41_res, n_reg_module_74_res,
         n_reg_module_75_res, n_and_module_42_res, n_reg_module_76_res,
         n_reg_module_77_res, n_xor_module_103_res, n_xor_module_104_res,
         n_reg_module_78_res, n_not_module_15_res, n_and_module_43_res,
         n_xor_module_105_res, n_not_module_16_res, n_and_module_44_res,
         n_xor_module_106_res, n_reg_module_79_res, n_and_module_45_res,
         n_reg_module_80_res, n_reg_module_81_res, n_and_module_46_res,
         n_reg_module_82_res, n_reg_module_83_res, n_xor_module_107_res,
         n_xor_module_108_res, n_reg_module_84_res, n_and_module_47_res,
         n_reg_module_85_res, n_reg_module_86_res, n_and_module_48_res,
         n_reg_module_87_res, n_reg_module_88_res, n_xor_module_109_res,
         n_xor_module_110_res, n_xor_module_111_res, n_xor_module_112_res,
         n_reg_module_89_res, n_not_module_17_res, n_and_module_49_res,
         n_xor_module_113_res, n_not_module_18_res, n_and_module_50_res,
         n_xor_module_114_res, n_reg_module_90_res, n_and_module_51_res,
         n_reg_module_91_res, n_reg_module_92_res, n_and_module_52_res,
         n_reg_module_93_res, n_reg_module_94_res, n_xor_module_115_res,
         n_xor_module_116_res, n_reg_module_95_res, n_and_module_53_res,
         n_reg_module_96_res, n_reg_module_97_res, n_and_module_54_res,
         n_reg_module_98_res, n_reg_module_99_res, n_xor_module_117_res,
         n_xor_module_118_res, n_xor_module_119_res, n_xor_module_120_res,
         n_xor_module_121_res, n_xor_module_122_res, n_xor_module_123_res,
         n_xor_module_124_res, n_xor_module_125_res, n_xor_module_126_res,
         n_xor_module_127_res, n_xor_module_128_res, n_xor_module_129_res,
         n_xor_module_130_res, n_xor_module_131_res, n_xor_module_132_res,
         n_xor_module_133_res, n_xor_module_134_res, n_xor_module_135_res,
         n_xor_module_136_res, n_xor_module_137_res, n_xor_module_138_res,
         n_reg_module_100_res, n_not_module_19_res, n_and_module_55_res,
         n_xor_module_139_res, n_not_module_20_res, n_and_module_56_res,
         n_xor_module_140_res, n_reg_module_101_res, n_and_module_57_res,
         n_reg_module_102_res, n_reg_module_103_res, n_and_module_58_res,
         n_reg_module_104_res, n_reg_module_105_res, n_xor_module_141_res,
         n_xor_module_142_res, n_reg_module_106_res, n_and_module_59_res,
         n_reg_module_107_res, n_reg_module_108_res, n_and_module_60_res,
         n_reg_module_109_res, n_reg_module_110_res, n_xor_module_143_res,
         n_xor_module_144_res, n_xor_module_145_res, n_xor_module_146_res,
         n_xor_module_147_res, n_xor_module_148_res, n_xor_module_149_res,
         n_xor_module_150_res, n_reg_module_111_res, n_not_module_21_res,
         n_and_module_61_res, n_xor_module_151_res, n_not_module_22_res,
         n_and_module_62_res, n_xor_module_152_res, n_reg_module_112_res,
         n_and_module_63_res, n_reg_module_113_res, n_reg_module_114_res,
         n_and_module_64_res, n_reg_module_115_res, n_reg_module_116_res,
         n_xor_module_153_res, n_xor_module_154_res, n_reg_module_117_res,
         n_and_module_65_res, n_reg_module_118_res, n_reg_module_119_res,
         n_and_module_66_res, n_reg_module_120_res, n_reg_module_121_res,
         n_xor_module_155_res, n_xor_module_156_res, n_reg_module_122_res,
         n_not_module_23_res, n_and_module_67_res, n_xor_module_157_res,
         n_not_module_24_res, n_and_module_68_res, n_xor_module_158_res,
         n_reg_module_123_res, n_and_module_69_res, n_reg_module_124_res,
         n_reg_module_125_res, n_and_module_70_res, n_reg_module_126_res,
         n_reg_module_127_res, n_xor_module_159_res, n_xor_module_160_res,
         n_reg_module_128_res, n_and_module_71_res, n_reg_module_129_res,
         n_reg_module_130_res, n_and_module_72_res, n_reg_module_131_res,
         n_reg_module_132_res, n_xor_module_161_res, n_xor_module_162_res,
         n_reg_module_133_res, n_not_module_25_res, n_and_module_73_res,
         n_xor_module_163_res, n_not_module_26_res, n_and_module_74_res,
         n_xor_module_164_res, n_reg_module_134_res, n_and_module_75_res,
         n_reg_module_135_res, n_reg_module_136_res, n_and_module_76_res,
         n_reg_module_137_res, n_reg_module_138_res, n_xor_module_165_res,
         n_xor_module_166_res, n_reg_module_139_res, n_and_module_77_res,
         n_reg_module_140_res, n_reg_module_141_res, n_and_module_78_res,
         n_reg_module_142_res, n_reg_module_143_res, n_xor_module_167_res,
         n_xor_module_168_res, n_reg_module_144_res, n_not_module_27_res,
         n_and_module_79_res, n_xor_module_169_res, n_not_module_28_res,
         n_and_module_80_res, n_xor_module_170_res, n_reg_module_145_res,
         n_and_module_81_res, n_reg_module_146_res, n_reg_module_147_res,
         n_and_module_82_res, n_reg_module_148_res, n_reg_module_149_res,
         n_xor_module_171_res, n_xor_module_172_res, n_reg_module_150_res,
         n_and_module_83_res, n_reg_module_151_res, n_reg_module_152_res,
         n_and_module_84_res, n_reg_module_153_res, n_reg_module_154_res,
         n_xor_module_173_res, n_xor_module_174_res, n_xor_module_175_res,
         n_xor_module_176_res, n_reg_module_155_res, n_not_module_29_res,
         n_and_module_85_res, n_xor_module_177_res, n_not_module_30_res,
         n_and_module_86_res, n_xor_module_178_res, n_reg_module_156_res,
         n_and_module_87_res, n_reg_module_157_res, n_reg_module_158_res,
         n_and_module_88_res, n_reg_module_159_res, n_reg_module_160_res,
         n_xor_module_179_res, n_xor_module_180_res, n_reg_module_161_res,
         n_and_module_89_res, n_reg_module_162_res, n_reg_module_163_res,
         n_and_module_90_res, n_reg_module_164_res, n_reg_module_165_res,
         n_xor_module_181_res, n_xor_module_182_res, n_reg_module_166_res,
         n_not_module_31_res, n_and_module_91_res, n_xor_module_183_res,
         n_not_module_32_res, n_and_module_92_res, n_xor_module_184_res,
         n_reg_module_167_res, n_and_module_93_res, n_reg_module_168_res,
         n_reg_module_169_res, n_and_module_94_res, n_reg_module_170_res,
         n_reg_module_171_res, n_xor_module_185_res, n_xor_module_186_res,
         n_reg_module_172_res, n_and_module_95_res, n_reg_module_173_res,
         n_reg_module_174_res, n_and_module_96_res, n_reg_module_175_res,
         n_reg_module_176_res, n_xor_module_187_res, n_xor_module_188_res,
         n_xor_module_189_res, n_xor_module_190_res, n_xor_module_191_res,
         n_xor_module_192_res, n_xor_module_193_res, n_xor_module_194_res,
         n_xor_module_195_res, n_xor_module_196_res, n_xor_module_197_res,
         n_xor_module_198_res, n_xor_module_199_res, n_xor_module_200_res,
         n_xor_module_201_res, n_xor_module_202_res, n_xor_module_203_res,
         n_xor_module_204_res, n_xor_module_205_res, n_xor_module_206_res,
         n_xor_module_207_res, n_xor_module_208_res, n_reg_module_177_res,
         n_not_module_33_res, n_and_module_97_res, n_xor_module_209_res,
         n_not_module_34_res, n_and_module_98_res, n_xor_module_210_res,
         n_reg_module_178_res, n_and_module_99_res, n_reg_module_179_res,
         n_reg_module_180_res, n_and_module_100_res, n_reg_module_181_res,
         n_reg_module_182_res, n_xor_module_211_res, n_xor_module_212_res,
         n_reg_module_183_res, n_and_module_101_res, n_reg_module_184_res,
         n_reg_module_185_res, n_and_module_102_res, n_reg_module_186_res,
         n_reg_module_187_res, n_xor_module_213_res, n_xor_module_214_res,
         n_reg_module_188_res, n_not_module_35_res, n_and_module_103_res,
         n_xor_module_215_res, n_not_module_36_res, n_and_module_104_res,
         n_xor_module_216_res, n_reg_module_189_res, n_and_module_105_res,
         n_reg_module_190_res, n_reg_module_191_res, n_and_module_106_res,
         n_reg_module_192_res, n_reg_module_193_res, n_xor_module_217_res,
         n_xor_module_218_res, n_reg_module_194_res, n_and_module_107_res,
         n_reg_module_195_res, n_reg_module_196_res, n_and_module_108_res,
         n_reg_module_197_res, n_reg_module_198_res, n_xor_module_219_res,
         n_xor_module_220_res, n_reg_module_199_res, n_not_module_37_res,
         n_and_module_109_res, n_xor_module_221_res, n_not_module_38_res,
         n_and_module_110_res, n_xor_module_222_res, n_reg_module_200_res,
         n_and_module_111_res, n_reg_module_201_res, n_reg_module_202_res,
         n_and_module_112_res, n_reg_module_203_res, n_reg_module_204_res,
         n_xor_module_223_res, n_xor_module_224_res, n_reg_module_205_res,
         n_and_module_113_res, n_reg_module_206_res, n_reg_module_207_res,
         n_and_module_114_res, n_reg_module_208_res, n_reg_module_209_res,
         n_xor_module_225_res, n_xor_module_226_res, n_reg_module_210_res,
         n_not_module_39_res, n_and_module_115_res, n_xor_module_227_res,
         n_not_module_40_res, n_and_module_116_res, n_xor_module_228_res,
         n_reg_module_211_res, n_and_module_117_res, n_reg_module_212_res,
         n_reg_module_213_res, n_and_module_118_res, n_reg_module_214_res,
         n_reg_module_215_res, n_xor_module_229_res, n_xor_module_230_res,
         n_reg_module_216_res, n_and_module_119_res, n_reg_module_217_res,
         n_reg_module_218_res, n_and_module_120_res, n_reg_module_219_res,
         n_reg_module_220_res, n_xor_module_231_res, n_xor_module_232_res,
         n_reg_module_221_res, n_not_module_41_res, n_and_module_121_res,
         n_xor_module_233_res, n_not_module_42_res, n_and_module_122_res,
         n_xor_module_234_res, n_reg_module_222_res, n_and_module_123_res,
         n_reg_module_223_res, n_reg_module_224_res, n_and_module_124_res,
         n_reg_module_225_res, n_reg_module_226_res, n_xor_module_235_res,
         n_xor_module_236_res, n_reg_module_227_res, n_and_module_125_res,
         n_reg_module_228_res, n_reg_module_229_res, n_and_module_126_res,
         n_reg_module_230_res, n_reg_module_231_res, n_xor_module_237_res,
         n_xor_module_238_res, n_reg_module_232_res, n_not_module_43_res,
         n_and_module_127_res, n_xor_module_239_res, n_not_module_44_res,
         n_and_module_128_res, n_xor_module_240_res, n_reg_module_233_res,
         n_and_module_129_res, n_reg_module_234_res, n_reg_module_235_res,
         n_and_module_130_res, n_reg_module_236_res, n_reg_module_237_res,
         n_xor_module_241_res, n_xor_module_242_res, n_reg_module_238_res,
         n_and_module_131_res, n_reg_module_239_res, n_reg_module_240_res,
         n_and_module_132_res, n_reg_module_241_res, n_reg_module_242_res,
         n_xor_module_243_res, n_xor_module_244_res, n_reg_module_243_res,
         n_not_module_45_res, n_and_module_133_res, n_xor_module_245_res,
         n_not_module_46_res, n_and_module_134_res, n_xor_module_246_res,
         n_reg_module_244_res, n_and_module_135_res, n_reg_module_245_res,
         n_reg_module_246_res, n_and_module_136_res, n_reg_module_247_res,
         n_reg_module_248_res, n_xor_module_247_res, n_xor_module_248_res,
         n_reg_module_249_res, n_and_module_137_res, n_reg_module_250_res,
         n_reg_module_251_res, n_and_module_138_res, n_reg_module_252_res,
         n_reg_module_253_res, n_xor_module_249_res, n_xor_module_250_res,
         n_reg_module_254_res, n_not_module_47_res, n_and_module_139_res,
         n_xor_module_251_res, n_not_module_48_res, n_and_module_140_res,
         n_xor_module_252_res, n_reg_module_255_res, n_and_module_141_res,
         n_reg_module_256_res, n_reg_module_257_res, n_and_module_142_res,
         n_reg_module_258_res, n_reg_module_259_res, n_xor_module_253_res,
         n_xor_module_254_res, n_reg_module_260_res, n_and_module_143_res,
         n_reg_module_261_res, n_reg_module_262_res, n_and_module_144_res,
         n_reg_module_263_res, n_reg_module_264_res, n_xor_module_255_res,
         n_xor_module_256_res, n_reg_module_265_res, n_not_module_49_res,
         n_and_module_145_res, n_xor_module_257_res, n_not_module_50_res,
         n_and_module_146_res, n_xor_module_258_res, n_reg_module_266_res,
         n_and_module_147_res, n_reg_module_267_res, n_reg_module_268_res,
         n_and_module_148_res, n_reg_module_269_res, n_reg_module_270_res,
         n_xor_module_259_res, n_xor_module_260_res, n_reg_module_271_res,
         n_and_module_149_res, n_reg_module_272_res, n_reg_module_273_res,
         n_and_module_150_res, n_reg_module_274_res, n_reg_module_275_res,
         n_xor_module_261_res, n_xor_module_262_res, n_reg_module_276_res,
         n_not_module_51_res, n_and_module_151_res, n_xor_module_263_res,
         n_not_module_52_res, n_and_module_152_res, n_xor_module_264_res,
         n_reg_module_277_res, n_and_module_153_res, n_reg_module_278_res,
         n_reg_module_279_res, n_and_module_154_res, n_reg_module_280_res,
         n_reg_module_281_res, n_xor_module_265_res, n_xor_module_266_res,
         n_reg_module_282_res, n_and_module_155_res, n_reg_module_283_res,
         n_reg_module_284_res, n_and_module_156_res, n_reg_module_285_res,
         n_reg_module_286_res, n_xor_module_267_res, n_xor_module_268_res,
         n_reg_module_287_res, n_not_module_53_res, n_and_module_157_res,
         n_xor_module_269_res, n_not_module_54_res, n_and_module_158_res,
         n_xor_module_270_res, n_reg_module_288_res, n_and_module_159_res,
         n_reg_module_289_res, n_reg_module_290_res, n_and_module_160_res,
         n_reg_module_291_res, n_reg_module_292_res, n_xor_module_271_res,
         n_xor_module_272_res, n_reg_module_293_res, n_and_module_161_res,
         n_reg_module_294_res, n_reg_module_295_res, n_and_module_162_res,
         n_reg_module_296_res, n_reg_module_297_res, n_xor_module_273_res,
         n_xor_module_274_res, n_reg_module_298_res, n_not_module_55_res,
         n_and_module_163_res, n_xor_module_275_res, n_not_module_56_res,
         n_and_module_164_res, n_xor_module_276_res, n_reg_module_299_res,
         n_and_module_165_res, n_reg_module_300_res, n_reg_module_301_res,
         n_and_module_166_res, n_reg_module_302_res, n_reg_module_303_res,
         n_xor_module_277_res, n_xor_module_278_res, n_reg_module_304_res,
         n_and_module_167_res, n_reg_module_305_res, n_reg_module_306_res,
         n_and_module_168_res, n_reg_module_307_res, n_reg_module_308_res,
         n_xor_module_279_res, n_xor_module_280_res, n_reg_module_309_res,
         n_not_module_57_res, n_and_module_169_res, n_xor_module_281_res,
         n_not_module_58_res, n_and_module_170_res, n_xor_module_282_res,
         n_reg_module_310_res, n_and_module_171_res, n_reg_module_311_res,
         n_reg_module_312_res, n_and_module_172_res, n_reg_module_313_res,
         n_reg_module_314_res, n_xor_module_283_res, n_xor_module_284_res,
         n_reg_module_315_res, n_and_module_173_res, n_reg_module_316_res,
         n_reg_module_317_res, n_and_module_174_res, n_reg_module_318_res,
         n_reg_module_319_res, n_xor_module_285_res, n_xor_module_286_res,
         n_reg_module_320_res, n_not_module_59_res, n_and_module_175_res,
         n_xor_module_287_res, n_not_module_60_res, n_and_module_176_res,
         n_xor_module_288_res, n_reg_module_321_res, n_and_module_177_res,
         n_reg_module_322_res, n_reg_module_323_res, n_and_module_178_res,
         n_reg_module_324_res, n_reg_module_325_res, n_xor_module_289_res,
         n_xor_module_290_res, n_reg_module_326_res, n_and_module_179_res,
         n_reg_module_327_res, n_reg_module_328_res, n_and_module_180_res,
         n_reg_module_329_res, n_reg_module_330_res, n_xor_module_291_res,
         n_xor_module_292_res, n_reg_module_331_res, n_not_module_61_res,
         n_and_module_181_res, n_xor_module_293_res, n_not_module_62_res,
         n_and_module_182_res, n_xor_module_294_res, n_reg_module_332_res,
         n_and_module_183_res, n_reg_module_333_res, n_reg_module_334_res,
         n_and_module_184_res, n_reg_module_335_res, n_reg_module_336_res,
         n_xor_module_295_res, n_xor_module_296_res, n_reg_module_337_res,
         n_and_module_185_res, n_reg_module_338_res, n_reg_module_339_res,
         n_and_module_186_res, n_reg_module_340_res, n_reg_module_341_res,
         n_xor_module_297_res, n_xor_module_298_res, n_reg_module_342_res,
         n_not_module_63_res, n_and_module_187_res, n_xor_module_299_res,
         n_not_module_64_res, n_and_module_188_res, n_xor_module_300_res,
         n_reg_module_343_res, n_and_module_189_res, n_reg_module_344_res,
         n_reg_module_345_res, n_and_module_190_res, n_reg_module_346_res,
         n_reg_module_347_res, n_xor_module_301_res, n_xor_module_302_res,
         n_reg_module_348_res, n_and_module_191_res, n_reg_module_349_res,
         n_reg_module_350_res, n_and_module_192_res, n_reg_module_351_res,
         n_reg_module_352_res, n_xor_module_303_res, n_xor_module_304_res,
         n_reg_module_353_res, n_not_module_65_res, n_and_module_193_res,
         n_xor_module_305_res, n_not_module_66_res, n_and_module_194_res,
         n_xor_module_306_res, n_reg_module_354_res, n_and_module_195_res,
         n_reg_module_355_res, n_reg_module_356_res, n_and_module_196_res,
         n_reg_module_357_res, n_reg_module_358_res, n_xor_module_307_res,
         n_xor_module_308_res, n_reg_module_359_res, n_and_module_197_res,
         n_reg_module_360_res, n_reg_module_361_res, n_and_module_198_res,
         n_reg_module_362_res, n_reg_module_363_res, n_xor_module_309_res,
         n_xor_module_310_res, n_reg_module_364_res, n_not_module_67_res,
         n_and_module_199_res, n_xor_module_311_res, n_not_module_68_res,
         n_and_module_200_res, n_xor_module_312_res, n_reg_module_365_res,
         n_and_module_201_res, n_reg_module_366_res, n_reg_module_367_res,
         n_and_module_202_res, n_reg_module_368_res, n_reg_module_369_res,
         n_xor_module_313_res, n_xor_module_314_res, n_reg_module_370_res,
         n_and_module_203_res, n_reg_module_371_res, n_reg_module_372_res,
         n_and_module_204_res, n_reg_module_373_res, n_reg_module_374_res,
         n_xor_module_315_res, n_xor_module_316_res, n_xor_module_317_res,
         n_xor_module_318_res, n_xor_module_319_res, n_xor_module_320_res,
         n_xor_module_321_res, n_xor_module_322_res, n_xor_module_323_res,
         n_xor_module_324_res, n_xor_module_325_res, n_xor_module_326_res,
         n_xor_module_327_res, n_xor_module_328_res, n_xor_module_329_res,
         n_xor_module_330_res, n_xor_module_331_res, n_xor_module_332_res,
         n_xor_module_333_res, n_xor_module_334_res, n_xor_module_335_res,
         n_xor_module_336_res, n_xor_module_337_res, n_xor_module_338_res,
         n_xor_module_339_res, n_xor_module_340_res, n_xor_module_341_res,
         n_xor_module_342_res, n_xor_module_343_res, n_xor_module_344_res,
         n_xor_module_345_res, n_xor_module_346_res, n_xor_module_347_res,
         n_xor_module_348_res, n_xor_module_349_res, n_xor_module_350_res,
         n_xor_module_351_res, n_xor_module_352_res, n_xor_module_353_res,
         n_xor_module_354_res, n_xor_module_355_res, n_xor_module_356_res,
         n_xor_module_357_res, n_xor_module_358_res, n_xor_module_359_res,
         n_xor_module_360_res, n_xor_module_361_res, n_xor_module_362_res,
         n_xor_module_363_res, n_xor_module_364_res, n_xor_module_365_res,
         n_xor_module_366_res, n_xor_module_367_res, n_xor_module_368_res,
         n_xor_module_369_res, n_xor_module_370_res, n_xor_module_371_res,
         n_xor_module_372_res, n_xor_module_373_res, n_xor_module_374_res,
         n_xor_module_375_res, n_xor_module_376_res, n_xor_module_377_res,
         n_xor_module_378_res, n_xor_module_379_res, n_xor_module_380_res,
         n_not_module_69_res, n_xor_module_381_res, n_xor_module_382_res,
         n_not_module_70_res, n_xor_module_383_res, n_xor_module_384_res,
         n_xor_module_385_res, n_xor_module_386_res, n_xor_module_387_res,
         n_xor_module_388_res, n_xor_module_389_res, n_xor_module_390_res,
         n_not_module_71_res, n_xor_module_391_res, n_xor_module_392_res,
         n_not_module_72_res;

  XOR2_X1 u_xor_module_1_U1 ( .A(io_i3_s0), .B(io_i0_s0), .Z(
        n_xor_module_1_res) );
  XOR2_X1 u_xor_module_2_U1 ( .A(io_i3_s1), .B(io_i0_s1), .Z(
        n_xor_module_2_res) );
  XOR2_X1 u_xor_module_3_U1 ( .A(io_i5_s0), .B(io_i0_s0), .Z(
        n_xor_module_3_res) );
  XOR2_X1 u_xor_module_4_U1 ( .A(io_i5_s1), .B(io_i0_s1), .Z(
        n_xor_module_4_res) );
  XOR2_X1 u_xor_module_5_U1 ( .A(io_i6_s0), .B(io_i0_s0), .Z(
        n_xor_module_5_res) );
  XOR2_X1 u_xor_module_6_U1 ( .A(io_i6_s1), .B(io_i0_s1), .Z(
        n_xor_module_6_res) );
  XOR2_X1 u_xor_module_7_U1 ( .A(io_i5_s0), .B(io_i3_s0), .Z(
        n_xor_module_7_res) );
  XOR2_X1 u_xor_module_8_U1 ( .A(io_i5_s1), .B(io_i3_s1), .Z(
        n_xor_module_8_res) );
  XOR2_X1 u_xor_module_9_U1 ( .A(io_i6_s0), .B(io_i4_s0), .Z(
        n_xor_module_9_res) );
  XOR2_X1 u_xor_module_10_U1 ( .A(io_i6_s1), .B(io_i4_s1), .Z(
        n_xor_module_10_res) );
  XOR2_X1 u_xor_module_11_U1 ( .A(n_xor_module_9_res), .B(n_xor_module_1_res), 
        .Z(n_xor_module_11_res) );
  XOR2_X1 u_xor_module_12_U1 ( .A(n_xor_module_10_res), .B(n_xor_module_2_res), 
        .Z(n_xor_module_12_res) );
  XOR2_X1 u_xor_module_13_U1 ( .A(io_i2_s0), .B(io_i1_s0), .Z(
        n_xor_module_13_res) );
  XOR2_X1 u_xor_module_14_U1 ( .A(io_i2_s1), .B(io_i1_s1), .Z(
        n_xor_module_14_res) );
  XOR2_X1 u_xor_module_15_U1 ( .A(n_xor_module_11_res), .B(io_i7_s0), .Z(
        n_xor_module_15_res) );
  XOR2_X1 u_xor_module_16_U1 ( .A(n_xor_module_12_res), .B(io_i7_s1), .Z(
        n_xor_module_16_res) );
  XOR2_X1 u_xor_module_17_U1 ( .A(n_xor_module_13_res), .B(io_i7_s0), .Z(
        n_xor_module_17_res) );
  XOR2_X1 u_xor_module_18_U1 ( .A(n_xor_module_14_res), .B(io_i7_s1), .Z(
        n_xor_module_18_res) );
  XOR2_X1 u_xor_module_19_U1 ( .A(n_xor_module_13_res), .B(n_xor_module_11_res), .Z(n_xor_module_19_res) );
  XOR2_X1 u_xor_module_20_U1 ( .A(n_xor_module_14_res), .B(n_xor_module_12_res), .Z(n_xor_module_20_res) );
  XOR2_X1 u_xor_module_21_U1 ( .A(io_i5_s0), .B(io_i1_s0), .Z(
        n_xor_module_21_res) );
  XOR2_X1 u_xor_module_22_U1 ( .A(io_i5_s1), .B(io_i1_s1), .Z(
        n_xor_module_22_res) );
  XOR2_X1 u_xor_module_23_U1 ( .A(io_i5_s0), .B(io_i2_s0), .Z(
        n_xor_module_23_res) );
  XOR2_X1 u_xor_module_24_U1 ( .A(io_i5_s1), .B(io_i2_s1), .Z(
        n_xor_module_24_res) );
  XOR2_X1 u_xor_module_25_U1 ( .A(n_xor_module_7_res), .B(n_xor_module_5_res), 
        .Z(n_xor_module_25_res) );
  XOR2_X1 u_xor_module_26_U1 ( .A(n_xor_module_8_res), .B(n_xor_module_6_res), 
        .Z(n_xor_module_26_res) );
  XOR2_X1 u_xor_module_27_U1 ( .A(n_xor_module_21_res), .B(n_xor_module_11_res), .Z(n_xor_module_27_res) );
  XOR2_X1 u_xor_module_28_U1 ( .A(n_xor_module_22_res), .B(n_xor_module_12_res), .Z(n_xor_module_28_res) );
  XOR2_X1 u_xor_module_29_U1 ( .A(n_xor_module_21_res), .B(n_xor_module_9_res), 
        .Z(n_xor_module_29_res) );
  XOR2_X1 u_xor_module_30_U1 ( .A(n_xor_module_22_res), .B(n_xor_module_10_res), .Z(n_xor_module_30_res) );
  XOR2_X1 u_xor_module_31_U1 ( .A(n_xor_module_23_res), .B(n_xor_module_9_res), 
        .Z(n_xor_module_31_res) );
  XOR2_X1 u_xor_module_32_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_10_res), .Z(n_xor_module_32_res) );
  XOR2_X1 u_xor_module_33_U1 ( .A(n_xor_module_31_res), .B(n_xor_module_17_res), .Z(n_xor_module_33_res) );
  XOR2_X1 u_xor_module_34_U1 ( .A(n_xor_module_32_res), .B(n_xor_module_18_res), .Z(n_xor_module_34_res) );
  XOR2_X1 u_xor_module_35_U1 ( .A(io_i7_s0), .B(io_i3_s0), .Z(
        n_xor_module_35_res) );
  XOR2_X1 u_xor_module_36_U1 ( .A(io_i7_s1), .B(io_i3_s1), .Z(
        n_xor_module_36_res) );
  XOR2_X1 u_xor_module_37_U1 ( .A(n_xor_module_35_res), .B(n_xor_module_13_res), .Z(n_xor_module_37_res) );
  XOR2_X1 u_xor_module_38_U1 ( .A(n_xor_module_36_res), .B(n_xor_module_14_res), .Z(n_xor_module_38_res) );
  XOR2_X1 u_xor_module_39_U1 ( .A(n_xor_module_37_res), .B(n_xor_module_1_res), 
        .Z(n_xor_module_39_res) );
  XOR2_X1 u_xor_module_40_U1 ( .A(n_xor_module_38_res), .B(n_xor_module_2_res), 
        .Z(n_xor_module_40_res) );
  XOR2_X1 u_xor_module_41_U1 ( .A(io_i7_s0), .B(io_i6_s0), .Z(
        n_xor_module_41_res) );
  XOR2_X1 u_xor_module_42_U1 ( .A(io_i7_s1), .B(io_i6_s1), .Z(
        n_xor_module_42_res) );
  XOR2_X1 u_xor_module_43_U1 ( .A(n_xor_module_41_res), .B(n_xor_module_13_res), .Z(n_xor_module_43_res) );
  XOR2_X1 u_xor_module_44_U1 ( .A(n_xor_module_42_res), .B(n_xor_module_14_res), .Z(n_xor_module_44_res) );
  XOR2_X1 u_xor_module_45_U1 ( .A(n_xor_module_43_res), .B(n_xor_module_3_res), 
        .Z(n_xor_module_45_res) );
  XOR2_X1 u_xor_module_46_U1 ( .A(n_xor_module_44_res), .B(n_xor_module_4_res), 
        .Z(n_xor_module_46_res) );
  XOR2_X1 u_xor_module_47_U1 ( .A(n_xor_module_19_res), .B(n_xor_module_3_res), 
        .Z(n_xor_module_47_res) );
  XOR2_X1 u_xor_module_48_U1 ( .A(n_xor_module_20_res), .B(n_xor_module_4_res), 
        .Z(n_xor_module_48_res) );
  XOR2_X1 u_xor_module_49_U1 ( .A(n_xor_module_33_res), .B(n_xor_module_39_res), .Z(n_xor_module_49_res) );
  XOR2_X1 u_xor_module_50_U1 ( .A(n_xor_module_34_res), .B(n_xor_module_40_res), .Z(n_xor_module_50_res) );
  XOR2_X1 u_xor_module_51_U1 ( .A(n_xor_module_31_res), .B(n_xor_module_5_res), 
        .Z(n_xor_module_51_res) );
  XOR2_X1 u_xor_module_52_U1 ( .A(n_xor_module_32_res), .B(n_xor_module_6_res), 
        .Z(n_xor_module_52_res) );
  XOR2_X1 u_xor_module_53_U1 ( .A(n_xor_module_23_res), .B(n_xor_module_1_res), 
        .Z(n_xor_module_53_res) );
  XOR2_X1 u_xor_module_54_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_2_res), 
        .Z(n_xor_module_54_res) );
  DFF_X1 u_reg_module_1__hpc_r0_reg ( .D(p_rand_0), .CK(clock_0), .Q(
        n_reg_module_1_res), .QN() );
  INV_X1 u_not_module_1_U1 ( .A(n_xor_module_25_res), .ZN(n_not_module_1_res)
         );
  AND2_X1 u_and_module_1_U1 ( .A1(n_not_module_1_res), .A2(n_reg_module_1_res), 
        .ZN(n_and_module_1_res) );
  XOR2_X1 u_xor_module_55_U1 ( .A(p_rand_0), .B(n_xor_module_12_res), .Z(
        n_xor_module_55_res) );
  INV_X1 u_not_module_2_U1 ( .A(n_xor_module_26_res), .ZN(n_not_module_2_res)
         );
  AND2_X1 u_and_module_2_U1 ( .A1(n_not_module_2_res), .A2(n_reg_module_1_res), 
        .ZN(n_and_module_2_res) );
  XOR2_X1 u_xor_module_56_U1 ( .A(p_rand_0), .B(n_xor_module_11_res), .Z(
        n_xor_module_56_res) );
  DFF_X1 u_reg_module_2__hpc_r0_reg ( .D(n_xor_module_11_res), .CK(clock_0), 
        .Q(n_reg_module_2_res), .QN() );
  AND2_X1 u_and_module_3_U1 ( .A1(n_reg_module_2_res), .A2(n_xor_module_25_res), .ZN(n_and_module_3_res) );
  DFF_X1 u_reg_module_3__hpc_r0_reg ( .D(n_and_module_3_res), .CK(clock_0), 
        .Q(n_reg_module_3_res), .QN() );
  DFF_X1 u_reg_module_4__hpc_r0_reg ( .D(n_xor_module_55_res), .CK(clock_0), 
        .Q(n_reg_module_4_res), .QN() );
  AND2_X1 u_and_module_4_U1 ( .A1(n_reg_module_4_res), .A2(n_xor_module_25_res), .ZN(n_and_module_4_res) );
  DFF_X1 u_reg_module_5__hpc_r0_reg ( .D(n_and_module_4_res), .CK(clock_0), 
        .Q(n_reg_module_5_res), .QN() );
  DFF_X1 u_reg_module_6__hpc_r0_reg ( .D(n_and_module_1_res), .CK(clock_0), 
        .Q(n_reg_module_6_res), .QN() );
  XOR2_X1 u_xor_module_57_U1 ( .A(n_reg_module_6_res), .B(n_reg_module_5_res), 
        .Z(n_xor_module_57_res) );
  XOR2_X1 u_xor_module_58_U1 ( .A(n_xor_module_57_res), .B(n_reg_module_3_res), 
        .Z(n_xor_module_58_res) );
  DFF_X1 u_reg_module_7__hpc_r0_reg ( .D(n_xor_module_12_res), .CK(clock_0), 
        .Q(n_reg_module_7_res), .QN() );
  AND2_X1 u_and_module_5_U1 ( .A1(n_reg_module_7_res), .A2(n_xor_module_26_res), .ZN(n_and_module_5_res) );
  DFF_X1 u_reg_module_8__hpc_r0_reg ( .D(n_and_module_5_res), .CK(clock_0), 
        .Q(n_reg_module_8_res), .QN() );
  DFF_X1 u_reg_module_9__hpc_r0_reg ( .D(n_xor_module_56_res), .CK(clock_0), 
        .Q(n_reg_module_9_res), .QN() );
  AND2_X1 u_and_module_6_U1 ( .A1(n_reg_module_9_res), .A2(n_xor_module_26_res), .ZN(n_and_module_6_res) );
  DFF_X1 u_reg_module_10__hpc_r0_reg ( .D(n_and_module_6_res), .CK(clock_0), 
        .Q(n_reg_module_10_res), .QN() );
  DFF_X1 u_reg_module_11__hpc_r0_reg ( .D(n_and_module_2_res), .CK(clock_0), 
        .Q(n_reg_module_11_res), .QN() );
  XOR2_X1 u_xor_module_59_U1 ( .A(n_reg_module_11_res), .B(n_reg_module_10_res), .Z(n_xor_module_59_res) );
  XOR2_X1 u_xor_module_60_U1 ( .A(n_xor_module_59_res), .B(n_reg_module_8_res), 
        .Z(n_xor_module_60_res) );
  DFF_X1 u_reg_module_12__hpc_r0_reg ( .D(p_rand_1), .CK(clock_0), .Q(
        n_reg_module_12_res), .QN() );
  INV_X1 u_not_module_3_U1 ( .A(n_xor_module_45_res), .ZN(n_not_module_3_res)
         );
  AND2_X1 u_and_module_7_U1 ( .A1(n_not_module_3_res), .A2(n_reg_module_12_res), .ZN(n_and_module_7_res) );
  XOR2_X1 u_xor_module_61_U1 ( .A(p_rand_1), .B(n_xor_module_16_res), .Z(
        n_xor_module_61_res) );
  INV_X1 u_not_module_4_U1 ( .A(n_xor_module_46_res), .ZN(n_not_module_4_res)
         );
  AND2_X1 u_and_module_8_U1 ( .A1(n_not_module_4_res), .A2(n_reg_module_12_res), .ZN(n_and_module_8_res) );
  XOR2_X1 u_xor_module_62_U1 ( .A(p_rand_1), .B(n_xor_module_15_res), .Z(
        n_xor_module_62_res) );
  DFF_X1 u_reg_module_13__hpc_r0_reg ( .D(n_xor_module_15_res), .CK(clock_0), 
        .Q(n_reg_module_13_res), .QN() );
  AND2_X1 u_and_module_9_U1 ( .A1(n_reg_module_13_res), .A2(
        n_xor_module_45_res), .ZN(n_and_module_9_res) );
  DFF_X1 u_reg_module_14__hpc_r0_reg ( .D(n_and_module_9_res), .CK(clock_0), 
        .Q(n_reg_module_14_res), .QN() );
  DFF_X1 u_reg_module_15__hpc_r0_reg ( .D(n_xor_module_61_res), .CK(clock_0), 
        .Q(n_reg_module_15_res), .QN() );
  AND2_X1 u_and_module_10_U1 ( .A1(n_reg_module_15_res), .A2(
        n_xor_module_45_res), .ZN(n_and_module_10_res) );
  DFF_X1 u_reg_module_16__hpc_r0_reg ( .D(n_and_module_10_res), .CK(clock_0), 
        .Q(n_reg_module_16_res), .QN() );
  DFF_X1 u_reg_module_17__hpc_r0_reg ( .D(n_and_module_7_res), .CK(clock_0), 
        .Q(n_reg_module_17_res), .QN() );
  XOR2_X1 u_xor_module_63_U1 ( .A(n_reg_module_17_res), .B(n_reg_module_16_res), .Z(n_xor_module_63_res) );
  XOR2_X1 u_xor_module_64_U1 ( .A(n_xor_module_63_res), .B(n_reg_module_14_res), .Z(n_xor_module_64_res) );
  DFF_X1 u_reg_module_18__hpc_r0_reg ( .D(n_xor_module_16_res), .CK(clock_0), 
        .Q(n_reg_module_18_res), .QN() );
  AND2_X1 u_and_module_11_U1 ( .A1(n_reg_module_18_res), .A2(
        n_xor_module_46_res), .ZN(n_and_module_11_res) );
  DFF_X1 u_reg_module_19__hpc_r0_reg ( .D(n_and_module_11_res), .CK(clock_0), 
        .Q(n_reg_module_19_res), .QN() );
  DFF_X1 u_reg_module_20__hpc_r0_reg ( .D(n_xor_module_62_res), .CK(clock_0), 
        .Q(n_reg_module_20_res), .QN() );
  AND2_X1 u_and_module_12_U1 ( .A1(n_reg_module_20_res), .A2(
        n_xor_module_46_res), .ZN(n_and_module_12_res) );
  DFF_X1 u_reg_module_21__hpc_r0_reg ( .D(n_and_module_12_res), .CK(clock_0), 
        .Q(n_reg_module_21_res), .QN() );
  DFF_X1 u_reg_module_22__hpc_r0_reg ( .D(n_and_module_8_res), .CK(clock_0), 
        .Q(n_reg_module_22_res), .QN() );
  XOR2_X1 u_xor_module_65_U1 ( .A(n_reg_module_22_res), .B(n_reg_module_21_res), .Z(n_xor_module_65_res) );
  XOR2_X1 u_xor_module_66_U1 ( .A(n_xor_module_65_res), .B(n_reg_module_19_res), .Z(n_xor_module_66_res) );
  XOR2_X1 u_xor_module_67_U1 ( .A(n_xor_module_58_res), .B(n_xor_module_27_res), .Z(n_xor_module_67_res) );
  XOR2_X1 u_xor_module_68_U1 ( .A(n_xor_module_60_res), .B(n_xor_module_28_res), .Z(n_xor_module_68_res) );
  DFF_X1 u_reg_module_23__hpc_r0_reg ( .D(p_rand_2), .CK(clock_0), .Q(
        n_reg_module_23_res), .QN() );
  INV_X1 u_not_module_5_U1 ( .A(n_xor_module_37_res), .ZN(n_not_module_5_res)
         );
  AND2_X1 u_and_module_13_U1 ( .A1(n_not_module_5_res), .A2(
        n_reg_module_23_res), .ZN(n_and_module_13_res) );
  XOR2_X1 u_xor_module_69_U1 ( .A(p_rand_2), .B(io_i7_s1), .Z(
        n_xor_module_69_res) );
  INV_X1 u_not_module_6_U1 ( .A(n_xor_module_38_res), .ZN(n_not_module_6_res)
         );
  AND2_X1 u_and_module_14_U1 ( .A1(n_not_module_6_res), .A2(
        n_reg_module_23_res), .ZN(n_and_module_14_res) );
  XOR2_X1 u_xor_module_70_U1 ( .A(p_rand_2), .B(io_i7_s0), .Z(
        n_xor_module_70_res) );
  DFF_X1 u_reg_module_24__hpc_r0_reg ( .D(io_i7_s0), .CK(clock_0), .Q(
        n_reg_module_24_res), .QN() );
  AND2_X1 u_and_module_15_U1 ( .A1(n_reg_module_24_res), .A2(
        n_xor_module_37_res), .ZN(n_and_module_15_res) );
  DFF_X1 u_reg_module_25__hpc_r0_reg ( .D(n_and_module_15_res), .CK(clock_0), 
        .Q(n_reg_module_25_res), .QN() );
  DFF_X1 u_reg_module_26__hpc_r0_reg ( .D(n_xor_module_69_res), .CK(clock_0), 
        .Q(n_reg_module_26_res), .QN() );
  AND2_X1 u_and_module_16_U1 ( .A1(n_reg_module_26_res), .A2(
        n_xor_module_37_res), .ZN(n_and_module_16_res) );
  DFF_X1 u_reg_module_27__hpc_r0_reg ( .D(n_and_module_16_res), .CK(clock_0), 
        .Q(n_reg_module_27_res), .QN() );
  DFF_X1 u_reg_module_28__hpc_r0_reg ( .D(n_and_module_13_res), .CK(clock_0), 
        .Q(n_reg_module_28_res), .QN() );
  XOR2_X1 u_xor_module_71_U1 ( .A(n_reg_module_28_res), .B(n_reg_module_27_res), .Z(n_xor_module_71_res) );
  XOR2_X1 u_xor_module_72_U1 ( .A(n_xor_module_71_res), .B(n_reg_module_25_res), .Z(n_xor_module_72_res) );
  DFF_X1 u_reg_module_29__hpc_r0_reg ( .D(io_i7_s1), .CK(clock_0), .Q(
        n_reg_module_29_res), .QN() );
  AND2_X1 u_and_module_17_U1 ( .A1(n_reg_module_29_res), .A2(
        n_xor_module_38_res), .ZN(n_and_module_17_res) );
  DFF_X1 u_reg_module_30__hpc_r0_reg ( .D(n_and_module_17_res), .CK(clock_0), 
        .Q(n_reg_module_30_res), .QN() );
  DFF_X1 u_reg_module_31__hpc_r0_reg ( .D(n_xor_module_70_res), .CK(clock_0), 
        .Q(n_reg_module_31_res), .QN() );
  AND2_X1 u_and_module_18_U1 ( .A1(n_reg_module_31_res), .A2(
        n_xor_module_38_res), .ZN(n_and_module_18_res) );
  DFF_X1 u_reg_module_32__hpc_r0_reg ( .D(n_and_module_18_res), .CK(clock_0), 
        .Q(n_reg_module_32_res), .QN() );
  DFF_X1 u_reg_module_33__hpc_r0_reg ( .D(n_and_module_14_res), .CK(clock_0), 
        .Q(n_reg_module_33_res), .QN() );
  XOR2_X1 u_xor_module_73_U1 ( .A(n_reg_module_33_res), .B(n_reg_module_32_res), .Z(n_xor_module_73_res) );
  XOR2_X1 u_xor_module_74_U1 ( .A(n_xor_module_73_res), .B(n_reg_module_30_res), .Z(n_xor_module_74_res) );
  XOR2_X1 u_xor_module_75_U1 ( .A(n_xor_module_58_res), .B(n_xor_module_72_res), .Z(n_xor_module_75_res) );
  XOR2_X1 u_xor_module_76_U1 ( .A(n_xor_module_60_res), .B(n_xor_module_74_res), .Z(n_xor_module_76_res) );
  DFF_X1 u_reg_module_34__hpc_r0_reg ( .D(p_rand_3), .CK(clock_0), .Q(
        n_reg_module_34_res), .QN() );
  INV_X1 u_not_module_7_U1 ( .A(n_xor_module_5_res), .ZN(n_not_module_7_res)
         );
  AND2_X1 u_and_module_19_U1 ( .A1(n_not_module_7_res), .A2(
        n_reg_module_34_res), .ZN(n_and_module_19_res) );
  XOR2_X1 u_xor_module_77_U1 ( .A(p_rand_3), .B(n_xor_module_32_res), .Z(
        n_xor_module_77_res) );
  INV_X1 u_not_module_8_U1 ( .A(n_xor_module_6_res), .ZN(n_not_module_8_res)
         );
  AND2_X1 u_and_module_20_U1 ( .A1(n_not_module_8_res), .A2(
        n_reg_module_34_res), .ZN(n_and_module_20_res) );
  XOR2_X1 u_xor_module_78_U1 ( .A(p_rand_3), .B(n_xor_module_31_res), .Z(
        n_xor_module_78_res) );
  DFF_X1 u_reg_module_35__hpc_r0_reg ( .D(n_xor_module_31_res), .CK(clock_0), 
        .Q(n_reg_module_35_res), .QN() );
  AND2_X1 u_and_module_21_U1 ( .A1(n_reg_module_35_res), .A2(
        n_xor_module_5_res), .ZN(n_and_module_21_res) );
  DFF_X1 u_reg_module_36__hpc_r0_reg ( .D(n_and_module_21_res), .CK(clock_0), 
        .Q(n_reg_module_36_res), .QN() );
  DFF_X1 u_reg_module_37__hpc_r0_reg ( .D(n_xor_module_77_res), .CK(clock_0), 
        .Q(n_reg_module_37_res), .QN() );
  AND2_X1 u_and_module_22_U1 ( .A1(n_reg_module_37_res), .A2(
        n_xor_module_5_res), .ZN(n_and_module_22_res) );
  DFF_X1 u_reg_module_38__hpc_r0_reg ( .D(n_and_module_22_res), .CK(clock_0), 
        .Q(n_reg_module_38_res), .QN() );
  DFF_X1 u_reg_module_39__hpc_r0_reg ( .D(n_and_module_19_res), .CK(clock_0), 
        .Q(n_reg_module_39_res), .QN() );
  XOR2_X1 u_xor_module_79_U1 ( .A(n_reg_module_39_res), .B(n_reg_module_38_res), .Z(n_xor_module_79_res) );
  XOR2_X1 u_xor_module_80_U1 ( .A(n_xor_module_79_res), .B(n_reg_module_36_res), .Z(n_xor_module_80_res) );
  DFF_X1 u_reg_module_40__hpc_r0_reg ( .D(n_xor_module_32_res), .CK(clock_0), 
        .Q(n_reg_module_40_res), .QN() );
  AND2_X1 u_and_module_23_U1 ( .A1(n_reg_module_40_res), .A2(
        n_xor_module_6_res), .ZN(n_and_module_23_res) );
  DFF_X1 u_reg_module_41__hpc_r0_reg ( .D(n_and_module_23_res), .CK(clock_0), 
        .Q(n_reg_module_41_res), .QN() );
  DFF_X1 u_reg_module_42__hpc_r0_reg ( .D(n_xor_module_78_res), .CK(clock_0), 
        .Q(n_reg_module_42_res), .QN() );
  AND2_X1 u_and_module_24_U1 ( .A1(n_reg_module_42_res), .A2(
        n_xor_module_6_res), .ZN(n_and_module_24_res) );
  DFF_X1 u_reg_module_43__hpc_r0_reg ( .D(n_and_module_24_res), .CK(clock_0), 
        .Q(n_reg_module_43_res), .QN() );
  DFF_X1 u_reg_module_44__hpc_r0_reg ( .D(n_and_module_20_res), .CK(clock_0), 
        .Q(n_reg_module_44_res), .QN() );
  XOR2_X1 u_xor_module_81_U1 ( .A(n_reg_module_44_res), .B(n_reg_module_43_res), .Z(n_xor_module_81_res) );
  XOR2_X1 u_xor_module_82_U1 ( .A(n_xor_module_81_res), .B(n_reg_module_41_res), .Z(n_xor_module_82_res) );
  DFF_X1 u_reg_module_45__hpc_r0_reg ( .D(p_rand_4), .CK(clock_0), .Q(
        n_reg_module_45_res), .QN() );
  INV_X1 u_not_module_9_U1 ( .A(n_xor_module_43_res), .ZN(n_not_module_9_res)
         );
  AND2_X1 u_and_module_25_U1 ( .A1(n_not_module_9_res), .A2(
        n_reg_module_45_res), .ZN(n_and_module_25_res) );
  XOR2_X1 u_xor_module_83_U1 ( .A(p_rand_4), .B(n_xor_module_18_res), .Z(
        n_xor_module_83_res) );
  INV_X1 u_not_module_10_U1 ( .A(n_xor_module_44_res), .ZN(n_not_module_10_res) );
  AND2_X1 u_and_module_26_U1 ( .A1(n_not_module_10_res), .A2(
        n_reg_module_45_res), .ZN(n_and_module_26_res) );
  XOR2_X1 u_xor_module_84_U1 ( .A(p_rand_4), .B(n_xor_module_17_res), .Z(
        n_xor_module_84_res) );
  DFF_X1 u_reg_module_46__hpc_r0_reg ( .D(n_xor_module_17_res), .CK(clock_0), 
        .Q(n_reg_module_46_res), .QN() );
  AND2_X1 u_and_module_27_U1 ( .A1(n_reg_module_46_res), .A2(
        n_xor_module_43_res), .ZN(n_and_module_27_res) );
  DFF_X1 u_reg_module_47__hpc_r0_reg ( .D(n_and_module_27_res), .CK(clock_0), 
        .Q(n_reg_module_47_res), .QN() );
  DFF_X1 u_reg_module_48__hpc_r0_reg ( .D(n_xor_module_83_res), .CK(clock_0), 
        .Q(n_reg_module_48_res), .QN() );
  AND2_X1 u_and_module_28_U1 ( .A1(n_reg_module_48_res), .A2(
        n_xor_module_43_res), .ZN(n_and_module_28_res) );
  DFF_X1 u_reg_module_49__hpc_r0_reg ( .D(n_and_module_28_res), .CK(clock_0), 
        .Q(n_reg_module_49_res), .QN() );
  DFF_X1 u_reg_module_50__hpc_r0_reg ( .D(n_and_module_25_res), .CK(clock_0), 
        .Q(n_reg_module_50_res), .QN() );
  XOR2_X1 u_xor_module_85_U1 ( .A(n_reg_module_50_res), .B(n_reg_module_49_res), .Z(n_xor_module_85_res) );
  XOR2_X1 u_xor_module_86_U1 ( .A(n_xor_module_85_res), .B(n_reg_module_47_res), .Z(n_xor_module_86_res) );
  DFF_X1 u_reg_module_51__hpc_r0_reg ( .D(n_xor_module_18_res), .CK(clock_0), 
        .Q(n_reg_module_51_res), .QN() );
  AND2_X1 u_and_module_29_U1 ( .A1(n_reg_module_51_res), .A2(
        n_xor_module_44_res), .ZN(n_and_module_29_res) );
  DFF_X1 u_reg_module_52__hpc_r0_reg ( .D(n_and_module_29_res), .CK(clock_0), 
        .Q(n_reg_module_52_res), .QN() );
  DFF_X1 u_reg_module_53__hpc_r0_reg ( .D(n_xor_module_84_res), .CK(clock_0), 
        .Q(n_reg_module_53_res), .QN() );
  AND2_X1 u_and_module_30_U1 ( .A1(n_reg_module_53_res), .A2(
        n_xor_module_44_res), .ZN(n_and_module_30_res) );
  DFF_X1 u_reg_module_54__hpc_r0_reg ( .D(n_and_module_30_res), .CK(clock_0), 
        .Q(n_reg_module_54_res), .QN() );
  DFF_X1 u_reg_module_55__hpc_r0_reg ( .D(n_and_module_26_res), .CK(clock_0), 
        .Q(n_reg_module_55_res), .QN() );
  XOR2_X1 u_xor_module_87_U1 ( .A(n_reg_module_55_res), .B(n_reg_module_54_res), .Z(n_xor_module_87_res) );
  XOR2_X1 u_xor_module_88_U1 ( .A(n_xor_module_87_res), .B(n_reg_module_52_res), .Z(n_xor_module_88_res) );
  XOR2_X1 u_xor_module_89_U1 ( .A(n_xor_module_80_res), .B(n_xor_module_51_res), .Z(n_xor_module_89_res) );
  XOR2_X1 u_xor_module_90_U1 ( .A(n_xor_module_82_res), .B(n_xor_module_52_res), .Z(n_xor_module_90_res) );
  DFF_X1 u_reg_module_56__hpc_r0_reg ( .D(p_rand_5), .CK(clock_0), .Q(
        n_reg_module_56_res), .QN() );
  INV_X1 u_not_module_11_U1 ( .A(n_xor_module_39_res), .ZN(n_not_module_11_res) );
  AND2_X1 u_and_module_31_U1 ( .A1(n_not_module_11_res), .A2(
        n_reg_module_56_res), .ZN(n_and_module_31_res) );
  XOR2_X1 u_xor_module_91_U1 ( .A(p_rand_5), .B(n_xor_module_34_res), .Z(
        n_xor_module_91_res) );
  INV_X1 u_not_module_12_U1 ( .A(n_xor_module_40_res), .ZN(n_not_module_12_res) );
  AND2_X1 u_and_module_32_U1 ( .A1(n_not_module_12_res), .A2(
        n_reg_module_56_res), .ZN(n_and_module_32_res) );
  XOR2_X1 u_xor_module_92_U1 ( .A(p_rand_5), .B(n_xor_module_33_res), .Z(
        n_xor_module_92_res) );
  DFF_X1 u_reg_module_57__hpc_r0_reg ( .D(n_xor_module_33_res), .CK(clock_0), 
        .Q(n_reg_module_57_res), .QN() );
  AND2_X1 u_and_module_33_U1 ( .A1(n_reg_module_57_res), .A2(
        n_xor_module_39_res), .ZN(n_and_module_33_res) );
  DFF_X1 u_reg_module_58__hpc_r0_reg ( .D(n_and_module_33_res), .CK(clock_0), 
        .Q(n_reg_module_58_res), .QN() );
  DFF_X1 u_reg_module_59__hpc_r0_reg ( .D(n_xor_module_91_res), .CK(clock_0), 
        .Q(n_reg_module_59_res), .QN() );
  AND2_X1 u_and_module_34_U1 ( .A1(n_reg_module_59_res), .A2(
        n_xor_module_39_res), .ZN(n_and_module_34_res) );
  DFF_X1 u_reg_module_60__hpc_r0_reg ( .D(n_and_module_34_res), .CK(clock_0), 
        .Q(n_reg_module_60_res), .QN() );
  DFF_X1 u_reg_module_61__hpc_r0_reg ( .D(n_and_module_31_res), .CK(clock_0), 
        .Q(n_reg_module_61_res), .QN() );
  XOR2_X1 u_xor_module_93_U1 ( .A(n_reg_module_61_res), .B(n_reg_module_60_res), .Z(n_xor_module_93_res) );
  XOR2_X1 u_xor_module_94_U1 ( .A(n_xor_module_93_res), .B(n_reg_module_58_res), .Z(n_xor_module_94_res) );
  DFF_X1 u_reg_module_62__hpc_r0_reg ( .D(n_xor_module_34_res), .CK(clock_0), 
        .Q(n_reg_module_62_res), .QN() );
  AND2_X1 u_and_module_35_U1 ( .A1(n_reg_module_62_res), .A2(
        n_xor_module_40_res), .ZN(n_and_module_35_res) );
  DFF_X1 u_reg_module_63__hpc_r0_reg ( .D(n_and_module_35_res), .CK(clock_0), 
        .Q(n_reg_module_63_res), .QN() );
  DFF_X1 u_reg_module_64__hpc_r0_reg ( .D(n_xor_module_92_res), .CK(clock_0), 
        .Q(n_reg_module_64_res), .QN() );
  AND2_X1 u_and_module_36_U1 ( .A1(n_reg_module_64_res), .A2(
        n_xor_module_40_res), .ZN(n_and_module_36_res) );
  DFF_X1 u_reg_module_65__hpc_r0_reg ( .D(n_and_module_36_res), .CK(clock_0), 
        .Q(n_reg_module_65_res), .QN() );
  DFF_X1 u_reg_module_66__hpc_r0_reg ( .D(n_and_module_32_res), .CK(clock_0), 
        .Q(n_reg_module_66_res), .QN() );
  XOR2_X1 u_xor_module_95_U1 ( .A(n_reg_module_66_res), .B(n_reg_module_65_res), .Z(n_xor_module_95_res) );
  XOR2_X1 u_xor_module_96_U1 ( .A(n_xor_module_95_res), .B(n_reg_module_63_res), .Z(n_xor_module_96_res) );
  XOR2_X1 u_xor_module_97_U1 ( .A(n_xor_module_80_res), .B(n_xor_module_94_res), .Z(n_xor_module_97_res) );
  XOR2_X1 u_xor_module_98_U1 ( .A(n_xor_module_82_res), .B(n_xor_module_96_res), .Z(n_xor_module_98_res) );
  DFF_X1 u_reg_module_67__hpc_r0_reg ( .D(p_rand_6), .CK(clock_0), .Q(
        n_reg_module_67_res), .QN() );
  INV_X1 u_not_module_13_U1 ( .A(n_xor_module_1_res), .ZN(n_not_module_13_res)
         );
  AND2_X1 u_and_module_37_U1 ( .A1(n_not_module_13_res), .A2(
        n_reg_module_67_res), .ZN(n_and_module_37_res) );
  XOR2_X1 u_xor_module_99_U1 ( .A(p_rand_6), .B(n_xor_module_30_res), .Z(
        n_xor_module_99_res) );
  INV_X1 u_not_module_14_U1 ( .A(n_xor_module_2_res), .ZN(n_not_module_14_res)
         );
  AND2_X1 u_and_module_38_U1 ( .A1(n_not_module_14_res), .A2(
        n_reg_module_67_res), .ZN(n_and_module_38_res) );
  XOR2_X1 u_xor_module_100_U1 ( .A(p_rand_6), .B(n_xor_module_29_res), .Z(
        n_xor_module_100_res) );
  DFF_X1 u_reg_module_68__hpc_r0_reg ( .D(n_xor_module_29_res), .CK(clock_0), 
        .Q(n_reg_module_68_res), .QN() );
  AND2_X1 u_and_module_39_U1 ( .A1(n_reg_module_68_res), .A2(
        n_xor_module_1_res), .ZN(n_and_module_39_res) );
  DFF_X1 u_reg_module_69__hpc_r0_reg ( .D(n_and_module_39_res), .CK(clock_0), 
        .Q(n_reg_module_69_res), .QN() );
  DFF_X1 u_reg_module_70__hpc_r0_reg ( .D(n_xor_module_99_res), .CK(clock_0), 
        .Q(n_reg_module_70_res), .QN() );
  AND2_X1 u_and_module_40_U1 ( .A1(n_reg_module_70_res), .A2(
        n_xor_module_1_res), .ZN(n_and_module_40_res) );
  DFF_X1 u_reg_module_71__hpc_r0_reg ( .D(n_and_module_40_res), .CK(clock_0), 
        .Q(n_reg_module_71_res), .QN() );
  DFF_X1 u_reg_module_72__hpc_r0_reg ( .D(n_and_module_37_res), .CK(clock_0), 
        .Q(n_reg_module_72_res), .QN() );
  XOR2_X1 u_xor_module_101_U1 ( .A(n_reg_module_72_res), .B(
        n_reg_module_71_res), .Z(n_xor_module_101_res) );
  XOR2_X1 u_xor_module_102_U1 ( .A(n_xor_module_101_res), .B(
        n_reg_module_69_res), .Z(n_xor_module_102_res) );
  DFF_X1 u_reg_module_73__hpc_r0_reg ( .D(n_xor_module_30_res), .CK(clock_0), 
        .Q(n_reg_module_73_res), .QN() );
  AND2_X1 u_and_module_41_U1 ( .A1(n_reg_module_73_res), .A2(
        n_xor_module_2_res), .ZN(n_and_module_41_res) );
  DFF_X1 u_reg_module_74__hpc_r0_reg ( .D(n_and_module_41_res), .CK(clock_0), 
        .Q(n_reg_module_74_res), .QN() );
  DFF_X1 u_reg_module_75__hpc_r0_reg ( .D(n_xor_module_100_res), .CK(clock_0), 
        .Q(n_reg_module_75_res), .QN() );
  AND2_X1 u_and_module_42_U1 ( .A1(n_reg_module_75_res), .A2(
        n_xor_module_2_res), .ZN(n_and_module_42_res) );
  DFF_X1 u_reg_module_76__hpc_r0_reg ( .D(n_and_module_42_res), .CK(clock_0), 
        .Q(n_reg_module_76_res), .QN() );
  DFF_X1 u_reg_module_77__hpc_r0_reg ( .D(n_and_module_38_res), .CK(clock_0), 
        .Q(n_reg_module_77_res), .QN() );
  XOR2_X1 u_xor_module_103_U1 ( .A(n_reg_module_77_res), .B(
        n_reg_module_76_res), .Z(n_xor_module_103_res) );
  XOR2_X1 u_xor_module_104_U1 ( .A(n_xor_module_103_res), .B(
        n_reg_module_74_res), .Z(n_xor_module_104_res) );
  DFF_X1 u_reg_module_78__hpc_r0_reg ( .D(p_rand_7), .CK(clock_0), .Q(
        n_reg_module_78_res), .QN() );
  INV_X1 u_not_module_15_U1 ( .A(n_xor_module_7_res), .ZN(n_not_module_15_res)
         );
  AND2_X1 u_and_module_43_U1 ( .A1(n_not_module_15_res), .A2(
        n_reg_module_78_res), .ZN(n_and_module_43_res) );
  XOR2_X1 u_xor_module_105_U1 ( .A(p_rand_7), .B(n_xor_module_54_res), .Z(
        n_xor_module_105_res) );
  INV_X1 u_not_module_16_U1 ( .A(n_xor_module_8_res), .ZN(n_not_module_16_res)
         );
  AND2_X1 u_and_module_44_U1 ( .A1(n_not_module_16_res), .A2(
        n_reg_module_78_res), .ZN(n_and_module_44_res) );
  XOR2_X1 u_xor_module_106_U1 ( .A(p_rand_7), .B(n_xor_module_53_res), .Z(
        n_xor_module_106_res) );
  DFF_X1 u_reg_module_79__hpc_r0_reg ( .D(n_xor_module_53_res), .CK(clock_0), 
        .Q(n_reg_module_79_res), .QN() );
  AND2_X1 u_and_module_45_U1 ( .A1(n_reg_module_79_res), .A2(
        n_xor_module_7_res), .ZN(n_and_module_45_res) );
  DFF_X1 u_reg_module_80__hpc_r0_reg ( .D(n_and_module_45_res), .CK(clock_0), 
        .Q(n_reg_module_80_res), .QN() );
  DFF_X1 u_reg_module_81__hpc_r0_reg ( .D(n_xor_module_105_res), .CK(clock_0), 
        .Q(n_reg_module_81_res), .QN() );
  AND2_X1 u_and_module_46_U1 ( .A1(n_reg_module_81_res), .A2(
        n_xor_module_7_res), .ZN(n_and_module_46_res) );
  DFF_X1 u_reg_module_82__hpc_r0_reg ( .D(n_and_module_46_res), .CK(clock_0), 
        .Q(n_reg_module_82_res), .QN() );
  DFF_X1 u_reg_module_83__hpc_r0_reg ( .D(n_and_module_43_res), .CK(clock_0), 
        .Q(n_reg_module_83_res), .QN() );
  XOR2_X1 u_xor_module_107_U1 ( .A(n_reg_module_83_res), .B(
        n_reg_module_82_res), .Z(n_xor_module_107_res) );
  XOR2_X1 u_xor_module_108_U1 ( .A(n_xor_module_107_res), .B(
        n_reg_module_80_res), .Z(n_xor_module_108_res) );
  DFF_X1 u_reg_module_84__hpc_r0_reg ( .D(n_xor_module_54_res), .CK(clock_0), 
        .Q(n_reg_module_84_res), .QN() );
  AND2_X1 u_and_module_47_U1 ( .A1(n_reg_module_84_res), .A2(
        n_xor_module_8_res), .ZN(n_and_module_47_res) );
  DFF_X1 u_reg_module_85__hpc_r0_reg ( .D(n_and_module_47_res), .CK(clock_0), 
        .Q(n_reg_module_85_res), .QN() );
  DFF_X1 u_reg_module_86__hpc_r0_reg ( .D(n_xor_module_106_res), .CK(clock_0), 
        .Q(n_reg_module_86_res), .QN() );
  AND2_X1 u_and_module_48_U1 ( .A1(n_reg_module_86_res), .A2(
        n_xor_module_8_res), .ZN(n_and_module_48_res) );
  DFF_X1 u_reg_module_87__hpc_r0_reg ( .D(n_and_module_48_res), .CK(clock_0), 
        .Q(n_reg_module_87_res), .QN() );
  DFF_X1 u_reg_module_88__hpc_r0_reg ( .D(n_and_module_44_res), .CK(clock_0), 
        .Q(n_reg_module_88_res), .QN() );
  XOR2_X1 u_xor_module_109_U1 ( .A(n_reg_module_88_res), .B(
        n_reg_module_87_res), .Z(n_xor_module_109_res) );
  XOR2_X1 u_xor_module_110_U1 ( .A(n_xor_module_109_res), .B(
        n_reg_module_85_res), .Z(n_xor_module_110_res) );
  XOR2_X1 u_xor_module_111_U1 ( .A(n_xor_module_102_res), .B(
        n_xor_module_108_res), .Z(n_xor_module_111_res) );
  XOR2_X1 u_xor_module_112_U1 ( .A(n_xor_module_104_res), .B(
        n_xor_module_110_res), .Z(n_xor_module_112_res) );
  DFF_X1 u_reg_module_89__hpc_r0_reg ( .D(p_rand_8), .CK(clock_0), .Q(
        n_reg_module_89_res), .QN() );
  INV_X1 u_not_module_17_U1 ( .A(n_xor_module_3_res), .ZN(n_not_module_17_res)
         );
  AND2_X1 u_and_module_49_U1 ( .A1(n_not_module_17_res), .A2(
        n_reg_module_89_res), .ZN(n_and_module_49_res) );
  XOR2_X1 u_xor_module_113_U1 ( .A(p_rand_8), .B(n_xor_module_20_res), .Z(
        n_xor_module_113_res) );
  INV_X1 u_not_module_18_U1 ( .A(n_xor_module_4_res), .ZN(n_not_module_18_res)
         );
  AND2_X1 u_and_module_50_U1 ( .A1(n_not_module_18_res), .A2(
        n_reg_module_89_res), .ZN(n_and_module_50_res) );
  XOR2_X1 u_xor_module_114_U1 ( .A(p_rand_8), .B(n_xor_module_19_res), .Z(
        n_xor_module_114_res) );
  DFF_X1 u_reg_module_90__hpc_r0_reg ( .D(n_xor_module_19_res), .CK(clock_0), 
        .Q(n_reg_module_90_res), .QN() );
  AND2_X1 u_and_module_51_U1 ( .A1(n_reg_module_90_res), .A2(
        n_xor_module_3_res), .ZN(n_and_module_51_res) );
  DFF_X1 u_reg_module_91__hpc_r0_reg ( .D(n_and_module_51_res), .CK(clock_0), 
        .Q(n_reg_module_91_res), .QN() );
  DFF_X1 u_reg_module_92__hpc_r0_reg ( .D(n_xor_module_113_res), .CK(clock_0), 
        .Q(n_reg_module_92_res), .QN() );
  AND2_X1 u_and_module_52_U1 ( .A1(n_reg_module_92_res), .A2(
        n_xor_module_3_res), .ZN(n_and_module_52_res) );
  DFF_X1 u_reg_module_93__hpc_r0_reg ( .D(n_and_module_52_res), .CK(clock_0), 
        .Q(n_reg_module_93_res), .QN() );
  DFF_X1 u_reg_module_94__hpc_r0_reg ( .D(n_and_module_49_res), .CK(clock_0), 
        .Q(n_reg_module_94_res), .QN() );
  XOR2_X1 u_xor_module_115_U1 ( .A(n_reg_module_94_res), .B(
        n_reg_module_93_res), .Z(n_xor_module_115_res) );
  XOR2_X1 u_xor_module_116_U1 ( .A(n_xor_module_115_res), .B(
        n_reg_module_91_res), .Z(n_xor_module_116_res) );
  DFF_X1 u_reg_module_95__hpc_r0_reg ( .D(n_xor_module_20_res), .CK(clock_0), 
        .Q(n_reg_module_95_res), .QN() );
  AND2_X1 u_and_module_53_U1 ( .A1(n_reg_module_95_res), .A2(
        n_xor_module_4_res), .ZN(n_and_module_53_res) );
  DFF_X1 u_reg_module_96__hpc_r0_reg ( .D(n_and_module_53_res), .CK(clock_0), 
        .Q(n_reg_module_96_res), .QN() );
  DFF_X1 u_reg_module_97__hpc_r0_reg ( .D(n_xor_module_114_res), .CK(clock_0), 
        .Q(n_reg_module_97_res), .QN() );
  AND2_X1 u_and_module_54_U1 ( .A1(n_reg_module_97_res), .A2(
        n_xor_module_4_res), .ZN(n_and_module_54_res) );
  DFF_X1 u_reg_module_98__hpc_r0_reg ( .D(n_and_module_54_res), .CK(clock_0), 
        .Q(n_reg_module_98_res), .QN() );
  DFF_X1 u_reg_module_99__hpc_r0_reg ( .D(n_and_module_50_res), .CK(clock_0), 
        .Q(n_reg_module_99_res), .QN() );
  XOR2_X1 u_xor_module_117_U1 ( .A(n_reg_module_99_res), .B(
        n_reg_module_98_res), .Z(n_xor_module_117_res) );
  XOR2_X1 u_xor_module_118_U1 ( .A(n_xor_module_117_res), .B(
        n_reg_module_96_res), .Z(n_xor_module_118_res) );
  XOR2_X1 u_xor_module_119_U1 ( .A(n_xor_module_102_res), .B(
        n_xor_module_116_res), .Z(n_xor_module_119_res) );
  XOR2_X1 u_xor_module_120_U1 ( .A(n_xor_module_104_res), .B(
        n_xor_module_118_res), .Z(n_xor_module_120_res) );
  XOR2_X1 u_xor_module_121_U1 ( .A(n_xor_module_64_res), .B(
        n_xor_module_67_res), .Z(n_xor_module_121_res) );
  XOR2_X1 u_xor_module_122_U1 ( .A(n_xor_module_66_res), .B(
        n_xor_module_68_res), .Z(n_xor_module_122_res) );
  XOR2_X1 u_xor_module_123_U1 ( .A(n_xor_module_47_res), .B(
        n_xor_module_75_res), .Z(n_xor_module_123_res) );
  XOR2_X1 u_xor_module_124_U1 ( .A(n_xor_module_48_res), .B(
        n_xor_module_76_res), .Z(n_xor_module_124_res) );
  XOR2_X1 u_xor_module_125_U1 ( .A(n_xor_module_86_res), .B(
        n_xor_module_89_res), .Z(n_xor_module_125_res) );
  XOR2_X1 u_xor_module_126_U1 ( .A(n_xor_module_88_res), .B(
        n_xor_module_90_res), .Z(n_xor_module_126_res) );
  XOR2_X1 u_xor_module_127_U1 ( .A(n_xor_module_119_res), .B(
        n_xor_module_97_res), .Z(n_xor_module_127_res) );
  XOR2_X1 u_xor_module_128_U1 ( .A(n_xor_module_120_res), .B(
        n_xor_module_98_res), .Z(n_xor_module_128_res) );
  XOR2_X1 u_xor_module_129_U1 ( .A(n_xor_module_111_res), .B(
        n_xor_module_121_res), .Z(n_xor_module_129_res) );
  XOR2_X1 u_xor_module_130_U1 ( .A(n_xor_module_112_res), .B(
        n_xor_module_122_res), .Z(n_xor_module_130_res) );
  XOR2_X1 u_xor_module_131_U1 ( .A(n_xor_module_119_res), .B(
        n_xor_module_123_res), .Z(n_xor_module_131_res) );
  XOR2_X1 u_xor_module_132_U1 ( .A(n_xor_module_120_res), .B(
        n_xor_module_124_res), .Z(n_xor_module_132_res) );
  XOR2_X1 u_xor_module_133_U1 ( .A(n_xor_module_111_res), .B(
        n_xor_module_125_res), .Z(n_xor_module_133_res) );
  XOR2_X1 u_xor_module_134_U1 ( .A(n_xor_module_112_res), .B(
        n_xor_module_126_res), .Z(n_xor_module_134_res) );
  XOR2_X1 u_xor_module_135_U1 ( .A(n_xor_module_49_res), .B(
        n_xor_module_127_res), .Z(n_xor_module_135_res) );
  XOR2_X1 u_xor_module_136_U1 ( .A(n_xor_module_50_res), .B(
        n_xor_module_128_res), .Z(n_xor_module_136_res) );
  XOR2_X1 u_xor_module_137_U1 ( .A(n_xor_module_135_res), .B(
        n_xor_module_133_res), .Z(n_xor_module_137_res) );
  XOR2_X1 u_xor_module_138_U1 ( .A(n_xor_module_136_res), .B(
        n_xor_module_134_res), .Z(n_xor_module_138_res) );
  DFF_X1 u_reg_module_100__hpc_r0_reg ( .D(p_rand_9), .CK(clock_0), .Q(
        n_reg_module_100_res), .QN() );
  INV_X1 u_not_module_19_U1 ( .A(n_xor_module_133_res), .ZN(
        n_not_module_19_res) );
  AND2_X1 u_and_module_55_U1 ( .A1(n_not_module_19_res), .A2(
        n_reg_module_100_res), .ZN(n_and_module_55_res) );
  XOR2_X1 u_xor_module_139_U1 ( .A(p_rand_9), .B(n_xor_module_130_res), .Z(
        n_xor_module_139_res) );
  INV_X1 u_not_module_20_U1 ( .A(n_xor_module_134_res), .ZN(
        n_not_module_20_res) );
  AND2_X1 u_and_module_56_U1 ( .A1(n_not_module_20_res), .A2(
        n_reg_module_100_res), .ZN(n_and_module_56_res) );
  XOR2_X1 u_xor_module_140_U1 ( .A(p_rand_9), .B(n_xor_module_129_res), .Z(
        n_xor_module_140_res) );
  DFF_X1 u_reg_module_101__hpc_r0_reg ( .D(n_xor_module_129_res), .CK(clock_0), 
        .Q(n_reg_module_101_res), .QN() );
  AND2_X1 u_and_module_57_U1 ( .A1(n_reg_module_101_res), .A2(
        n_xor_module_133_res), .ZN(n_and_module_57_res) );
  DFF_X1 u_reg_module_102__hpc_r0_reg ( .D(n_and_module_57_res), .CK(clock_0), 
        .Q(n_reg_module_102_res), .QN() );
  DFF_X1 u_reg_module_103__hpc_r0_reg ( .D(n_xor_module_139_res), .CK(clock_0), 
        .Q(n_reg_module_103_res), .QN() );
  AND2_X1 u_and_module_58_U1 ( .A1(n_reg_module_103_res), .A2(
        n_xor_module_133_res), .ZN(n_and_module_58_res) );
  DFF_X1 u_reg_module_104__hpc_r0_reg ( .D(n_and_module_58_res), .CK(clock_0), 
        .Q(n_reg_module_104_res), .QN() );
  DFF_X1 u_reg_module_105__hpc_r0_reg ( .D(n_and_module_55_res), .CK(clock_0), 
        .Q(n_reg_module_105_res), .QN() );
  XOR2_X1 u_xor_module_141_U1 ( .A(n_reg_module_105_res), .B(
        n_reg_module_104_res), .Z(n_xor_module_141_res) );
  XOR2_X1 u_xor_module_142_U1 ( .A(n_xor_module_141_res), .B(
        n_reg_module_102_res), .Z(n_xor_module_142_res) );
  DFF_X1 u_reg_module_106__hpc_r0_reg ( .D(n_xor_module_130_res), .CK(clock_0), 
        .Q(n_reg_module_106_res), .QN() );
  AND2_X1 u_and_module_59_U1 ( .A1(n_reg_module_106_res), .A2(
        n_xor_module_134_res), .ZN(n_and_module_59_res) );
  DFF_X1 u_reg_module_107__hpc_r0_reg ( .D(n_and_module_59_res), .CK(clock_0), 
        .Q(n_reg_module_107_res), .QN() );
  DFF_X1 u_reg_module_108__hpc_r0_reg ( .D(n_xor_module_140_res), .CK(clock_0), 
        .Q(n_reg_module_108_res), .QN() );
  AND2_X1 u_and_module_60_U1 ( .A1(n_reg_module_108_res), .A2(
        n_xor_module_134_res), .ZN(n_and_module_60_res) );
  DFF_X1 u_reg_module_109__hpc_r0_reg ( .D(n_and_module_60_res), .CK(clock_0), 
        .Q(n_reg_module_109_res), .QN() );
  DFF_X1 u_reg_module_110__hpc_r0_reg ( .D(n_and_module_56_res), .CK(clock_0), 
        .Q(n_reg_module_110_res), .QN() );
  XOR2_X1 u_xor_module_143_U1 ( .A(n_reg_module_110_res), .B(
        n_reg_module_109_res), .Z(n_xor_module_143_res) );
  XOR2_X1 u_xor_module_144_U1 ( .A(n_xor_module_143_res), .B(
        n_reg_module_107_res), .Z(n_xor_module_144_res) );
  XOR2_X1 u_xor_module_145_U1 ( .A(n_xor_module_142_res), .B(
        n_xor_module_131_res), .Z(n_xor_module_145_res) );
  XOR2_X1 u_xor_module_146_U1 ( .A(n_xor_module_144_res), .B(
        n_xor_module_132_res), .Z(n_xor_module_146_res) );
  XOR2_X1 u_xor_module_147_U1 ( .A(n_xor_module_131_res), .B(
        n_xor_module_129_res), .Z(n_xor_module_147_res) );
  XOR2_X1 u_xor_module_148_U1 ( .A(n_xor_module_132_res), .B(
        n_xor_module_130_res), .Z(n_xor_module_148_res) );
  XOR2_X1 u_xor_module_149_U1 ( .A(n_xor_module_142_res), .B(
        n_xor_module_135_res), .Z(n_xor_module_149_res) );
  XOR2_X1 u_xor_module_150_U1 ( .A(n_xor_module_144_res), .B(
        n_xor_module_136_res), .Z(n_xor_module_150_res) );
  DFF_X1 u_reg_module_111__hpc_r0_reg ( .D(p_rand_10), .CK(clock_0), .Q(
        n_reg_module_111_res), .QN() );
  INV_X1 u_not_module_21_U1 ( .A(n_xor_module_149_res), .ZN(
        n_not_module_21_res) );
  AND2_X1 u_and_module_61_U1 ( .A1(n_not_module_21_res), .A2(
        n_reg_module_111_res), .ZN(n_and_module_61_res) );
  XOR2_X1 u_xor_module_151_U1 ( .A(p_rand_10), .B(n_xor_module_148_res), .Z(
        n_xor_module_151_res) );
  INV_X1 u_not_module_22_U1 ( .A(n_xor_module_150_res), .ZN(
        n_not_module_22_res) );
  AND2_X1 u_and_module_62_U1 ( .A1(n_not_module_22_res), .A2(
        n_reg_module_111_res), .ZN(n_and_module_62_res) );
  XOR2_X1 u_xor_module_152_U1 ( .A(p_rand_10), .B(n_xor_module_147_res), .Z(
        n_xor_module_152_res) );
  DFF_X1 u_reg_module_112__hpc_r0_reg ( .D(n_xor_module_147_res), .CK(clock_0), 
        .Q(n_reg_module_112_res), .QN() );
  AND2_X1 u_and_module_63_U1 ( .A1(n_reg_module_112_res), .A2(
        n_xor_module_149_res), .ZN(n_and_module_63_res) );
  DFF_X1 u_reg_module_113__hpc_r0_reg ( .D(n_and_module_63_res), .CK(clock_0), 
        .Q(n_reg_module_113_res), .QN() );
  DFF_X1 u_reg_module_114__hpc_r0_reg ( .D(n_xor_module_151_res), .CK(clock_0), 
        .Q(n_reg_module_114_res), .QN() );
  AND2_X1 u_and_module_64_U1 ( .A1(n_reg_module_114_res), .A2(
        n_xor_module_149_res), .ZN(n_and_module_64_res) );
  DFF_X1 u_reg_module_115__hpc_r0_reg ( .D(n_and_module_64_res), .CK(clock_0), 
        .Q(n_reg_module_115_res), .QN() );
  DFF_X1 u_reg_module_116__hpc_r0_reg ( .D(n_and_module_61_res), .CK(clock_0), 
        .Q(n_reg_module_116_res), .QN() );
  XOR2_X1 u_xor_module_153_U1 ( .A(n_reg_module_116_res), .B(
        n_reg_module_115_res), .Z(n_xor_module_153_res) );
  XOR2_X1 u_xor_module_154_U1 ( .A(n_xor_module_153_res), .B(
        n_reg_module_113_res), .Z(n_xor_module_154_res) );
  DFF_X1 u_reg_module_117__hpc_r0_reg ( .D(n_xor_module_148_res), .CK(clock_0), 
        .Q(n_reg_module_117_res), .QN() );
  AND2_X1 u_and_module_65_U1 ( .A1(n_reg_module_117_res), .A2(
        n_xor_module_150_res), .ZN(n_and_module_65_res) );
  DFF_X1 u_reg_module_118__hpc_r0_reg ( .D(n_and_module_65_res), .CK(clock_0), 
        .Q(n_reg_module_118_res), .QN() );
  DFF_X1 u_reg_module_119__hpc_r0_reg ( .D(n_xor_module_152_res), .CK(clock_0), 
        .Q(n_reg_module_119_res), .QN() );
  AND2_X1 u_and_module_66_U1 ( .A1(n_reg_module_119_res), .A2(
        n_xor_module_150_res), .ZN(n_and_module_66_res) );
  DFF_X1 u_reg_module_120__hpc_r0_reg ( .D(n_and_module_66_res), .CK(clock_0), 
        .Q(n_reg_module_120_res), .QN() );
  DFF_X1 u_reg_module_121__hpc_r0_reg ( .D(n_and_module_62_res), .CK(clock_0), 
        .Q(n_reg_module_121_res), .QN() );
  XOR2_X1 u_xor_module_155_U1 ( .A(n_reg_module_121_res), .B(
        n_reg_module_120_res), .Z(n_xor_module_155_res) );
  XOR2_X1 u_xor_module_156_U1 ( .A(n_xor_module_155_res), .B(
        n_reg_module_118_res), .Z(n_xor_module_156_res) );
  DFF_X1 u_reg_module_122__hpc_r0_reg ( .D(p_rand_11), .CK(clock_0), .Q(
        n_reg_module_122_res), .QN() );
  INV_X1 u_not_module_23_U1 ( .A(n_xor_module_145_res), .ZN(
        n_not_module_23_res) );
  AND2_X1 u_and_module_67_U1 ( .A1(n_not_module_23_res), .A2(
        n_reg_module_122_res), .ZN(n_and_module_67_res) );
  XOR2_X1 u_xor_module_157_U1 ( .A(p_rand_11), .B(n_xor_module_138_res), .Z(
        n_xor_module_157_res) );
  INV_X1 u_not_module_24_U1 ( .A(n_xor_module_146_res), .ZN(
        n_not_module_24_res) );
  AND2_X1 u_and_module_68_U1 ( .A1(n_not_module_24_res), .A2(
        n_reg_module_122_res), .ZN(n_and_module_68_res) );
  XOR2_X1 u_xor_module_158_U1 ( .A(p_rand_11), .B(n_xor_module_137_res), .Z(
        n_xor_module_158_res) );
  DFF_X1 u_reg_module_123__hpc_r0_reg ( .D(n_xor_module_137_res), .CK(clock_0), 
        .Q(n_reg_module_123_res), .QN() );
  AND2_X1 u_and_module_69_U1 ( .A1(n_reg_module_123_res), .A2(
        n_xor_module_145_res), .ZN(n_and_module_69_res) );
  DFF_X1 u_reg_module_124__hpc_r0_reg ( .D(n_and_module_69_res), .CK(clock_0), 
        .Q(n_reg_module_124_res), .QN() );
  DFF_X1 u_reg_module_125__hpc_r0_reg ( .D(n_xor_module_157_res), .CK(clock_0), 
        .Q(n_reg_module_125_res), .QN() );
  AND2_X1 u_and_module_70_U1 ( .A1(n_reg_module_125_res), .A2(
        n_xor_module_145_res), .ZN(n_and_module_70_res) );
  DFF_X1 u_reg_module_126__hpc_r0_reg ( .D(n_and_module_70_res), .CK(clock_0), 
        .Q(n_reg_module_126_res), .QN() );
  DFF_X1 u_reg_module_127__hpc_r0_reg ( .D(n_and_module_67_res), .CK(clock_0), 
        .Q(n_reg_module_127_res), .QN() );
  XOR2_X1 u_xor_module_159_U1 ( .A(n_reg_module_127_res), .B(
        n_reg_module_126_res), .Z(n_xor_module_159_res) );
  XOR2_X1 u_xor_module_160_U1 ( .A(n_xor_module_159_res), .B(
        n_reg_module_124_res), .Z(n_xor_module_160_res) );
  DFF_X1 u_reg_module_128__hpc_r0_reg ( .D(n_xor_module_138_res), .CK(clock_0), 
        .Q(n_reg_module_128_res), .QN() );
  AND2_X1 u_and_module_71_U1 ( .A1(n_reg_module_128_res), .A2(
        n_xor_module_146_res), .ZN(n_and_module_71_res) );
  DFF_X1 u_reg_module_129__hpc_r0_reg ( .D(n_and_module_71_res), .CK(clock_0), 
        .Q(n_reg_module_129_res), .QN() );
  DFF_X1 u_reg_module_130__hpc_r0_reg ( .D(n_xor_module_158_res), .CK(clock_0), 
        .Q(n_reg_module_130_res), .QN() );
  AND2_X1 u_and_module_72_U1 ( .A1(n_reg_module_130_res), .A2(
        n_xor_module_146_res), .ZN(n_and_module_72_res) );
  DFF_X1 u_reg_module_131__hpc_r0_reg ( .D(n_and_module_72_res), .CK(clock_0), 
        .Q(n_reg_module_131_res), .QN() );
  DFF_X1 u_reg_module_132__hpc_r0_reg ( .D(n_and_module_68_res), .CK(clock_0), 
        .Q(n_reg_module_132_res), .QN() );
  XOR2_X1 u_xor_module_161_U1 ( .A(n_reg_module_132_res), .B(
        n_reg_module_131_res), .Z(n_xor_module_161_res) );
  XOR2_X1 u_xor_module_162_U1 ( .A(n_xor_module_161_res), .B(
        n_reg_module_129_res), .Z(n_xor_module_162_res) );
  DFF_X1 u_reg_module_133__hpc_r0_reg ( .D(p_rand_12), .CK(clock_0), .Q(
        n_reg_module_133_res), .QN() );
  INV_X1 u_not_module_25_U1 ( .A(n_xor_module_129_res), .ZN(
        n_not_module_25_res) );
  AND2_X1 u_and_module_73_U1 ( .A1(n_not_module_25_res), .A2(
        n_reg_module_133_res), .ZN(n_and_module_73_res) );
  XOR2_X1 u_xor_module_163_U1 ( .A(p_rand_12), .B(n_xor_module_136_res), .Z(
        n_xor_module_163_res) );
  INV_X1 u_not_module_26_U1 ( .A(n_xor_module_130_res), .ZN(
        n_not_module_26_res) );
  AND2_X1 u_and_module_74_U1 ( .A1(n_not_module_26_res), .A2(
        n_reg_module_133_res), .ZN(n_and_module_74_res) );
  XOR2_X1 u_xor_module_164_U1 ( .A(p_rand_12), .B(n_xor_module_135_res), .Z(
        n_xor_module_164_res) );
  DFF_X1 u_reg_module_134__hpc_r0_reg ( .D(n_xor_module_135_res), .CK(clock_0), 
        .Q(n_reg_module_134_res), .QN() );
  AND2_X1 u_and_module_75_U1 ( .A1(n_reg_module_134_res), .A2(
        n_xor_module_129_res), .ZN(n_and_module_75_res) );
  DFF_X1 u_reg_module_135__hpc_r0_reg ( .D(n_and_module_75_res), .CK(clock_0), 
        .Q(n_reg_module_135_res), .QN() );
  DFF_X1 u_reg_module_136__hpc_r0_reg ( .D(n_xor_module_163_res), .CK(clock_0), 
        .Q(n_reg_module_136_res), .QN() );
  AND2_X1 u_and_module_76_U1 ( .A1(n_reg_module_136_res), .A2(
        n_xor_module_129_res), .ZN(n_and_module_76_res) );
  DFF_X1 u_reg_module_137__hpc_r0_reg ( .D(n_and_module_76_res), .CK(clock_0), 
        .Q(n_reg_module_137_res), .QN() );
  DFF_X1 u_reg_module_138__hpc_r0_reg ( .D(n_and_module_73_res), .CK(clock_0), 
        .Q(n_reg_module_138_res), .QN() );
  XOR2_X1 u_xor_module_165_U1 ( .A(n_reg_module_138_res), .B(
        n_reg_module_137_res), .Z(n_xor_module_165_res) );
  XOR2_X1 u_xor_module_166_U1 ( .A(n_xor_module_165_res), .B(
        n_reg_module_135_res), .Z(n_xor_module_166_res) );
  DFF_X1 u_reg_module_139__hpc_r0_reg ( .D(n_xor_module_136_res), .CK(clock_0), 
        .Q(n_reg_module_139_res), .QN() );
  AND2_X1 u_and_module_77_U1 ( .A1(n_reg_module_139_res), .A2(
        n_xor_module_130_res), .ZN(n_and_module_77_res) );
  DFF_X1 u_reg_module_140__hpc_r0_reg ( .D(n_and_module_77_res), .CK(clock_0), 
        .Q(n_reg_module_140_res), .QN() );
  DFF_X1 u_reg_module_141__hpc_r0_reg ( .D(n_xor_module_164_res), .CK(clock_0), 
        .Q(n_reg_module_141_res), .QN() );
  AND2_X1 u_and_module_78_U1 ( .A1(n_reg_module_141_res), .A2(
        n_xor_module_130_res), .ZN(n_and_module_78_res) );
  DFF_X1 u_reg_module_142__hpc_r0_reg ( .D(n_and_module_78_res), .CK(clock_0), 
        .Q(n_reg_module_142_res), .QN() );
  DFF_X1 u_reg_module_143__hpc_r0_reg ( .D(n_and_module_74_res), .CK(clock_0), 
        .Q(n_reg_module_143_res), .QN() );
  XOR2_X1 u_xor_module_167_U1 ( .A(n_reg_module_143_res), .B(
        n_reg_module_142_res), .Z(n_xor_module_167_res) );
  XOR2_X1 u_xor_module_168_U1 ( .A(n_xor_module_167_res), .B(
        n_reg_module_140_res), .Z(n_xor_module_168_res) );
  DFF_X1 u_reg_module_144__hpc_r0_reg ( .D(p_rand_13), .CK(clock_0), .Q(
        n_reg_module_144_res), .QN() );
  INV_X1 u_not_module_27_U1 ( .A(n_xor_module_147_res), .ZN(
        n_not_module_27_res) );
  AND2_X1 u_and_module_79_U1 ( .A1(n_not_module_27_res), .A2(
        n_reg_module_144_res), .ZN(n_and_module_79_res) );
  XOR2_X1 u_xor_module_169_U1 ( .A(p_rand_13), .B(n_xor_module_168_res), .Z(
        n_xor_module_169_res) );
  INV_X1 u_not_module_28_U1 ( .A(n_xor_module_148_res), .ZN(
        n_not_module_28_res) );
  AND2_X1 u_and_module_80_U1 ( .A1(n_not_module_28_res), .A2(
        n_reg_module_144_res), .ZN(n_and_module_80_res) );
  XOR2_X1 u_xor_module_170_U1 ( .A(p_rand_13), .B(n_xor_module_166_res), .Z(
        n_xor_module_170_res) );
  DFF_X1 u_reg_module_145__hpc_r0_reg ( .D(n_xor_module_166_res), .CK(clock_0), 
        .Q(n_reg_module_145_res), .QN() );
  AND2_X1 u_and_module_81_U1 ( .A1(n_reg_module_145_res), .A2(
        n_xor_module_147_res), .ZN(n_and_module_81_res) );
  DFF_X1 u_reg_module_146__hpc_r0_reg ( .D(n_and_module_81_res), .CK(clock_0), 
        .Q(n_reg_module_146_res), .QN() );
  DFF_X1 u_reg_module_147__hpc_r0_reg ( .D(n_xor_module_169_res), .CK(clock_0), 
        .Q(n_reg_module_147_res), .QN() );
  AND2_X1 u_and_module_82_U1 ( .A1(n_reg_module_147_res), .A2(
        n_xor_module_147_res), .ZN(n_and_module_82_res) );
  DFF_X1 u_reg_module_148__hpc_r0_reg ( .D(n_and_module_82_res), .CK(clock_0), 
        .Q(n_reg_module_148_res), .QN() );
  DFF_X1 u_reg_module_149__hpc_r0_reg ( .D(n_and_module_79_res), .CK(clock_0), 
        .Q(n_reg_module_149_res), .QN() );
  XOR2_X1 u_xor_module_171_U1 ( .A(n_reg_module_149_res), .B(
        n_reg_module_148_res), .Z(n_xor_module_171_res) );
  XOR2_X1 u_xor_module_172_U1 ( .A(n_xor_module_171_res), .B(
        n_reg_module_146_res), .Z(n_xor_module_172_res) );
  DFF_X1 u_reg_module_150__hpc_r0_reg ( .D(n_xor_module_168_res), .CK(clock_0), 
        .Q(n_reg_module_150_res), .QN() );
  AND2_X1 u_and_module_83_U1 ( .A1(n_reg_module_150_res), .A2(
        n_xor_module_148_res), .ZN(n_and_module_83_res) );
  DFF_X1 u_reg_module_151__hpc_r0_reg ( .D(n_and_module_83_res), .CK(clock_0), 
        .Q(n_reg_module_151_res), .QN() );
  DFF_X1 u_reg_module_152__hpc_r0_reg ( .D(n_xor_module_170_res), .CK(clock_0), 
        .Q(n_reg_module_152_res), .QN() );
  AND2_X1 u_and_module_84_U1 ( .A1(n_reg_module_152_res), .A2(
        n_xor_module_148_res), .ZN(n_and_module_84_res) );
  DFF_X1 u_reg_module_153__hpc_r0_reg ( .D(n_and_module_84_res), .CK(clock_0), 
        .Q(n_reg_module_153_res), .QN() );
  DFF_X1 u_reg_module_154__hpc_r0_reg ( .D(n_and_module_80_res), .CK(clock_0), 
        .Q(n_reg_module_154_res), .QN() );
  XOR2_X1 u_xor_module_173_U1 ( .A(n_reg_module_154_res), .B(
        n_reg_module_153_res), .Z(n_xor_module_173_res) );
  XOR2_X1 u_xor_module_174_U1 ( .A(n_xor_module_173_res), .B(
        n_reg_module_151_res), .Z(n_xor_module_174_res) );
  XOR2_X1 u_xor_module_175_U1 ( .A(n_xor_module_142_res), .B(
        n_xor_module_147_res), .Z(n_xor_module_175_res) );
  XOR2_X1 u_xor_module_176_U1 ( .A(n_xor_module_144_res), .B(
        n_xor_module_148_res), .Z(n_xor_module_176_res) );
  DFF_X1 u_reg_module_155__hpc_r0_reg ( .D(p_rand_14), .CK(clock_0), .Q(
        n_reg_module_155_res), .QN() );
  INV_X1 u_not_module_29_U1 ( .A(n_xor_module_131_res), .ZN(
        n_not_module_29_res) );
  AND2_X1 u_and_module_85_U1 ( .A1(n_not_module_29_res), .A2(
        n_reg_module_155_res), .ZN(n_and_module_85_res) );
  XOR2_X1 u_xor_module_177_U1 ( .A(p_rand_14), .B(n_xor_module_134_res), .Z(
        n_xor_module_177_res) );
  INV_X1 u_not_module_30_U1 ( .A(n_xor_module_132_res), .ZN(
        n_not_module_30_res) );
  AND2_X1 u_and_module_86_U1 ( .A1(n_not_module_30_res), .A2(
        n_reg_module_155_res), .ZN(n_and_module_86_res) );
  XOR2_X1 u_xor_module_178_U1 ( .A(p_rand_14), .B(n_xor_module_133_res), .Z(
        n_xor_module_178_res) );
  DFF_X1 u_reg_module_156__hpc_r0_reg ( .D(n_xor_module_133_res), .CK(clock_0), 
        .Q(n_reg_module_156_res), .QN() );
  AND2_X1 u_and_module_87_U1 ( .A1(n_reg_module_156_res), .A2(
        n_xor_module_131_res), .ZN(n_and_module_87_res) );
  DFF_X1 u_reg_module_157__hpc_r0_reg ( .D(n_and_module_87_res), .CK(clock_0), 
        .Q(n_reg_module_157_res), .QN() );
  DFF_X1 u_reg_module_158__hpc_r0_reg ( .D(n_xor_module_177_res), .CK(clock_0), 
        .Q(n_reg_module_158_res), .QN() );
  AND2_X1 u_and_module_88_U1 ( .A1(n_reg_module_158_res), .A2(
        n_xor_module_131_res), .ZN(n_and_module_88_res) );
  DFF_X1 u_reg_module_159__hpc_r0_reg ( .D(n_and_module_88_res), .CK(clock_0), 
        .Q(n_reg_module_159_res), .QN() );
  DFF_X1 u_reg_module_160__hpc_r0_reg ( .D(n_and_module_85_res), .CK(clock_0), 
        .Q(n_reg_module_160_res), .QN() );
  XOR2_X1 u_xor_module_179_U1 ( .A(n_reg_module_160_res), .B(
        n_reg_module_159_res), .Z(n_xor_module_179_res) );
  XOR2_X1 u_xor_module_180_U1 ( .A(n_xor_module_179_res), .B(
        n_reg_module_157_res), .Z(n_xor_module_180_res) );
  DFF_X1 u_reg_module_161__hpc_r0_reg ( .D(n_xor_module_134_res), .CK(clock_0), 
        .Q(n_reg_module_161_res), .QN() );
  AND2_X1 u_and_module_89_U1 ( .A1(n_reg_module_161_res), .A2(
        n_xor_module_132_res), .ZN(n_and_module_89_res) );
  DFF_X1 u_reg_module_162__hpc_r0_reg ( .D(n_and_module_89_res), .CK(clock_0), 
        .Q(n_reg_module_162_res), .QN() );
  DFF_X1 u_reg_module_163__hpc_r0_reg ( .D(n_xor_module_178_res), .CK(clock_0), 
        .Q(n_reg_module_163_res), .QN() );
  AND2_X1 u_and_module_90_U1 ( .A1(n_reg_module_163_res), .A2(
        n_xor_module_132_res), .ZN(n_and_module_90_res) );
  DFF_X1 u_reg_module_164__hpc_r0_reg ( .D(n_and_module_90_res), .CK(clock_0), 
        .Q(n_reg_module_164_res), .QN() );
  DFF_X1 u_reg_module_165__hpc_r0_reg ( .D(n_and_module_86_res), .CK(clock_0), 
        .Q(n_reg_module_165_res), .QN() );
  XOR2_X1 u_xor_module_181_U1 ( .A(n_reg_module_165_res), .B(
        n_reg_module_164_res), .Z(n_xor_module_181_res) );
  XOR2_X1 u_xor_module_182_U1 ( .A(n_xor_module_181_res), .B(
        n_reg_module_162_res), .Z(n_xor_module_182_res) );
  DFF_X1 u_reg_module_166__hpc_r0_reg ( .D(p_rand_15), .CK(clock_0), .Q(
        n_reg_module_166_res), .QN() );
  INV_X1 u_not_module_31_U1 ( .A(n_xor_module_137_res), .ZN(
        n_not_module_31_res) );
  AND2_X1 u_and_module_91_U1 ( .A1(n_not_module_31_res), .A2(
        n_reg_module_166_res), .ZN(n_and_module_91_res) );
  XOR2_X1 u_xor_module_183_U1 ( .A(p_rand_15), .B(n_xor_module_182_res), .Z(
        n_xor_module_183_res) );
  INV_X1 u_not_module_32_U1 ( .A(n_xor_module_138_res), .ZN(
        n_not_module_32_res) );
  AND2_X1 u_and_module_92_U1 ( .A1(n_not_module_32_res), .A2(
        n_reg_module_166_res), .ZN(n_and_module_92_res) );
  XOR2_X1 u_xor_module_184_U1 ( .A(p_rand_15), .B(n_xor_module_180_res), .Z(
        n_xor_module_184_res) );
  DFF_X1 u_reg_module_167__hpc_r0_reg ( .D(n_xor_module_180_res), .CK(clock_0), 
        .Q(n_reg_module_167_res), .QN() );
  AND2_X1 u_and_module_93_U1 ( .A1(n_reg_module_167_res), .A2(
        n_xor_module_137_res), .ZN(n_and_module_93_res) );
  DFF_X1 u_reg_module_168__hpc_r0_reg ( .D(n_and_module_93_res), .CK(clock_0), 
        .Q(n_reg_module_168_res), .QN() );
  DFF_X1 u_reg_module_169__hpc_r0_reg ( .D(n_xor_module_183_res), .CK(clock_0), 
        .Q(n_reg_module_169_res), .QN() );
  AND2_X1 u_and_module_94_U1 ( .A1(n_reg_module_169_res), .A2(
        n_xor_module_137_res), .ZN(n_and_module_94_res) );
  DFF_X1 u_reg_module_170__hpc_r0_reg ( .D(n_and_module_94_res), .CK(clock_0), 
        .Q(n_reg_module_170_res), .QN() );
  DFF_X1 u_reg_module_171__hpc_r0_reg ( .D(n_and_module_91_res), .CK(clock_0), 
        .Q(n_reg_module_171_res), .QN() );
  XOR2_X1 u_xor_module_185_U1 ( .A(n_reg_module_171_res), .B(
        n_reg_module_170_res), .Z(n_xor_module_185_res) );
  XOR2_X1 u_xor_module_186_U1 ( .A(n_xor_module_185_res), .B(
        n_reg_module_168_res), .Z(n_xor_module_186_res) );
  DFF_X1 u_reg_module_172__hpc_r0_reg ( .D(n_xor_module_182_res), .CK(clock_0), 
        .Q(n_reg_module_172_res), .QN() );
  AND2_X1 u_and_module_95_U1 ( .A1(n_reg_module_172_res), .A2(
        n_xor_module_138_res), .ZN(n_and_module_95_res) );
  DFF_X1 u_reg_module_173__hpc_r0_reg ( .D(n_and_module_95_res), .CK(clock_0), 
        .Q(n_reg_module_173_res), .QN() );
  DFF_X1 u_reg_module_174__hpc_r0_reg ( .D(n_xor_module_184_res), .CK(clock_0), 
        .Q(n_reg_module_174_res), .QN() );
  AND2_X1 u_and_module_96_U1 ( .A1(n_reg_module_174_res), .A2(
        n_xor_module_138_res), .ZN(n_and_module_96_res) );
  DFF_X1 u_reg_module_175__hpc_r0_reg ( .D(n_and_module_96_res), .CK(clock_0), 
        .Q(n_reg_module_175_res), .QN() );
  DFF_X1 u_reg_module_176__hpc_r0_reg ( .D(n_and_module_92_res), .CK(clock_0), 
        .Q(n_reg_module_176_res), .QN() );
  XOR2_X1 u_xor_module_187_U1 ( .A(n_reg_module_176_res), .B(
        n_reg_module_175_res), .Z(n_xor_module_187_res) );
  XOR2_X1 u_xor_module_188_U1 ( .A(n_xor_module_187_res), .B(
        n_reg_module_173_res), .Z(n_xor_module_188_res) );
  XOR2_X1 u_xor_module_189_U1 ( .A(n_xor_module_142_res), .B(
        n_xor_module_137_res), .Z(n_xor_module_189_res) );
  XOR2_X1 u_xor_module_190_U1 ( .A(n_xor_module_144_res), .B(
        n_xor_module_138_res), .Z(n_xor_module_190_res) );
  XOR2_X1 u_xor_module_191_U1 ( .A(n_xor_module_154_res), .B(
        n_xor_module_131_res), .Z(n_xor_module_191_res) );
  XOR2_X1 u_xor_module_192_U1 ( .A(n_xor_module_156_res), .B(
        n_xor_module_132_res), .Z(n_xor_module_192_res) );
  XOR2_X1 u_xor_module_193_U1 ( .A(n_xor_module_175_res), .B(
        n_xor_module_172_res), .Z(n_xor_module_193_res) );
  XOR2_X1 u_xor_module_194_U1 ( .A(n_xor_module_176_res), .B(
        n_xor_module_174_res), .Z(n_xor_module_194_res) );
  XOR2_X1 u_xor_module_195_U1 ( .A(n_xor_module_160_res), .B(
        n_xor_module_135_res), .Z(n_xor_module_195_res) );
  XOR2_X1 u_xor_module_196_U1 ( .A(n_xor_module_162_res), .B(
        n_xor_module_136_res), .Z(n_xor_module_196_res) );
  XOR2_X1 u_xor_module_197_U1 ( .A(n_xor_module_189_res), .B(
        n_xor_module_186_res), .Z(n_xor_module_197_res) );
  XOR2_X1 u_xor_module_198_U1 ( .A(n_xor_module_190_res), .B(
        n_xor_module_188_res), .Z(n_xor_module_198_res) );
  XOR2_X1 u_xor_module_199_U1 ( .A(n_xor_module_197_res), .B(
        n_xor_module_193_res), .Z(n_xor_module_199_res) );
  XOR2_X1 u_xor_module_200_U1 ( .A(n_xor_module_198_res), .B(
        n_xor_module_194_res), .Z(n_xor_module_200_res) );
  XOR2_X1 u_xor_module_201_U1 ( .A(n_xor_module_195_res), .B(
        n_xor_module_191_res), .Z(n_xor_module_201_res) );
  XOR2_X1 u_xor_module_202_U1 ( .A(n_xor_module_196_res), .B(
        n_xor_module_192_res), .Z(n_xor_module_202_res) );
  XOR2_X1 u_xor_module_203_U1 ( .A(n_xor_module_193_res), .B(
        n_xor_module_191_res), .Z(n_xor_module_203_res) );
  XOR2_X1 u_xor_module_204_U1 ( .A(n_xor_module_194_res), .B(
        n_xor_module_192_res), .Z(n_xor_module_204_res) );
  XOR2_X1 u_xor_module_205_U1 ( .A(n_xor_module_197_res), .B(
        n_xor_module_195_res), .Z(n_xor_module_205_res) );
  XOR2_X1 u_xor_module_206_U1 ( .A(n_xor_module_198_res), .B(
        n_xor_module_196_res), .Z(n_xor_module_206_res) );
  XOR2_X1 u_xor_module_207_U1 ( .A(n_xor_module_199_res), .B(
        n_xor_module_201_res), .Z(n_xor_module_207_res) );
  XOR2_X1 u_xor_module_208_U1 ( .A(n_xor_module_200_res), .B(
        n_xor_module_202_res), .Z(n_xor_module_208_res) );
  DFF_X1 u_reg_module_177__hpc_r0_reg ( .D(p_rand_16), .CK(clock_0), .Q(
        n_reg_module_177_res), .QN() );
  INV_X1 u_not_module_33_U1 ( .A(n_xor_module_205_res), .ZN(
        n_not_module_33_res) );
  AND2_X1 u_and_module_97_U1 ( .A1(n_not_module_33_res), .A2(
        n_reg_module_177_res), .ZN(n_and_module_97_res) );
  XOR2_X1 u_xor_module_209_U1 ( .A(p_rand_16), .B(n_xor_module_12_res), .Z(
        n_xor_module_209_res) );
  INV_X1 u_not_module_34_U1 ( .A(n_xor_module_206_res), .ZN(
        n_not_module_34_res) );
  AND2_X1 u_and_module_98_U1 ( .A1(n_not_module_34_res), .A2(
        n_reg_module_177_res), .ZN(n_and_module_98_res) );
  XOR2_X1 u_xor_module_210_U1 ( .A(p_rand_16), .B(n_xor_module_11_res), .Z(
        n_xor_module_210_res) );
  DFF_X1 u_reg_module_178__hpc_r0_reg ( .D(n_xor_module_11_res), .CK(clock_0), 
        .Q(n_reg_module_178_res), .QN() );
  AND2_X1 u_and_module_99_U1 ( .A1(n_reg_module_178_res), .A2(
        n_xor_module_205_res), .ZN(n_and_module_99_res) );
  DFF_X1 u_reg_module_179__hpc_r0_reg ( .D(n_and_module_99_res), .CK(clock_0), 
        .Q(n_reg_module_179_res), .QN() );
  DFF_X1 u_reg_module_180__hpc_r0_reg ( .D(n_xor_module_209_res), .CK(clock_0), 
        .Q(n_reg_module_180_res), .QN() );
  AND2_X1 u_and_module_100_U1 ( .A1(n_reg_module_180_res), .A2(
        n_xor_module_205_res), .ZN(n_and_module_100_res) );
  DFF_X1 u_reg_module_181__hpc_r0_reg ( .D(n_and_module_100_res), .CK(clock_0), 
        .Q(n_reg_module_181_res), .QN() );
  DFF_X1 u_reg_module_182__hpc_r0_reg ( .D(n_and_module_97_res), .CK(clock_0), 
        .Q(n_reg_module_182_res), .QN() );
  XOR2_X1 u_xor_module_211_U1 ( .A(n_reg_module_182_res), .B(
        n_reg_module_181_res), .Z(n_xor_module_211_res) );
  XOR2_X1 u_xor_module_212_U1 ( .A(n_xor_module_211_res), .B(
        n_reg_module_179_res), .Z(n_xor_module_212_res) );
  DFF_X1 u_reg_module_183__hpc_r0_reg ( .D(n_xor_module_12_res), .CK(clock_0), 
        .Q(n_reg_module_183_res), .QN() );
  AND2_X1 u_and_module_101_U1 ( .A1(n_reg_module_183_res), .A2(
        n_xor_module_206_res), .ZN(n_and_module_101_res) );
  DFF_X1 u_reg_module_184__hpc_r0_reg ( .D(n_and_module_101_res), .CK(clock_0), 
        .Q(n_reg_module_184_res), .QN() );
  DFF_X1 u_reg_module_185__hpc_r0_reg ( .D(n_xor_module_210_res), .CK(clock_0), 
        .Q(n_reg_module_185_res), .QN() );
  AND2_X1 u_and_module_102_U1 ( .A1(n_reg_module_185_res), .A2(
        n_xor_module_206_res), .ZN(n_and_module_102_res) );
  DFF_X1 u_reg_module_186__hpc_r0_reg ( .D(n_and_module_102_res), .CK(clock_0), 
        .Q(n_reg_module_186_res), .QN() );
  DFF_X1 u_reg_module_187__hpc_r0_reg ( .D(n_and_module_98_res), .CK(clock_0), 
        .Q(n_reg_module_187_res), .QN() );
  XOR2_X1 u_xor_module_213_U1 ( .A(n_reg_module_187_res), .B(
        n_reg_module_186_res), .Z(n_xor_module_213_res) );
  XOR2_X1 u_xor_module_214_U1 ( .A(n_xor_module_213_res), .B(
        n_reg_module_184_res), .Z(n_xor_module_214_res) );
  DFF_X1 u_reg_module_188__hpc_r0_reg ( .D(p_rand_17), .CK(clock_0), .Q(
        n_reg_module_188_res), .QN() );
  INV_X1 u_not_module_35_U1 ( .A(n_xor_module_197_res), .ZN(
        n_not_module_35_res) );
  AND2_X1 u_and_module_103_U1 ( .A1(n_not_module_35_res), .A2(
        n_reg_module_188_res), .ZN(n_and_module_103_res) );
  XOR2_X1 u_xor_module_215_U1 ( .A(p_rand_17), .B(n_xor_module_16_res), .Z(
        n_xor_module_215_res) );
  INV_X1 u_not_module_36_U1 ( .A(n_xor_module_198_res), .ZN(
        n_not_module_36_res) );
  AND2_X1 u_and_module_104_U1 ( .A1(n_not_module_36_res), .A2(
        n_reg_module_188_res), .ZN(n_and_module_104_res) );
  XOR2_X1 u_xor_module_216_U1 ( .A(p_rand_17), .B(n_xor_module_15_res), .Z(
        n_xor_module_216_res) );
  DFF_X1 u_reg_module_189__hpc_r0_reg ( .D(n_xor_module_15_res), .CK(clock_0), 
        .Q(n_reg_module_189_res), .QN() );
  AND2_X1 u_and_module_105_U1 ( .A1(n_reg_module_189_res), .A2(
        n_xor_module_197_res), .ZN(n_and_module_105_res) );
  DFF_X1 u_reg_module_190__hpc_r0_reg ( .D(n_and_module_105_res), .CK(clock_0), 
        .Q(n_reg_module_190_res), .QN() );
  DFF_X1 u_reg_module_191__hpc_r0_reg ( .D(n_xor_module_215_res), .CK(clock_0), 
        .Q(n_reg_module_191_res), .QN() );
  AND2_X1 u_and_module_106_U1 ( .A1(n_reg_module_191_res), .A2(
        n_xor_module_197_res), .ZN(n_and_module_106_res) );
  DFF_X1 u_reg_module_192__hpc_r0_reg ( .D(n_and_module_106_res), .CK(clock_0), 
        .Q(n_reg_module_192_res), .QN() );
  DFF_X1 u_reg_module_193__hpc_r0_reg ( .D(n_and_module_103_res), .CK(clock_0), 
        .Q(n_reg_module_193_res), .QN() );
  XOR2_X1 u_xor_module_217_U1 ( .A(n_reg_module_193_res), .B(
        n_reg_module_192_res), .Z(n_xor_module_217_res) );
  XOR2_X1 u_xor_module_218_U1 ( .A(n_xor_module_217_res), .B(
        n_reg_module_190_res), .Z(n_xor_module_218_res) );
  DFF_X1 u_reg_module_194__hpc_r0_reg ( .D(n_xor_module_16_res), .CK(clock_0), 
        .Q(n_reg_module_194_res), .QN() );
  AND2_X1 u_and_module_107_U1 ( .A1(n_reg_module_194_res), .A2(
        n_xor_module_198_res), .ZN(n_and_module_107_res) );
  DFF_X1 u_reg_module_195__hpc_r0_reg ( .D(n_and_module_107_res), .CK(clock_0), 
        .Q(n_reg_module_195_res), .QN() );
  DFF_X1 u_reg_module_196__hpc_r0_reg ( .D(n_xor_module_216_res), .CK(clock_0), 
        .Q(n_reg_module_196_res), .QN() );
  AND2_X1 u_and_module_108_U1 ( .A1(n_reg_module_196_res), .A2(
        n_xor_module_198_res), .ZN(n_and_module_108_res) );
  DFF_X1 u_reg_module_197__hpc_r0_reg ( .D(n_and_module_108_res), .CK(clock_0), 
        .Q(n_reg_module_197_res), .QN() );
  DFF_X1 u_reg_module_198__hpc_r0_reg ( .D(n_and_module_104_res), .CK(clock_0), 
        .Q(n_reg_module_198_res), .QN() );
  XOR2_X1 u_xor_module_219_U1 ( .A(n_reg_module_198_res), .B(
        n_reg_module_197_res), .Z(n_xor_module_219_res) );
  XOR2_X1 u_xor_module_220_U1 ( .A(n_xor_module_219_res), .B(
        n_reg_module_195_res), .Z(n_xor_module_220_res) );
  DFF_X1 u_reg_module_199__hpc_r0_reg ( .D(p_rand_18), .CK(clock_0), .Q(
        n_reg_module_199_res), .QN() );
  INV_X1 u_not_module_37_U1 ( .A(n_xor_module_195_res), .ZN(
        n_not_module_37_res) );
  AND2_X1 u_and_module_109_U1 ( .A1(n_not_module_37_res), .A2(
        n_reg_module_199_res), .ZN(n_and_module_109_res) );
  XOR2_X1 u_xor_module_221_U1 ( .A(p_rand_18), .B(io_i7_s1), .Z(
        n_xor_module_221_res) );
  INV_X1 u_not_module_38_U1 ( .A(n_xor_module_196_res), .ZN(
        n_not_module_38_res) );
  AND2_X1 u_and_module_110_U1 ( .A1(n_not_module_38_res), .A2(
        n_reg_module_199_res), .ZN(n_and_module_110_res) );
  XOR2_X1 u_xor_module_222_U1 ( .A(p_rand_18), .B(io_i7_s0), .Z(
        n_xor_module_222_res) );
  DFF_X1 u_reg_module_200__hpc_r0_reg ( .D(io_i7_s0), .CK(clock_0), .Q(
        n_reg_module_200_res), .QN() );
  AND2_X1 u_and_module_111_U1 ( .A1(n_reg_module_200_res), .A2(
        n_xor_module_195_res), .ZN(n_and_module_111_res) );
  DFF_X1 u_reg_module_201__hpc_r0_reg ( .D(n_and_module_111_res), .CK(clock_0), 
        .Q(n_reg_module_201_res), .QN() );
  DFF_X1 u_reg_module_202__hpc_r0_reg ( .D(n_xor_module_221_res), .CK(clock_0), 
        .Q(n_reg_module_202_res), .QN() );
  AND2_X1 u_and_module_112_U1 ( .A1(n_reg_module_202_res), .A2(
        n_xor_module_195_res), .ZN(n_and_module_112_res) );
  DFF_X1 u_reg_module_203__hpc_r0_reg ( .D(n_and_module_112_res), .CK(clock_0), 
        .Q(n_reg_module_203_res), .QN() );
  DFF_X1 u_reg_module_204__hpc_r0_reg ( .D(n_and_module_109_res), .CK(clock_0), 
        .Q(n_reg_module_204_res), .QN() );
  XOR2_X1 u_xor_module_223_U1 ( .A(n_reg_module_204_res), .B(
        n_reg_module_203_res), .Z(n_xor_module_223_res) );
  XOR2_X1 u_xor_module_224_U1 ( .A(n_xor_module_223_res), .B(
        n_reg_module_201_res), .Z(n_xor_module_224_res) );
  DFF_X1 u_reg_module_205__hpc_r0_reg ( .D(io_i7_s1), .CK(clock_0), .Q(
        n_reg_module_205_res), .QN() );
  AND2_X1 u_and_module_113_U1 ( .A1(n_reg_module_205_res), .A2(
        n_xor_module_196_res), .ZN(n_and_module_113_res) );
  DFF_X1 u_reg_module_206__hpc_r0_reg ( .D(n_and_module_113_res), .CK(clock_0), 
        .Q(n_reg_module_206_res), .QN() );
  DFF_X1 u_reg_module_207__hpc_r0_reg ( .D(n_xor_module_222_res), .CK(clock_0), 
        .Q(n_reg_module_207_res), .QN() );
  AND2_X1 u_and_module_114_U1 ( .A1(n_reg_module_207_res), .A2(
        n_xor_module_196_res), .ZN(n_and_module_114_res) );
  DFF_X1 u_reg_module_208__hpc_r0_reg ( .D(n_and_module_114_res), .CK(clock_0), 
        .Q(n_reg_module_208_res), .QN() );
  DFF_X1 u_reg_module_209__hpc_r0_reg ( .D(n_and_module_110_res), .CK(clock_0), 
        .Q(n_reg_module_209_res), .QN() );
  XOR2_X1 u_xor_module_225_U1 ( .A(n_reg_module_209_res), .B(
        n_reg_module_208_res), .Z(n_xor_module_225_res) );
  XOR2_X1 u_xor_module_226_U1 ( .A(n_xor_module_225_res), .B(
        n_reg_module_206_res), .Z(n_xor_module_226_res) );
  DFF_X1 u_reg_module_210__hpc_r0_reg ( .D(p_rand_19), .CK(clock_0), .Q(
        n_reg_module_210_res), .QN() );
  INV_X1 u_not_module_39_U1 ( .A(n_xor_module_203_res), .ZN(
        n_not_module_39_res) );
  AND2_X1 u_and_module_115_U1 ( .A1(n_not_module_39_res), .A2(
        n_reg_module_210_res), .ZN(n_and_module_115_res) );
  XOR2_X1 u_xor_module_227_U1 ( .A(p_rand_19), .B(n_xor_module_32_res), .Z(
        n_xor_module_227_res) );
  INV_X1 u_not_module_40_U1 ( .A(n_xor_module_204_res), .ZN(
        n_not_module_40_res) );
  AND2_X1 u_and_module_116_U1 ( .A1(n_not_module_40_res), .A2(
        n_reg_module_210_res), .ZN(n_and_module_116_res) );
  XOR2_X1 u_xor_module_228_U1 ( .A(p_rand_19), .B(n_xor_module_31_res), .Z(
        n_xor_module_228_res) );
  DFF_X1 u_reg_module_211__hpc_r0_reg ( .D(n_xor_module_31_res), .CK(clock_0), 
        .Q(n_reg_module_211_res), .QN() );
  AND2_X1 u_and_module_117_U1 ( .A1(n_reg_module_211_res), .A2(
        n_xor_module_203_res), .ZN(n_and_module_117_res) );
  DFF_X1 u_reg_module_212__hpc_r0_reg ( .D(n_and_module_117_res), .CK(clock_0), 
        .Q(n_reg_module_212_res), .QN() );
  DFF_X1 u_reg_module_213__hpc_r0_reg ( .D(n_xor_module_227_res), .CK(clock_0), 
        .Q(n_reg_module_213_res), .QN() );
  AND2_X1 u_and_module_118_U1 ( .A1(n_reg_module_213_res), .A2(
        n_xor_module_203_res), .ZN(n_and_module_118_res) );
  DFF_X1 u_reg_module_214__hpc_r0_reg ( .D(n_and_module_118_res), .CK(clock_0), 
        .Q(n_reg_module_214_res), .QN() );
  DFF_X1 u_reg_module_215__hpc_r0_reg ( .D(n_and_module_115_res), .CK(clock_0), 
        .Q(n_reg_module_215_res), .QN() );
  XOR2_X1 u_xor_module_229_U1 ( .A(n_reg_module_215_res), .B(
        n_reg_module_214_res), .Z(n_xor_module_229_res) );
  XOR2_X1 u_xor_module_230_U1 ( .A(n_xor_module_229_res), .B(
        n_reg_module_212_res), .Z(n_xor_module_230_res) );
  DFF_X1 u_reg_module_216__hpc_r0_reg ( .D(n_xor_module_32_res), .CK(clock_0), 
        .Q(n_reg_module_216_res), .QN() );
  AND2_X1 u_and_module_119_U1 ( .A1(n_reg_module_216_res), .A2(
        n_xor_module_204_res), .ZN(n_and_module_119_res) );
  DFF_X1 u_reg_module_217__hpc_r0_reg ( .D(n_and_module_119_res), .CK(clock_0), 
        .Q(n_reg_module_217_res), .QN() );
  DFF_X1 u_reg_module_218__hpc_r0_reg ( .D(n_xor_module_228_res), .CK(clock_0), 
        .Q(n_reg_module_218_res), .QN() );
  AND2_X1 u_and_module_120_U1 ( .A1(n_reg_module_218_res), .A2(
        n_xor_module_204_res), .ZN(n_and_module_120_res) );
  DFF_X1 u_reg_module_219__hpc_r0_reg ( .D(n_and_module_120_res), .CK(clock_0), 
        .Q(n_reg_module_219_res), .QN() );
  DFF_X1 u_reg_module_220__hpc_r0_reg ( .D(n_and_module_116_res), .CK(clock_0), 
        .Q(n_reg_module_220_res), .QN() );
  XOR2_X1 u_xor_module_231_U1 ( .A(n_reg_module_220_res), .B(
        n_reg_module_219_res), .Z(n_xor_module_231_res) );
  XOR2_X1 u_xor_module_232_U1 ( .A(n_xor_module_231_res), .B(
        n_reg_module_217_res), .Z(n_xor_module_232_res) );
  DFF_X1 u_reg_module_221__hpc_r0_reg ( .D(p_rand_20), .CK(clock_0), .Q(
        n_reg_module_221_res), .QN() );
  INV_X1 u_not_module_41_U1 ( .A(n_xor_module_193_res), .ZN(
        n_not_module_41_res) );
  AND2_X1 u_and_module_121_U1 ( .A1(n_not_module_41_res), .A2(
        n_reg_module_221_res), .ZN(n_and_module_121_res) );
  XOR2_X1 u_xor_module_233_U1 ( .A(p_rand_20), .B(n_xor_module_18_res), .Z(
        n_xor_module_233_res) );
  INV_X1 u_not_module_42_U1 ( .A(n_xor_module_194_res), .ZN(
        n_not_module_42_res) );
  AND2_X1 u_and_module_122_U1 ( .A1(n_not_module_42_res), .A2(
        n_reg_module_221_res), .ZN(n_and_module_122_res) );
  XOR2_X1 u_xor_module_234_U1 ( .A(p_rand_20), .B(n_xor_module_17_res), .Z(
        n_xor_module_234_res) );
  DFF_X1 u_reg_module_222__hpc_r0_reg ( .D(n_xor_module_17_res), .CK(clock_0), 
        .Q(n_reg_module_222_res), .QN() );
  AND2_X1 u_and_module_123_U1 ( .A1(n_reg_module_222_res), .A2(
        n_xor_module_193_res), .ZN(n_and_module_123_res) );
  DFF_X1 u_reg_module_223__hpc_r0_reg ( .D(n_and_module_123_res), .CK(clock_0), 
        .Q(n_reg_module_223_res), .QN() );
  DFF_X1 u_reg_module_224__hpc_r0_reg ( .D(n_xor_module_233_res), .CK(clock_0), 
        .Q(n_reg_module_224_res), .QN() );
  AND2_X1 u_and_module_124_U1 ( .A1(n_reg_module_224_res), .A2(
        n_xor_module_193_res), .ZN(n_and_module_124_res) );
  DFF_X1 u_reg_module_225__hpc_r0_reg ( .D(n_and_module_124_res), .CK(clock_0), 
        .Q(n_reg_module_225_res), .QN() );
  DFF_X1 u_reg_module_226__hpc_r0_reg ( .D(n_and_module_121_res), .CK(clock_0), 
        .Q(n_reg_module_226_res), .QN() );
  XOR2_X1 u_xor_module_235_U1 ( .A(n_reg_module_226_res), .B(
        n_reg_module_225_res), .Z(n_xor_module_235_res) );
  XOR2_X1 u_xor_module_236_U1 ( .A(n_xor_module_235_res), .B(
        n_reg_module_223_res), .Z(n_xor_module_236_res) );
  DFF_X1 u_reg_module_227__hpc_r0_reg ( .D(n_xor_module_18_res), .CK(clock_0), 
        .Q(n_reg_module_227_res), .QN() );
  AND2_X1 u_and_module_125_U1 ( .A1(n_reg_module_227_res), .A2(
        n_xor_module_194_res), .ZN(n_and_module_125_res) );
  DFF_X1 u_reg_module_228__hpc_r0_reg ( .D(n_and_module_125_res), .CK(clock_0), 
        .Q(n_reg_module_228_res), .QN() );
  DFF_X1 u_reg_module_229__hpc_r0_reg ( .D(n_xor_module_234_res), .CK(clock_0), 
        .Q(n_reg_module_229_res), .QN() );
  AND2_X1 u_and_module_126_U1 ( .A1(n_reg_module_229_res), .A2(
        n_xor_module_194_res), .ZN(n_and_module_126_res) );
  DFF_X1 u_reg_module_230__hpc_r0_reg ( .D(n_and_module_126_res), .CK(clock_0), 
        .Q(n_reg_module_230_res), .QN() );
  DFF_X1 u_reg_module_231__hpc_r0_reg ( .D(n_and_module_122_res), .CK(clock_0), 
        .Q(n_reg_module_231_res), .QN() );
  XOR2_X1 u_xor_module_237_U1 ( .A(n_reg_module_231_res), .B(
        n_reg_module_230_res), .Z(n_xor_module_237_res) );
  XOR2_X1 u_xor_module_238_U1 ( .A(n_xor_module_237_res), .B(
        n_reg_module_228_res), .Z(n_xor_module_238_res) );
  DFF_X1 u_reg_module_232__hpc_r0_reg ( .D(p_rand_21), .CK(clock_0), .Q(
        n_reg_module_232_res), .QN() );
  INV_X1 u_not_module_43_U1 ( .A(n_xor_module_191_res), .ZN(
        n_not_module_43_res) );
  AND2_X1 u_and_module_127_U1 ( .A1(n_not_module_43_res), .A2(
        n_reg_module_232_res), .ZN(n_and_module_127_res) );
  XOR2_X1 u_xor_module_239_U1 ( .A(p_rand_21), .B(n_xor_module_34_res), .Z(
        n_xor_module_239_res) );
  INV_X1 u_not_module_44_U1 ( .A(n_xor_module_192_res), .ZN(
        n_not_module_44_res) );
  AND2_X1 u_and_module_128_U1 ( .A1(n_not_module_44_res), .A2(
        n_reg_module_232_res), .ZN(n_and_module_128_res) );
  XOR2_X1 u_xor_module_240_U1 ( .A(p_rand_21), .B(n_xor_module_33_res), .Z(
        n_xor_module_240_res) );
  DFF_X1 u_reg_module_233__hpc_r0_reg ( .D(n_xor_module_33_res), .CK(clock_0), 
        .Q(n_reg_module_233_res), .QN() );
  AND2_X1 u_and_module_129_U1 ( .A1(n_reg_module_233_res), .A2(
        n_xor_module_191_res), .ZN(n_and_module_129_res) );
  DFF_X1 u_reg_module_234__hpc_r0_reg ( .D(n_and_module_129_res), .CK(clock_0), 
        .Q(n_reg_module_234_res), .QN() );
  DFF_X1 u_reg_module_235__hpc_r0_reg ( .D(n_xor_module_239_res), .CK(clock_0), 
        .Q(n_reg_module_235_res), .QN() );
  AND2_X1 u_and_module_130_U1 ( .A1(n_reg_module_235_res), .A2(
        n_xor_module_191_res), .ZN(n_and_module_130_res) );
  DFF_X1 u_reg_module_236__hpc_r0_reg ( .D(n_and_module_130_res), .CK(clock_0), 
        .Q(n_reg_module_236_res), .QN() );
  DFF_X1 u_reg_module_237__hpc_r0_reg ( .D(n_and_module_127_res), .CK(clock_0), 
        .Q(n_reg_module_237_res), .QN() );
  XOR2_X1 u_xor_module_241_U1 ( .A(n_reg_module_237_res), .B(
        n_reg_module_236_res), .Z(n_xor_module_241_res) );
  XOR2_X1 u_xor_module_242_U1 ( .A(n_xor_module_241_res), .B(
        n_reg_module_234_res), .Z(n_xor_module_242_res) );
  DFF_X1 u_reg_module_238__hpc_r0_reg ( .D(n_xor_module_34_res), .CK(clock_0), 
        .Q(n_reg_module_238_res), .QN() );
  AND2_X1 u_and_module_131_U1 ( .A1(n_reg_module_238_res), .A2(
        n_xor_module_192_res), .ZN(n_and_module_131_res) );
  DFF_X1 u_reg_module_239__hpc_r0_reg ( .D(n_and_module_131_res), .CK(clock_0), 
        .Q(n_reg_module_239_res), .QN() );
  DFF_X1 u_reg_module_240__hpc_r0_reg ( .D(n_xor_module_240_res), .CK(clock_0), 
        .Q(n_reg_module_240_res), .QN() );
  AND2_X1 u_and_module_132_U1 ( .A1(n_reg_module_240_res), .A2(
        n_xor_module_192_res), .ZN(n_and_module_132_res) );
  DFF_X1 u_reg_module_241__hpc_r0_reg ( .D(n_and_module_132_res), .CK(clock_0), 
        .Q(n_reg_module_241_res), .QN() );
  DFF_X1 u_reg_module_242__hpc_r0_reg ( .D(n_and_module_128_res), .CK(clock_0), 
        .Q(n_reg_module_242_res), .QN() );
  XOR2_X1 u_xor_module_243_U1 ( .A(n_reg_module_242_res), .B(
        n_reg_module_241_res), .Z(n_xor_module_243_res) );
  XOR2_X1 u_xor_module_244_U1 ( .A(n_xor_module_243_res), .B(
        n_reg_module_239_res), .Z(n_xor_module_244_res) );
  DFF_X1 u_reg_module_243__hpc_r0_reg ( .D(p_rand_22), .CK(clock_0), .Q(
        n_reg_module_243_res), .QN() );
  INV_X1 u_not_module_45_U1 ( .A(n_xor_module_201_res), .ZN(
        n_not_module_45_res) );
  AND2_X1 u_and_module_133_U1 ( .A1(n_not_module_45_res), .A2(
        n_reg_module_243_res), .ZN(n_and_module_133_res) );
  XOR2_X1 u_xor_module_245_U1 ( .A(p_rand_22), .B(n_xor_module_30_res), .Z(
        n_xor_module_245_res) );
  INV_X1 u_not_module_46_U1 ( .A(n_xor_module_202_res), .ZN(
        n_not_module_46_res) );
  AND2_X1 u_and_module_134_U1 ( .A1(n_not_module_46_res), .A2(
        n_reg_module_243_res), .ZN(n_and_module_134_res) );
  XOR2_X1 u_xor_module_246_U1 ( .A(p_rand_22), .B(n_xor_module_29_res), .Z(
        n_xor_module_246_res) );
  DFF_X1 u_reg_module_244__hpc_r0_reg ( .D(n_xor_module_29_res), .CK(clock_0), 
        .Q(n_reg_module_244_res), .QN() );
  AND2_X1 u_and_module_135_U1 ( .A1(n_reg_module_244_res), .A2(
        n_xor_module_201_res), .ZN(n_and_module_135_res) );
  DFF_X1 u_reg_module_245__hpc_r0_reg ( .D(n_and_module_135_res), .CK(clock_0), 
        .Q(n_reg_module_245_res), .QN() );
  DFF_X1 u_reg_module_246__hpc_r0_reg ( .D(n_xor_module_245_res), .CK(clock_0), 
        .Q(n_reg_module_246_res), .QN() );
  AND2_X1 u_and_module_136_U1 ( .A1(n_reg_module_246_res), .A2(
        n_xor_module_201_res), .ZN(n_and_module_136_res) );
  DFF_X1 u_reg_module_247__hpc_r0_reg ( .D(n_and_module_136_res), .CK(clock_0), 
        .Q(n_reg_module_247_res), .QN() );
  DFF_X1 u_reg_module_248__hpc_r0_reg ( .D(n_and_module_133_res), .CK(clock_0), 
        .Q(n_reg_module_248_res), .QN() );
  XOR2_X1 u_xor_module_247_U1 ( .A(n_reg_module_248_res), .B(
        n_reg_module_247_res), .Z(n_xor_module_247_res) );
  XOR2_X1 u_xor_module_248_U1 ( .A(n_xor_module_247_res), .B(
        n_reg_module_245_res), .Z(n_xor_module_248_res) );
  DFF_X1 u_reg_module_249__hpc_r0_reg ( .D(n_xor_module_30_res), .CK(clock_0), 
        .Q(n_reg_module_249_res), .QN() );
  AND2_X1 u_and_module_137_U1 ( .A1(n_reg_module_249_res), .A2(
        n_xor_module_202_res), .ZN(n_and_module_137_res) );
  DFF_X1 u_reg_module_250__hpc_r0_reg ( .D(n_and_module_137_res), .CK(clock_0), 
        .Q(n_reg_module_250_res), .QN() );
  DFF_X1 u_reg_module_251__hpc_r0_reg ( .D(n_xor_module_246_res), .CK(clock_0), 
        .Q(n_reg_module_251_res), .QN() );
  AND2_X1 u_and_module_138_U1 ( .A1(n_reg_module_251_res), .A2(
        n_xor_module_202_res), .ZN(n_and_module_138_res) );
  DFF_X1 u_reg_module_252__hpc_r0_reg ( .D(n_and_module_138_res), .CK(clock_0), 
        .Q(n_reg_module_252_res), .QN() );
  DFF_X1 u_reg_module_253__hpc_r0_reg ( .D(n_and_module_134_res), .CK(clock_0), 
        .Q(n_reg_module_253_res), .QN() );
  XOR2_X1 u_xor_module_249_U1 ( .A(n_reg_module_253_res), .B(
        n_reg_module_252_res), .Z(n_xor_module_249_res) );
  XOR2_X1 u_xor_module_250_U1 ( .A(n_xor_module_249_res), .B(
        n_reg_module_250_res), .Z(n_xor_module_250_res) );
  DFF_X1 u_reg_module_254__hpc_r0_reg ( .D(p_rand_23), .CK(clock_0), .Q(
        n_reg_module_254_res), .QN() );
  INV_X1 u_not_module_47_U1 ( .A(n_xor_module_207_res), .ZN(
        n_not_module_47_res) );
  AND2_X1 u_and_module_139_U1 ( .A1(n_not_module_47_res), .A2(
        n_reg_module_254_res), .ZN(n_and_module_139_res) );
  XOR2_X1 u_xor_module_251_U1 ( .A(p_rand_23), .B(n_xor_module_54_res), .Z(
        n_xor_module_251_res) );
  INV_X1 u_not_module_48_U1 ( .A(n_xor_module_208_res), .ZN(
        n_not_module_48_res) );
  AND2_X1 u_and_module_140_U1 ( .A1(n_not_module_48_res), .A2(
        n_reg_module_254_res), .ZN(n_and_module_140_res) );
  XOR2_X1 u_xor_module_252_U1 ( .A(p_rand_23), .B(n_xor_module_53_res), .Z(
        n_xor_module_252_res) );
  DFF_X1 u_reg_module_255__hpc_r0_reg ( .D(n_xor_module_53_res), .CK(clock_0), 
        .Q(n_reg_module_255_res), .QN() );
  AND2_X1 u_and_module_141_U1 ( .A1(n_reg_module_255_res), .A2(
        n_xor_module_207_res), .ZN(n_and_module_141_res) );
  DFF_X1 u_reg_module_256__hpc_r0_reg ( .D(n_and_module_141_res), .CK(clock_0), 
        .Q(n_reg_module_256_res), .QN() );
  DFF_X1 u_reg_module_257__hpc_r0_reg ( .D(n_xor_module_251_res), .CK(clock_0), 
        .Q(n_reg_module_257_res), .QN() );
  AND2_X1 u_and_module_142_U1 ( .A1(n_reg_module_257_res), .A2(
        n_xor_module_207_res), .ZN(n_and_module_142_res) );
  DFF_X1 u_reg_module_258__hpc_r0_reg ( .D(n_and_module_142_res), .CK(clock_0), 
        .Q(n_reg_module_258_res), .QN() );
  DFF_X1 u_reg_module_259__hpc_r0_reg ( .D(n_and_module_139_res), .CK(clock_0), 
        .Q(n_reg_module_259_res), .QN() );
  XOR2_X1 u_xor_module_253_U1 ( .A(n_reg_module_259_res), .B(
        n_reg_module_258_res), .Z(n_xor_module_253_res) );
  XOR2_X1 u_xor_module_254_U1 ( .A(n_xor_module_253_res), .B(
        n_reg_module_256_res), .Z(n_xor_module_254_res) );
  DFF_X1 u_reg_module_260__hpc_r0_reg ( .D(n_xor_module_54_res), .CK(clock_0), 
        .Q(n_reg_module_260_res), .QN() );
  AND2_X1 u_and_module_143_U1 ( .A1(n_reg_module_260_res), .A2(
        n_xor_module_208_res), .ZN(n_and_module_143_res) );
  DFF_X1 u_reg_module_261__hpc_r0_reg ( .D(n_and_module_143_res), .CK(clock_0), 
        .Q(n_reg_module_261_res), .QN() );
  DFF_X1 u_reg_module_262__hpc_r0_reg ( .D(n_xor_module_252_res), .CK(clock_0), 
        .Q(n_reg_module_262_res), .QN() );
  AND2_X1 u_and_module_144_U1 ( .A1(n_reg_module_262_res), .A2(
        n_xor_module_208_res), .ZN(n_and_module_144_res) );
  DFF_X1 u_reg_module_263__hpc_r0_reg ( .D(n_and_module_144_res), .CK(clock_0), 
        .Q(n_reg_module_263_res), .QN() );
  DFF_X1 u_reg_module_264__hpc_r0_reg ( .D(n_and_module_140_res), .CK(clock_0), 
        .Q(n_reg_module_264_res), .QN() );
  XOR2_X1 u_xor_module_255_U1 ( .A(n_reg_module_264_res), .B(
        n_reg_module_263_res), .Z(n_xor_module_255_res) );
  XOR2_X1 u_xor_module_256_U1 ( .A(n_xor_module_255_res), .B(
        n_reg_module_261_res), .Z(n_xor_module_256_res) );
  DFF_X1 u_reg_module_265__hpc_r0_reg ( .D(p_rand_24), .CK(clock_0), .Q(
        n_reg_module_265_res), .QN() );
  INV_X1 u_not_module_49_U1 ( .A(n_xor_module_199_res), .ZN(
        n_not_module_49_res) );
  AND2_X1 u_and_module_145_U1 ( .A1(n_not_module_49_res), .A2(
        n_reg_module_265_res), .ZN(n_and_module_145_res) );
  XOR2_X1 u_xor_module_257_U1 ( .A(p_rand_24), .B(n_xor_module_20_res), .Z(
        n_xor_module_257_res) );
  INV_X1 u_not_module_50_U1 ( .A(n_xor_module_200_res), .ZN(
        n_not_module_50_res) );
  AND2_X1 u_and_module_146_U1 ( .A1(n_not_module_50_res), .A2(
        n_reg_module_265_res), .ZN(n_and_module_146_res) );
  XOR2_X1 u_xor_module_258_U1 ( .A(p_rand_24), .B(n_xor_module_19_res), .Z(
        n_xor_module_258_res) );
  DFF_X1 u_reg_module_266__hpc_r0_reg ( .D(n_xor_module_19_res), .CK(clock_0), 
        .Q(n_reg_module_266_res), .QN() );
  AND2_X1 u_and_module_147_U1 ( .A1(n_reg_module_266_res), .A2(
        n_xor_module_199_res), .ZN(n_and_module_147_res) );
  DFF_X1 u_reg_module_267__hpc_r0_reg ( .D(n_and_module_147_res), .CK(clock_0), 
        .Q(n_reg_module_267_res), .QN() );
  DFF_X1 u_reg_module_268__hpc_r0_reg ( .D(n_xor_module_257_res), .CK(clock_0), 
        .Q(n_reg_module_268_res), .QN() );
  AND2_X1 u_and_module_148_U1 ( .A1(n_reg_module_268_res), .A2(
        n_xor_module_199_res), .ZN(n_and_module_148_res) );
  DFF_X1 u_reg_module_269__hpc_r0_reg ( .D(n_and_module_148_res), .CK(clock_0), 
        .Q(n_reg_module_269_res), .QN() );
  DFF_X1 u_reg_module_270__hpc_r0_reg ( .D(n_and_module_145_res), .CK(clock_0), 
        .Q(n_reg_module_270_res), .QN() );
  XOR2_X1 u_xor_module_259_U1 ( .A(n_reg_module_270_res), .B(
        n_reg_module_269_res), .Z(n_xor_module_259_res) );
  XOR2_X1 u_xor_module_260_U1 ( .A(n_xor_module_259_res), .B(
        n_reg_module_267_res), .Z(n_xor_module_260_res) );
  DFF_X1 u_reg_module_271__hpc_r0_reg ( .D(n_xor_module_20_res), .CK(clock_0), 
        .Q(n_reg_module_271_res), .QN() );
  AND2_X1 u_and_module_149_U1 ( .A1(n_reg_module_271_res), .A2(
        n_xor_module_200_res), .ZN(n_and_module_149_res) );
  DFF_X1 u_reg_module_272__hpc_r0_reg ( .D(n_and_module_149_res), .CK(clock_0), 
        .Q(n_reg_module_272_res), .QN() );
  DFF_X1 u_reg_module_273__hpc_r0_reg ( .D(n_xor_module_258_res), .CK(clock_0), 
        .Q(n_reg_module_273_res), .QN() );
  AND2_X1 u_and_module_150_U1 ( .A1(n_reg_module_273_res), .A2(
        n_xor_module_200_res), .ZN(n_and_module_150_res) );
  DFF_X1 u_reg_module_274__hpc_r0_reg ( .D(n_and_module_150_res), .CK(clock_0), 
        .Q(n_reg_module_274_res), .QN() );
  DFF_X1 u_reg_module_275__hpc_r0_reg ( .D(n_and_module_146_res), .CK(clock_0), 
        .Q(n_reg_module_275_res), .QN() );
  XOR2_X1 u_xor_module_261_U1 ( .A(n_reg_module_275_res), .B(
        n_reg_module_274_res), .Z(n_xor_module_261_res) );
  XOR2_X1 u_xor_module_262_U1 ( .A(n_xor_module_261_res), .B(
        n_reg_module_272_res), .Z(n_xor_module_262_res) );
  DFF_X1 u_reg_module_276__hpc_r0_reg ( .D(p_rand_25), .CK(clock_0), .Q(
        n_reg_module_276_res), .QN() );
  INV_X1 u_not_module_51_U1 ( .A(n_xor_module_205_res), .ZN(
        n_not_module_51_res) );
  AND2_X1 u_and_module_151_U1 ( .A1(n_not_module_51_res), .A2(
        n_reg_module_276_res), .ZN(n_and_module_151_res) );
  XOR2_X1 u_xor_module_263_U1 ( .A(p_rand_25), .B(n_xor_module_26_res), .Z(
        n_xor_module_263_res) );
  INV_X1 u_not_module_52_U1 ( .A(n_xor_module_206_res), .ZN(
        n_not_module_52_res) );
  AND2_X1 u_and_module_152_U1 ( .A1(n_not_module_52_res), .A2(
        n_reg_module_276_res), .ZN(n_and_module_152_res) );
  XOR2_X1 u_xor_module_264_U1 ( .A(p_rand_25), .B(n_xor_module_25_res), .Z(
        n_xor_module_264_res) );
  DFF_X1 u_reg_module_277__hpc_r0_reg ( .D(n_xor_module_25_res), .CK(clock_0), 
        .Q(n_reg_module_277_res), .QN() );
  AND2_X1 u_and_module_153_U1 ( .A1(n_reg_module_277_res), .A2(
        n_xor_module_205_res), .ZN(n_and_module_153_res) );
  DFF_X1 u_reg_module_278__hpc_r0_reg ( .D(n_and_module_153_res), .CK(clock_0), 
        .Q(n_reg_module_278_res), .QN() );
  DFF_X1 u_reg_module_279__hpc_r0_reg ( .D(n_xor_module_263_res), .CK(clock_0), 
        .Q(n_reg_module_279_res), .QN() );
  AND2_X1 u_and_module_154_U1 ( .A1(n_reg_module_279_res), .A2(
        n_xor_module_205_res), .ZN(n_and_module_154_res) );
  DFF_X1 u_reg_module_280__hpc_r0_reg ( .D(n_and_module_154_res), .CK(clock_0), 
        .Q(n_reg_module_280_res), .QN() );
  DFF_X1 u_reg_module_281__hpc_r0_reg ( .D(n_and_module_151_res), .CK(clock_0), 
        .Q(n_reg_module_281_res), .QN() );
  XOR2_X1 u_xor_module_265_U1 ( .A(n_reg_module_281_res), .B(
        n_reg_module_280_res), .Z(n_xor_module_265_res) );
  XOR2_X1 u_xor_module_266_U1 ( .A(n_xor_module_265_res), .B(
        n_reg_module_278_res), .Z(n_xor_module_266_res) );
  DFF_X1 u_reg_module_282__hpc_r0_reg ( .D(n_xor_module_26_res), .CK(clock_0), 
        .Q(n_reg_module_282_res), .QN() );
  AND2_X1 u_and_module_155_U1 ( .A1(n_reg_module_282_res), .A2(
        n_xor_module_206_res), .ZN(n_and_module_155_res) );
  DFF_X1 u_reg_module_283__hpc_r0_reg ( .D(n_and_module_155_res), .CK(clock_0), 
        .Q(n_reg_module_283_res), .QN() );
  DFF_X1 u_reg_module_284__hpc_r0_reg ( .D(n_xor_module_264_res), .CK(clock_0), 
        .Q(n_reg_module_284_res), .QN() );
  AND2_X1 u_and_module_156_U1 ( .A1(n_reg_module_284_res), .A2(
        n_xor_module_206_res), .ZN(n_and_module_156_res) );
  DFF_X1 u_reg_module_285__hpc_r0_reg ( .D(n_and_module_156_res), .CK(clock_0), 
        .Q(n_reg_module_285_res), .QN() );
  DFF_X1 u_reg_module_286__hpc_r0_reg ( .D(n_and_module_152_res), .CK(clock_0), 
        .Q(n_reg_module_286_res), .QN() );
  XOR2_X1 u_xor_module_267_U1 ( .A(n_reg_module_286_res), .B(
        n_reg_module_285_res), .Z(n_xor_module_267_res) );
  XOR2_X1 u_xor_module_268_U1 ( .A(n_xor_module_267_res), .B(
        n_reg_module_283_res), .Z(n_xor_module_268_res) );
  DFF_X1 u_reg_module_287__hpc_r0_reg ( .D(p_rand_26), .CK(clock_0), .Q(
        n_reg_module_287_res), .QN() );
  INV_X1 u_not_module_53_U1 ( .A(n_xor_module_197_res), .ZN(
        n_not_module_53_res) );
  AND2_X1 u_and_module_157_U1 ( .A1(n_not_module_53_res), .A2(
        n_reg_module_287_res), .ZN(n_and_module_157_res) );
  XOR2_X1 u_xor_module_269_U1 ( .A(p_rand_26), .B(n_xor_module_46_res), .Z(
        n_xor_module_269_res) );
  INV_X1 u_not_module_54_U1 ( .A(n_xor_module_198_res), .ZN(
        n_not_module_54_res) );
  AND2_X1 u_and_module_158_U1 ( .A1(n_not_module_54_res), .A2(
        n_reg_module_287_res), .ZN(n_and_module_158_res) );
  XOR2_X1 u_xor_module_270_U1 ( .A(p_rand_26), .B(n_xor_module_45_res), .Z(
        n_xor_module_270_res) );
  DFF_X1 u_reg_module_288__hpc_r0_reg ( .D(n_xor_module_45_res), .CK(clock_0), 
        .Q(n_reg_module_288_res), .QN() );
  AND2_X1 u_and_module_159_U1 ( .A1(n_reg_module_288_res), .A2(
        n_xor_module_197_res), .ZN(n_and_module_159_res) );
  DFF_X1 u_reg_module_289__hpc_r0_reg ( .D(n_and_module_159_res), .CK(clock_0), 
        .Q(n_reg_module_289_res), .QN() );
  DFF_X1 u_reg_module_290__hpc_r0_reg ( .D(n_xor_module_269_res), .CK(clock_0), 
        .Q(n_reg_module_290_res), .QN() );
  AND2_X1 u_and_module_160_U1 ( .A1(n_reg_module_290_res), .A2(
        n_xor_module_197_res), .ZN(n_and_module_160_res) );
  DFF_X1 u_reg_module_291__hpc_r0_reg ( .D(n_and_module_160_res), .CK(clock_0), 
        .Q(n_reg_module_291_res), .QN() );
  DFF_X1 u_reg_module_292__hpc_r0_reg ( .D(n_and_module_157_res), .CK(clock_0), 
        .Q(n_reg_module_292_res), .QN() );
  XOR2_X1 u_xor_module_271_U1 ( .A(n_reg_module_292_res), .B(
        n_reg_module_291_res), .Z(n_xor_module_271_res) );
  XOR2_X1 u_xor_module_272_U1 ( .A(n_xor_module_271_res), .B(
        n_reg_module_289_res), .Z(n_xor_module_272_res) );
  DFF_X1 u_reg_module_293__hpc_r0_reg ( .D(n_xor_module_46_res), .CK(clock_0), 
        .Q(n_reg_module_293_res), .QN() );
  AND2_X1 u_and_module_161_U1 ( .A1(n_reg_module_293_res), .A2(
        n_xor_module_198_res), .ZN(n_and_module_161_res) );
  DFF_X1 u_reg_module_294__hpc_r0_reg ( .D(n_and_module_161_res), .CK(clock_0), 
        .Q(n_reg_module_294_res), .QN() );
  DFF_X1 u_reg_module_295__hpc_r0_reg ( .D(n_xor_module_270_res), .CK(clock_0), 
        .Q(n_reg_module_295_res), .QN() );
  AND2_X1 u_and_module_162_U1 ( .A1(n_reg_module_295_res), .A2(
        n_xor_module_198_res), .ZN(n_and_module_162_res) );
  DFF_X1 u_reg_module_296__hpc_r0_reg ( .D(n_and_module_162_res), .CK(clock_0), 
        .Q(n_reg_module_296_res), .QN() );
  DFF_X1 u_reg_module_297__hpc_r0_reg ( .D(n_and_module_158_res), .CK(clock_0), 
        .Q(n_reg_module_297_res), .QN() );
  XOR2_X1 u_xor_module_273_U1 ( .A(n_reg_module_297_res), .B(
        n_reg_module_296_res), .Z(n_xor_module_273_res) );
  XOR2_X1 u_xor_module_274_U1 ( .A(n_xor_module_273_res), .B(
        n_reg_module_294_res), .Z(n_xor_module_274_res) );
  DFF_X1 u_reg_module_298__hpc_r0_reg ( .D(p_rand_27), .CK(clock_0), .Q(
        n_reg_module_298_res), .QN() );
  INV_X1 u_not_module_55_U1 ( .A(n_xor_module_195_res), .ZN(
        n_not_module_55_res) );
  AND2_X1 u_and_module_163_U1 ( .A1(n_not_module_55_res), .A2(
        n_reg_module_298_res), .ZN(n_and_module_163_res) );
  XOR2_X1 u_xor_module_275_U1 ( .A(p_rand_27), .B(n_xor_module_38_res), .Z(
        n_xor_module_275_res) );
  INV_X1 u_not_module_56_U1 ( .A(n_xor_module_196_res), .ZN(
        n_not_module_56_res) );
  AND2_X1 u_and_module_164_U1 ( .A1(n_not_module_56_res), .A2(
        n_reg_module_298_res), .ZN(n_and_module_164_res) );
  XOR2_X1 u_xor_module_276_U1 ( .A(p_rand_27), .B(n_xor_module_37_res), .Z(
        n_xor_module_276_res) );
  DFF_X1 u_reg_module_299__hpc_r0_reg ( .D(n_xor_module_37_res), .CK(clock_0), 
        .Q(n_reg_module_299_res), .QN() );
  AND2_X1 u_and_module_165_U1 ( .A1(n_reg_module_299_res), .A2(
        n_xor_module_195_res), .ZN(n_and_module_165_res) );
  DFF_X1 u_reg_module_300__hpc_r0_reg ( .D(n_and_module_165_res), .CK(clock_0), 
        .Q(n_reg_module_300_res), .QN() );
  DFF_X1 u_reg_module_301__hpc_r0_reg ( .D(n_xor_module_275_res), .CK(clock_0), 
        .Q(n_reg_module_301_res), .QN() );
  AND2_X1 u_and_module_166_U1 ( .A1(n_reg_module_301_res), .A2(
        n_xor_module_195_res), .ZN(n_and_module_166_res) );
  DFF_X1 u_reg_module_302__hpc_r0_reg ( .D(n_and_module_166_res), .CK(clock_0), 
        .Q(n_reg_module_302_res), .QN() );
  DFF_X1 u_reg_module_303__hpc_r0_reg ( .D(n_and_module_163_res), .CK(clock_0), 
        .Q(n_reg_module_303_res), .QN() );
  XOR2_X1 u_xor_module_277_U1 ( .A(n_reg_module_303_res), .B(
        n_reg_module_302_res), .Z(n_xor_module_277_res) );
  XOR2_X1 u_xor_module_278_U1 ( .A(n_xor_module_277_res), .B(
        n_reg_module_300_res), .Z(n_xor_module_278_res) );
  DFF_X1 u_reg_module_304__hpc_r0_reg ( .D(n_xor_module_38_res), .CK(clock_0), 
        .Q(n_reg_module_304_res), .QN() );
  AND2_X1 u_and_module_167_U1 ( .A1(n_reg_module_304_res), .A2(
        n_xor_module_196_res), .ZN(n_and_module_167_res) );
  DFF_X1 u_reg_module_305__hpc_r0_reg ( .D(n_and_module_167_res), .CK(clock_0), 
        .Q(n_reg_module_305_res), .QN() );
  DFF_X1 u_reg_module_306__hpc_r0_reg ( .D(n_xor_module_276_res), .CK(clock_0), 
        .Q(n_reg_module_306_res), .QN() );
  AND2_X1 u_and_module_168_U1 ( .A1(n_reg_module_306_res), .A2(
        n_xor_module_196_res), .ZN(n_and_module_168_res) );
  DFF_X1 u_reg_module_307__hpc_r0_reg ( .D(n_and_module_168_res), .CK(clock_0), 
        .Q(n_reg_module_307_res), .QN() );
  DFF_X1 u_reg_module_308__hpc_r0_reg ( .D(n_and_module_164_res), .CK(clock_0), 
        .Q(n_reg_module_308_res), .QN() );
  XOR2_X1 u_xor_module_279_U1 ( .A(n_reg_module_308_res), .B(
        n_reg_module_307_res), .Z(n_xor_module_279_res) );
  XOR2_X1 u_xor_module_280_U1 ( .A(n_xor_module_279_res), .B(
        n_reg_module_305_res), .Z(n_xor_module_280_res) );
  DFF_X1 u_reg_module_309__hpc_r0_reg ( .D(p_rand_28), .CK(clock_0), .Q(
        n_reg_module_309_res), .QN() );
  INV_X1 u_not_module_57_U1 ( .A(n_xor_module_203_res), .ZN(
        n_not_module_57_res) );
  AND2_X1 u_and_module_169_U1 ( .A1(n_not_module_57_res), .A2(
        n_reg_module_309_res), .ZN(n_and_module_169_res) );
  XOR2_X1 u_xor_module_281_U1 ( .A(p_rand_28), .B(n_xor_module_6_res), .Z(
        n_xor_module_281_res) );
  INV_X1 u_not_module_58_U1 ( .A(n_xor_module_204_res), .ZN(
        n_not_module_58_res) );
  AND2_X1 u_and_module_170_U1 ( .A1(n_not_module_58_res), .A2(
        n_reg_module_309_res), .ZN(n_and_module_170_res) );
  XOR2_X1 u_xor_module_282_U1 ( .A(p_rand_28), .B(n_xor_module_5_res), .Z(
        n_xor_module_282_res) );
  DFF_X1 u_reg_module_310__hpc_r0_reg ( .D(n_xor_module_5_res), .CK(clock_0), 
        .Q(n_reg_module_310_res), .QN() );
  AND2_X1 u_and_module_171_U1 ( .A1(n_reg_module_310_res), .A2(
        n_xor_module_203_res), .ZN(n_and_module_171_res) );
  DFF_X1 u_reg_module_311__hpc_r0_reg ( .D(n_and_module_171_res), .CK(clock_0), 
        .Q(n_reg_module_311_res), .QN() );
  DFF_X1 u_reg_module_312__hpc_r0_reg ( .D(n_xor_module_281_res), .CK(clock_0), 
        .Q(n_reg_module_312_res), .QN() );
  AND2_X1 u_and_module_172_U1 ( .A1(n_reg_module_312_res), .A2(
        n_xor_module_203_res), .ZN(n_and_module_172_res) );
  DFF_X1 u_reg_module_313__hpc_r0_reg ( .D(n_and_module_172_res), .CK(clock_0), 
        .Q(n_reg_module_313_res), .QN() );
  DFF_X1 u_reg_module_314__hpc_r0_reg ( .D(n_and_module_169_res), .CK(clock_0), 
        .Q(n_reg_module_314_res), .QN() );
  XOR2_X1 u_xor_module_283_U1 ( .A(n_reg_module_314_res), .B(
        n_reg_module_313_res), .Z(n_xor_module_283_res) );
  XOR2_X1 u_xor_module_284_U1 ( .A(n_xor_module_283_res), .B(
        n_reg_module_311_res), .Z(n_xor_module_284_res) );
  DFF_X1 u_reg_module_315__hpc_r0_reg ( .D(n_xor_module_6_res), .CK(clock_0), 
        .Q(n_reg_module_315_res), .QN() );
  AND2_X1 u_and_module_173_U1 ( .A1(n_reg_module_315_res), .A2(
        n_xor_module_204_res), .ZN(n_and_module_173_res) );
  DFF_X1 u_reg_module_316__hpc_r0_reg ( .D(n_and_module_173_res), .CK(clock_0), 
        .Q(n_reg_module_316_res), .QN() );
  DFF_X1 u_reg_module_317__hpc_r0_reg ( .D(n_xor_module_282_res), .CK(clock_0), 
        .Q(n_reg_module_317_res), .QN() );
  AND2_X1 u_and_module_174_U1 ( .A1(n_reg_module_317_res), .A2(
        n_xor_module_204_res), .ZN(n_and_module_174_res) );
  DFF_X1 u_reg_module_318__hpc_r0_reg ( .D(n_and_module_174_res), .CK(clock_0), 
        .Q(n_reg_module_318_res), .QN() );
  DFF_X1 u_reg_module_319__hpc_r0_reg ( .D(n_and_module_170_res), .CK(clock_0), 
        .Q(n_reg_module_319_res), .QN() );
  XOR2_X1 u_xor_module_285_U1 ( .A(n_reg_module_319_res), .B(
        n_reg_module_318_res), .Z(n_xor_module_285_res) );
  XOR2_X1 u_xor_module_286_U1 ( .A(n_xor_module_285_res), .B(
        n_reg_module_316_res), .Z(n_xor_module_286_res) );
  DFF_X1 u_reg_module_320__hpc_r0_reg ( .D(p_rand_29), .CK(clock_0), .Q(
        n_reg_module_320_res), .QN() );
  INV_X1 u_not_module_59_U1 ( .A(n_xor_module_193_res), .ZN(
        n_not_module_59_res) );
  AND2_X1 u_and_module_175_U1 ( .A1(n_not_module_59_res), .A2(
        n_reg_module_320_res), .ZN(n_and_module_175_res) );
  XOR2_X1 u_xor_module_287_U1 ( .A(p_rand_29), .B(n_xor_module_44_res), .Z(
        n_xor_module_287_res) );
  INV_X1 u_not_module_60_U1 ( .A(n_xor_module_194_res), .ZN(
        n_not_module_60_res) );
  AND2_X1 u_and_module_176_U1 ( .A1(n_not_module_60_res), .A2(
        n_reg_module_320_res), .ZN(n_and_module_176_res) );
  XOR2_X1 u_xor_module_288_U1 ( .A(p_rand_29), .B(n_xor_module_43_res), .Z(
        n_xor_module_288_res) );
  DFF_X1 u_reg_module_321__hpc_r0_reg ( .D(n_xor_module_43_res), .CK(clock_0), 
        .Q(n_reg_module_321_res), .QN() );
  AND2_X1 u_and_module_177_U1 ( .A1(n_reg_module_321_res), .A2(
        n_xor_module_193_res), .ZN(n_and_module_177_res) );
  DFF_X1 u_reg_module_322__hpc_r0_reg ( .D(n_and_module_177_res), .CK(clock_0), 
        .Q(n_reg_module_322_res), .QN() );
  DFF_X1 u_reg_module_323__hpc_r0_reg ( .D(n_xor_module_287_res), .CK(clock_0), 
        .Q(n_reg_module_323_res), .QN() );
  AND2_X1 u_and_module_178_U1 ( .A1(n_reg_module_323_res), .A2(
        n_xor_module_193_res), .ZN(n_and_module_178_res) );
  DFF_X1 u_reg_module_324__hpc_r0_reg ( .D(n_and_module_178_res), .CK(clock_0), 
        .Q(n_reg_module_324_res), .QN() );
  DFF_X1 u_reg_module_325__hpc_r0_reg ( .D(n_and_module_175_res), .CK(clock_0), 
        .Q(n_reg_module_325_res), .QN() );
  XOR2_X1 u_xor_module_289_U1 ( .A(n_reg_module_325_res), .B(
        n_reg_module_324_res), .Z(n_xor_module_289_res) );
  XOR2_X1 u_xor_module_290_U1 ( .A(n_xor_module_289_res), .B(
        n_reg_module_322_res), .Z(n_xor_module_290_res) );
  DFF_X1 u_reg_module_326__hpc_r0_reg ( .D(n_xor_module_44_res), .CK(clock_0), 
        .Q(n_reg_module_326_res), .QN() );
  AND2_X1 u_and_module_179_U1 ( .A1(n_reg_module_326_res), .A2(
        n_xor_module_194_res), .ZN(n_and_module_179_res) );
  DFF_X1 u_reg_module_327__hpc_r0_reg ( .D(n_and_module_179_res), .CK(clock_0), 
        .Q(n_reg_module_327_res), .QN() );
  DFF_X1 u_reg_module_328__hpc_r0_reg ( .D(n_xor_module_288_res), .CK(clock_0), 
        .Q(n_reg_module_328_res), .QN() );
  AND2_X1 u_and_module_180_U1 ( .A1(n_reg_module_328_res), .A2(
        n_xor_module_194_res), .ZN(n_and_module_180_res) );
  DFF_X1 u_reg_module_329__hpc_r0_reg ( .D(n_and_module_180_res), .CK(clock_0), 
        .Q(n_reg_module_329_res), .QN() );
  DFF_X1 u_reg_module_330__hpc_r0_reg ( .D(n_and_module_176_res), .CK(clock_0), 
        .Q(n_reg_module_330_res), .QN() );
  XOR2_X1 u_xor_module_291_U1 ( .A(n_reg_module_330_res), .B(
        n_reg_module_329_res), .Z(n_xor_module_291_res) );
  XOR2_X1 u_xor_module_292_U1 ( .A(n_xor_module_291_res), .B(
        n_reg_module_327_res), .Z(n_xor_module_292_res) );
  DFF_X1 u_reg_module_331__hpc_r0_reg ( .D(p_rand_30), .CK(clock_0), .Q(
        n_reg_module_331_res), .QN() );
  INV_X1 u_not_module_61_U1 ( .A(n_xor_module_191_res), .ZN(
        n_not_module_61_res) );
  AND2_X1 u_and_module_181_U1 ( .A1(n_not_module_61_res), .A2(
        n_reg_module_331_res), .ZN(n_and_module_181_res) );
  XOR2_X1 u_xor_module_293_U1 ( .A(p_rand_30), .B(n_xor_module_40_res), .Z(
        n_xor_module_293_res) );
  INV_X1 u_not_module_62_U1 ( .A(n_xor_module_192_res), .ZN(
        n_not_module_62_res) );
  AND2_X1 u_and_module_182_U1 ( .A1(n_not_module_62_res), .A2(
        n_reg_module_331_res), .ZN(n_and_module_182_res) );
  XOR2_X1 u_xor_module_294_U1 ( .A(p_rand_30), .B(n_xor_module_39_res), .Z(
        n_xor_module_294_res) );
  DFF_X1 u_reg_module_332__hpc_r0_reg ( .D(n_xor_module_39_res), .CK(clock_0), 
        .Q(n_reg_module_332_res), .QN() );
  AND2_X1 u_and_module_183_U1 ( .A1(n_reg_module_332_res), .A2(
        n_xor_module_191_res), .ZN(n_and_module_183_res) );
  DFF_X1 u_reg_module_333__hpc_r0_reg ( .D(n_and_module_183_res), .CK(clock_0), 
        .Q(n_reg_module_333_res), .QN() );
  DFF_X1 u_reg_module_334__hpc_r0_reg ( .D(n_xor_module_293_res), .CK(clock_0), 
        .Q(n_reg_module_334_res), .QN() );
  AND2_X1 u_and_module_184_U1 ( .A1(n_reg_module_334_res), .A2(
        n_xor_module_191_res), .ZN(n_and_module_184_res) );
  DFF_X1 u_reg_module_335__hpc_r0_reg ( .D(n_and_module_184_res), .CK(clock_0), 
        .Q(n_reg_module_335_res), .QN() );
  DFF_X1 u_reg_module_336__hpc_r0_reg ( .D(n_and_module_181_res), .CK(clock_0), 
        .Q(n_reg_module_336_res), .QN() );
  XOR2_X1 u_xor_module_295_U1 ( .A(n_reg_module_336_res), .B(
        n_reg_module_335_res), .Z(n_xor_module_295_res) );
  XOR2_X1 u_xor_module_296_U1 ( .A(n_xor_module_295_res), .B(
        n_reg_module_333_res), .Z(n_xor_module_296_res) );
  DFF_X1 u_reg_module_337__hpc_r0_reg ( .D(n_xor_module_40_res), .CK(clock_0), 
        .Q(n_reg_module_337_res), .QN() );
  AND2_X1 u_and_module_185_U1 ( .A1(n_reg_module_337_res), .A2(
        n_xor_module_192_res), .ZN(n_and_module_185_res) );
  DFF_X1 u_reg_module_338__hpc_r0_reg ( .D(n_and_module_185_res), .CK(clock_0), 
        .Q(n_reg_module_338_res), .QN() );
  DFF_X1 u_reg_module_339__hpc_r0_reg ( .D(n_xor_module_294_res), .CK(clock_0), 
        .Q(n_reg_module_339_res), .QN() );
  AND2_X1 u_and_module_186_U1 ( .A1(n_reg_module_339_res), .A2(
        n_xor_module_192_res), .ZN(n_and_module_186_res) );
  DFF_X1 u_reg_module_340__hpc_r0_reg ( .D(n_and_module_186_res), .CK(clock_0), 
        .Q(n_reg_module_340_res), .QN() );
  DFF_X1 u_reg_module_341__hpc_r0_reg ( .D(n_and_module_182_res), .CK(clock_0), 
        .Q(n_reg_module_341_res), .QN() );
  XOR2_X1 u_xor_module_297_U1 ( .A(n_reg_module_341_res), .B(
        n_reg_module_340_res), .Z(n_xor_module_297_res) );
  XOR2_X1 u_xor_module_298_U1 ( .A(n_xor_module_297_res), .B(
        n_reg_module_338_res), .Z(n_xor_module_298_res) );
  DFF_X1 u_reg_module_342__hpc_r0_reg ( .D(p_rand_31), .CK(clock_0), .Q(
        n_reg_module_342_res), .QN() );
  INV_X1 u_not_module_63_U1 ( .A(n_xor_module_201_res), .ZN(
        n_not_module_63_res) );
  AND2_X1 u_and_module_187_U1 ( .A1(n_not_module_63_res), .A2(
        n_reg_module_342_res), .ZN(n_and_module_187_res) );
  XOR2_X1 u_xor_module_299_U1 ( .A(p_rand_31), .B(n_xor_module_2_res), .Z(
        n_xor_module_299_res) );
  INV_X1 u_not_module_64_U1 ( .A(n_xor_module_202_res), .ZN(
        n_not_module_64_res) );
  AND2_X1 u_and_module_188_U1 ( .A1(n_not_module_64_res), .A2(
        n_reg_module_342_res), .ZN(n_and_module_188_res) );
  XOR2_X1 u_xor_module_300_U1 ( .A(p_rand_31), .B(n_xor_module_1_res), .Z(
        n_xor_module_300_res) );
  DFF_X1 u_reg_module_343__hpc_r0_reg ( .D(n_xor_module_1_res), .CK(clock_0), 
        .Q(n_reg_module_343_res), .QN() );
  AND2_X1 u_and_module_189_U1 ( .A1(n_reg_module_343_res), .A2(
        n_xor_module_201_res), .ZN(n_and_module_189_res) );
  DFF_X1 u_reg_module_344__hpc_r0_reg ( .D(n_and_module_189_res), .CK(clock_0), 
        .Q(n_reg_module_344_res), .QN() );
  DFF_X1 u_reg_module_345__hpc_r0_reg ( .D(n_xor_module_299_res), .CK(clock_0), 
        .Q(n_reg_module_345_res), .QN() );
  AND2_X1 u_and_module_190_U1 ( .A1(n_reg_module_345_res), .A2(
        n_xor_module_201_res), .ZN(n_and_module_190_res) );
  DFF_X1 u_reg_module_346__hpc_r0_reg ( .D(n_and_module_190_res), .CK(clock_0), 
        .Q(n_reg_module_346_res), .QN() );
  DFF_X1 u_reg_module_347__hpc_r0_reg ( .D(n_and_module_187_res), .CK(clock_0), 
        .Q(n_reg_module_347_res), .QN() );
  XOR2_X1 u_xor_module_301_U1 ( .A(n_reg_module_347_res), .B(
        n_reg_module_346_res), .Z(n_xor_module_301_res) );
  XOR2_X1 u_xor_module_302_U1 ( .A(n_xor_module_301_res), .B(
        n_reg_module_344_res), .Z(n_xor_module_302_res) );
  DFF_X1 u_reg_module_348__hpc_r0_reg ( .D(n_xor_module_2_res), .CK(clock_0), 
        .Q(n_reg_module_348_res), .QN() );
  AND2_X1 u_and_module_191_U1 ( .A1(n_reg_module_348_res), .A2(
        n_xor_module_202_res), .ZN(n_and_module_191_res) );
  DFF_X1 u_reg_module_349__hpc_r0_reg ( .D(n_and_module_191_res), .CK(clock_0), 
        .Q(n_reg_module_349_res), .QN() );
  DFF_X1 u_reg_module_350__hpc_r0_reg ( .D(n_xor_module_300_res), .CK(clock_0), 
        .Q(n_reg_module_350_res), .QN() );
  AND2_X1 u_and_module_192_U1 ( .A1(n_reg_module_350_res), .A2(
        n_xor_module_202_res), .ZN(n_and_module_192_res) );
  DFF_X1 u_reg_module_351__hpc_r0_reg ( .D(n_and_module_192_res), .CK(clock_0), 
        .Q(n_reg_module_351_res), .QN() );
  DFF_X1 u_reg_module_352__hpc_r0_reg ( .D(n_and_module_188_res), .CK(clock_0), 
        .Q(n_reg_module_352_res), .QN() );
  XOR2_X1 u_xor_module_303_U1 ( .A(n_reg_module_352_res), .B(
        n_reg_module_351_res), .Z(n_xor_module_303_res) );
  XOR2_X1 u_xor_module_304_U1 ( .A(n_xor_module_303_res), .B(
        n_reg_module_349_res), .Z(n_xor_module_304_res) );
  DFF_X1 u_reg_module_353__hpc_r0_reg ( .D(p_rand_32), .CK(clock_0), .Q(
        n_reg_module_353_res), .QN() );
  INV_X1 u_not_module_65_U1 ( .A(n_xor_module_207_res), .ZN(
        n_not_module_65_res) );
  AND2_X1 u_and_module_193_U1 ( .A1(n_not_module_65_res), .A2(
        n_reg_module_353_res), .ZN(n_and_module_193_res) );
  XOR2_X1 u_xor_module_305_U1 ( .A(p_rand_32), .B(n_xor_module_8_res), .Z(
        n_xor_module_305_res) );
  INV_X1 u_not_module_66_U1 ( .A(n_xor_module_208_res), .ZN(
        n_not_module_66_res) );
  AND2_X1 u_and_module_194_U1 ( .A1(n_not_module_66_res), .A2(
        n_reg_module_353_res), .ZN(n_and_module_194_res) );
  XOR2_X1 u_xor_module_306_U1 ( .A(p_rand_32), .B(n_xor_module_7_res), .Z(
        n_xor_module_306_res) );
  DFF_X1 u_reg_module_354__hpc_r0_reg ( .D(n_xor_module_7_res), .CK(clock_0), 
        .Q(n_reg_module_354_res), .QN() );
  AND2_X1 u_and_module_195_U1 ( .A1(n_reg_module_354_res), .A2(
        n_xor_module_207_res), .ZN(n_and_module_195_res) );
  DFF_X1 u_reg_module_355__hpc_r0_reg ( .D(n_and_module_195_res), .CK(clock_0), 
        .Q(n_reg_module_355_res), .QN() );
  DFF_X1 u_reg_module_356__hpc_r0_reg ( .D(n_xor_module_305_res), .CK(clock_0), 
        .Q(n_reg_module_356_res), .QN() );
  AND2_X1 u_and_module_196_U1 ( .A1(n_reg_module_356_res), .A2(
        n_xor_module_207_res), .ZN(n_and_module_196_res) );
  DFF_X1 u_reg_module_357__hpc_r0_reg ( .D(n_and_module_196_res), .CK(clock_0), 
        .Q(n_reg_module_357_res), .QN() );
  DFF_X1 u_reg_module_358__hpc_r0_reg ( .D(n_and_module_193_res), .CK(clock_0), 
        .Q(n_reg_module_358_res), .QN() );
  XOR2_X1 u_xor_module_307_U1 ( .A(n_reg_module_358_res), .B(
        n_reg_module_357_res), .Z(n_xor_module_307_res) );
  XOR2_X1 u_xor_module_308_U1 ( .A(n_xor_module_307_res), .B(
        n_reg_module_355_res), .Z(n_xor_module_308_res) );
  DFF_X1 u_reg_module_359__hpc_r0_reg ( .D(n_xor_module_8_res), .CK(clock_0), 
        .Q(n_reg_module_359_res), .QN() );
  AND2_X1 u_and_module_197_U1 ( .A1(n_reg_module_359_res), .A2(
        n_xor_module_208_res), .ZN(n_and_module_197_res) );
  DFF_X1 u_reg_module_360__hpc_r0_reg ( .D(n_and_module_197_res), .CK(clock_0), 
        .Q(n_reg_module_360_res), .QN() );
  DFF_X1 u_reg_module_361__hpc_r0_reg ( .D(n_xor_module_306_res), .CK(clock_0), 
        .Q(n_reg_module_361_res), .QN() );
  AND2_X1 u_and_module_198_U1 ( .A1(n_reg_module_361_res), .A2(
        n_xor_module_208_res), .ZN(n_and_module_198_res) );
  DFF_X1 u_reg_module_362__hpc_r0_reg ( .D(n_and_module_198_res), .CK(clock_0), 
        .Q(n_reg_module_362_res), .QN() );
  DFF_X1 u_reg_module_363__hpc_r0_reg ( .D(n_and_module_194_res), .CK(clock_0), 
        .Q(n_reg_module_363_res), .QN() );
  XOR2_X1 u_xor_module_309_U1 ( .A(n_reg_module_363_res), .B(
        n_reg_module_362_res), .Z(n_xor_module_309_res) );
  XOR2_X1 u_xor_module_310_U1 ( .A(n_xor_module_309_res), .B(
        n_reg_module_360_res), .Z(n_xor_module_310_res) );
  DFF_X1 u_reg_module_364__hpc_r0_reg ( .D(p_rand_33), .CK(clock_0), .Q(
        n_reg_module_364_res), .QN() );
  INV_X1 u_not_module_67_U1 ( .A(n_xor_module_199_res), .ZN(
        n_not_module_67_res) );
  AND2_X1 u_and_module_199_U1 ( .A1(n_not_module_67_res), .A2(
        n_reg_module_364_res), .ZN(n_and_module_199_res) );
  XOR2_X1 u_xor_module_311_U1 ( .A(p_rand_33), .B(n_xor_module_4_res), .Z(
        n_xor_module_311_res) );
  INV_X1 u_not_module_68_U1 ( .A(n_xor_module_200_res), .ZN(
        n_not_module_68_res) );
  AND2_X1 u_and_module_200_U1 ( .A1(n_not_module_68_res), .A2(
        n_reg_module_364_res), .ZN(n_and_module_200_res) );
  XOR2_X1 u_xor_module_312_U1 ( .A(p_rand_33), .B(n_xor_module_3_res), .Z(
        n_xor_module_312_res) );
  DFF_X1 u_reg_module_365__hpc_r0_reg ( .D(n_xor_module_3_res), .CK(clock_0), 
        .Q(n_reg_module_365_res), .QN() );
  AND2_X1 u_and_module_201_U1 ( .A1(n_reg_module_365_res), .A2(
        n_xor_module_199_res), .ZN(n_and_module_201_res) );
  DFF_X1 u_reg_module_366__hpc_r0_reg ( .D(n_and_module_201_res), .CK(clock_0), 
        .Q(n_reg_module_366_res), .QN() );
  DFF_X1 u_reg_module_367__hpc_r0_reg ( .D(n_xor_module_311_res), .CK(clock_0), 
        .Q(n_reg_module_367_res), .QN() );
  AND2_X1 u_and_module_202_U1 ( .A1(n_reg_module_367_res), .A2(
        n_xor_module_199_res), .ZN(n_and_module_202_res) );
  DFF_X1 u_reg_module_368__hpc_r0_reg ( .D(n_and_module_202_res), .CK(clock_0), 
        .Q(n_reg_module_368_res), .QN() );
  DFF_X1 u_reg_module_369__hpc_r0_reg ( .D(n_and_module_199_res), .CK(clock_0), 
        .Q(n_reg_module_369_res), .QN() );
  XOR2_X1 u_xor_module_313_U1 ( .A(n_reg_module_369_res), .B(
        n_reg_module_368_res), .Z(n_xor_module_313_res) );
  XOR2_X1 u_xor_module_314_U1 ( .A(n_xor_module_313_res), .B(
        n_reg_module_366_res), .Z(n_xor_module_314_res) );
  DFF_X1 u_reg_module_370__hpc_r0_reg ( .D(n_xor_module_4_res), .CK(clock_0), 
        .Q(n_reg_module_370_res), .QN() );
  AND2_X1 u_and_module_203_U1 ( .A1(n_reg_module_370_res), .A2(
        n_xor_module_200_res), .ZN(n_and_module_203_res) );
  DFF_X1 u_reg_module_371__hpc_r0_reg ( .D(n_and_module_203_res), .CK(clock_0), 
        .Q(n_reg_module_371_res), .QN() );
  DFF_X1 u_reg_module_372__hpc_r0_reg ( .D(n_xor_module_312_res), .CK(clock_0), 
        .Q(n_reg_module_372_res), .QN() );
  AND2_X1 u_and_module_204_U1 ( .A1(n_reg_module_372_res), .A2(
        n_xor_module_200_res), .ZN(n_and_module_204_res) );
  DFF_X1 u_reg_module_373__hpc_r0_reg ( .D(n_and_module_204_res), .CK(clock_0), 
        .Q(n_reg_module_373_res), .QN() );
  DFF_X1 u_reg_module_374__hpc_r0_reg ( .D(n_and_module_200_res), .CK(clock_0), 
        .Q(n_reg_module_374_res), .QN() );
  XOR2_X1 u_xor_module_315_U1 ( .A(n_reg_module_374_res), .B(
        n_reg_module_373_res), .Z(n_xor_module_315_res) );
  XOR2_X1 u_xor_module_316_U1 ( .A(n_xor_module_315_res), .B(
        n_reg_module_371_res), .Z(n_xor_module_316_res) );
  XOR2_X1 u_xor_module_317_U1 ( .A(n_xor_module_308_res), .B(
        n_xor_module_302_res), .Z(n_xor_module_317_res) );
  XOR2_X1 u_xor_module_318_U1 ( .A(n_xor_module_310_res), .B(
        n_xor_module_304_res), .Z(n_xor_module_318_res) );
  XOR2_X1 u_xor_module_319_U1 ( .A(n_xor_module_272_res), .B(
        n_xor_module_236_res), .Z(n_xor_module_319_res) );
  XOR2_X1 u_xor_module_320_U1 ( .A(n_xor_module_274_res), .B(
        n_xor_module_238_res), .Z(n_xor_module_320_res) );
  XOR2_X1 u_xor_module_321_U1 ( .A(n_xor_module_224_res), .B(
        n_xor_module_212_res), .Z(n_xor_module_321_res) );
  XOR2_X1 u_xor_module_322_U1 ( .A(n_xor_module_226_res), .B(
        n_xor_module_214_res), .Z(n_xor_module_322_res) );
  XOR2_X1 u_xor_module_323_U1 ( .A(n_xor_module_266_res), .B(
        n_xor_module_218_res), .Z(n_xor_module_323_res) );
  XOR2_X1 u_xor_module_324_U1 ( .A(n_xor_module_268_res), .B(
        n_xor_module_220_res), .Z(n_xor_module_324_res) );
  XOR2_X1 u_xor_module_325_U1 ( .A(n_xor_module_284_res), .B(
        n_xor_module_260_res), .Z(n_xor_module_325_res) );
  XOR2_X1 u_xor_module_326_U1 ( .A(n_xor_module_286_res), .B(
        n_xor_module_262_res), .Z(n_xor_module_326_res) );
  XOR2_X1 u_xor_module_327_U1 ( .A(n_xor_module_302_res), .B(
        n_xor_module_230_res), .Z(n_xor_module_327_res) );
  XOR2_X1 u_xor_module_328_U1 ( .A(n_xor_module_304_res), .B(
        n_xor_module_232_res), .Z(n_xor_module_328_res) );
  XOR2_X1 u_xor_module_329_U1 ( .A(n_xor_module_327_res), .B(
        n_xor_module_308_res), .Z(n_xor_module_329_res) );
  XOR2_X1 u_xor_module_330_U1 ( .A(n_xor_module_328_res), .B(
        n_xor_module_310_res), .Z(n_xor_module_330_res) );
  XOR2_X1 u_xor_module_331_U1 ( .A(n_xor_module_323_res), .B(
        n_xor_module_212_res), .Z(n_xor_module_331_res) );
  XOR2_X1 u_xor_module_332_U1 ( .A(n_xor_module_324_res), .B(
        n_xor_module_214_res), .Z(n_xor_module_332_res) );
  XOR2_X1 u_xor_module_333_U1 ( .A(n_xor_module_290_res), .B(
        n_xor_module_242_res), .Z(n_xor_module_333_res) );
  XOR2_X1 u_xor_module_334_U1 ( .A(n_xor_module_292_res), .B(
        n_xor_module_244_res), .Z(n_xor_module_334_res) );
  XOR2_X1 u_xor_module_335_U1 ( .A(n_xor_module_254_res), .B(
        n_xor_module_248_res), .Z(n_xor_module_335_res) );
  XOR2_X1 u_xor_module_336_U1 ( .A(n_xor_module_256_res), .B(
        n_xor_module_250_res), .Z(n_xor_module_336_res) );
  XOR2_X1 u_xor_module_337_U1 ( .A(n_xor_module_325_res), .B(
        n_xor_module_254_res), .Z(n_xor_module_337_res) );
  XOR2_X1 u_xor_module_338_U1 ( .A(n_xor_module_326_res), .B(
        n_xor_module_256_res), .Z(n_xor_module_338_res) );
  XOR2_X1 u_xor_module_339_U1 ( .A(n_xor_module_321_res), .B(
        n_xor_module_296_res), .Z(n_xor_module_339_res) );
  XOR2_X1 u_xor_module_340_U1 ( .A(n_xor_module_322_res), .B(
        n_xor_module_298_res), .Z(n_xor_module_340_res) );
  XOR2_X1 u_xor_module_341_U1 ( .A(n_xor_module_242_res), .B(
        n_xor_module_224_res), .Z(n_xor_module_341_res) );
  XOR2_X1 u_xor_module_342_U1 ( .A(n_xor_module_244_res), .B(
        n_xor_module_226_res), .Z(n_xor_module_342_res) );
  XOR2_X1 u_xor_module_343_U1 ( .A(n_xor_module_317_res), .B(
        n_xor_module_236_res), .Z(n_xor_module_343_res) );
  XOR2_X1 u_xor_module_344_U1 ( .A(n_xor_module_318_res), .B(
        n_xor_module_238_res), .Z(n_xor_module_344_res) );
  XOR2_X1 u_xor_module_345_U1 ( .A(n_xor_module_302_res), .B(
        n_xor_module_248_res), .Z(n_xor_module_345_res) );
  XOR2_X1 u_xor_module_346_U1 ( .A(n_xor_module_304_res), .B(
        n_xor_module_250_res), .Z(n_xor_module_346_res) );
  XOR2_X1 u_xor_module_347_U1 ( .A(n_xor_module_319_res), .B(
        n_xor_module_266_res), .Z(n_xor_module_347_res) );
  XOR2_X1 u_xor_module_348_U1 ( .A(n_xor_module_320_res), .B(
        n_xor_module_268_res), .Z(n_xor_module_348_res) );
  XOR2_X1 u_xor_module_349_U1 ( .A(n_xor_module_317_res), .B(
        n_xor_module_272_res), .Z(n_xor_module_349_res) );
  XOR2_X1 u_xor_module_350_U1 ( .A(n_xor_module_318_res), .B(
        n_xor_module_274_res), .Z(n_xor_module_350_res) );
  XOR2_X1 u_xor_module_351_U1 ( .A(n_xor_module_319_res), .B(
        n_xor_module_278_res), .Z(n_xor_module_351_res) );
  XOR2_X1 u_xor_module_352_U1 ( .A(n_xor_module_320_res), .B(
        n_xor_module_280_res), .Z(n_xor_module_352_res) );
  XOR2_X1 u_xor_module_353_U1 ( .A(n_xor_module_333_res), .B(
        n_xor_module_284_res), .Z(n_xor_module_353_res) );
  XOR2_X1 u_xor_module_354_U1 ( .A(n_xor_module_334_res), .B(
        n_xor_module_286_res), .Z(n_xor_module_354_res) );
  XOR2_X1 u_xor_module_355_U1 ( .A(n_xor_module_325_res), .B(
        n_xor_module_314_res), .Z(n_xor_module_355_res) );
  XOR2_X1 u_xor_module_356_U1 ( .A(n_xor_module_326_res), .B(
        n_xor_module_316_res), .Z(n_xor_module_356_res) );
  XOR2_X1 u_xor_module_357_U1 ( .A(n_xor_module_319_res), .B(
        n_xor_module_317_res), .Z(n_xor_module_357_res) );
  XOR2_X1 u_xor_module_358_U1 ( .A(n_xor_module_320_res), .B(
        n_xor_module_318_res), .Z(n_xor_module_358_res) );
  XOR2_X1 u_xor_module_359_U1 ( .A(n_xor_module_331_res), .B(
        n_xor_module_319_res), .Z(n_xor_module_359_res) );
  XOR2_X1 u_xor_module_360_U1 ( .A(n_xor_module_332_res), .B(
        n_xor_module_320_res), .Z(n_xor_module_360_res) );
  XOR2_X1 u_xor_module_361_U1 ( .A(n_xor_module_341_res), .B(
        n_xor_module_323_res), .Z(n_xor_module_361_res) );
  XOR2_X1 u_xor_module_362_U1 ( .A(n_xor_module_342_res), .B(
        n_xor_module_324_res), .Z(n_xor_module_362_res) );
  XOR2_X1 u_xor_module_363_U1 ( .A(n_xor_module_321_res), .B(
        n_xor_module_353_res), .Z(n_xor_module_363_res) );
  XOR2_X1 u_xor_module_364_U1 ( .A(n_xor_module_322_res), .B(
        n_xor_module_354_res), .Z(n_xor_module_364_res) );
  XOR2_X1 u_xor_module_365_U1 ( .A(n_xor_module_335_res), .B(
        n_xor_module_347_res), .Z(n_xor_module_365_res) );
  XOR2_X1 u_xor_module_366_U1 ( .A(n_xor_module_336_res), .B(
        n_xor_module_348_res), .Z(n_xor_module_366_res) );
  XOR2_X1 u_xor_module_367_U1 ( .A(n_xor_module_337_res), .B(
        n_xor_module_329_res), .Z(n_xor_module_367_res) );
  XOR2_X1 u_xor_module_368_U1 ( .A(n_xor_module_338_res), .B(
        n_xor_module_330_res), .Z(n_xor_module_368_res) );
  XOR2_X1 u_xor_module_369_U1 ( .A(n_xor_module_335_res), .B(
        n_xor_module_331_res), .Z(n_xor_module_369_res) );
  XOR2_X1 u_xor_module_370_U1 ( .A(n_xor_module_336_res), .B(
        n_xor_module_332_res), .Z(n_xor_module_370_res) );
  XOR2_X1 u_xor_module_371_U1 ( .A(n_xor_module_337_res), .B(
        n_xor_module_333_res), .Z(n_xor_module_371_res) );
  XOR2_X1 u_xor_module_372_U1 ( .A(n_xor_module_338_res), .B(
        n_xor_module_334_res), .Z(n_xor_module_372_res) );
  XOR2_X1 u_xor_module_373_U1 ( .A(n_xor_module_345_res), .B(
        n_xor_module_339_res), .Z(n_xor_module_373_res) );
  XOR2_X1 u_xor_module_374_U1 ( .A(n_xor_module_346_res), .B(
        n_xor_module_340_res), .Z(n_xor_module_374_res) );
  XOR2_X1 u_xor_module_375_U1 ( .A(n_xor_module_351_res), .B(
        n_xor_module_339_res), .Z(n_xor_module_375_res) );
  XOR2_X1 u_xor_module_376_U1 ( .A(n_xor_module_352_res), .B(
        n_xor_module_340_res), .Z(n_xor_module_376_res) );
  XOR2_X1 u_xor_module_377_U1 ( .A(n_xor_module_365_res), .B(
        n_xor_module_329_res), .Z(n_xor_module_377_res) );
  XOR2_X1 u_xor_module_378_U1 ( .A(n_xor_module_366_res), .B(
        n_xor_module_330_res), .Z(n_xor_module_378_res) );
  XOR2_X1 u_xor_module_379_U1 ( .A(n_xor_module_369_res), .B(
        n_xor_module_349_res), .Z(n_xor_module_379_res) );
  XOR2_X1 u_xor_module_380_U1 ( .A(n_xor_module_370_res), .B(
        n_xor_module_350_res), .Z(n_xor_module_380_res) );
  INV_X1 u_not_module_69_U1 ( .A(n_xor_module_379_res), .ZN(
        n_not_module_69_res) );
  XOR2_X1 u_xor_module_381_U1 ( .A(n_xor_module_373_res), .B(
        n_xor_module_355_res), .Z(n_xor_module_381_res) );
  XOR2_X1 u_xor_module_382_U1 ( .A(n_xor_module_374_res), .B(
        n_xor_module_356_res), .Z(n_xor_module_382_res) );
  INV_X1 u_not_module_70_U1 ( .A(n_xor_module_381_res), .ZN(
        n_not_module_70_res) );
  XOR2_X1 u_xor_module_383_U1 ( .A(n_xor_module_359_res), .B(
        n_xor_module_329_res), .Z(n_xor_module_383_res) );
  XOR2_X1 u_xor_module_384_U1 ( .A(n_xor_module_360_res), .B(
        n_xor_module_330_res), .Z(n_xor_module_384_res) );
  XOR2_X1 u_xor_module_385_U1 ( .A(n_xor_module_361_res), .B(
        n_xor_module_357_res), .Z(n_xor_module_385_res) );
  XOR2_X1 u_xor_module_386_U1 ( .A(n_xor_module_362_res), .B(
        n_xor_module_358_res), .Z(n_xor_module_386_res) );
  XOR2_X1 u_xor_module_387_U1 ( .A(n_xor_module_375_res), .B(
        n_xor_module_367_res), .Z(n_xor_module_387_res) );
  XOR2_X1 u_xor_module_388_U1 ( .A(n_xor_module_376_res), .B(
        n_xor_module_368_res), .Z(n_xor_module_388_res) );
  XOR2_X1 u_xor_module_389_U1 ( .A(n_xor_module_371_res), .B(
        n_xor_module_343_res), .Z(n_xor_module_389_res) );
  XOR2_X1 u_xor_module_390_U1 ( .A(n_xor_module_372_res), .B(
        n_xor_module_344_res), .Z(n_xor_module_390_res) );
  INV_X1 u_not_module_71_U1 ( .A(n_xor_module_389_res), .ZN(
        n_not_module_71_res) );
  XOR2_X1 u_xor_module_391_U1 ( .A(n_xor_module_363_res), .B(
        n_xor_module_329_res), .Z(n_xor_module_391_res) );
  XOR2_X1 u_xor_module_392_U1 ( .A(n_xor_module_364_res), .B(
        n_xor_module_330_res), .Z(n_xor_module_392_res) );
  INV_X1 u_not_module_72_U1 ( .A(n_xor_module_391_res), .ZN(
        n_not_module_72_res) );
  XOR2_X1 u_xor_module_393_U1 ( .A(io_k0_s0), .B(n_xor_module_377_res), .Z(
        io_o0_s0) );
  XOR2_X1 u_xor_module_394_U1 ( .A(io_k0_s1), .B(n_xor_module_378_res), .Z(
        io_o0_s1) );
  XOR2_X1 u_xor_module_395_U1 ( .A(io_k1_s0), .B(n_not_module_69_res), .Z(
        io_o1_s0) );
  XOR2_X1 u_xor_module_396_U1 ( .A(io_k1_s1), .B(n_xor_module_380_res), .Z(
        io_o1_s1) );
  XOR2_X1 u_xor_module_397_U1 ( .A(io_k2_s0), .B(n_not_module_70_res), .Z(
        io_o2_s0) );
  XOR2_X1 u_xor_module_398_U1 ( .A(io_k2_s1), .B(n_xor_module_382_res), .Z(
        io_o2_s1) );
  XOR2_X1 u_xor_module_399_U1 ( .A(io_k3_s0), .B(n_xor_module_383_res), .Z(
        io_o3_s0) );
  XOR2_X1 u_xor_module_400_U1 ( .A(io_k3_s1), .B(n_xor_module_384_res), .Z(
        io_o3_s1) );
  XOR2_X1 u_xor_module_401_U1 ( .A(io_k4_s0), .B(n_xor_module_385_res), .Z(
        io_o4_s0) );
  XOR2_X1 u_xor_module_402_U1 ( .A(io_k4_s1), .B(n_xor_module_386_res), .Z(
        io_o4_s1) );
  XOR2_X1 u_xor_module_403_U1 ( .A(io_k5_s0), .B(n_xor_module_387_res), .Z(
        io_o5_s0) );
  XOR2_X1 u_xor_module_404_U1 ( .A(io_k5_s1), .B(n_xor_module_388_res), .Z(
        io_o5_s1) );
  XOR2_X1 u_xor_module_405_U1 ( .A(io_k6_s0), .B(n_not_module_71_res), .Z(
        io_o6_s0) );
  XOR2_X1 u_xor_module_406_U1 ( .A(io_k6_s1), .B(n_xor_module_390_res), .Z(
        io_o6_s1) );
  XOR2_X1 u_xor_module_407_U1 ( .A(io_k7_s0), .B(n_not_module_72_res), .Z(
        io_o7_s0) );
  XOR2_X1 u_xor_module_408_U1 ( .A(io_k7_s1), .B(n_xor_module_392_res), .Z(
        io_o7_s1) );
endmodule

