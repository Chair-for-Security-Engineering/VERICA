
module CINI ( io_a_0, io_a_1, io_a_2, io_a_3, io_b_0, io_b_1, io_b_2, io_b_3, 
        io_c_0, io_c_1, io_c_2, io_c_3, io_rand, clk, reset );
  input [6:0] io_a_0;
  input [6:0] io_a_1;
  input [6:0] io_a_2;
  input [6:0] io_a_3;
  input [6:0] io_b_0;
  input [6:0] io_b_1;
  input [6:0] io_b_2;
  input [6:0] io_b_3;
  output [6:0] io_c_0;
  output [6:0] io_c_1;
  output [6:0] io_c_2;
  output [6:0] io_c_3;
  input [5:0] io_rand;
  input clk, reset;
  wire   simpleNot_84_port_z, simpleNot_85_port_z, simpleNot_86_port_z,
         simpleNot_87_port_z, simpleNot_88_port_z, simpleNot_89_port_z,
         simpleNot_90_port_z, simpleNot_91_port_z, simpleNot_92_port_z,
         simpleNot_93_port_z, simpleNot_94_port_z, simpleNot_95_port_z,
         simpleNot_96_port_z, simpleNot_97_port_z, simpleNot_98_port_z,
         simpleNot_99_port_z, simpleNot_100_port_z, simpleNot_101_port_z,
         simpleNot_102_port_z, simpleNot_103_port_z, simpleNot_104_port_z,
         simpleNot_105_port_z, simpleNot_106_port_z, simpleNot_107_port_z,
         simpleNot_108_port_z, simpleNot_109_port_z, simpleNot_110_port_z,
         simpleNot_111_port_z, simpleNot_112_port_z, simpleNot_113_port_z,
         simpleNot_114_port_z, simpleNot_115_port_z, simpleNot_116_port_z,
         simpleNot_117_port_z, simpleNot_118_port_z, simpleNot_119_port_z,
         simpleNot_120_port_z, simpleNot_121_port_z, simpleNot_122_port_z,
         simpleNot_123_port_z, simpleNot_124_port_z, simpleNot_125_port_z,
         simpleNot_126_port_z, simpleNot_127_port_z, simpleNot_128_port_z,
         simpleNot_129_port_z, simpleNot_130_port_z, simpleNot_131_port_z,
         simpleNot_132_port_z, simpleNot_133_port_z, simpleNot_134_port_z,
         simpleNot_135_port_z, simpleNot_136_port_z, simpleNot_137_port_z,
         simpleNot_138_port_z, simpleNot_139_port_z, simpleNot_140_port_z,
         simpleNot_141_port_z, simpleNot_142_port_z, simpleNot_143_port_z,
         simpleNot_144_port_z, simpleNot_145_port_z, simpleNot_146_port_z,
         simpleNot_147_port_z, simpleNot_148_port_z, simpleNot_149_port_z,
         simpleNot_150_port_z, simpleNot_151_port_z, simpleNot_152_port_z,
         simpleNot_153_port_z, simpleNot_154_port_z, simpleNot_155_port_z,
         simpleNot_156_port_z, simpleNot_157_port_z, simpleNot_158_port_z,
         simpleNot_159_port_z, simpleNot_160_port_z, simpleNot_161_port_z,
         simpleNot_162_port_z, simpleNot_163_port_z, simpleNot_164_port_z,
         simpleNot_165_port_z, simpleNot_166_port_z, simpleNot_167_port_z,
         simpleXor_84_port_z, simpleXor_85_port_z, simpleXor_86_port_z,
         simpleXor_87_port_z, simpleXor_88_port_z, simpleXor_89_port_z,
         simpleXor_90_port_z, simpleXor_91_port_z, simpleXor_92_port_z,
         simpleXor_93_port_z, simpleXor_94_port_z, simpleXor_95_port_z,
         simpleXor_96_port_z, simpleXor_97_port_z, simpleXor_98_port_z,
         simpleXor_99_port_z, simpleXor_100_port_z, simpleXor_101_port_z,
         simpleXor_102_port_z, simpleXor_103_port_z, simpleXor_104_port_z,
         simpleXor_105_port_z, simpleXor_106_port_z, simpleXor_107_port_z,
         simpleXor_108_port_z, simpleXor_109_port_z, simpleXor_110_port_z,
         simpleXor_111_port_z, simpleXor_112_port_z, simpleXor_113_port_z,
         simpleXor_114_port_z, simpleXor_115_port_z, simpleXor_116_port_z,
         simpleXor_117_port_z, simpleXor_118_port_z, simpleXor_119_port_z,
         simpleXor_120_port_z, simpleXor_121_port_z, simpleXor_122_port_z,
         simpleXor_123_port_z, simpleXor_124_port_z, simpleXor_125_port_z,
         simpleXor_126_port_z, simpleXor_127_port_z, simpleXor_128_port_z,
         simpleXor_129_port_z, simpleXor_130_port_z, simpleXor_131_port_z,
         simpleXor_132_port_z, simpleXor_133_port_z, simpleXor_134_port_z,
         simpleXor_135_port_z, simpleXor_136_port_z, simpleXor_137_port_z,
         simpleXor_138_port_z, simpleXor_139_port_z, simpleXor_140_port_z,
         simpleXor_141_port_z, simpleXor_142_port_z, simpleXor_143_port_z,
         simpleXor_144_port_z, simpleXor_145_port_z, simpleXor_146_port_z,
         simpleXor_147_port_z, simpleXor_148_port_z, simpleXor_149_port_z,
         simpleXor_150_port_z, simpleXor_151_port_z, simpleXor_152_port_z,
         simpleXor_153_port_z, simpleXor_154_port_z, simpleXor_155_port_z,
         simpleXor_156_port_z, simpleXor_157_port_z, simpleXor_158_port_z,
         simpleXor_159_port_z, simpleXor_160_port_z, simpleXor_161_port_z,
         simpleXor_162_port_z, simpleXor_163_port_z, simpleXor_164_port_z,
         simpleXor_165_port_z, simpleXor_166_port_z, simpleXor_167_port_z,
         n_zz_io_c_0_0_, n_zz_io_c_1_0_, n_zz_io_c_2_0_, n_zz_io_c_3_0_,
         n_zz_io_c_0_5_0_, n_zz_io_c_1_5_0_, n_zz_io_c_2_5_0_,
         n_zz_io_c_3_5_0_, n_zz_io_c_0_10_0_, n_zz_io_c_1_10_0_,
         n_zz_io_c_2_10_0_, n_zz_io_c_3_10_0_, n_zz_io_c_0_15_0_,
         n_zz_io_c_1_15_0_, n_zz_io_c_2_15_0_, n_zz_io_c_3_15_0_,
         n_zz_io_c_0_20_0_, n_zz_io_c_1_20_0_, n_zz_io_c_2_20_0_,
         n_zz_io_c_3_20_0_, n_zz_io_c_0_25_0_, n_zz_io_c_1_25_0_,
         n_zz_io_c_2_25_0_, n_zz_io_c_3_25_0_, n_zz_io_c_0_30_0_,
         n_zz_io_c_1_30_0_, n_zz_io_c_2_30_0_, n_zz_io_c_3_30_0_, N0, N1, N2,
         N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, cor_maj_167_port_o,
         cor_maj_166_port_o, cor_maj_165_port_o, cor_maj_164_port_o,
         cor_maj_163_port_o, cor_maj_162_port_o, cor_maj_161_port_o,
         cor_maj_160_port_o, cor_maj_159_port_o, cor_maj_158_port_o,
         cor_maj_157_port_o, cor_maj_156_port_o, cor_maj_155_port_o,
         cor_maj_154_port_o, cor_maj_153_port_o, cor_maj_152_port_o,
         cor_maj_151_port_o, cor_maj_150_port_o, cor_maj_149_port_o,
         cor_maj_148_port_o, cor_maj_147_port_o, cor_maj_146_port_o,
         cor_maj_145_port_o, cor_maj_144_port_o, cor_maj_143_port_o,
         cor_maj_142_port_o, cor_maj_141_port_o, cor_maj_140_port_o,
         cor_maj_139_port_o, cor_maj_138_port_o, cor_maj_137_port_o,
         cor_maj_136_port_o, cor_maj_135_port_o, cor_maj_134_port_o,
         cor_maj_133_port_o, cor_maj_132_port_o, cor_maj_131_port_o,
         cor_maj_130_port_o, cor_maj_129_port_o, cor_maj_128_port_o,
         cor_maj_127_port_o, cor_maj_126_port_o, cor_maj_125_port_o,
         cor_maj_124_port_o, cor_maj_123_port_o, cor_maj_122_port_o,
         cor_maj_121_port_o, cor_maj_120_port_o, cor_maj_119_port_o,
         cor_maj_118_port_o, cor_maj_117_port_o, cor_maj_116_port_o,
         cor_maj_115_port_o, cor_maj_114_port_o, cor_maj_113_port_o,
         cor_maj_112_port_o, cor_maj_111_port_o, cor_maj_110_port_o,
         cor_maj_109_port_o, cor_maj_108_port_o, cor_maj_107_port_o,
         cor_maj_106_port_o, cor_maj_105_port_o, cor_maj_104_port_o,
         cor_maj_103_port_o, cor_maj_102_port_o, cor_maj_101_port_o,
         cor_maj_100_port_o, cor_maj_99_port_o, cor_maj_98_port_o,
         cor_maj_97_port_o, cor_maj_96_port_o, cor_maj_95_port_o,
         cor_maj_94_port_o, cor_maj_93_port_o, cor_maj_92_port_o,
         cor_maj_91_port_o, cor_maj_90_port_o, cor_maj_89_port_o,
         cor_maj_88_port_o, cor_maj_87_port_o, cor_maj_86_port_o,
         cor_maj_85_port_o, cor_maj_84_port_o, cor_maj_84_n17, cor_maj_84_n16,
         cor_maj_84_n15, cor_maj_84_n14, cor_maj_84_n13, cor_maj_84_n12,
         cor_maj_84_n11, cor_maj_84_n10, cor_maj_84_n9, cor_maj_84_n8,
         cor_maj_84_n7, cor_maj_84_n6, cor_maj_84_n5, cor_maj_84_n4,
         cor_maj_84_n3, cor_maj_84_n2, cor_maj_84_n1, cor_maj_85_n34,
         cor_maj_85_n33, cor_maj_85_n32, cor_maj_85_n31, cor_maj_85_n30,
         cor_maj_85_n29, cor_maj_85_n28, cor_maj_85_n27, cor_maj_85_n26,
         cor_maj_85_n25, cor_maj_85_n24, cor_maj_85_n23, cor_maj_85_n22,
         cor_maj_85_n21, cor_maj_85_n20, cor_maj_85_n19, cor_maj_85_n18,
         cor_maj_86_n34, cor_maj_86_n33, cor_maj_86_n32, cor_maj_86_n31,
         cor_maj_86_n30, cor_maj_86_n29, cor_maj_86_n28, cor_maj_86_n27,
         cor_maj_86_n26, cor_maj_86_n25, cor_maj_86_n24, cor_maj_86_n23,
         cor_maj_86_n22, cor_maj_86_n21, cor_maj_86_n20, cor_maj_86_n19,
         cor_maj_86_n18, cor_maj_87_n34, cor_maj_87_n33, cor_maj_87_n32,
         cor_maj_87_n31, cor_maj_87_n30, cor_maj_87_n29, cor_maj_87_n28,
         cor_maj_87_n27, cor_maj_87_n26, cor_maj_87_n25, cor_maj_87_n24,
         cor_maj_87_n23, cor_maj_87_n22, cor_maj_87_n21, cor_maj_87_n20,
         cor_maj_87_n19, cor_maj_87_n18, cor_maj_88_n34, cor_maj_88_n33,
         cor_maj_88_n32, cor_maj_88_n31, cor_maj_88_n30, cor_maj_88_n29,
         cor_maj_88_n28, cor_maj_88_n27, cor_maj_88_n26, cor_maj_88_n25,
         cor_maj_88_n24, cor_maj_88_n23, cor_maj_88_n22, cor_maj_88_n21,
         cor_maj_88_n20, cor_maj_88_n19, cor_maj_88_n18, cor_maj_89_n34,
         cor_maj_89_n33, cor_maj_89_n32, cor_maj_89_n31, cor_maj_89_n30,
         cor_maj_89_n29, cor_maj_89_n28, cor_maj_89_n27, cor_maj_89_n26,
         cor_maj_89_n25, cor_maj_89_n24, cor_maj_89_n23, cor_maj_89_n22,
         cor_maj_89_n21, cor_maj_89_n20, cor_maj_89_n19, cor_maj_89_n18,
         cor_maj_90_n34, cor_maj_90_n33, cor_maj_90_n32, cor_maj_90_n31,
         cor_maj_90_n30, cor_maj_90_n29, cor_maj_90_n28, cor_maj_90_n27,
         cor_maj_90_n26, cor_maj_90_n25, cor_maj_90_n24, cor_maj_90_n23,
         cor_maj_90_n22, cor_maj_90_n21, cor_maj_90_n20, cor_maj_90_n19,
         cor_maj_90_n18, cor_maj_91_n34, cor_maj_91_n33, cor_maj_91_n32,
         cor_maj_91_n31, cor_maj_91_n30, cor_maj_91_n29, cor_maj_91_n28,
         cor_maj_91_n27, cor_maj_91_n26, cor_maj_91_n25, cor_maj_91_n24,
         cor_maj_91_n23, cor_maj_91_n22, cor_maj_91_n21, cor_maj_91_n20,
         cor_maj_91_n19, cor_maj_91_n18, cor_maj_92_n34, cor_maj_92_n33,
         cor_maj_92_n32, cor_maj_92_n31, cor_maj_92_n30, cor_maj_92_n29,
         cor_maj_92_n28, cor_maj_92_n27, cor_maj_92_n26, cor_maj_92_n25,
         cor_maj_92_n24, cor_maj_92_n23, cor_maj_92_n22, cor_maj_92_n21,
         cor_maj_92_n20, cor_maj_92_n19, cor_maj_92_n18, cor_maj_93_n34,
         cor_maj_93_n33, cor_maj_93_n32, cor_maj_93_n31, cor_maj_93_n30,
         cor_maj_93_n29, cor_maj_93_n28, cor_maj_93_n27, cor_maj_93_n26,
         cor_maj_93_n25, cor_maj_93_n24, cor_maj_93_n23, cor_maj_93_n22,
         cor_maj_93_n21, cor_maj_93_n20, cor_maj_93_n19, cor_maj_93_n18,
         cor_maj_94_n34, cor_maj_94_n33, cor_maj_94_n32, cor_maj_94_n31,
         cor_maj_94_n30, cor_maj_94_n29, cor_maj_94_n28, cor_maj_94_n27,
         cor_maj_94_n26, cor_maj_94_n25, cor_maj_94_n24, cor_maj_94_n23,
         cor_maj_94_n22, cor_maj_94_n21, cor_maj_94_n20, cor_maj_94_n19,
         cor_maj_94_n18, cor_maj_95_n34, cor_maj_95_n33, cor_maj_95_n32,
         cor_maj_95_n31, cor_maj_95_n30, cor_maj_95_n29, cor_maj_95_n28,
         cor_maj_95_n27, cor_maj_95_n26, cor_maj_95_n25, cor_maj_95_n24,
         cor_maj_95_n23, cor_maj_95_n22, cor_maj_95_n21, cor_maj_95_n20,
         cor_maj_95_n19, cor_maj_95_n18, cor_maj_96_n34, cor_maj_96_n33,
         cor_maj_96_n32, cor_maj_96_n31, cor_maj_96_n30, cor_maj_96_n29,
         cor_maj_96_n28, cor_maj_96_n27, cor_maj_96_n26, cor_maj_96_n25,
         cor_maj_96_n24, cor_maj_96_n23, cor_maj_96_n22, cor_maj_96_n21,
         cor_maj_96_n20, cor_maj_96_n19, cor_maj_96_n18, cor_maj_97_n34,
         cor_maj_97_n33, cor_maj_97_n32, cor_maj_97_n31, cor_maj_97_n30,
         cor_maj_97_n29, cor_maj_97_n28, cor_maj_97_n27, cor_maj_97_n26,
         cor_maj_97_n25, cor_maj_97_n24, cor_maj_97_n23, cor_maj_97_n22,
         cor_maj_97_n21, cor_maj_97_n20, cor_maj_97_n19, cor_maj_97_n18,
         cor_maj_98_n34, cor_maj_98_n33, cor_maj_98_n32, cor_maj_98_n31,
         cor_maj_98_n30, cor_maj_98_n29, cor_maj_98_n28, cor_maj_98_n27,
         cor_maj_98_n26, cor_maj_98_n25, cor_maj_98_n24, cor_maj_98_n23,
         cor_maj_98_n22, cor_maj_98_n21, cor_maj_98_n20, cor_maj_98_n19,
         cor_maj_98_n18, cor_maj_99_n34, cor_maj_99_n33, cor_maj_99_n32,
         cor_maj_99_n31, cor_maj_99_n30, cor_maj_99_n29, cor_maj_99_n28,
         cor_maj_99_n27, cor_maj_99_n26, cor_maj_99_n25, cor_maj_99_n24,
         cor_maj_99_n23, cor_maj_99_n22, cor_maj_99_n21, cor_maj_99_n20,
         cor_maj_99_n19, cor_maj_99_n18, cor_maj_100_n34, cor_maj_100_n33,
         cor_maj_100_n32, cor_maj_100_n31, cor_maj_100_n30, cor_maj_100_n29,
         cor_maj_100_n28, cor_maj_100_n27, cor_maj_100_n26, cor_maj_100_n25,
         cor_maj_100_n24, cor_maj_100_n23, cor_maj_100_n22, cor_maj_100_n21,
         cor_maj_100_n20, cor_maj_100_n19, cor_maj_100_n18, cor_maj_101_n34,
         cor_maj_101_n33, cor_maj_101_n32, cor_maj_101_n31, cor_maj_101_n30,
         cor_maj_101_n29, cor_maj_101_n28, cor_maj_101_n27, cor_maj_101_n26,
         cor_maj_101_n25, cor_maj_101_n24, cor_maj_101_n23, cor_maj_101_n22,
         cor_maj_101_n21, cor_maj_101_n20, cor_maj_101_n19, cor_maj_101_n18,
         cor_maj_102_n34, cor_maj_102_n33, cor_maj_102_n32, cor_maj_102_n31,
         cor_maj_102_n30, cor_maj_102_n29, cor_maj_102_n28, cor_maj_102_n27,
         cor_maj_102_n26, cor_maj_102_n25, cor_maj_102_n24, cor_maj_102_n23,
         cor_maj_102_n22, cor_maj_102_n21, cor_maj_102_n20, cor_maj_102_n19,
         cor_maj_102_n18, cor_maj_103_n34, cor_maj_103_n33, cor_maj_103_n32,
         cor_maj_103_n31, cor_maj_103_n30, cor_maj_103_n29, cor_maj_103_n28,
         cor_maj_103_n27, cor_maj_103_n26, cor_maj_103_n25, cor_maj_103_n24,
         cor_maj_103_n23, cor_maj_103_n22, cor_maj_103_n21, cor_maj_103_n20,
         cor_maj_103_n19, cor_maj_103_n18, cor_maj_104_n34, cor_maj_104_n33,
         cor_maj_104_n32, cor_maj_104_n31, cor_maj_104_n30, cor_maj_104_n29,
         cor_maj_104_n28, cor_maj_104_n27, cor_maj_104_n26, cor_maj_104_n25,
         cor_maj_104_n24, cor_maj_104_n23, cor_maj_104_n22, cor_maj_104_n21,
         cor_maj_104_n20, cor_maj_104_n19, cor_maj_104_n18, cor_maj_105_n34,
         cor_maj_105_n33, cor_maj_105_n32, cor_maj_105_n31, cor_maj_105_n30,
         cor_maj_105_n29, cor_maj_105_n28, cor_maj_105_n27, cor_maj_105_n26,
         cor_maj_105_n25, cor_maj_105_n24, cor_maj_105_n23, cor_maj_105_n22,
         cor_maj_105_n21, cor_maj_105_n20, cor_maj_105_n19, cor_maj_105_n18,
         cor_maj_106_n34, cor_maj_106_n33, cor_maj_106_n32, cor_maj_106_n31,
         cor_maj_106_n30, cor_maj_106_n29, cor_maj_106_n28, cor_maj_106_n27,
         cor_maj_106_n26, cor_maj_106_n25, cor_maj_106_n24, cor_maj_106_n23,
         cor_maj_106_n22, cor_maj_106_n21, cor_maj_106_n20, cor_maj_106_n19,
         cor_maj_106_n18, cor_maj_107_n34, cor_maj_107_n33, cor_maj_107_n32,
         cor_maj_107_n31, cor_maj_107_n30, cor_maj_107_n29, cor_maj_107_n28,
         cor_maj_107_n27, cor_maj_107_n26, cor_maj_107_n25, cor_maj_107_n24,
         cor_maj_107_n23, cor_maj_107_n22, cor_maj_107_n21, cor_maj_107_n20,
         cor_maj_107_n19, cor_maj_107_n18, cor_maj_108_n34, cor_maj_108_n33,
         cor_maj_108_n32, cor_maj_108_n31, cor_maj_108_n30, cor_maj_108_n29,
         cor_maj_108_n28, cor_maj_108_n27, cor_maj_108_n26, cor_maj_108_n25,
         cor_maj_108_n24, cor_maj_108_n23, cor_maj_108_n22, cor_maj_108_n21,
         cor_maj_108_n20, cor_maj_108_n19, cor_maj_108_n18, cor_maj_109_n34,
         cor_maj_109_n33, cor_maj_109_n32, cor_maj_109_n31, cor_maj_109_n30,
         cor_maj_109_n29, cor_maj_109_n28, cor_maj_109_n27, cor_maj_109_n26,
         cor_maj_109_n25, cor_maj_109_n24, cor_maj_109_n23, cor_maj_109_n22,
         cor_maj_109_n21, cor_maj_109_n20, cor_maj_109_n19, cor_maj_109_n18,
         cor_maj_110_n34, cor_maj_110_n33, cor_maj_110_n32, cor_maj_110_n31,
         cor_maj_110_n30, cor_maj_110_n29, cor_maj_110_n28, cor_maj_110_n27,
         cor_maj_110_n26, cor_maj_110_n25, cor_maj_110_n24, cor_maj_110_n23,
         cor_maj_110_n22, cor_maj_110_n21, cor_maj_110_n20, cor_maj_110_n19,
         cor_maj_110_n18, cor_maj_111_n34, cor_maj_111_n33, cor_maj_111_n32,
         cor_maj_111_n31, cor_maj_111_n30, cor_maj_111_n29, cor_maj_111_n28,
         cor_maj_111_n27, cor_maj_111_n26, cor_maj_111_n25, cor_maj_111_n24,
         cor_maj_111_n23, cor_maj_111_n22, cor_maj_111_n21, cor_maj_111_n20,
         cor_maj_111_n19, cor_maj_111_n18, cor_maj_112_n34, cor_maj_112_n33,
         cor_maj_112_n32, cor_maj_112_n31, cor_maj_112_n30, cor_maj_112_n29,
         cor_maj_112_n28, cor_maj_112_n27, cor_maj_112_n26, cor_maj_112_n25,
         cor_maj_112_n24, cor_maj_112_n23, cor_maj_112_n22, cor_maj_112_n21,
         cor_maj_112_n20, cor_maj_112_n19, cor_maj_112_n18, cor_maj_113_n34,
         cor_maj_113_n33, cor_maj_113_n32, cor_maj_113_n31, cor_maj_113_n30,
         cor_maj_113_n29, cor_maj_113_n28, cor_maj_113_n27, cor_maj_113_n26,
         cor_maj_113_n25, cor_maj_113_n24, cor_maj_113_n23, cor_maj_113_n22,
         cor_maj_113_n21, cor_maj_113_n20, cor_maj_113_n19, cor_maj_113_n18,
         cor_maj_114_n34, cor_maj_114_n33, cor_maj_114_n32, cor_maj_114_n31,
         cor_maj_114_n30, cor_maj_114_n29, cor_maj_114_n28, cor_maj_114_n27,
         cor_maj_114_n26, cor_maj_114_n25, cor_maj_114_n24, cor_maj_114_n23,
         cor_maj_114_n22, cor_maj_114_n21, cor_maj_114_n20, cor_maj_114_n19,
         cor_maj_114_n18, cor_maj_115_n34, cor_maj_115_n33, cor_maj_115_n32,
         cor_maj_115_n31, cor_maj_115_n30, cor_maj_115_n29, cor_maj_115_n28,
         cor_maj_115_n27, cor_maj_115_n26, cor_maj_115_n25, cor_maj_115_n24,
         cor_maj_115_n23, cor_maj_115_n22, cor_maj_115_n21, cor_maj_115_n20,
         cor_maj_115_n19, cor_maj_115_n18, cor_maj_116_n34, cor_maj_116_n33,
         cor_maj_116_n32, cor_maj_116_n31, cor_maj_116_n30, cor_maj_116_n29,
         cor_maj_116_n28, cor_maj_116_n27, cor_maj_116_n26, cor_maj_116_n25,
         cor_maj_116_n24, cor_maj_116_n23, cor_maj_116_n22, cor_maj_116_n21,
         cor_maj_116_n20, cor_maj_116_n19, cor_maj_116_n18, cor_maj_117_n34,
         cor_maj_117_n33, cor_maj_117_n32, cor_maj_117_n31, cor_maj_117_n30,
         cor_maj_117_n29, cor_maj_117_n28, cor_maj_117_n27, cor_maj_117_n26,
         cor_maj_117_n25, cor_maj_117_n24, cor_maj_117_n23, cor_maj_117_n22,
         cor_maj_117_n21, cor_maj_117_n20, cor_maj_117_n19, cor_maj_117_n18,
         cor_maj_118_n34, cor_maj_118_n33, cor_maj_118_n32, cor_maj_118_n31,
         cor_maj_118_n30, cor_maj_118_n29, cor_maj_118_n28, cor_maj_118_n27,
         cor_maj_118_n26, cor_maj_118_n25, cor_maj_118_n24, cor_maj_118_n23,
         cor_maj_118_n22, cor_maj_118_n21, cor_maj_118_n20, cor_maj_118_n19,
         cor_maj_118_n18, cor_maj_119_n34, cor_maj_119_n33, cor_maj_119_n32,
         cor_maj_119_n31, cor_maj_119_n30, cor_maj_119_n29, cor_maj_119_n28,
         cor_maj_119_n27, cor_maj_119_n26, cor_maj_119_n25, cor_maj_119_n24,
         cor_maj_119_n23, cor_maj_119_n22, cor_maj_119_n21, cor_maj_119_n20,
         cor_maj_119_n19, cor_maj_119_n18, cor_maj_120_n34, cor_maj_120_n33,
         cor_maj_120_n32, cor_maj_120_n31, cor_maj_120_n30, cor_maj_120_n29,
         cor_maj_120_n28, cor_maj_120_n27, cor_maj_120_n26, cor_maj_120_n25,
         cor_maj_120_n24, cor_maj_120_n23, cor_maj_120_n22, cor_maj_120_n21,
         cor_maj_120_n20, cor_maj_120_n19, cor_maj_120_n18, cor_maj_121_n34,
         cor_maj_121_n33, cor_maj_121_n32, cor_maj_121_n31, cor_maj_121_n30,
         cor_maj_121_n29, cor_maj_121_n28, cor_maj_121_n27, cor_maj_121_n26,
         cor_maj_121_n25, cor_maj_121_n24, cor_maj_121_n23, cor_maj_121_n22,
         cor_maj_121_n21, cor_maj_121_n20, cor_maj_121_n19, cor_maj_121_n18,
         cor_maj_122_n34, cor_maj_122_n33, cor_maj_122_n32, cor_maj_122_n31,
         cor_maj_122_n30, cor_maj_122_n29, cor_maj_122_n28, cor_maj_122_n27,
         cor_maj_122_n26, cor_maj_122_n25, cor_maj_122_n24, cor_maj_122_n23,
         cor_maj_122_n22, cor_maj_122_n21, cor_maj_122_n20, cor_maj_122_n19,
         cor_maj_122_n18, cor_maj_123_n34, cor_maj_123_n33, cor_maj_123_n32,
         cor_maj_123_n31, cor_maj_123_n30, cor_maj_123_n29, cor_maj_123_n28,
         cor_maj_123_n27, cor_maj_123_n26, cor_maj_123_n25, cor_maj_123_n24,
         cor_maj_123_n23, cor_maj_123_n22, cor_maj_123_n21, cor_maj_123_n20,
         cor_maj_123_n19, cor_maj_123_n18, cor_maj_124_n34, cor_maj_124_n33,
         cor_maj_124_n32, cor_maj_124_n31, cor_maj_124_n30, cor_maj_124_n29,
         cor_maj_124_n28, cor_maj_124_n27, cor_maj_124_n26, cor_maj_124_n25,
         cor_maj_124_n24, cor_maj_124_n23, cor_maj_124_n22, cor_maj_124_n21,
         cor_maj_124_n20, cor_maj_124_n19, cor_maj_124_n18, cor_maj_125_n34,
         cor_maj_125_n33, cor_maj_125_n32, cor_maj_125_n31, cor_maj_125_n30,
         cor_maj_125_n29, cor_maj_125_n28, cor_maj_125_n27, cor_maj_125_n26,
         cor_maj_125_n25, cor_maj_125_n24, cor_maj_125_n23, cor_maj_125_n22,
         cor_maj_125_n21, cor_maj_125_n20, cor_maj_125_n19, cor_maj_125_n18,
         cor_maj_126_n34, cor_maj_126_n33, cor_maj_126_n32, cor_maj_126_n31,
         cor_maj_126_n30, cor_maj_126_n29, cor_maj_126_n28, cor_maj_126_n27,
         cor_maj_126_n26, cor_maj_126_n25, cor_maj_126_n24, cor_maj_126_n23,
         cor_maj_126_n22, cor_maj_126_n21, cor_maj_126_n20, cor_maj_126_n19,
         cor_maj_126_n18, cor_maj_127_n34, cor_maj_127_n33, cor_maj_127_n32,
         cor_maj_127_n31, cor_maj_127_n30, cor_maj_127_n29, cor_maj_127_n28,
         cor_maj_127_n27, cor_maj_127_n26, cor_maj_127_n25, cor_maj_127_n24,
         cor_maj_127_n23, cor_maj_127_n22, cor_maj_127_n21, cor_maj_127_n20,
         cor_maj_127_n19, cor_maj_127_n18, cor_maj_128_n34, cor_maj_128_n33,
         cor_maj_128_n32, cor_maj_128_n31, cor_maj_128_n30, cor_maj_128_n29,
         cor_maj_128_n28, cor_maj_128_n27, cor_maj_128_n26, cor_maj_128_n25,
         cor_maj_128_n24, cor_maj_128_n23, cor_maj_128_n22, cor_maj_128_n21,
         cor_maj_128_n20, cor_maj_128_n19, cor_maj_128_n18, cor_maj_129_n34,
         cor_maj_129_n33, cor_maj_129_n32, cor_maj_129_n31, cor_maj_129_n30,
         cor_maj_129_n29, cor_maj_129_n28, cor_maj_129_n27, cor_maj_129_n26,
         cor_maj_129_n25, cor_maj_129_n24, cor_maj_129_n23, cor_maj_129_n22,
         cor_maj_129_n21, cor_maj_129_n20, cor_maj_129_n19, cor_maj_129_n18,
         cor_maj_130_n34, cor_maj_130_n33, cor_maj_130_n32, cor_maj_130_n31,
         cor_maj_130_n30, cor_maj_130_n29, cor_maj_130_n28, cor_maj_130_n27,
         cor_maj_130_n26, cor_maj_130_n25, cor_maj_130_n24, cor_maj_130_n23,
         cor_maj_130_n22, cor_maj_130_n21, cor_maj_130_n20, cor_maj_130_n19,
         cor_maj_130_n18, cor_maj_131_n34, cor_maj_131_n33, cor_maj_131_n32,
         cor_maj_131_n31, cor_maj_131_n30, cor_maj_131_n29, cor_maj_131_n28,
         cor_maj_131_n27, cor_maj_131_n26, cor_maj_131_n25, cor_maj_131_n24,
         cor_maj_131_n23, cor_maj_131_n22, cor_maj_131_n21, cor_maj_131_n20,
         cor_maj_131_n19, cor_maj_131_n18, cor_maj_132_n34, cor_maj_132_n33,
         cor_maj_132_n32, cor_maj_132_n31, cor_maj_132_n30, cor_maj_132_n29,
         cor_maj_132_n28, cor_maj_132_n27, cor_maj_132_n26, cor_maj_132_n25,
         cor_maj_132_n24, cor_maj_132_n23, cor_maj_132_n22, cor_maj_132_n21,
         cor_maj_132_n20, cor_maj_132_n19, cor_maj_132_n18, cor_maj_133_n34,
         cor_maj_133_n33, cor_maj_133_n32, cor_maj_133_n31, cor_maj_133_n30,
         cor_maj_133_n29, cor_maj_133_n28, cor_maj_133_n27, cor_maj_133_n26,
         cor_maj_133_n25, cor_maj_133_n24, cor_maj_133_n23, cor_maj_133_n22,
         cor_maj_133_n21, cor_maj_133_n20, cor_maj_133_n19, cor_maj_133_n18,
         cor_maj_134_n34, cor_maj_134_n33, cor_maj_134_n32, cor_maj_134_n31,
         cor_maj_134_n30, cor_maj_134_n29, cor_maj_134_n28, cor_maj_134_n27,
         cor_maj_134_n26, cor_maj_134_n25, cor_maj_134_n24, cor_maj_134_n23,
         cor_maj_134_n22, cor_maj_134_n21, cor_maj_134_n20, cor_maj_134_n19,
         cor_maj_134_n18, cor_maj_135_n34, cor_maj_135_n33, cor_maj_135_n32,
         cor_maj_135_n31, cor_maj_135_n30, cor_maj_135_n29, cor_maj_135_n28,
         cor_maj_135_n27, cor_maj_135_n26, cor_maj_135_n25, cor_maj_135_n24,
         cor_maj_135_n23, cor_maj_135_n22, cor_maj_135_n21, cor_maj_135_n20,
         cor_maj_135_n19, cor_maj_135_n18, cor_maj_136_n34, cor_maj_136_n33,
         cor_maj_136_n32, cor_maj_136_n31, cor_maj_136_n30, cor_maj_136_n29,
         cor_maj_136_n28, cor_maj_136_n27, cor_maj_136_n26, cor_maj_136_n25,
         cor_maj_136_n24, cor_maj_136_n23, cor_maj_136_n22, cor_maj_136_n21,
         cor_maj_136_n20, cor_maj_136_n19, cor_maj_136_n18, cor_maj_137_n34,
         cor_maj_137_n33, cor_maj_137_n32, cor_maj_137_n31, cor_maj_137_n30,
         cor_maj_137_n29, cor_maj_137_n28, cor_maj_137_n27, cor_maj_137_n26,
         cor_maj_137_n25, cor_maj_137_n24, cor_maj_137_n23, cor_maj_137_n22,
         cor_maj_137_n21, cor_maj_137_n20, cor_maj_137_n19, cor_maj_137_n18,
         cor_maj_138_n34, cor_maj_138_n33, cor_maj_138_n32, cor_maj_138_n31,
         cor_maj_138_n30, cor_maj_138_n29, cor_maj_138_n28, cor_maj_138_n27,
         cor_maj_138_n26, cor_maj_138_n25, cor_maj_138_n24, cor_maj_138_n23,
         cor_maj_138_n22, cor_maj_138_n21, cor_maj_138_n20, cor_maj_138_n19,
         cor_maj_138_n18, cor_maj_139_n34, cor_maj_139_n33, cor_maj_139_n32,
         cor_maj_139_n31, cor_maj_139_n30, cor_maj_139_n29, cor_maj_139_n28,
         cor_maj_139_n27, cor_maj_139_n26, cor_maj_139_n25, cor_maj_139_n24,
         cor_maj_139_n23, cor_maj_139_n22, cor_maj_139_n21, cor_maj_139_n20,
         cor_maj_139_n19, cor_maj_139_n18, cor_maj_140_n34, cor_maj_140_n33,
         cor_maj_140_n32, cor_maj_140_n31, cor_maj_140_n30, cor_maj_140_n29,
         cor_maj_140_n28, cor_maj_140_n27, cor_maj_140_n26, cor_maj_140_n25,
         cor_maj_140_n24, cor_maj_140_n23, cor_maj_140_n22, cor_maj_140_n21,
         cor_maj_140_n20, cor_maj_140_n19, cor_maj_140_n18, cor_maj_141_n34,
         cor_maj_141_n33, cor_maj_141_n32, cor_maj_141_n31, cor_maj_141_n30,
         cor_maj_141_n29, cor_maj_141_n28, cor_maj_141_n27, cor_maj_141_n26,
         cor_maj_141_n25, cor_maj_141_n24, cor_maj_141_n23, cor_maj_141_n22,
         cor_maj_141_n21, cor_maj_141_n20, cor_maj_141_n19, cor_maj_141_n18,
         cor_maj_142_n34, cor_maj_142_n33, cor_maj_142_n32, cor_maj_142_n31,
         cor_maj_142_n30, cor_maj_142_n29, cor_maj_142_n28, cor_maj_142_n27,
         cor_maj_142_n26, cor_maj_142_n25, cor_maj_142_n24, cor_maj_142_n23,
         cor_maj_142_n22, cor_maj_142_n21, cor_maj_142_n20, cor_maj_142_n19,
         cor_maj_142_n18, cor_maj_143_n34, cor_maj_143_n33, cor_maj_143_n32,
         cor_maj_143_n31, cor_maj_143_n30, cor_maj_143_n29, cor_maj_143_n28,
         cor_maj_143_n27, cor_maj_143_n26, cor_maj_143_n25, cor_maj_143_n24,
         cor_maj_143_n23, cor_maj_143_n22, cor_maj_143_n21, cor_maj_143_n20,
         cor_maj_143_n19, cor_maj_143_n18, cor_maj_144_n34, cor_maj_144_n33,
         cor_maj_144_n32, cor_maj_144_n31, cor_maj_144_n30, cor_maj_144_n29,
         cor_maj_144_n28, cor_maj_144_n27, cor_maj_144_n26, cor_maj_144_n25,
         cor_maj_144_n24, cor_maj_144_n23, cor_maj_144_n22, cor_maj_144_n21,
         cor_maj_144_n20, cor_maj_144_n19, cor_maj_144_n18, cor_maj_145_n34,
         cor_maj_145_n33, cor_maj_145_n32, cor_maj_145_n31, cor_maj_145_n30,
         cor_maj_145_n29, cor_maj_145_n28, cor_maj_145_n27, cor_maj_145_n26,
         cor_maj_145_n25, cor_maj_145_n24, cor_maj_145_n23, cor_maj_145_n22,
         cor_maj_145_n21, cor_maj_145_n20, cor_maj_145_n19, cor_maj_145_n18,
         cor_maj_146_n34, cor_maj_146_n33, cor_maj_146_n32, cor_maj_146_n31,
         cor_maj_146_n30, cor_maj_146_n29, cor_maj_146_n28, cor_maj_146_n27,
         cor_maj_146_n26, cor_maj_146_n25, cor_maj_146_n24, cor_maj_146_n23,
         cor_maj_146_n22, cor_maj_146_n21, cor_maj_146_n20, cor_maj_146_n19,
         cor_maj_146_n18, cor_maj_147_n34, cor_maj_147_n33, cor_maj_147_n32,
         cor_maj_147_n31, cor_maj_147_n30, cor_maj_147_n29, cor_maj_147_n28,
         cor_maj_147_n27, cor_maj_147_n26, cor_maj_147_n25, cor_maj_147_n24,
         cor_maj_147_n23, cor_maj_147_n22, cor_maj_147_n21, cor_maj_147_n20,
         cor_maj_147_n19, cor_maj_147_n18, cor_maj_148_n34, cor_maj_148_n33,
         cor_maj_148_n32, cor_maj_148_n31, cor_maj_148_n30, cor_maj_148_n29,
         cor_maj_148_n28, cor_maj_148_n27, cor_maj_148_n26, cor_maj_148_n25,
         cor_maj_148_n24, cor_maj_148_n23, cor_maj_148_n22, cor_maj_148_n21,
         cor_maj_148_n20, cor_maj_148_n19, cor_maj_148_n18, cor_maj_149_n34,
         cor_maj_149_n33, cor_maj_149_n32, cor_maj_149_n31, cor_maj_149_n30,
         cor_maj_149_n29, cor_maj_149_n28, cor_maj_149_n27, cor_maj_149_n26,
         cor_maj_149_n25, cor_maj_149_n24, cor_maj_149_n23, cor_maj_149_n22,
         cor_maj_149_n21, cor_maj_149_n20, cor_maj_149_n19, cor_maj_149_n18,
         cor_maj_150_n34, cor_maj_150_n33, cor_maj_150_n32, cor_maj_150_n31,
         cor_maj_150_n30, cor_maj_150_n29, cor_maj_150_n28, cor_maj_150_n27,
         cor_maj_150_n26, cor_maj_150_n25, cor_maj_150_n24, cor_maj_150_n23,
         cor_maj_150_n22, cor_maj_150_n21, cor_maj_150_n20, cor_maj_150_n19,
         cor_maj_150_n18, cor_maj_151_n34, cor_maj_151_n33, cor_maj_151_n32,
         cor_maj_151_n31, cor_maj_151_n30, cor_maj_151_n29, cor_maj_151_n28,
         cor_maj_151_n27, cor_maj_151_n26, cor_maj_151_n25, cor_maj_151_n24,
         cor_maj_151_n23, cor_maj_151_n22, cor_maj_151_n21, cor_maj_151_n20,
         cor_maj_151_n19, cor_maj_151_n18, cor_maj_152_n34, cor_maj_152_n33,
         cor_maj_152_n32, cor_maj_152_n31, cor_maj_152_n30, cor_maj_152_n29,
         cor_maj_152_n28, cor_maj_152_n27, cor_maj_152_n26, cor_maj_152_n25,
         cor_maj_152_n24, cor_maj_152_n23, cor_maj_152_n22, cor_maj_152_n21,
         cor_maj_152_n20, cor_maj_152_n19, cor_maj_152_n18, cor_maj_153_n34,
         cor_maj_153_n33, cor_maj_153_n32, cor_maj_153_n31, cor_maj_153_n30,
         cor_maj_153_n29, cor_maj_153_n28, cor_maj_153_n27, cor_maj_153_n26,
         cor_maj_153_n25, cor_maj_153_n24, cor_maj_153_n23, cor_maj_153_n22,
         cor_maj_153_n21, cor_maj_153_n20, cor_maj_153_n19, cor_maj_153_n18,
         cor_maj_154_n34, cor_maj_154_n33, cor_maj_154_n32, cor_maj_154_n31,
         cor_maj_154_n30, cor_maj_154_n29, cor_maj_154_n28, cor_maj_154_n27,
         cor_maj_154_n26, cor_maj_154_n25, cor_maj_154_n24, cor_maj_154_n23,
         cor_maj_154_n22, cor_maj_154_n21, cor_maj_154_n20, cor_maj_154_n19,
         cor_maj_154_n18, cor_maj_155_n34, cor_maj_155_n33, cor_maj_155_n32,
         cor_maj_155_n31, cor_maj_155_n30, cor_maj_155_n29, cor_maj_155_n28,
         cor_maj_155_n27, cor_maj_155_n26, cor_maj_155_n25, cor_maj_155_n24,
         cor_maj_155_n23, cor_maj_155_n22, cor_maj_155_n21, cor_maj_155_n20,
         cor_maj_155_n19, cor_maj_155_n18, cor_maj_156_n34, cor_maj_156_n33,
         cor_maj_156_n32, cor_maj_156_n31, cor_maj_156_n30, cor_maj_156_n29,
         cor_maj_156_n28, cor_maj_156_n27, cor_maj_156_n26, cor_maj_156_n25,
         cor_maj_156_n24, cor_maj_156_n23, cor_maj_156_n22, cor_maj_156_n21,
         cor_maj_156_n20, cor_maj_156_n19, cor_maj_156_n18, cor_maj_157_n34,
         cor_maj_157_n33, cor_maj_157_n32, cor_maj_157_n31, cor_maj_157_n30,
         cor_maj_157_n29, cor_maj_157_n28, cor_maj_157_n27, cor_maj_157_n26,
         cor_maj_157_n25, cor_maj_157_n24, cor_maj_157_n23, cor_maj_157_n22,
         cor_maj_157_n21, cor_maj_157_n20, cor_maj_157_n19, cor_maj_157_n18,
         cor_maj_158_n34, cor_maj_158_n33, cor_maj_158_n32, cor_maj_158_n31,
         cor_maj_158_n30, cor_maj_158_n29, cor_maj_158_n28, cor_maj_158_n27,
         cor_maj_158_n26, cor_maj_158_n25, cor_maj_158_n24, cor_maj_158_n23,
         cor_maj_158_n22, cor_maj_158_n21, cor_maj_158_n20, cor_maj_158_n19,
         cor_maj_158_n18, cor_maj_159_n34, cor_maj_159_n33, cor_maj_159_n32,
         cor_maj_159_n31, cor_maj_159_n30, cor_maj_159_n29, cor_maj_159_n28,
         cor_maj_159_n27, cor_maj_159_n26, cor_maj_159_n25, cor_maj_159_n24,
         cor_maj_159_n23, cor_maj_159_n22, cor_maj_159_n21, cor_maj_159_n20,
         cor_maj_159_n19, cor_maj_159_n18, cor_maj_160_n34, cor_maj_160_n33,
         cor_maj_160_n32, cor_maj_160_n31, cor_maj_160_n30, cor_maj_160_n29,
         cor_maj_160_n28, cor_maj_160_n27, cor_maj_160_n26, cor_maj_160_n25,
         cor_maj_160_n24, cor_maj_160_n23, cor_maj_160_n22, cor_maj_160_n21,
         cor_maj_160_n20, cor_maj_160_n19, cor_maj_160_n18, cor_maj_161_n34,
         cor_maj_161_n33, cor_maj_161_n32, cor_maj_161_n31, cor_maj_161_n30,
         cor_maj_161_n29, cor_maj_161_n28, cor_maj_161_n27, cor_maj_161_n26,
         cor_maj_161_n25, cor_maj_161_n24, cor_maj_161_n23, cor_maj_161_n22,
         cor_maj_161_n21, cor_maj_161_n20, cor_maj_161_n19, cor_maj_161_n18,
         cor_maj_162_n34, cor_maj_162_n33, cor_maj_162_n32, cor_maj_162_n31,
         cor_maj_162_n30, cor_maj_162_n29, cor_maj_162_n28, cor_maj_162_n27,
         cor_maj_162_n26, cor_maj_162_n25, cor_maj_162_n24, cor_maj_162_n23,
         cor_maj_162_n22, cor_maj_162_n21, cor_maj_162_n20, cor_maj_162_n19,
         cor_maj_162_n18, cor_maj_163_n34, cor_maj_163_n33, cor_maj_163_n32,
         cor_maj_163_n31, cor_maj_163_n30, cor_maj_163_n29, cor_maj_163_n28,
         cor_maj_163_n27, cor_maj_163_n26, cor_maj_163_n25, cor_maj_163_n24,
         cor_maj_163_n23, cor_maj_163_n22, cor_maj_163_n21, cor_maj_163_n20,
         cor_maj_163_n19, cor_maj_163_n18, cor_maj_164_n34, cor_maj_164_n33,
         cor_maj_164_n32, cor_maj_164_n31, cor_maj_164_n30, cor_maj_164_n29,
         cor_maj_164_n28, cor_maj_164_n27, cor_maj_164_n26, cor_maj_164_n25,
         cor_maj_164_n24, cor_maj_164_n23, cor_maj_164_n22, cor_maj_164_n21,
         cor_maj_164_n20, cor_maj_164_n19, cor_maj_164_n18, cor_maj_165_n34,
         cor_maj_165_n33, cor_maj_165_n32, cor_maj_165_n31, cor_maj_165_n30,
         cor_maj_165_n29, cor_maj_165_n28, cor_maj_165_n27, cor_maj_165_n26,
         cor_maj_165_n25, cor_maj_165_n24, cor_maj_165_n23, cor_maj_165_n22,
         cor_maj_165_n21, cor_maj_165_n20, cor_maj_165_n19, cor_maj_165_n18,
         cor_maj_166_n34, cor_maj_166_n33, cor_maj_166_n32, cor_maj_166_n31,
         cor_maj_166_n30, cor_maj_166_n29, cor_maj_166_n28, cor_maj_166_n27,
         cor_maj_166_n26, cor_maj_166_n25, cor_maj_166_n24, cor_maj_166_n23,
         cor_maj_166_n22, cor_maj_166_n21, cor_maj_166_n20, cor_maj_166_n19,
         cor_maj_166_n18, cor_maj_167_n34, cor_maj_167_n33, cor_maj_167_n32,
         cor_maj_167_n31, cor_maj_167_n30, cor_maj_167_n29, cor_maj_167_n28,
         cor_maj_167_n27, cor_maj_167_n26, cor_maj_167_n25, cor_maj_167_n24,
         cor_maj_167_n23, cor_maj_167_n22, cor_maj_167_n21, cor_maj_167_n20,
         cor_maj_167_n19, cor_maj_167_n18;
  wire   [6:0] v_1_0_1;
  wire   [6:0] v_1_0_2;
  wire   [6:0] v_1_0_3;
  wire   [6:0] v_1_1_0;
  wire   [6:0] v_1_1_2;
  wire   [6:0] v_1_1_3;
  wire   [6:0] v_1_2_0;
  wire   [6:0] v_1_2_1;
  wire   [6:0] v_1_2_3;
  wire   [6:0] v_1_3_0;
  wire   [6:0] v_1_3_1;
  wire   [6:0] v_1_3_2;
  wire   [6:0] cor_port_v_0_1;
  wire   [6:0] cor_port_v_0_2;
  wire   [6:0] cor_port_v_0_3;
  wire   [6:0] cor_port_v_1_0;
  wire   [6:0] cor_port_v_1_2;
  wire   [6:0] cor_port_v_1_3;
  wire   [6:0] cor_port_v_2_0;
  wire   [6:0] cor_port_v_2_1;
  wire   [6:0] cor_port_v_2_3;
  wire   [6:0] cor_port_v_3_0;
  wire   [6:0] cor_port_v_3_1;
  wire   [6:0] cor_port_v_3_2;
  wire   [3:1] n_zz_io_c_0_4;
  wire   [6:0] u_0_1;
  wire   [6:0] u_0_2;
  wire   [6:0] u_0_3;
  wire   [3:1] n_zz_io_c_1_4;
  wire   [6:0] u_1_0;
  wire   [6:0] u_1_2;
  wire   [6:0] u_1_3;
  wire   [3:1] n_zz_io_c_2_4;
  wire   [6:0] u_2_0;
  wire   [6:0] u_2_1;
  wire   [6:0] u_2_3;
  wire   [3:1] n_zz_io_c_3_4;
  wire   [6:0] u_3_0;
  wire   [6:0] u_3_1;
  wire   [6:0] u_3_2;
  wire   [3:1] n_zz_io_c_0_9;
  wire   [3:1] n_zz_io_c_1_9;
  wire   [3:1] n_zz_io_c_2_9;
  wire   [3:1] n_zz_io_c_3_9;
  wire   [3:1] n_zz_io_c_0_14;
  wire   [3:1] n_zz_io_c_1_14;
  wire   [3:1] n_zz_io_c_2_14;
  wire   [3:1] n_zz_io_c_3_14;
  wire   [3:1] n_zz_io_c_0_19;
  wire   [3:1] n_zz_io_c_1_19;
  wire   [3:1] n_zz_io_c_2_19;
  wire   [3:1] n_zz_io_c_3_19;
  wire   [3:1] n_zz_io_c_0_24;
  wire   [3:1] n_zz_io_c_1_24;
  wire   [3:1] n_zz_io_c_2_24;
  wire   [3:1] n_zz_io_c_3_24;
  wire   [3:1] n_zz_io_c_0_29;
  wire   [3:1] n_zz_io_c_1_29;
  wire   [3:1] n_zz_io_c_2_29;
  wire   [3:1] n_zz_io_c_3_29;
  wire   [3:1] n_zz_io_c_0_34;
  wire   [3:1] n_zz_io_c_1_34;
  wire   [3:1] n_zz_io_c_2_34;
  wire   [3:1] n_zz_io_c_3_34;
  wire   [6:0] rand_reg_0;
  wire   [6:0] rand_reg_1;
  wire   [6:0] rand_reg_2;
  wire   [6:0] rand_reg_6;
  wire   [6:0] rand_reg_3;
  wire   [6:0] rand_reg_4;
  wire   [6:0] rand_reg_7;
  wire   [6:0] rand_reg_9;
  wire   [6:0] rand_reg_5;
  wire   [6:0] rand_reg_8;
  wire   [6:0] rand_reg_10;
  wire   [6:0] rand_reg_11;
  wire   [6:0] b_reg_0;
  wire   [6:0] b_reg_1;
  wire   [6:0] b_reg_2;
  wire   [6:0] b_reg_3;

  DFF_X1 b_reg_1_reg_6_ ( .D(io_b_1[6]), .CK(clk), .Q(b_reg_1[6]), .QN() );
  DFF_X1 b_reg_1_reg_5_ ( .D(io_b_1[5]), .CK(clk), .Q(b_reg_1[5]), .QN() );
  DFF_X1 b_reg_1_reg_4_ ( .D(io_b_1[4]), .CK(clk), .Q(b_reg_1[4]), .QN() );
  DFF_X1 b_reg_1_reg_3_ ( .D(io_b_1[3]), .CK(clk), .Q(b_reg_1[3]), .QN() );
  DFF_X1 b_reg_1_reg_2_ ( .D(io_b_1[2]), .CK(clk), .Q(b_reg_1[2]), .QN() );
  DFF_X1 b_reg_1_reg_1_ ( .D(io_b_1[1]), .CK(clk), .Q(b_reg_1[1]), .QN() );
  DFF_X1 b_reg_1_reg_0_ ( .D(io_b_1[0]), .CK(clk), .Q(b_reg_1[0]), .QN() );
  DFF_X1 b_reg_2_reg_6_ ( .D(io_b_2[6]), .CK(clk), .Q(b_reg_2[6]), .QN() );
  DFF_X1 b_reg_2_reg_5_ ( .D(io_b_2[5]), .CK(clk), .Q(b_reg_2[5]), .QN() );
  DFF_X1 b_reg_2_reg_4_ ( .D(io_b_2[4]), .CK(clk), .Q(b_reg_2[4]), .QN() );
  DFF_X1 b_reg_2_reg_3_ ( .D(io_b_2[3]), .CK(clk), .Q(b_reg_2[3]), .QN() );
  DFF_X1 b_reg_2_reg_2_ ( .D(io_b_2[2]), .CK(clk), .Q(b_reg_2[2]), .QN() );
  DFF_X1 b_reg_2_reg_1_ ( .D(io_b_2[1]), .CK(clk), .Q(b_reg_2[1]), .QN() );
  DFF_X1 b_reg_2_reg_0_ ( .D(io_b_2[0]), .CK(clk), .Q(b_reg_2[0]), .QN() );
  DFF_X1 b_reg_3_reg_6_ ( .D(io_b_3[6]), .CK(clk), .Q(b_reg_3[6]), .QN() );
  DFF_X1 b_reg_3_reg_5_ ( .D(io_b_3[5]), .CK(clk), .Q(b_reg_3[5]), .QN() );
  DFF_X1 b_reg_3_reg_4_ ( .D(io_b_3[4]), .CK(clk), .Q(b_reg_3[4]), .QN() );
  DFF_X1 b_reg_3_reg_3_ ( .D(io_b_3[3]), .CK(clk), .Q(b_reg_3[3]), .QN() );
  DFF_X1 b_reg_3_reg_2_ ( .D(io_b_3[2]), .CK(clk), .Q(b_reg_3[2]), .QN() );
  DFF_X1 b_reg_3_reg_1_ ( .D(io_b_3[1]), .CK(clk), .Q(b_reg_3[1]), .QN() );
  DFF_X1 b_reg_3_reg_0_ ( .D(io_b_3[0]), .CK(clk), .Q(b_reg_3[0]), .QN() );
  DFF_X1 u_zz_io_c_3_34_reg_3_ ( .D(N195), .CK(clk), .Q(n_zz_io_c_3_34[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_34_reg_2_ ( .D(N194), .CK(clk), .Q(n_zz_io_c_3_34[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_34_reg_1_ ( .D(N193), .CK(clk), .Q(n_zz_io_c_3_34[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_34_reg_0_ ( .D(N192), .CK(clk), .Q(n_zz_io_c_3_30_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_34_reg_3_ ( .D(N191), .CK(clk), .Q(n_zz_io_c_2_34[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_34_reg_2_ ( .D(N190), .CK(clk), .Q(n_zz_io_c_2_34[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_34_reg_1_ ( .D(N189), .CK(clk), .Q(n_zz_io_c_2_34[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_34_reg_0_ ( .D(N188), .CK(clk), .Q(n_zz_io_c_2_30_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_34_reg_3_ ( .D(N187), .CK(clk), .Q(n_zz_io_c_1_34[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_34_reg_2_ ( .D(N186), .CK(clk), .Q(n_zz_io_c_1_34[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_34_reg_1_ ( .D(N185), .CK(clk), .Q(n_zz_io_c_1_34[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_34_reg_0_ ( .D(N184), .CK(clk), .Q(n_zz_io_c_1_30_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_34_reg_3_ ( .D(N183), .CK(clk), .Q(n_zz_io_c_0_34[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_34_reg_2_ ( .D(N182), .CK(clk), .Q(n_zz_io_c_0_34[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_34_reg_1_ ( .D(N181), .CK(clk), .Q(n_zz_io_c_0_34[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_29_reg_3_ ( .D(N179), .CK(clk), .Q(n_zz_io_c_3_29[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_29_reg_2_ ( .D(N178), .CK(clk), .Q(n_zz_io_c_3_29[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_29_reg_1_ ( .D(N177), .CK(clk), .Q(n_zz_io_c_3_29[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_29_reg_0_ ( .D(N176), .CK(clk), .Q(n_zz_io_c_3_25_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_29_reg_3_ ( .D(N175), .CK(clk), .Q(n_zz_io_c_2_29[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_29_reg_2_ ( .D(N174), .CK(clk), .Q(n_zz_io_c_2_29[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_29_reg_1_ ( .D(N173), .CK(clk), .Q(n_zz_io_c_2_29[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_29_reg_0_ ( .D(N172), .CK(clk), .Q(n_zz_io_c_2_25_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_29_reg_3_ ( .D(N171), .CK(clk), .Q(n_zz_io_c_1_29[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_29_reg_2_ ( .D(N170), .CK(clk), .Q(n_zz_io_c_1_29[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_29_reg_1_ ( .D(N169), .CK(clk), .Q(n_zz_io_c_1_29[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_29_reg_0_ ( .D(N168), .CK(clk), .Q(n_zz_io_c_1_25_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_29_reg_3_ ( .D(N167), .CK(clk), .Q(n_zz_io_c_0_29[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_29_reg_2_ ( .D(N166), .CK(clk), .Q(n_zz_io_c_0_29[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_29_reg_1_ ( .D(N165), .CK(clk), .Q(n_zz_io_c_0_29[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_3_ ( .D(N163), .CK(clk), .Q(n_zz_io_c_3_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_2_ ( .D(N162), .CK(clk), .Q(n_zz_io_c_3_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_1_ ( .D(N161), .CK(clk), .Q(n_zz_io_c_3_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_0_ ( .D(N160), .CK(clk), .Q(n_zz_io_c_3_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_3_ ( .D(N159), .CK(clk), .Q(n_zz_io_c_2_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_2_ ( .D(N158), .CK(clk), .Q(n_zz_io_c_2_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_1_ ( .D(N157), .CK(clk), .Q(n_zz_io_c_2_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_0_ ( .D(N156), .CK(clk), .Q(n_zz_io_c_2_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_3_ ( .D(N155), .CK(clk), .Q(n_zz_io_c_1_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_2_ ( .D(N154), .CK(clk), .Q(n_zz_io_c_1_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_1_ ( .D(N153), .CK(clk), .Q(n_zz_io_c_1_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_0_ ( .D(N152), .CK(clk), .Q(n_zz_io_c_1_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_3_ ( .D(N151), .CK(clk), .Q(n_zz_io_c_0_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_2_ ( .D(N150), .CK(clk), .Q(n_zz_io_c_0_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_1_ ( .D(N149), .CK(clk), .Q(n_zz_io_c_0_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_3_ ( .D(N147), .CK(clk), .Q(n_zz_io_c_3_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_2_ ( .D(N146), .CK(clk), .Q(n_zz_io_c_3_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_1_ ( .D(N145), .CK(clk), .Q(n_zz_io_c_3_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_0_ ( .D(N144), .CK(clk), .Q(n_zz_io_c_3_15_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_3_ ( .D(N143), .CK(clk), .Q(n_zz_io_c_2_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_2_ ( .D(N142), .CK(clk), .Q(n_zz_io_c_2_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_1_ ( .D(N141), .CK(clk), .Q(n_zz_io_c_2_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_0_ ( .D(N140), .CK(clk), .Q(n_zz_io_c_2_15_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_3_ ( .D(N139), .CK(clk), .Q(n_zz_io_c_1_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_2_ ( .D(N138), .CK(clk), .Q(n_zz_io_c_1_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_1_ ( .D(N137), .CK(clk), .Q(n_zz_io_c_1_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_0_ ( .D(N136), .CK(clk), .Q(n_zz_io_c_1_15_0_), 
        .QN() );
  DFF_X1 rand_reg_9_reg_6_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[6]), 
        .QN() );
  DFF_X1 u_2_1_reg_6_ ( .D(N79), .CK(clk), .Q(u_2_1[6]), .QN() );
  DFF_X1 rand_reg_9_reg_5_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[5]), 
        .QN() );
  DFF_X1 u_2_1_reg_5_ ( .D(N67), .CK(clk), .Q(u_2_1[5]), .QN() );
  DFF_X1 rand_reg_9_reg_4_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[4]), 
        .QN() );
  DFF_X1 u_2_1_reg_4_ ( .D(N55), .CK(clk), .Q(u_2_1[4]), .QN() );
  DFF_X1 rand_reg_9_reg_3_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[3]), 
        .QN() );
  DFF_X1 u_2_1_reg_3_ ( .D(N43), .CK(clk), .Q(u_2_1[3]), .QN() );
  DFF_X1 rand_reg_9_reg_2_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[2]), 
        .QN() );
  DFF_X1 u_2_1_reg_2_ ( .D(N31), .CK(clk), .Q(u_2_1[2]), .QN() );
  DFF_X1 rand_reg_9_reg_1_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[1]), 
        .QN() );
  DFF_X1 u_2_1_reg_1_ ( .D(N19), .CK(clk), .Q(u_2_1[1]), .QN() );
  DFF_X1 rand_reg_9_reg_0_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[0]), 
        .QN() );
  DFF_X1 u_2_1_reg_0_ ( .D(N7), .CK(clk), .Q(u_2_1[0]), .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_3_ ( .D(N135), .CK(clk), .Q(n_zz_io_c_0_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_2_ ( .D(N134), .CK(clk), .Q(n_zz_io_c_0_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_1_ ( .D(N133), .CK(clk), .Q(n_zz_io_c_0_19[1]), 
        .QN() );
  DFF_X1 rand_reg_1_reg_6_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[6]), 
        .QN() );
  DFF_X1 u_0_2_reg_6_ ( .D(N73), .CK(clk), .Q(u_0_2[6]), .QN() );
  DFF_X1 rand_reg_1_reg_5_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[5]), 
        .QN() );
  DFF_X1 u_0_2_reg_5_ ( .D(N61), .CK(clk), .Q(u_0_2[5]), .QN() );
  DFF_X1 rand_reg_1_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[4]), 
        .QN() );
  DFF_X1 u_0_2_reg_4_ ( .D(N49), .CK(clk), .Q(u_0_2[4]), .QN() );
  DFF_X1 rand_reg_1_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[3]), 
        .QN() );
  DFF_X1 u_0_2_reg_3_ ( .D(N37), .CK(clk), .Q(u_0_2[3]), .QN() );
  DFF_X1 rand_reg_1_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[2]), 
        .QN() );
  DFF_X1 u_0_2_reg_2_ ( .D(N25), .CK(clk), .Q(u_0_2[2]), .QN() );
  DFF_X1 rand_reg_1_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[1]), 
        .QN() );
  DFF_X1 u_0_2_reg_1_ ( .D(N13), .CK(clk), .Q(u_0_2[1]), .QN() );
  DFF_X1 rand_reg_1_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[0]), 
        .QN() );
  DFF_X1 u_0_2_reg_0_ ( .D(N1), .CK(clk), .Q(u_0_2[0]), .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_3_ ( .D(N131), .CK(clk), .Q(n_zz_io_c_3_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_2_ ( .D(N130), .CK(clk), .Q(n_zz_io_c_3_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_1_ ( .D(N129), .CK(clk), .Q(n_zz_io_c_3_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_0_ ( .D(N128), .CK(clk), .Q(n_zz_io_c_3_10_0_), 
        .QN() );
  DFF_X1 rand_reg_0_reg_6_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[6]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_5_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[5]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[4]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[3]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[2]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[1]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[0]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_6_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[6]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_5_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[5]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_4_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[4]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_3_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[3]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_2_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[2]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_1_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[1]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_0_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[0]), 
        .QN() );
  DFF_X1 rand_reg_6_reg_6_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[6]), 
        .QN() );
  DFF_X1 u_1_0_reg_6_ ( .D(N75), .CK(clk), .Q(u_1_0[6]), .QN() );
  DFF_X1 rand_reg_6_reg_5_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[5]), 
        .QN() );
  DFF_X1 u_1_0_reg_5_ ( .D(N63), .CK(clk), .Q(u_1_0[5]), .QN() );
  DFF_X1 rand_reg_6_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[4]), 
        .QN() );
  DFF_X1 u_1_0_reg_4_ ( .D(N51), .CK(clk), .Q(u_1_0[4]), .QN() );
  DFF_X1 rand_reg_6_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[3]), 
        .QN() );
  DFF_X1 u_1_0_reg_3_ ( .D(N39), .CK(clk), .Q(u_1_0[3]), .QN() );
  DFF_X1 rand_reg_6_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[2]), 
        .QN() );
  DFF_X1 u_1_0_reg_2_ ( .D(N27), .CK(clk), .Q(u_1_0[2]), .QN() );
  DFF_X1 rand_reg_6_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[1]), 
        .QN() );
  DFF_X1 u_1_0_reg_1_ ( .D(N15), .CK(clk), .Q(u_1_0[1]), .QN() );
  DFF_X1 rand_reg_6_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[0]), 
        .QN() );
  DFF_X1 u_1_0_reg_0_ ( .D(N3), .CK(clk), .Q(u_1_0[0]), .QN() );
  DFF_X1 rand_reg_7_reg_6_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[6]), 
        .QN() );
  DFF_X1 u_2_0_reg_6_ ( .D(N78), .CK(clk), .Q(u_2_0[6]), .QN() );
  DFF_X1 rand_reg_7_reg_5_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[5]), 
        .QN() );
  DFF_X1 u_2_0_reg_5_ ( .D(N66), .CK(clk), .Q(u_2_0[5]), .QN() );
  DFF_X1 rand_reg_7_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[4]), 
        .QN() );
  DFF_X1 u_2_0_reg_4_ ( .D(N54), .CK(clk), .Q(u_2_0[4]), .QN() );
  DFF_X1 rand_reg_7_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[3]), 
        .QN() );
  DFF_X1 u_2_0_reg_3_ ( .D(N42), .CK(clk), .Q(u_2_0[3]), .QN() );
  DFF_X1 rand_reg_7_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[2]), 
        .QN() );
  DFF_X1 u_2_0_reg_2_ ( .D(N30), .CK(clk), .Q(u_2_0[2]), .QN() );
  DFF_X1 rand_reg_7_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[1]), 
        .QN() );
  DFF_X1 u_2_0_reg_1_ ( .D(N18), .CK(clk), .Q(u_2_0[1]), .QN() );
  DFF_X1 rand_reg_7_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[0]), 
        .QN() );
  DFF_X1 u_2_0_reg_0_ ( .D(N6), .CK(clk), .Q(u_2_0[0]), .QN() );
  DFF_X1 u_0_1_reg_6_ ( .D(N72), .CK(clk), .Q(u_0_1[6]), .QN() );
  DFF_X1 u_0_1_reg_5_ ( .D(N60), .CK(clk), .Q(u_0_1[5]), .QN() );
  DFF_X1 u_0_1_reg_4_ ( .D(N48), .CK(clk), .Q(u_0_1[4]), .QN() );
  DFF_X1 u_0_1_reg_3_ ( .D(N36), .CK(clk), .Q(u_0_1[3]), .QN() );
  DFF_X1 u_0_1_reg_2_ ( .D(N24), .CK(clk), .Q(u_0_1[2]), .QN() );
  DFF_X1 u_0_1_reg_1_ ( .D(N12), .CK(clk), .Q(u_0_1[1]), .QN() );
  DFF_X1 u_0_1_reg_0_ ( .D(N0), .CK(clk), .Q(u_0_1[0]), .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_3_ ( .D(N127), .CK(clk), .Q(n_zz_io_c_2_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_2_ ( .D(N126), .CK(clk), .Q(n_zz_io_c_2_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_1_ ( .D(N125), .CK(clk), .Q(n_zz_io_c_2_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_0_ ( .D(N124), .CK(clk), .Q(n_zz_io_c_2_10_0_), 
        .QN() );
  DFF_X1 rand_reg_2_reg_6_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[6]), 
        .QN() );
  DFF_X1 u_0_3_reg_6_ ( .D(N74), .CK(clk), .Q(u_0_3[6]), .QN() );
  DFF_X1 rand_reg_2_reg_5_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[5]), 
        .QN() );
  DFF_X1 u_0_3_reg_5_ ( .D(N62), .CK(clk), .Q(u_0_3[5]), .QN() );
  DFF_X1 rand_reg_2_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[4]), 
        .QN() );
  DFF_X1 u_0_3_reg_4_ ( .D(N50), .CK(clk), .Q(u_0_3[4]), .QN() );
  DFF_X1 rand_reg_2_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[3]), 
        .QN() );
  DFF_X1 u_0_3_reg_3_ ( .D(N38), .CK(clk), .Q(u_0_3[3]), .QN() );
  DFF_X1 rand_reg_2_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[2]), 
        .QN() );
  DFF_X1 u_0_3_reg_2_ ( .D(N26), .CK(clk), .Q(u_0_3[2]), .QN() );
  DFF_X1 rand_reg_2_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[1]), 
        .QN() );
  DFF_X1 u_0_3_reg_1_ ( .D(N14), .CK(clk), .Q(u_0_3[1]), .QN() );
  DFF_X1 rand_reg_2_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[0]), 
        .QN() );
  DFF_X1 u_0_3_reg_0_ ( .D(N2), .CK(clk), .Q(u_0_3[0]), .QN() );
  DFF_X1 rand_reg_8_reg_6_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[6]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_5_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[5]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[4]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[3]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[2]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[1]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[0]), 
        .QN() );
  DFF_X1 rand_reg_3_reg_6_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[6]), 
        .QN() );
  DFF_X1 u_1_2_reg_6_ ( .D(N76), .CK(clk), .Q(u_1_2[6]), .QN() );
  DFF_X1 rand_reg_3_reg_5_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[5]), 
        .QN() );
  DFF_X1 u_1_2_reg_5_ ( .D(N64), .CK(clk), .Q(u_1_2[5]), .QN() );
  DFF_X1 rand_reg_3_reg_4_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[4]), 
        .QN() );
  DFF_X1 u_1_2_reg_4_ ( .D(N52), .CK(clk), .Q(u_1_2[4]), .QN() );
  DFF_X1 rand_reg_3_reg_3_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[3]), 
        .QN() );
  DFF_X1 u_1_2_reg_3_ ( .D(N40), .CK(clk), .Q(u_1_2[3]), .QN() );
  DFF_X1 rand_reg_3_reg_2_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[2]), 
        .QN() );
  DFF_X1 u_1_2_reg_2_ ( .D(N28), .CK(clk), .Q(u_1_2[2]), .QN() );
  DFF_X1 rand_reg_3_reg_1_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[1]), 
        .QN() );
  DFF_X1 u_1_2_reg_1_ ( .D(N16), .CK(clk), .Q(u_1_2[1]), .QN() );
  DFF_X1 rand_reg_3_reg_0_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[0]), 
        .QN() );
  DFF_X1 u_1_2_reg_0_ ( .D(N4), .CK(clk), .Q(u_1_2[0]), .QN() );
  DFF_X1 rand_reg_4_reg_6_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[6]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_5_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[5]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_4_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[4]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_3_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[3]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_2_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[2]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_1_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[1]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_0_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[0]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_3_ ( .D(N123), .CK(clk), .Q(n_zz_io_c_1_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_2_ ( .D(N122), .CK(clk), .Q(n_zz_io_c_1_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_1_ ( .D(N121), .CK(clk), .Q(n_zz_io_c_1_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_0_ ( .D(N120), .CK(clk), .Q(n_zz_io_c_1_10_0_), 
        .QN() );
  DFF_X1 rand_reg_10_reg_6_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[6]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_5_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[5]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_4_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[4]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_3_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[3]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_2_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[2]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_1_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[1]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_0_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[0]), 
        .QN() );
  DFF_X1 rand_reg_5_reg_6_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[6]), 
        .QN() );
  DFF_X1 u_2_3_reg_6_ ( .D(N80), .CK(clk), .Q(u_2_3[6]), .QN() );
  DFF_X1 rand_reg_5_reg_5_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[5]), 
        .QN() );
  DFF_X1 u_2_3_reg_5_ ( .D(N68), .CK(clk), .Q(u_2_3[5]), .QN() );
  DFF_X1 rand_reg_5_reg_4_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[4]), 
        .QN() );
  DFF_X1 u_2_3_reg_4_ ( .D(N56), .CK(clk), .Q(u_2_3[4]), .QN() );
  DFF_X1 rand_reg_5_reg_3_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[3]), 
        .QN() );
  DFF_X1 u_2_3_reg_3_ ( .D(N44), .CK(clk), .Q(u_2_3[3]), .QN() );
  DFF_X1 rand_reg_5_reg_2_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[2]), 
        .QN() );
  DFF_X1 u_2_3_reg_2_ ( .D(N32), .CK(clk), .Q(u_2_3[2]), .QN() );
  DFF_X1 rand_reg_5_reg_1_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[1]), 
        .QN() );
  DFF_X1 u_2_3_reg_1_ ( .D(N20), .CK(clk), .Q(u_2_3[1]), .QN() );
  DFF_X1 rand_reg_5_reg_0_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[0]), 
        .QN() );
  DFF_X1 u_2_3_reg_0_ ( .D(N8), .CK(clk), .Q(u_2_3[0]), .QN() );
  DFF_X1 b_reg_0_reg_6_ ( .D(io_b_0[6]), .CK(clk), .Q(b_reg_0[6]), .QN() );
  DFF_X1 u_zz_io_c_0_34_reg_0_ ( .D(N180), .CK(clk), .Q(n_zz_io_c_0_30_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_5_ ( .D(io_b_0[5]), .CK(clk), .Q(b_reg_0[5]), .QN() );
  DFF_X1 u_zz_io_c_0_29_reg_0_ ( .D(N164), .CK(clk), .Q(n_zz_io_c_0_25_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_4_ ( .D(io_b_0[4]), .CK(clk), .Q(b_reg_0[4]), .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_0_ ( .D(N148), .CK(clk), .Q(n_zz_io_c_0_20_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_3_ ( .D(io_b_0[3]), .CK(clk), .Q(b_reg_0[3]), .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_0_ ( .D(N132), .CK(clk), .Q(n_zz_io_c_0_15_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_2_ ( .D(io_b_0[2]), .CK(clk), .Q(b_reg_0[2]), .QN() );
  DFF_X1 b_reg_0_reg_1_ ( .D(io_b_0[1]), .CK(clk), .Q(b_reg_0[1]), .QN() );
  DFF_X1 b_reg_0_reg_0_ ( .D(io_b_0[0]), .CK(clk), .Q(b_reg_0[0]), .QN() );
  DFF_X1 u_1_3_reg_6_ ( .D(N77), .CK(clk), .Q(u_1_3[6]), .QN() );
  DFF_X1 u_1_3_reg_5_ ( .D(N65), .CK(clk), .Q(u_1_3[5]), .QN() );
  DFF_X1 u_1_3_reg_4_ ( .D(N53), .CK(clk), .Q(u_1_3[4]), .QN() );
  DFF_X1 u_1_3_reg_3_ ( .D(N41), .CK(clk), .Q(u_1_3[3]), .QN() );
  DFF_X1 u_1_3_reg_2_ ( .D(N29), .CK(clk), .Q(u_1_3[2]), .QN() );
  DFF_X1 u_1_3_reg_1_ ( .D(N17), .CK(clk), .Q(u_1_3[1]), .QN() );
  DFF_X1 u_1_3_reg_0_ ( .D(N5), .CK(clk), .Q(u_1_3[0]), .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_3_ ( .D(N119), .CK(clk), .Q(n_zz_io_c_0_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_2_ ( .D(N118), .CK(clk), .Q(n_zz_io_c_0_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_1_ ( .D(N117), .CK(clk), .Q(n_zz_io_c_0_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_0_ ( .D(N116), .CK(clk), .Q(n_zz_io_c_0_10_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_3_9_reg_3_ ( .D(N115), .CK(clk), .Q(n_zz_io_c_3_9[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_9_reg_2_ ( .D(N114), .CK(clk), .Q(n_zz_io_c_3_9[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_9_reg_1_ ( .D(N113), .CK(clk), .Q(n_zz_io_c_3_9[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_9_reg_0_ ( .D(N112), .CK(clk), .Q(n_zz_io_c_3_5_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_9_reg_3_ ( .D(N111), .CK(clk), .Q(n_zz_io_c_2_9[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_9_reg_2_ ( .D(N110), .CK(clk), .Q(n_zz_io_c_2_9[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_9_reg_1_ ( .D(N109), .CK(clk), .Q(n_zz_io_c_2_9[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_9_reg_0_ ( .D(N108), .CK(clk), .Q(n_zz_io_c_2_5_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_9_reg_3_ ( .D(N107), .CK(clk), .Q(n_zz_io_c_1_9[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_9_reg_2_ ( .D(N106), .CK(clk), .Q(n_zz_io_c_1_9[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_9_reg_1_ ( .D(N105), .CK(clk), .Q(n_zz_io_c_1_9[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_9_reg_0_ ( .D(N104), .CK(clk), .Q(n_zz_io_c_1_5_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_9_reg_3_ ( .D(N103), .CK(clk), .Q(n_zz_io_c_0_9[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_9_reg_2_ ( .D(N102), .CK(clk), .Q(n_zz_io_c_0_9[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_9_reg_1_ ( .D(N101), .CK(clk), .Q(n_zz_io_c_0_9[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_9_reg_0_ ( .D(N100), .CK(clk), .Q(n_zz_io_c_0_5_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_3_4_reg_3_ ( .D(N99), .CK(clk), .Q(n_zz_io_c_3_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_3_4_reg_2_ ( .D(N98), .CK(clk), .Q(n_zz_io_c_3_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_3_4_reg_1_ ( .D(N97), .CK(clk), .Q(n_zz_io_c_3_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_3_4_reg_0_ ( .D(N96), .CK(clk), .Q(n_zz_io_c_3_0_), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_3_ ( .D(N95), .CK(clk), .Q(n_zz_io_c_2_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_2_ ( .D(N94), .CK(clk), .Q(n_zz_io_c_2_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_1_ ( .D(N93), .CK(clk), .Q(n_zz_io_c_2_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_0_ ( .D(N92), .CK(clk), .Q(n_zz_io_c_2_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_3_ ( .D(N91), .CK(clk), .Q(n_zz_io_c_1_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_2_ ( .D(N90), .CK(clk), .Q(n_zz_io_c_1_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_1_ ( .D(N89), .CK(clk), .Q(n_zz_io_c_1_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_0_ ( .D(N88), .CK(clk), .Q(n_zz_io_c_1_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_3_ ( .D(N87), .CK(clk), .Q(n_zz_io_c_0_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_2_ ( .D(N86), .CK(clk), .Q(n_zz_io_c_0_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_1_ ( .D(N85), .CK(clk), .Q(n_zz_io_c_0_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_0_ ( .D(N84), .CK(clk), .Q(n_zz_io_c_0_0_), .QN()
         );
  DFF_X1 u_3_2_reg_6_ ( .D(N83), .CK(clk), .Q(u_3_2[6]), .QN() );
  DFF_X1 u_3_2_reg_5_ ( .D(N71), .CK(clk), .Q(u_3_2[5]), .QN() );
  DFF_X1 u_3_2_reg_4_ ( .D(N59), .CK(clk), .Q(u_3_2[4]), .QN() );
  DFF_X1 u_3_2_reg_3_ ( .D(N47), .CK(clk), .Q(u_3_2[3]), .QN() );
  DFF_X1 u_3_2_reg_2_ ( .D(N35), .CK(clk), .Q(u_3_2[2]), .QN() );
  DFF_X1 u_3_2_reg_1_ ( .D(N23), .CK(clk), .Q(u_3_2[1]), .QN() );
  DFF_X1 u_3_2_reg_0_ ( .D(N11), .CK(clk), .Q(u_3_2[0]), .QN() );
  DFF_X1 u_3_1_reg_6_ ( .D(N82), .CK(clk), .Q(u_3_1[6]), .QN() );
  DFF_X1 u_3_1_reg_5_ ( .D(N70), .CK(clk), .Q(u_3_1[5]), .QN() );
  DFF_X1 u_3_1_reg_4_ ( .D(N58), .CK(clk), .Q(u_3_1[4]), .QN() );
  DFF_X1 u_3_1_reg_3_ ( .D(N46), .CK(clk), .Q(u_3_1[3]), .QN() );
  DFF_X1 u_3_1_reg_2_ ( .D(N34), .CK(clk), .Q(u_3_1[2]), .QN() );
  DFF_X1 u_3_1_reg_1_ ( .D(N22), .CK(clk), .Q(u_3_1[1]), .QN() );
  DFF_X1 u_3_1_reg_0_ ( .D(N10), .CK(clk), .Q(u_3_1[0]), .QN() );
  DFF_X1 u_3_0_reg_6_ ( .D(N81), .CK(clk), .Q(u_3_0[6]), .QN() );
  DFF_X1 u_3_0_reg_5_ ( .D(N69), .CK(clk), .Q(u_3_0[5]), .QN() );
  DFF_X1 u_3_0_reg_4_ ( .D(N57), .CK(clk), .Q(u_3_0[4]), .QN() );
  DFF_X1 u_3_0_reg_3_ ( .D(N45), .CK(clk), .Q(u_3_0[3]), .QN() );
  DFF_X1 u_3_0_reg_2_ ( .D(N33), .CK(clk), .Q(u_3_0[2]), .QN() );
  DFF_X1 u_3_0_reg_1_ ( .D(N21), .CK(clk), .Q(u_3_0[1]), .QN() );
  DFF_X1 u_3_0_reg_0_ ( .D(N9), .CK(clk), .Q(u_3_0[0]), .QN() );
  XOR2_X2 U4 ( .A(io_rand[5]), .B(io_b_2[5]), .Z(v_1_3_2[5]) );
  XOR2_X2 U5 ( .A(io_rand[5]), .B(io_b_2[4]), .Z(v_1_3_2[4]) );
  XOR2_X2 U6 ( .A(io_rand[5]), .B(io_b_2[3]), .Z(v_1_3_2[3]) );
  XOR2_X2 U7 ( .A(io_rand[5]), .B(io_b_2[2]), .Z(v_1_3_2[2]) );
  XOR2_X2 U8 ( .A(io_rand[5]), .B(io_b_2[1]), .Z(v_1_3_2[1]) );
  XOR2_X2 U9 ( .A(io_rand[5]), .B(io_b_2[0]), .Z(v_1_3_2[0]) );
  XOR2_X2 U11 ( .A(io_rand[4]), .B(io_b_1[5]), .Z(v_1_3_1[5]) );
  XOR2_X2 U12 ( .A(io_rand[4]), .B(io_b_1[4]), .Z(v_1_3_1[4]) );
  XOR2_X2 U13 ( .A(io_rand[4]), .B(io_b_1[3]), .Z(v_1_3_1[3]) );
  XOR2_X2 U14 ( .A(io_rand[4]), .B(io_b_1[2]), .Z(v_1_3_1[2]) );
  XOR2_X2 U15 ( .A(io_rand[4]), .B(io_b_1[1]), .Z(v_1_3_1[1]) );
  XOR2_X2 U16 ( .A(io_rand[4]), .B(io_b_1[0]), .Z(v_1_3_1[0]) );
  XOR2_X2 U18 ( .A(io_rand[2]), .B(io_b_0[5]), .Z(v_1_3_0[5]) );
  XOR2_X2 U19 ( .A(io_rand[2]), .B(io_b_0[4]), .Z(v_1_3_0[4]) );
  XOR2_X2 U20 ( .A(io_rand[2]), .B(io_b_0[3]), .Z(v_1_3_0[3]) );
  XOR2_X2 U21 ( .A(io_rand[2]), .B(io_b_0[2]), .Z(v_1_3_0[2]) );
  XOR2_X2 U22 ( .A(io_rand[2]), .B(io_b_0[1]), .Z(v_1_3_0[1]) );
  XOR2_X2 U23 ( .A(io_rand[2]), .B(io_b_0[0]), .Z(v_1_3_0[0]) );
  XOR2_X2 U25 ( .A(io_rand[5]), .B(io_b_3[5]), .Z(v_1_2_3[5]) );
  XOR2_X2 U26 ( .A(io_rand[5]), .B(io_b_3[4]), .Z(v_1_2_3[4]) );
  XOR2_X2 U27 ( .A(io_rand[5]), .B(io_b_3[3]), .Z(v_1_2_3[3]) );
  XOR2_X2 U28 ( .A(io_rand[5]), .B(io_b_3[2]), .Z(v_1_2_3[2]) );
  XOR2_X2 U29 ( .A(io_rand[5]), .B(io_b_3[1]), .Z(v_1_2_3[1]) );
  XOR2_X2 U30 ( .A(io_rand[5]), .B(io_b_3[0]), .Z(v_1_2_3[0]) );
  XOR2_X2 U32 ( .A(io_rand[3]), .B(io_b_1[5]), .Z(v_1_2_1[5]) );
  XOR2_X2 U33 ( .A(io_rand[3]), .B(io_b_1[4]), .Z(v_1_2_1[4]) );
  XOR2_X2 U34 ( .A(io_rand[3]), .B(io_b_1[3]), .Z(v_1_2_1[3]) );
  XOR2_X2 U35 ( .A(io_rand[3]), .B(io_b_1[2]), .Z(v_1_2_1[2]) );
  XOR2_X2 U36 ( .A(io_rand[3]), .B(io_b_1[1]), .Z(v_1_2_1[1]) );
  XOR2_X2 U37 ( .A(io_rand[3]), .B(io_b_1[0]), .Z(v_1_2_1[0]) );
  XOR2_X2 U39 ( .A(io_rand[1]), .B(io_b_0[5]), .Z(v_1_2_0[5]) );
  XOR2_X2 U40 ( .A(io_rand[1]), .B(io_b_0[4]), .Z(v_1_2_0[4]) );
  XOR2_X2 U41 ( .A(io_rand[1]), .B(io_b_0[3]), .Z(v_1_2_0[3]) );
  XOR2_X2 U42 ( .A(io_rand[1]), .B(io_b_0[2]), .Z(v_1_2_0[2]) );
  XOR2_X2 U43 ( .A(io_rand[1]), .B(io_b_0[1]), .Z(v_1_2_0[1]) );
  XOR2_X2 U44 ( .A(io_rand[1]), .B(io_b_0[0]), .Z(v_1_2_0[0]) );
  XOR2_X2 U46 ( .A(io_rand[4]), .B(io_b_3[5]), .Z(v_1_1_3[5]) );
  XOR2_X2 U47 ( .A(io_rand[4]), .B(io_b_3[4]), .Z(v_1_1_3[4]) );
  XOR2_X2 U48 ( .A(io_rand[4]), .B(io_b_3[3]), .Z(v_1_1_3[3]) );
  XOR2_X2 U49 ( .A(io_rand[4]), .B(io_b_3[2]), .Z(v_1_1_3[2]) );
  XOR2_X2 U50 ( .A(io_rand[4]), .B(io_b_3[1]), .Z(v_1_1_3[1]) );
  XOR2_X2 U51 ( .A(io_rand[4]), .B(io_b_3[0]), .Z(v_1_1_3[0]) );
  XOR2_X2 U53 ( .A(io_rand[3]), .B(io_b_2[5]), .Z(v_1_1_2[5]) );
  XOR2_X2 U54 ( .A(io_rand[3]), .B(io_b_2[4]), .Z(v_1_1_2[4]) );
  XOR2_X2 U55 ( .A(io_rand[3]), .B(io_b_2[3]), .Z(v_1_1_2[3]) );
  XOR2_X2 U56 ( .A(io_rand[3]), .B(io_b_2[2]), .Z(v_1_1_2[2]) );
  XOR2_X2 U57 ( .A(io_rand[3]), .B(io_b_2[1]), .Z(v_1_1_2[1]) );
  XOR2_X2 U58 ( .A(io_rand[3]), .B(io_b_2[0]), .Z(v_1_1_2[0]) );
  XOR2_X2 U60 ( .A(io_rand[0]), .B(io_b_0[5]), .Z(v_1_1_0[5]) );
  XOR2_X2 U61 ( .A(io_rand[0]), .B(io_b_0[4]), .Z(v_1_1_0[4]) );
  XOR2_X2 U62 ( .A(io_rand[0]), .B(io_b_0[3]), .Z(v_1_1_0[3]) );
  XOR2_X2 U63 ( .A(io_rand[0]), .B(io_b_0[2]), .Z(v_1_1_0[2]) );
  XOR2_X2 U64 ( .A(io_rand[0]), .B(io_b_0[1]), .Z(v_1_1_0[1]) );
  XOR2_X2 U65 ( .A(io_rand[0]), .B(io_b_0[0]), .Z(v_1_1_0[0]) );
  XOR2_X2 U67 ( .A(io_rand[2]), .B(io_b_3[5]), .Z(v_1_0_3[5]) );
  XOR2_X2 U68 ( .A(io_rand[2]), .B(io_b_3[4]), .Z(v_1_0_3[4]) );
  XOR2_X2 U69 ( .A(io_rand[2]), .B(io_b_3[3]), .Z(v_1_0_3[3]) );
  XOR2_X2 U70 ( .A(io_rand[2]), .B(io_b_3[2]), .Z(v_1_0_3[2]) );
  XOR2_X2 U71 ( .A(io_rand[2]), .B(io_b_3[1]), .Z(v_1_0_3[1]) );
  XOR2_X2 U72 ( .A(io_rand[2]), .B(io_b_3[0]), .Z(v_1_0_3[0]) );
  XOR2_X2 U74 ( .A(io_rand[1]), .B(io_b_2[5]), .Z(v_1_0_2[5]) );
  XOR2_X2 U75 ( .A(io_rand[1]), .B(io_b_2[4]), .Z(v_1_0_2[4]) );
  XOR2_X2 U76 ( .A(io_rand[1]), .B(io_b_2[3]), .Z(v_1_0_2[3]) );
  XOR2_X2 U77 ( .A(io_rand[1]), .B(io_b_2[2]), .Z(v_1_0_2[2]) );
  XOR2_X2 U78 ( .A(io_rand[1]), .B(io_b_2[1]), .Z(v_1_0_2[1]) );
  XOR2_X2 U79 ( .A(io_rand[1]), .B(io_b_2[0]), .Z(v_1_0_2[0]) );
  XOR2_X2 U81 ( .A(io_rand[0]), .B(io_b_1[5]), .Z(v_1_0_1[5]) );
  XOR2_X2 U82 ( .A(io_rand[0]), .B(io_b_1[4]), .Z(v_1_0_1[4]) );
  XOR2_X2 U83 ( .A(io_rand[0]), .B(io_b_1[3]), .Z(v_1_0_1[3]) );
  XOR2_X2 U84 ( .A(io_rand[0]), .B(io_b_1[2]), .Z(v_1_0_1[2]) );
  XOR2_X2 U85 ( .A(io_rand[0]), .B(io_b_1[1]), .Z(v_1_0_1[1]) );
  XOR2_X2 U86 ( .A(io_rand[0]), .B(io_b_1[0]), .Z(v_1_0_1[0]) );
  XOR2_X1 U367 ( .A(io_rand[5]), .B(io_b_2[6]), .Z(v_1_3_2[6]) );
  XOR2_X1 U368 ( .A(io_rand[4]), .B(io_b_1[6]), .Z(v_1_3_1[6]) );
  XOR2_X1 U369 ( .A(io_rand[2]), .B(io_b_0[6]), .Z(v_1_3_0[6]) );
  XOR2_X1 U370 ( .A(io_rand[5]), .B(io_b_3[6]), .Z(v_1_2_3[6]) );
  XOR2_X1 U371 ( .A(io_rand[3]), .B(io_b_1[6]), .Z(v_1_2_1[6]) );
  XOR2_X1 U372 ( .A(io_rand[1]), .B(io_b_0[6]), .Z(v_1_2_0[6]) );
  XOR2_X1 U373 ( .A(io_rand[4]), .B(io_b_3[6]), .Z(v_1_1_3[6]) );
  XOR2_X1 U374 ( .A(io_rand[3]), .B(io_b_2[6]), .Z(v_1_1_2[6]) );
  XOR2_X1 U375 ( .A(io_rand[0]), .B(io_b_0[6]), .Z(v_1_1_0[6]) );
  XOR2_X1 U376 ( .A(io_rand[2]), .B(io_b_3[6]), .Z(v_1_0_3[6]) );
  XOR2_X1 U377 ( .A(io_rand[1]), .B(io_b_2[6]), .Z(v_1_0_2[6]) );
  XOR2_X1 U378 ( .A(io_rand[0]), .B(io_b_1[6]), .Z(v_1_0_1[6]) );
  AND2_X1 U379 ( .A1(b_reg_0[0]), .A2(io_a_0[0]), .ZN(N84) );
  AND2_X1 U380 ( .A1(cor_port_v_0_1[0]), .A2(io_a_0[0]), .ZN(N85) );
  AND2_X1 U381 ( .A1(cor_port_v_0_2[0]), .A2(io_a_0[0]), .ZN(N86) );
  AND2_X1 U382 ( .A1(b_reg_1[0]), .A2(io_a_1[0]), .ZN(N88) );
  AND2_X1 U383 ( .A1(cor_port_v_1_0[0]), .A2(io_a_1[0]), .ZN(N89) );
  AND2_X1 U384 ( .A1(cor_port_v_1_2[0]), .A2(io_a_1[0]), .ZN(N90) );
  AND2_X1 U385 ( .A1(b_reg_2[0]), .A2(io_a_2[0]), .ZN(N92) );
  AND2_X1 U386 ( .A1(cor_port_v_2_0[0]), .A2(io_a_2[0]), .ZN(N93) );
  AND2_X1 U387 ( .A1(cor_port_v_2_1[0]), .A2(io_a_2[0]), .ZN(N94) );
  AND2_X1 U388 ( .A1(b_reg_3[0]), .A2(io_a_3[0]), .ZN(N96) );
  AND2_X1 U389 ( .A1(cor_port_v_3_0[0]), .A2(io_a_3[0]), .ZN(N97) );
  AND2_X1 U390 ( .A1(cor_port_v_3_1[0]), .A2(io_a_3[0]), .ZN(N98) );
  AND2_X1 U391 ( .A1(b_reg_0[1]), .A2(io_a_0[1]), .ZN(N100) );
  AND2_X1 U392 ( .A1(cor_port_v_0_1[1]), .A2(io_a_0[1]), .ZN(N101) );
  AND2_X1 U393 ( .A1(cor_port_v_0_2[1]), .A2(io_a_0[1]), .ZN(N102) );
  AND2_X1 U394 ( .A1(b_reg_1[1]), .A2(io_a_1[1]), .ZN(N104) );
  AND2_X1 U395 ( .A1(cor_port_v_1_0[1]), .A2(io_a_1[1]), .ZN(N105) );
  AND2_X1 U396 ( .A1(cor_port_v_1_2[1]), .A2(io_a_1[1]), .ZN(N106) );
  AND2_X1 U397 ( .A1(b_reg_2[1]), .A2(io_a_2[1]), .ZN(N108) );
  AND2_X1 U398 ( .A1(cor_port_v_2_0[1]), .A2(io_a_2[1]), .ZN(N109) );
  AND2_X1 U399 ( .A1(cor_port_v_2_1[1]), .A2(io_a_2[1]), .ZN(N110) );
  AND2_X1 U400 ( .A1(b_reg_3[1]), .A2(io_a_3[1]), .ZN(N112) );
  AND2_X1 U401 ( .A1(cor_port_v_3_0[1]), .A2(io_a_3[1]), .ZN(N113) );
  AND2_X1 U402 ( .A1(cor_port_v_3_1[1]), .A2(io_a_3[1]), .ZN(N114) );
  AND2_X1 U403 ( .A1(b_reg_0[2]), .A2(io_a_0[2]), .ZN(N116) );
  AND2_X1 U404 ( .A1(cor_port_v_0_1[2]), .A2(io_a_0[2]), .ZN(N117) );
  AND2_X1 U405 ( .A1(cor_port_v_0_2[2]), .A2(io_a_0[2]), .ZN(N118) );
  AND2_X1 U406 ( .A1(b_reg_0[3]), .A2(io_a_0[3]), .ZN(N132) );
  AND2_X1 U407 ( .A1(b_reg_0[4]), .A2(io_a_0[4]), .ZN(N148) );
  AND2_X1 U408 ( .A1(b_reg_0[5]), .A2(io_a_0[5]), .ZN(N164) );
  AND2_X1 U409 ( .A1(b_reg_0[6]), .A2(io_a_0[6]), .ZN(N180) );
  AND2_X1 U410 ( .A1(b_reg_1[2]), .A2(io_a_1[2]), .ZN(N120) );
  AND2_X1 U411 ( .A1(cor_port_v_1_0[2]), .A2(io_a_1[2]), .ZN(N121) );
  AND2_X1 U412 ( .A1(cor_port_v_1_2[2]), .A2(io_a_1[2]), .ZN(N122) );
  AND2_X1 U413 ( .A1(b_reg_2[2]), .A2(io_a_2[2]), .ZN(N124) );
  AND2_X1 U414 ( .A1(cor_port_v_2_0[2]), .A2(io_a_2[2]), .ZN(N125) );
  AND2_X1 U415 ( .A1(cor_port_v_2_1[2]), .A2(io_a_2[2]), .ZN(N126) );
  AND2_X1 U416 ( .A1(b_reg_3[2]), .A2(io_a_3[2]), .ZN(N128) );
  AND2_X1 U417 ( .A1(cor_port_v_3_0[2]), .A2(io_a_3[2]), .ZN(N129) );
  AND2_X1 U418 ( .A1(cor_port_v_3_1[2]), .A2(io_a_3[2]), .ZN(N130) );
  AND2_X1 U419 ( .A1(cor_port_v_0_1[3]), .A2(io_a_0[3]), .ZN(N133) );
  AND2_X1 U420 ( .A1(cor_port_v_0_2[3]), .A2(io_a_0[3]), .ZN(N134) );
  AND2_X1 U421 ( .A1(b_reg_1[3]), .A2(io_a_1[3]), .ZN(N136) );
  AND2_X1 U422 ( .A1(cor_port_v_1_0[3]), .A2(io_a_1[3]), .ZN(N137) );
  AND2_X1 U423 ( .A1(cor_port_v_1_2[3]), .A2(io_a_1[3]), .ZN(N138) );
  AND2_X1 U424 ( .A1(b_reg_2[3]), .A2(io_a_2[3]), .ZN(N140) );
  AND2_X1 U425 ( .A1(cor_port_v_2_0[3]), .A2(io_a_2[3]), .ZN(N141) );
  AND2_X1 U426 ( .A1(cor_port_v_2_1[3]), .A2(io_a_2[3]), .ZN(N142) );
  AND2_X1 U427 ( .A1(b_reg_3[3]), .A2(io_a_3[3]), .ZN(N144) );
  AND2_X1 U428 ( .A1(cor_port_v_3_0[3]), .A2(io_a_3[3]), .ZN(N145) );
  AND2_X1 U429 ( .A1(cor_port_v_3_1[3]), .A2(io_a_3[3]), .ZN(N146) );
  AND2_X1 U430 ( .A1(cor_port_v_0_1[4]), .A2(io_a_0[4]), .ZN(N149) );
  AND2_X1 U431 ( .A1(cor_port_v_0_2[4]), .A2(io_a_0[4]), .ZN(N150) );
  AND2_X1 U432 ( .A1(b_reg_1[4]), .A2(io_a_1[4]), .ZN(N152) );
  AND2_X1 U433 ( .A1(cor_port_v_1_0[4]), .A2(io_a_1[4]), .ZN(N153) );
  AND2_X1 U434 ( .A1(cor_port_v_1_2[4]), .A2(io_a_1[4]), .ZN(N154) );
  AND2_X1 U435 ( .A1(b_reg_2[4]), .A2(io_a_2[4]), .ZN(N156) );
  AND2_X1 U436 ( .A1(cor_port_v_2_0[4]), .A2(io_a_2[4]), .ZN(N157) );
  AND2_X1 U437 ( .A1(cor_port_v_2_1[4]), .A2(io_a_2[4]), .ZN(N158) );
  AND2_X1 U438 ( .A1(b_reg_3[4]), .A2(io_a_3[4]), .ZN(N160) );
  AND2_X1 U439 ( .A1(cor_port_v_3_0[4]), .A2(io_a_3[4]), .ZN(N161) );
  AND2_X1 U440 ( .A1(cor_port_v_3_1[4]), .A2(io_a_3[4]), .ZN(N162) );
  AND2_X1 U441 ( .A1(cor_port_v_0_1[5]), .A2(io_a_0[5]), .ZN(N165) );
  AND2_X1 U442 ( .A1(cor_port_v_0_2[5]), .A2(io_a_0[5]), .ZN(N166) );
  AND2_X1 U443 ( .A1(b_reg_1[5]), .A2(io_a_1[5]), .ZN(N168) );
  AND2_X1 U444 ( .A1(cor_port_v_1_0[5]), .A2(io_a_1[5]), .ZN(N169) );
  AND2_X1 U445 ( .A1(cor_port_v_1_2[5]), .A2(io_a_1[5]), .ZN(N170) );
  AND2_X1 U446 ( .A1(b_reg_2[5]), .A2(io_a_2[5]), .ZN(N172) );
  AND2_X1 U447 ( .A1(cor_port_v_2_0[5]), .A2(io_a_2[5]), .ZN(N173) );
  AND2_X1 U448 ( .A1(cor_port_v_2_1[5]), .A2(io_a_2[5]), .ZN(N174) );
  AND2_X1 U449 ( .A1(b_reg_3[5]), .A2(io_a_3[5]), .ZN(N176) );
  AND2_X1 U450 ( .A1(cor_port_v_3_0[5]), .A2(io_a_3[5]), .ZN(N177) );
  AND2_X1 U451 ( .A1(cor_port_v_3_1[5]), .A2(io_a_3[5]), .ZN(N178) );
  AND2_X1 U452 ( .A1(cor_port_v_0_1[6]), .A2(io_a_0[6]), .ZN(N181) );
  AND2_X1 U453 ( .A1(cor_port_v_0_2[6]), .A2(io_a_0[6]), .ZN(N182) );
  AND2_X1 U454 ( .A1(b_reg_1[6]), .A2(io_a_1[6]), .ZN(N184) );
  AND2_X1 U455 ( .A1(cor_port_v_1_0[6]), .A2(io_a_1[6]), .ZN(N185) );
  AND2_X1 U456 ( .A1(cor_port_v_1_2[6]), .A2(io_a_1[6]), .ZN(N186) );
  AND2_X1 U457 ( .A1(b_reg_2[6]), .A2(io_a_2[6]), .ZN(N188) );
  AND2_X1 U458 ( .A1(cor_port_v_2_0[6]), .A2(io_a_2[6]), .ZN(N189) );
  AND2_X1 U459 ( .A1(cor_port_v_2_1[6]), .A2(io_a_2[6]), .ZN(N190) );
  AND2_X1 U460 ( .A1(b_reg_3[6]), .A2(io_a_3[6]), .ZN(N192) );
  AND2_X1 U461 ( .A1(cor_port_v_3_0[6]), .A2(io_a_3[6]), .ZN(N193) );
  AND2_X1 U462 ( .A1(cor_port_v_3_1[6]), .A2(io_a_3[6]), .ZN(N194) );
  AND2_X1 U463 ( .A1(simpleNot_93_port_z), .A2(rand_reg_8[0]), .ZN(N9) );
  AND2_X1 U464 ( .A1(simpleNot_105_port_z), .A2(rand_reg_8[1]), .ZN(N21) );
  AND2_X1 U465 ( .A1(simpleNot_117_port_z), .A2(rand_reg_8[2]), .ZN(N33) );
  AND2_X1 U466 ( .A1(simpleNot_129_port_z), .A2(rand_reg_8[3]), .ZN(N45) );
  AND2_X1 U467 ( .A1(simpleNot_141_port_z), .A2(rand_reg_8[4]), .ZN(N57) );
  AND2_X1 U468 ( .A1(simpleNot_153_port_z), .A2(rand_reg_8[5]), .ZN(N69) );
  AND2_X1 U469 ( .A1(simpleNot_165_port_z), .A2(rand_reg_8[6]), .ZN(N81) );
  AND2_X1 U470 ( .A1(simpleNot_94_port_z), .A2(rand_reg_10[0]), .ZN(N10) );
  AND2_X1 U471 ( .A1(simpleNot_106_port_z), .A2(rand_reg_10[1]), .ZN(N22) );
  AND2_X1 U472 ( .A1(simpleNot_118_port_z), .A2(rand_reg_10[2]), .ZN(N34) );
  AND2_X1 U473 ( .A1(simpleNot_130_port_z), .A2(rand_reg_10[3]), .ZN(N46) );
  AND2_X1 U474 ( .A1(simpleNot_142_port_z), .A2(rand_reg_10[4]), .ZN(N58) );
  AND2_X1 U475 ( .A1(simpleNot_154_port_z), .A2(rand_reg_10[5]), .ZN(N70) );
  AND2_X1 U476 ( .A1(simpleNot_166_port_z), .A2(rand_reg_10[6]), .ZN(N82) );
  AND2_X1 U477 ( .A1(simpleNot_95_port_z), .A2(rand_reg_11[0]), .ZN(N11) );
  AND2_X1 U478 ( .A1(simpleNot_107_port_z), .A2(rand_reg_11[1]), .ZN(N23) );
  AND2_X1 U479 ( .A1(simpleNot_119_port_z), .A2(rand_reg_11[2]), .ZN(N35) );
  AND2_X1 U480 ( .A1(simpleNot_131_port_z), .A2(rand_reg_11[3]), .ZN(N47) );
  AND2_X1 U481 ( .A1(simpleNot_143_port_z), .A2(rand_reg_11[4]), .ZN(N59) );
  AND2_X1 U482 ( .A1(simpleNot_155_port_z), .A2(rand_reg_11[5]), .ZN(N71) );
  AND2_X1 U483 ( .A1(simpleNot_167_port_z), .A2(rand_reg_11[6]), .ZN(N83) );
  AND2_X1 U484 ( .A1(io_a_0[0]), .A2(cor_port_v_0_3[0]), .ZN(N87) );
  AND2_X1 U485 ( .A1(io_a_1[0]), .A2(cor_port_v_1_3[0]), .ZN(N91) );
  AND2_X1 U486 ( .A1(io_a_2[0]), .A2(cor_port_v_2_3[0]), .ZN(N95) );
  AND2_X1 U487 ( .A1(io_a_3[0]), .A2(cor_port_v_3_2[0]), .ZN(N99) );
  AND2_X1 U488 ( .A1(io_a_0[1]), .A2(cor_port_v_0_3[1]), .ZN(N103) );
  AND2_X1 U489 ( .A1(io_a_1[1]), .A2(cor_port_v_1_3[1]), .ZN(N107) );
  AND2_X1 U490 ( .A1(io_a_2[1]), .A2(cor_port_v_2_3[1]), .ZN(N111) );
  AND2_X1 U491 ( .A1(io_a_3[1]), .A2(cor_port_v_3_2[1]), .ZN(N115) );
  AND2_X1 U492 ( .A1(io_a_0[2]), .A2(cor_port_v_0_3[2]), .ZN(N119) );
  AND2_X1 U493 ( .A1(simpleNot_89_port_z), .A2(rand_reg_4[0]), .ZN(N5) );
  AND2_X1 U494 ( .A1(simpleNot_101_port_z), .A2(rand_reg_4[1]), .ZN(N17) );
  AND2_X1 U495 ( .A1(simpleNot_113_port_z), .A2(rand_reg_4[2]), .ZN(N29) );
  AND2_X1 U496 ( .A1(simpleNot_125_port_z), .A2(rand_reg_4[3]), .ZN(N41) );
  AND2_X1 U497 ( .A1(simpleNot_137_port_z), .A2(rand_reg_4[4]), .ZN(N53) );
  AND2_X1 U498 ( .A1(simpleNot_149_port_z), .A2(rand_reg_4[5]), .ZN(N65) );
  AND2_X1 U499 ( .A1(simpleNot_161_port_z), .A2(rand_reg_4[6]), .ZN(N77) );
  AND2_X1 U500 ( .A1(simpleNot_92_port_z), .A2(rand_reg_5[0]), .ZN(N8) );
  AND2_X1 U501 ( .A1(simpleNot_104_port_z), .A2(rand_reg_5[1]), .ZN(N20) );
  AND2_X1 U502 ( .A1(simpleNot_116_port_z), .A2(rand_reg_5[2]), .ZN(N32) );
  AND2_X1 U503 ( .A1(simpleNot_128_port_z), .A2(rand_reg_5[3]), .ZN(N44) );
  AND2_X1 U504 ( .A1(simpleNot_140_port_z), .A2(rand_reg_5[4]), .ZN(N56) );
  AND2_X1 U505 ( .A1(simpleNot_152_port_z), .A2(rand_reg_5[5]), .ZN(N68) );
  AND2_X1 U506 ( .A1(simpleNot_164_port_z), .A2(rand_reg_5[6]), .ZN(N80) );
  AND2_X1 U507 ( .A1(io_a_1[2]), .A2(cor_port_v_1_3[2]), .ZN(N123) );
  AND2_X1 U508 ( .A1(simpleNot_88_port_z), .A2(rand_reg_3[0]), .ZN(N4) );
  AND2_X1 U509 ( .A1(simpleNot_100_port_z), .A2(rand_reg_3[1]), .ZN(N16) );
  AND2_X1 U510 ( .A1(simpleNot_112_port_z), .A2(rand_reg_3[2]), .ZN(N28) );
  AND2_X1 U511 ( .A1(simpleNot_124_port_z), .A2(rand_reg_3[3]), .ZN(N40) );
  AND2_X1 U512 ( .A1(simpleNot_136_port_z), .A2(rand_reg_3[4]), .ZN(N52) );
  AND2_X1 U513 ( .A1(simpleNot_148_port_z), .A2(rand_reg_3[5]), .ZN(N64) );
  AND2_X1 U514 ( .A1(simpleNot_160_port_z), .A2(rand_reg_3[6]), .ZN(N76) );
  AND2_X1 U515 ( .A1(simpleNot_86_port_z), .A2(rand_reg_2[0]), .ZN(N2) );
  AND2_X1 U516 ( .A1(simpleNot_98_port_z), .A2(rand_reg_2[1]), .ZN(N14) );
  AND2_X1 U517 ( .A1(simpleNot_110_port_z), .A2(rand_reg_2[2]), .ZN(N26) );
  AND2_X1 U518 ( .A1(simpleNot_122_port_z), .A2(rand_reg_2[3]), .ZN(N38) );
  AND2_X1 U519 ( .A1(simpleNot_134_port_z), .A2(rand_reg_2[4]), .ZN(N50) );
  AND2_X1 U520 ( .A1(simpleNot_146_port_z), .A2(rand_reg_2[5]), .ZN(N62) );
  AND2_X1 U521 ( .A1(simpleNot_158_port_z), .A2(rand_reg_2[6]), .ZN(N74) );
  AND2_X1 U522 ( .A1(io_a_2[2]), .A2(cor_port_v_2_3[2]), .ZN(N127) );
  AND2_X1 U523 ( .A1(simpleNot_84_port_z), .A2(rand_reg_0[0]), .ZN(N0) );
  AND2_X1 U524 ( .A1(simpleNot_96_port_z), .A2(rand_reg_0[1]), .ZN(N12) );
  AND2_X1 U525 ( .A1(simpleNot_108_port_z), .A2(rand_reg_0[2]), .ZN(N24) );
  AND2_X1 U526 ( .A1(simpleNot_120_port_z), .A2(rand_reg_0[3]), .ZN(N36) );
  AND2_X1 U527 ( .A1(simpleNot_132_port_z), .A2(rand_reg_0[4]), .ZN(N48) );
  AND2_X1 U528 ( .A1(simpleNot_144_port_z), .A2(rand_reg_0[5]), .ZN(N60) );
  AND2_X1 U529 ( .A1(simpleNot_156_port_z), .A2(rand_reg_0[6]), .ZN(N72) );
  AND2_X1 U530 ( .A1(simpleNot_90_port_z), .A2(rand_reg_7[0]), .ZN(N6) );
  AND2_X1 U531 ( .A1(simpleNot_102_port_z), .A2(rand_reg_7[1]), .ZN(N18) );
  AND2_X1 U532 ( .A1(simpleNot_114_port_z), .A2(rand_reg_7[2]), .ZN(N30) );
  AND2_X1 U533 ( .A1(simpleNot_126_port_z), .A2(rand_reg_7[3]), .ZN(N42) );
  AND2_X1 U534 ( .A1(simpleNot_138_port_z), .A2(rand_reg_7[4]), .ZN(N54) );
  AND2_X1 U535 ( .A1(simpleNot_150_port_z), .A2(rand_reg_7[5]), .ZN(N66) );
  AND2_X1 U536 ( .A1(simpleNot_162_port_z), .A2(rand_reg_7[6]), .ZN(N78) );
  AND2_X1 U537 ( .A1(simpleNot_87_port_z), .A2(rand_reg_6[0]), .ZN(N3) );
  AND2_X1 U538 ( .A1(simpleNot_99_port_z), .A2(rand_reg_6[1]), .ZN(N15) );
  AND2_X1 U539 ( .A1(simpleNot_111_port_z), .A2(rand_reg_6[2]), .ZN(N27) );
  AND2_X1 U540 ( .A1(simpleNot_123_port_z), .A2(rand_reg_6[3]), .ZN(N39) );
  AND2_X1 U541 ( .A1(simpleNot_135_port_z), .A2(rand_reg_6[4]), .ZN(N51) );
  AND2_X1 U542 ( .A1(simpleNot_147_port_z), .A2(rand_reg_6[5]), .ZN(N63) );
  AND2_X1 U543 ( .A1(simpleNot_159_port_z), .A2(rand_reg_6[6]), .ZN(N75) );
  AND2_X1 U544 ( .A1(io_a_3[2]), .A2(cor_port_v_3_2[2]), .ZN(N131) );
  AND2_X1 U545 ( .A1(simpleNot_85_port_z), .A2(rand_reg_1[0]), .ZN(N1) );
  AND2_X1 U546 ( .A1(simpleNot_97_port_z), .A2(rand_reg_1[1]), .ZN(N13) );
  AND2_X1 U547 ( .A1(simpleNot_109_port_z), .A2(rand_reg_1[2]), .ZN(N25) );
  AND2_X1 U548 ( .A1(simpleNot_121_port_z), .A2(rand_reg_1[3]), .ZN(N37) );
  AND2_X1 U549 ( .A1(simpleNot_133_port_z), .A2(rand_reg_1[4]), .ZN(N49) );
  AND2_X1 U550 ( .A1(simpleNot_145_port_z), .A2(rand_reg_1[5]), .ZN(N61) );
  AND2_X1 U551 ( .A1(simpleNot_157_port_z), .A2(rand_reg_1[6]), .ZN(N73) );
  AND2_X1 U552 ( .A1(io_a_0[3]), .A2(cor_port_v_0_3[3]), .ZN(N135) );
  AND2_X1 U553 ( .A1(simpleNot_91_port_z), .A2(rand_reg_9[0]), .ZN(N7) );
  AND2_X1 U554 ( .A1(simpleNot_103_port_z), .A2(rand_reg_9[1]), .ZN(N19) );
  AND2_X1 U555 ( .A1(simpleNot_115_port_z), .A2(rand_reg_9[2]), .ZN(N31) );
  AND2_X1 U556 ( .A1(simpleNot_127_port_z), .A2(rand_reg_9[3]), .ZN(N43) );
  AND2_X1 U557 ( .A1(simpleNot_139_port_z), .A2(rand_reg_9[4]), .ZN(N55) );
  AND2_X1 U558 ( .A1(simpleNot_151_port_z), .A2(rand_reg_9[5]), .ZN(N67) );
  AND2_X1 U559 ( .A1(simpleNot_163_port_z), .A2(rand_reg_9[6]), .ZN(N79) );
  AND2_X1 U560 ( .A1(io_a_1[3]), .A2(cor_port_v_1_3[3]), .ZN(N139) );
  AND2_X1 U561 ( .A1(io_a_2[3]), .A2(cor_port_v_2_3[3]), .ZN(N143) );
  AND2_X1 U562 ( .A1(io_a_3[3]), .A2(cor_port_v_3_2[3]), .ZN(N147) );
  AND2_X1 U563 ( .A1(io_a_0[4]), .A2(cor_port_v_0_3[4]), .ZN(N151) );
  AND2_X1 U564 ( .A1(io_a_1[4]), .A2(cor_port_v_1_3[4]), .ZN(N155) );
  AND2_X1 U565 ( .A1(io_a_2[4]), .A2(cor_port_v_2_3[4]), .ZN(N159) );
  AND2_X1 U566 ( .A1(io_a_3[4]), .A2(cor_port_v_3_2[4]), .ZN(N163) );
  AND2_X1 U567 ( .A1(io_a_0[5]), .A2(cor_port_v_0_3[5]), .ZN(N167) );
  AND2_X1 U568 ( .A1(io_a_1[5]), .A2(cor_port_v_1_3[5]), .ZN(N171) );
  AND2_X1 U569 ( .A1(io_a_2[5]), .A2(cor_port_v_2_3[5]), .ZN(N175) );
  AND2_X1 U570 ( .A1(io_a_3[5]), .A2(cor_port_v_3_2[5]), .ZN(N179) );
  AND2_X1 U571 ( .A1(io_a_0[6]), .A2(cor_port_v_0_3[6]), .ZN(N183) );
  AND2_X1 U572 ( .A1(io_a_1[6]), .A2(cor_port_v_1_3[6]), .ZN(N187) );
  AND2_X1 U573 ( .A1(io_a_2[6]), .A2(cor_port_v_2_3[6]), .ZN(N191) );
  AND2_X1 U574 ( .A1(io_a_3[6]), .A2(cor_port_v_3_2[6]), .ZN(N195) );
  XOR2_X1 U575 ( .A(n13), .B(n14), .Z(io_c_3[0]) );
  XNOR2_X1 U576 ( .A(simpleXor_95_port_z), .B(simpleXor_94_port_z), .ZN(n13)
         );
  XNOR2_X1 U577 ( .A(simpleXor_93_port_z), .B(n_zz_io_c_3_0_), .ZN(n14) );
  XOR2_X1 U578 ( .A(n11), .B(n12), .Z(io_c_3[1]) );
  XNOR2_X1 U579 ( .A(simpleXor_107_port_z), .B(simpleXor_106_port_z), .ZN(n11)
         );
  XNOR2_X1 U580 ( .A(simpleXor_105_port_z), .B(n_zz_io_c_3_5_0_), .ZN(n12) );
  XOR2_X1 U581 ( .A(n9), .B(n10), .Z(io_c_3[2]) );
  XNOR2_X1 U582 ( .A(simpleXor_119_port_z), .B(simpleXor_118_port_z), .ZN(n9)
         );
  XNOR2_X1 U583 ( .A(simpleXor_117_port_z), .B(n_zz_io_c_3_10_0_), .ZN(n10) );
  XOR2_X1 U584 ( .A(n7), .B(n8), .Z(io_c_3[3]) );
  XNOR2_X1 U585 ( .A(simpleXor_131_port_z), .B(simpleXor_130_port_z), .ZN(n7)
         );
  XNOR2_X1 U586 ( .A(simpleXor_129_port_z), .B(n_zz_io_c_3_15_0_), .ZN(n8) );
  XOR2_X1 U587 ( .A(n5), .B(n6), .Z(io_c_3[4]) );
  XNOR2_X1 U588 ( .A(simpleXor_143_port_z), .B(simpleXor_142_port_z), .ZN(n5)
         );
  XNOR2_X1 U589 ( .A(simpleXor_141_port_z), .B(n_zz_io_c_3_20_0_), .ZN(n6) );
  XOR2_X1 U590 ( .A(n3), .B(n4), .Z(io_c_3[5]) );
  XNOR2_X1 U591 ( .A(simpleXor_155_port_z), .B(simpleXor_154_port_z), .ZN(n3)
         );
  XNOR2_X1 U592 ( .A(simpleXor_153_port_z), .B(n_zz_io_c_3_25_0_), .ZN(n4) );
  XOR2_X1 U593 ( .A(n1), .B(n2), .Z(io_c_3[6]) );
  XNOR2_X1 U594 ( .A(simpleXor_167_port_z), .B(simpleXor_166_port_z), .ZN(n1)
         );
  XNOR2_X1 U595 ( .A(simpleXor_165_port_z), .B(n_zz_io_c_3_30_0_), .ZN(n2) );
  XOR2_X1 U596 ( .A(n27), .B(n28), .Z(io_c_2[0]) );
  XNOR2_X1 U597 ( .A(simpleXor_92_port_z), .B(simpleXor_91_port_z), .ZN(n27)
         );
  XNOR2_X1 U598 ( .A(simpleXor_90_port_z), .B(n_zz_io_c_2_0_), .ZN(n28) );
  XOR2_X1 U599 ( .A(n25), .B(n26), .Z(io_c_2[1]) );
  XNOR2_X1 U600 ( .A(simpleXor_104_port_z), .B(simpleXor_103_port_z), .ZN(n25)
         );
  XNOR2_X1 U601 ( .A(simpleXor_102_port_z), .B(n_zz_io_c_2_5_0_), .ZN(n26) );
  XOR2_X1 U602 ( .A(n23), .B(n24), .Z(io_c_2[2]) );
  XNOR2_X1 U603 ( .A(simpleXor_116_port_z), .B(simpleXor_115_port_z), .ZN(n23)
         );
  XNOR2_X1 U604 ( .A(simpleXor_114_port_z), .B(n_zz_io_c_2_10_0_), .ZN(n24) );
  XOR2_X1 U605 ( .A(n21), .B(n22), .Z(io_c_2[3]) );
  XNOR2_X1 U606 ( .A(simpleXor_128_port_z), .B(simpleXor_127_port_z), .ZN(n21)
         );
  XNOR2_X1 U607 ( .A(simpleXor_126_port_z), .B(n_zz_io_c_2_15_0_), .ZN(n22) );
  XOR2_X1 U608 ( .A(n19), .B(n20), .Z(io_c_2[4]) );
  XNOR2_X1 U609 ( .A(simpleXor_140_port_z), .B(simpleXor_139_port_z), .ZN(n19)
         );
  XNOR2_X1 U610 ( .A(simpleXor_138_port_z), .B(n_zz_io_c_2_20_0_), .ZN(n20) );
  XOR2_X1 U611 ( .A(n17), .B(n18), .Z(io_c_2[5]) );
  XNOR2_X1 U612 ( .A(simpleXor_152_port_z), .B(simpleXor_151_port_z), .ZN(n17)
         );
  XNOR2_X1 U613 ( .A(simpleXor_150_port_z), .B(n_zz_io_c_2_25_0_), .ZN(n18) );
  XOR2_X1 U614 ( .A(n15), .B(n16), .Z(io_c_2[6]) );
  XNOR2_X1 U615 ( .A(simpleXor_164_port_z), .B(simpleXor_163_port_z), .ZN(n15)
         );
  XNOR2_X1 U616 ( .A(simpleXor_162_port_z), .B(n_zz_io_c_2_30_0_), .ZN(n16) );
  XOR2_X1 U617 ( .A(n41), .B(n42), .Z(io_c_1[0]) );
  XNOR2_X1 U618 ( .A(simpleXor_89_port_z), .B(simpleXor_88_port_z), .ZN(n41)
         );
  XNOR2_X1 U619 ( .A(simpleXor_87_port_z), .B(n_zz_io_c_1_0_), .ZN(n42) );
  XOR2_X1 U620 ( .A(n39), .B(n40), .Z(io_c_1[1]) );
  XNOR2_X1 U621 ( .A(simpleXor_99_port_z), .B(simpleXor_101_port_z), .ZN(n39)
         );
  XNOR2_X1 U622 ( .A(simpleXor_100_port_z), .B(n_zz_io_c_1_5_0_), .ZN(n40) );
  XOR2_X1 U623 ( .A(n37), .B(n38), .Z(io_c_1[2]) );
  XNOR2_X1 U624 ( .A(simpleXor_113_port_z), .B(simpleXor_112_port_z), .ZN(n37)
         );
  XNOR2_X1 U625 ( .A(simpleXor_111_port_z), .B(n_zz_io_c_1_10_0_), .ZN(n38) );
  XOR2_X1 U626 ( .A(n35), .B(n36), .Z(io_c_1[3]) );
  XNOR2_X1 U627 ( .A(simpleXor_125_port_z), .B(simpleXor_124_port_z), .ZN(n35)
         );
  XNOR2_X1 U628 ( .A(simpleXor_123_port_z), .B(n_zz_io_c_1_15_0_), .ZN(n36) );
  XOR2_X1 U629 ( .A(n33), .B(n34), .Z(io_c_1[4]) );
  XNOR2_X1 U630 ( .A(simpleXor_137_port_z), .B(simpleXor_136_port_z), .ZN(n33)
         );
  XNOR2_X1 U631 ( .A(simpleXor_135_port_z), .B(n_zz_io_c_1_20_0_), .ZN(n34) );
  XOR2_X1 U632 ( .A(n31), .B(n32), .Z(io_c_1[5]) );
  XNOR2_X1 U633 ( .A(simpleXor_149_port_z), .B(simpleXor_148_port_z), .ZN(n31)
         );
  XNOR2_X1 U634 ( .A(simpleXor_147_port_z), .B(n_zz_io_c_1_25_0_), .ZN(n32) );
  XOR2_X1 U635 ( .A(n29), .B(n30), .Z(io_c_1[6]) );
  XNOR2_X1 U636 ( .A(simpleXor_161_port_z), .B(simpleXor_160_port_z), .ZN(n29)
         );
  XNOR2_X1 U637 ( .A(simpleXor_159_port_z), .B(n_zz_io_c_1_30_0_), .ZN(n30) );
  XOR2_X1 U638 ( .A(n55), .B(n56), .Z(io_c_0[0]) );
  XNOR2_X1 U639 ( .A(simpleXor_86_port_z), .B(simpleXor_85_port_z), .ZN(n55)
         );
  XNOR2_X1 U640 ( .A(simpleXor_84_port_z), .B(n_zz_io_c_0_0_), .ZN(n56) );
  XOR2_X1 U641 ( .A(n53), .B(n54), .Z(io_c_0[1]) );
  XNOR2_X1 U642 ( .A(simpleXor_98_port_z), .B(simpleXor_97_port_z), .ZN(n53)
         );
  XNOR2_X1 U643 ( .A(simpleXor_96_port_z), .B(n_zz_io_c_0_5_0_), .ZN(n54) );
  XOR2_X1 U644 ( .A(n51), .B(n52), .Z(io_c_0[2]) );
  XNOR2_X1 U645 ( .A(simpleXor_110_port_z), .B(simpleXor_109_port_z), .ZN(n51)
         );
  XNOR2_X1 U646 ( .A(simpleXor_108_port_z), .B(n_zz_io_c_0_10_0_), .ZN(n52) );
  XOR2_X1 U647 ( .A(n49), .B(n50), .Z(io_c_0[3]) );
  XNOR2_X1 U648 ( .A(simpleXor_122_port_z), .B(simpleXor_121_port_z), .ZN(n49)
         );
  XNOR2_X1 U649 ( .A(simpleXor_120_port_z), .B(n_zz_io_c_0_15_0_), .ZN(n50) );
  XOR2_X1 U650 ( .A(n47), .B(n48), .Z(io_c_0[4]) );
  XNOR2_X1 U651 ( .A(simpleXor_134_port_z), .B(simpleXor_133_port_z), .ZN(n47)
         );
  XNOR2_X1 U652 ( .A(simpleXor_132_port_z), .B(n_zz_io_c_0_20_0_), .ZN(n48) );
  XOR2_X1 U653 ( .A(n45), .B(n46), .Z(io_c_0[5]) );
  XNOR2_X1 U654 ( .A(simpleXor_146_port_z), .B(simpleXor_145_port_z), .ZN(n45)
         );
  XNOR2_X1 U655 ( .A(simpleXor_144_port_z), .B(n_zz_io_c_0_25_0_), .ZN(n46) );
  XOR2_X1 U656 ( .A(n43), .B(n44), .Z(io_c_0[6]) );
  XNOR2_X1 U657 ( .A(simpleXor_158_port_z), .B(simpleXor_157_port_z), .ZN(n43)
         );
  XNOR2_X1 U658 ( .A(simpleXor_156_port_z), .B(n_zz_io_c_0_30_0_), .ZN(n44) );
  INV_X1 simpleNot_84_U1 ( .A(io_a_0[0]), .ZN(simpleNot_84_port_z) );
  INV_X1 simpleNot_85_U1 ( .A(io_a_0[0]), .ZN(simpleNot_85_port_z) );
  INV_X1 simpleNot_86_U1 ( .A(io_a_0[0]), .ZN(simpleNot_86_port_z) );
  INV_X1 simpleNot_87_U1 ( .A(io_a_1[0]), .ZN(simpleNot_87_port_z) );
  INV_X1 simpleNot_88_U1 ( .A(io_a_1[0]), .ZN(simpleNot_88_port_z) );
  INV_X1 simpleNot_89_U1 ( .A(io_a_1[0]), .ZN(simpleNot_89_port_z) );
  INV_X1 simpleNot_90_U1 ( .A(io_a_2[0]), .ZN(simpleNot_90_port_z) );
  INV_X1 simpleNot_91_U1 ( .A(io_a_2[0]), .ZN(simpleNot_91_port_z) );
  INV_X1 simpleNot_92_U1 ( .A(io_a_2[0]), .ZN(simpleNot_92_port_z) );
  INV_X1 simpleNot_93_U1 ( .A(io_a_3[0]), .ZN(simpleNot_93_port_z) );
  INV_X1 simpleNot_94_U1 ( .A(io_a_3[0]), .ZN(simpleNot_94_port_z) );
  INV_X1 simpleNot_95_U1 ( .A(io_a_3[0]), .ZN(simpleNot_95_port_z) );
  INV_X1 simpleNot_96_U1 ( .A(io_a_0[1]), .ZN(simpleNot_96_port_z) );
  INV_X1 simpleNot_97_U1 ( .A(io_a_0[1]), .ZN(simpleNot_97_port_z) );
  INV_X1 simpleNot_98_U1 ( .A(io_a_0[1]), .ZN(simpleNot_98_port_z) );
  INV_X1 simpleNot_99_U1 ( .A(io_a_1[1]), .ZN(simpleNot_99_port_z) );
  INV_X1 simpleNot_100_U1 ( .A(io_a_1[1]), .ZN(simpleNot_100_port_z) );
  INV_X1 simpleNot_101_U1 ( .A(io_a_1[1]), .ZN(simpleNot_101_port_z) );
  INV_X1 simpleNot_102_U1 ( .A(io_a_2[1]), .ZN(simpleNot_102_port_z) );
  INV_X1 simpleNot_103_U1 ( .A(io_a_2[1]), .ZN(simpleNot_103_port_z) );
  INV_X1 simpleNot_104_U1 ( .A(io_a_2[1]), .ZN(simpleNot_104_port_z) );
  INV_X1 simpleNot_105_U1 ( .A(io_a_3[1]), .ZN(simpleNot_105_port_z) );
  INV_X1 simpleNot_106_U1 ( .A(io_a_3[1]), .ZN(simpleNot_106_port_z) );
  INV_X1 simpleNot_107_U1 ( .A(io_a_3[1]), .ZN(simpleNot_107_port_z) );
  INV_X1 simpleNot_108_U1 ( .A(io_a_0[2]), .ZN(simpleNot_108_port_z) );
  INV_X1 simpleNot_109_U1 ( .A(io_a_0[2]), .ZN(simpleNot_109_port_z) );
  INV_X1 simpleNot_110_U1 ( .A(io_a_0[2]), .ZN(simpleNot_110_port_z) );
  INV_X1 simpleNot_111_U1 ( .A(io_a_1[2]), .ZN(simpleNot_111_port_z) );
  INV_X1 simpleNot_112_U1 ( .A(io_a_1[2]), .ZN(simpleNot_112_port_z) );
  INV_X1 simpleNot_113_U1 ( .A(io_a_1[2]), .ZN(simpleNot_113_port_z) );
  INV_X1 simpleNot_114_U1 ( .A(io_a_2[2]), .ZN(simpleNot_114_port_z) );
  INV_X1 simpleNot_115_U1 ( .A(io_a_2[2]), .ZN(simpleNot_115_port_z) );
  INV_X1 simpleNot_116_U1 ( .A(io_a_2[2]), .ZN(simpleNot_116_port_z) );
  INV_X1 simpleNot_117_U1 ( .A(io_a_3[2]), .ZN(simpleNot_117_port_z) );
  INV_X1 simpleNot_118_U1 ( .A(io_a_3[2]), .ZN(simpleNot_118_port_z) );
  INV_X1 simpleNot_119_U1 ( .A(io_a_3[2]), .ZN(simpleNot_119_port_z) );
  INV_X1 simpleNot_120_U1 ( .A(io_a_0[3]), .ZN(simpleNot_120_port_z) );
  INV_X1 simpleNot_121_U1 ( .A(io_a_0[3]), .ZN(simpleNot_121_port_z) );
  INV_X1 simpleNot_122_U1 ( .A(io_a_0[3]), .ZN(simpleNot_122_port_z) );
  INV_X1 simpleNot_123_U1 ( .A(io_a_1[3]), .ZN(simpleNot_123_port_z) );
  INV_X1 simpleNot_124_U1 ( .A(io_a_1[3]), .ZN(simpleNot_124_port_z) );
  INV_X1 simpleNot_125_U1 ( .A(io_a_1[3]), .ZN(simpleNot_125_port_z) );
  INV_X1 simpleNot_126_U1 ( .A(io_a_2[3]), .ZN(simpleNot_126_port_z) );
  INV_X1 simpleNot_127_U1 ( .A(io_a_2[3]), .ZN(simpleNot_127_port_z) );
  INV_X1 simpleNot_128_U1 ( .A(io_a_2[3]), .ZN(simpleNot_128_port_z) );
  INV_X1 simpleNot_129_U1 ( .A(io_a_3[3]), .ZN(simpleNot_129_port_z) );
  INV_X1 simpleNot_130_U1 ( .A(io_a_3[3]), .ZN(simpleNot_130_port_z) );
  INV_X1 simpleNot_131_U1 ( .A(io_a_3[3]), .ZN(simpleNot_131_port_z) );
  INV_X1 simpleNot_132_U1 ( .A(io_a_0[4]), .ZN(simpleNot_132_port_z) );
  INV_X1 simpleNot_133_U1 ( .A(io_a_0[4]), .ZN(simpleNot_133_port_z) );
  INV_X1 simpleNot_134_U1 ( .A(io_a_0[4]), .ZN(simpleNot_134_port_z) );
  INV_X1 simpleNot_135_U1 ( .A(io_a_1[4]), .ZN(simpleNot_135_port_z) );
  INV_X1 simpleNot_136_U1 ( .A(io_a_1[4]), .ZN(simpleNot_136_port_z) );
  INV_X1 simpleNot_137_U1 ( .A(io_a_1[4]), .ZN(simpleNot_137_port_z) );
  INV_X1 simpleNot_138_U1 ( .A(io_a_2[4]), .ZN(simpleNot_138_port_z) );
  INV_X1 simpleNot_139_U1 ( .A(io_a_2[4]), .ZN(simpleNot_139_port_z) );
  INV_X1 simpleNot_140_U1 ( .A(io_a_2[4]), .ZN(simpleNot_140_port_z) );
  INV_X1 simpleNot_141_U1 ( .A(io_a_3[4]), .ZN(simpleNot_141_port_z) );
  INV_X1 simpleNot_142_U1 ( .A(io_a_3[4]), .ZN(simpleNot_142_port_z) );
  INV_X1 simpleNot_143_U1 ( .A(io_a_3[4]), .ZN(simpleNot_143_port_z) );
  INV_X1 simpleNot_144_U1 ( .A(io_a_0[5]), .ZN(simpleNot_144_port_z) );
  INV_X1 simpleNot_145_U1 ( .A(io_a_0[5]), .ZN(simpleNot_145_port_z) );
  INV_X1 simpleNot_146_U1 ( .A(io_a_0[5]), .ZN(simpleNot_146_port_z) );
  INV_X1 simpleNot_147_U1 ( .A(io_a_1[5]), .ZN(simpleNot_147_port_z) );
  INV_X1 simpleNot_148_U1 ( .A(io_a_1[5]), .ZN(simpleNot_148_port_z) );
  INV_X1 simpleNot_149_U1 ( .A(io_a_1[5]), .ZN(simpleNot_149_port_z) );
  INV_X1 simpleNot_150_U1 ( .A(io_a_2[5]), .ZN(simpleNot_150_port_z) );
  INV_X1 simpleNot_151_U1 ( .A(io_a_2[5]), .ZN(simpleNot_151_port_z) );
  INV_X1 simpleNot_152_U1 ( .A(io_a_2[5]), .ZN(simpleNot_152_port_z) );
  INV_X1 simpleNot_153_U1 ( .A(io_a_3[5]), .ZN(simpleNot_153_port_z) );
  INV_X1 simpleNot_154_U1 ( .A(io_a_3[5]), .ZN(simpleNot_154_port_z) );
  INV_X1 simpleNot_155_U1 ( .A(io_a_3[5]), .ZN(simpleNot_155_port_z) );
  INV_X1 simpleNot_156_U1 ( .A(io_a_0[6]), .ZN(simpleNot_156_port_z) );
  INV_X1 simpleNot_157_U1 ( .A(io_a_0[6]), .ZN(simpleNot_157_port_z) );
  INV_X1 simpleNot_158_U1 ( .A(io_a_0[6]), .ZN(simpleNot_158_port_z) );
  INV_X1 simpleNot_159_U1 ( .A(io_a_1[6]), .ZN(simpleNot_159_port_z) );
  INV_X1 simpleNot_160_U1 ( .A(io_a_1[6]), .ZN(simpleNot_160_port_z) );
  INV_X1 simpleNot_161_U1 ( .A(io_a_1[6]), .ZN(simpleNot_161_port_z) );
  INV_X1 simpleNot_162_U1 ( .A(io_a_2[6]), .ZN(simpleNot_162_port_z) );
  INV_X1 simpleNot_163_U1 ( .A(io_a_2[6]), .ZN(simpleNot_163_port_z) );
  INV_X1 simpleNot_164_U1 ( .A(io_a_2[6]), .ZN(simpleNot_164_port_z) );
  INV_X1 simpleNot_165_U1 ( .A(io_a_3[6]), .ZN(simpleNot_165_port_z) );
  INV_X1 simpleNot_166_U1 ( .A(io_a_3[6]), .ZN(simpleNot_166_port_z) );
  INV_X1 simpleNot_167_U1 ( .A(io_a_3[6]), .ZN(simpleNot_167_port_z) );
  DFF_X1 cor_m_3_2_reg_0_ ( .D(cor_maj_161_port_o), .CK(clk), .Q(
        cor_port_v_3_2[0]), .QN() );
  DFF_X1 cor_m_3_2_reg_1_ ( .D(cor_maj_162_port_o), .CK(clk), .Q(
        cor_port_v_3_2[1]), .QN() );
  DFF_X1 cor_m_3_2_reg_2_ ( .D(cor_maj_163_port_o), .CK(clk), .Q(
        cor_port_v_3_2[2]), .QN() );
  DFF_X1 cor_m_3_2_reg_3_ ( .D(cor_maj_164_port_o), .CK(clk), .Q(
        cor_port_v_3_2[3]), .QN() );
  DFF_X1 cor_m_3_2_reg_4_ ( .D(cor_maj_165_port_o), .CK(clk), .Q(
        cor_port_v_3_2[4]), .QN() );
  DFF_X1 cor_m_3_2_reg_5_ ( .D(cor_maj_166_port_o), .CK(clk), .Q(
        cor_port_v_3_2[5]), .QN() );
  DFF_X1 cor_m_3_2_reg_6_ ( .D(cor_maj_167_port_o), .CK(clk), .Q(
        cor_port_v_3_2[6]), .QN() );
  DFF_X1 cor_m_3_1_reg_0_ ( .D(cor_maj_154_port_o), .CK(clk), .Q(
        cor_port_v_3_1[0]), .QN() );
  DFF_X1 cor_m_3_1_reg_1_ ( .D(cor_maj_155_port_o), .CK(clk), .Q(
        cor_port_v_3_1[1]), .QN() );
  DFF_X1 cor_m_3_1_reg_2_ ( .D(cor_maj_156_port_o), .CK(clk), .Q(
        cor_port_v_3_1[2]), .QN() );
  DFF_X1 cor_m_3_1_reg_3_ ( .D(cor_maj_157_port_o), .CK(clk), .Q(
        cor_port_v_3_1[3]), .QN() );
  DFF_X1 cor_m_3_1_reg_4_ ( .D(cor_maj_158_port_o), .CK(clk), .Q(
        cor_port_v_3_1[4]), .QN() );
  DFF_X1 cor_m_3_1_reg_5_ ( .D(cor_maj_159_port_o), .CK(clk), .Q(
        cor_port_v_3_1[5]), .QN() );
  DFF_X1 cor_m_3_1_reg_6_ ( .D(cor_maj_160_port_o), .CK(clk), .Q(
        cor_port_v_3_1[6]), .QN() );
  DFF_X1 cor_m_3_0_reg_0_ ( .D(cor_maj_147_port_o), .CK(clk), .Q(
        cor_port_v_3_0[0]), .QN() );
  DFF_X1 cor_m_3_0_reg_1_ ( .D(cor_maj_148_port_o), .CK(clk), .Q(
        cor_port_v_3_0[1]), .QN() );
  DFF_X1 cor_m_3_0_reg_2_ ( .D(cor_maj_149_port_o), .CK(clk), .Q(
        cor_port_v_3_0[2]), .QN() );
  DFF_X1 cor_m_3_0_reg_3_ ( .D(cor_maj_150_port_o), .CK(clk), .Q(
        cor_port_v_3_0[3]), .QN() );
  DFF_X1 cor_m_3_0_reg_4_ ( .D(cor_maj_151_port_o), .CK(clk), .Q(
        cor_port_v_3_0[4]), .QN() );
  DFF_X1 cor_m_3_0_reg_5_ ( .D(cor_maj_152_port_o), .CK(clk), .Q(
        cor_port_v_3_0[5]), .QN() );
  DFF_X1 cor_m_3_0_reg_6_ ( .D(cor_maj_153_port_o), .CK(clk), .Q(
        cor_port_v_3_0[6]), .QN() );
  DFF_X1 cor_m_2_3_reg_0_ ( .D(cor_maj_140_port_o), .CK(clk), .Q(
        cor_port_v_2_3[0]), .QN() );
  DFF_X1 cor_m_2_3_reg_1_ ( .D(cor_maj_141_port_o), .CK(clk), .Q(
        cor_port_v_2_3[1]), .QN() );
  DFF_X1 cor_m_2_3_reg_2_ ( .D(cor_maj_142_port_o), .CK(clk), .Q(
        cor_port_v_2_3[2]), .QN() );
  DFF_X1 cor_m_2_3_reg_3_ ( .D(cor_maj_143_port_o), .CK(clk), .Q(
        cor_port_v_2_3[3]), .QN() );
  DFF_X1 cor_m_2_3_reg_4_ ( .D(cor_maj_144_port_o), .CK(clk), .Q(
        cor_port_v_2_3[4]), .QN() );
  DFF_X1 cor_m_2_3_reg_5_ ( .D(cor_maj_145_port_o), .CK(clk), .Q(
        cor_port_v_2_3[5]), .QN() );
  DFF_X1 cor_m_2_3_reg_6_ ( .D(cor_maj_146_port_o), .CK(clk), .Q(
        cor_port_v_2_3[6]), .QN() );
  DFF_X1 cor_m_2_1_reg_0_ ( .D(cor_maj_133_port_o), .CK(clk), .Q(
        cor_port_v_2_1[0]), .QN() );
  DFF_X1 cor_m_2_1_reg_1_ ( .D(cor_maj_134_port_o), .CK(clk), .Q(
        cor_port_v_2_1[1]), .QN() );
  DFF_X1 cor_m_2_1_reg_2_ ( .D(cor_maj_135_port_o), .CK(clk), .Q(
        cor_port_v_2_1[2]), .QN() );
  DFF_X1 cor_m_2_1_reg_3_ ( .D(cor_maj_136_port_o), .CK(clk), .Q(
        cor_port_v_2_1[3]), .QN() );
  DFF_X1 cor_m_2_1_reg_4_ ( .D(cor_maj_137_port_o), .CK(clk), .Q(
        cor_port_v_2_1[4]), .QN() );
  DFF_X1 cor_m_2_1_reg_5_ ( .D(cor_maj_138_port_o), .CK(clk), .Q(
        cor_port_v_2_1[5]), .QN() );
  DFF_X1 cor_m_2_1_reg_6_ ( .D(cor_maj_139_port_o), .CK(clk), .Q(
        cor_port_v_2_1[6]), .QN() );
  DFF_X1 cor_m_2_0_reg_0_ ( .D(cor_maj_126_port_o), .CK(clk), .Q(
        cor_port_v_2_0[0]), .QN() );
  DFF_X1 cor_m_2_0_reg_1_ ( .D(cor_maj_127_port_o), .CK(clk), .Q(
        cor_port_v_2_0[1]), .QN() );
  DFF_X1 cor_m_2_0_reg_2_ ( .D(cor_maj_128_port_o), .CK(clk), .Q(
        cor_port_v_2_0[2]), .QN() );
  DFF_X1 cor_m_2_0_reg_3_ ( .D(cor_maj_129_port_o), .CK(clk), .Q(
        cor_port_v_2_0[3]), .QN() );
  DFF_X1 cor_m_2_0_reg_4_ ( .D(cor_maj_130_port_o), .CK(clk), .Q(
        cor_port_v_2_0[4]), .QN() );
  DFF_X1 cor_m_2_0_reg_5_ ( .D(cor_maj_131_port_o), .CK(clk), .Q(
        cor_port_v_2_0[5]), .QN() );
  DFF_X1 cor_m_2_0_reg_6_ ( .D(cor_maj_132_port_o), .CK(clk), .Q(
        cor_port_v_2_0[6]), .QN() );
  DFF_X1 cor_m_1_3_reg_0_ ( .D(cor_maj_119_port_o), .CK(clk), .Q(
        cor_port_v_1_3[0]), .QN() );
  DFF_X1 cor_m_1_3_reg_1_ ( .D(cor_maj_120_port_o), .CK(clk), .Q(
        cor_port_v_1_3[1]), .QN() );
  DFF_X1 cor_m_1_3_reg_2_ ( .D(cor_maj_121_port_o), .CK(clk), .Q(
        cor_port_v_1_3[2]), .QN() );
  DFF_X1 cor_m_1_3_reg_3_ ( .D(cor_maj_122_port_o), .CK(clk), .Q(
        cor_port_v_1_3[3]), .QN() );
  DFF_X1 cor_m_1_3_reg_4_ ( .D(cor_maj_123_port_o), .CK(clk), .Q(
        cor_port_v_1_3[4]), .QN() );
  DFF_X1 cor_m_1_3_reg_5_ ( .D(cor_maj_124_port_o), .CK(clk), .Q(
        cor_port_v_1_3[5]), .QN() );
  DFF_X1 cor_m_1_3_reg_6_ ( .D(cor_maj_125_port_o), .CK(clk), .Q(
        cor_port_v_1_3[6]), .QN() );
  DFF_X1 cor_m_1_2_reg_0_ ( .D(cor_maj_112_port_o), .CK(clk), .Q(
        cor_port_v_1_2[0]), .QN() );
  DFF_X1 cor_m_1_2_reg_1_ ( .D(cor_maj_113_port_o), .CK(clk), .Q(
        cor_port_v_1_2[1]), .QN() );
  DFF_X1 cor_m_1_2_reg_2_ ( .D(cor_maj_114_port_o), .CK(clk), .Q(
        cor_port_v_1_2[2]), .QN() );
  DFF_X1 cor_m_1_2_reg_3_ ( .D(cor_maj_115_port_o), .CK(clk), .Q(
        cor_port_v_1_2[3]), .QN() );
  DFF_X1 cor_m_1_2_reg_4_ ( .D(cor_maj_116_port_o), .CK(clk), .Q(
        cor_port_v_1_2[4]), .QN() );
  DFF_X1 cor_m_1_2_reg_5_ ( .D(cor_maj_117_port_o), .CK(clk), .Q(
        cor_port_v_1_2[5]), .QN() );
  DFF_X1 cor_m_1_2_reg_6_ ( .D(cor_maj_118_port_o), .CK(clk), .Q(
        cor_port_v_1_2[6]), .QN() );
  DFF_X1 cor_m_1_0_reg_0_ ( .D(cor_maj_105_port_o), .CK(clk), .Q(
        cor_port_v_1_0[0]), .QN() );
  DFF_X1 cor_m_1_0_reg_1_ ( .D(cor_maj_106_port_o), .CK(clk), .Q(
        cor_port_v_1_0[1]), .QN() );
  DFF_X1 cor_m_1_0_reg_2_ ( .D(cor_maj_107_port_o), .CK(clk), .Q(
        cor_port_v_1_0[2]), .QN() );
  DFF_X1 cor_m_1_0_reg_3_ ( .D(cor_maj_108_port_o), .CK(clk), .Q(
        cor_port_v_1_0[3]), .QN() );
  DFF_X1 cor_m_1_0_reg_4_ ( .D(cor_maj_109_port_o), .CK(clk), .Q(
        cor_port_v_1_0[4]), .QN() );
  DFF_X1 cor_m_1_0_reg_5_ ( .D(cor_maj_110_port_o), .CK(clk), .Q(
        cor_port_v_1_0[5]), .QN() );
  DFF_X1 cor_m_1_0_reg_6_ ( .D(cor_maj_111_port_o), .CK(clk), .Q(
        cor_port_v_1_0[6]), .QN() );
  DFF_X1 cor_m_0_3_reg_0_ ( .D(cor_maj_98_port_o), .CK(clk), .Q(
        cor_port_v_0_3[0]), .QN() );
  DFF_X1 cor_m_0_3_reg_1_ ( .D(cor_maj_99_port_o), .CK(clk), .Q(
        cor_port_v_0_3[1]), .QN() );
  DFF_X1 cor_m_0_3_reg_2_ ( .D(cor_maj_100_port_o), .CK(clk), .Q(
        cor_port_v_0_3[2]), .QN() );
  DFF_X1 cor_m_0_3_reg_3_ ( .D(cor_maj_101_port_o), .CK(clk), .Q(
        cor_port_v_0_3[3]), .QN() );
  DFF_X1 cor_m_0_3_reg_4_ ( .D(cor_maj_102_port_o), .CK(clk), .Q(
        cor_port_v_0_3[4]), .QN() );
  DFF_X1 cor_m_0_3_reg_5_ ( .D(cor_maj_103_port_o), .CK(clk), .Q(
        cor_port_v_0_3[5]), .QN() );
  DFF_X1 cor_m_0_3_reg_6_ ( .D(cor_maj_104_port_o), .CK(clk), .Q(
        cor_port_v_0_3[6]), .QN() );
  DFF_X1 cor_m_0_2_reg_0_ ( .D(cor_maj_91_port_o), .CK(clk), .Q(
        cor_port_v_0_2[0]), .QN() );
  DFF_X1 cor_m_0_2_reg_1_ ( .D(cor_maj_92_port_o), .CK(clk), .Q(
        cor_port_v_0_2[1]), .QN() );
  DFF_X1 cor_m_0_2_reg_2_ ( .D(cor_maj_93_port_o), .CK(clk), .Q(
        cor_port_v_0_2[2]), .QN() );
  DFF_X1 cor_m_0_2_reg_3_ ( .D(cor_maj_94_port_o), .CK(clk), .Q(
        cor_port_v_0_2[3]), .QN() );
  DFF_X1 cor_m_0_2_reg_4_ ( .D(cor_maj_95_port_o), .CK(clk), .Q(
        cor_port_v_0_2[4]), .QN() );
  DFF_X1 cor_m_0_2_reg_5_ ( .D(cor_maj_96_port_o), .CK(clk), .Q(
        cor_port_v_0_2[5]), .QN() );
  DFF_X1 cor_m_0_2_reg_6_ ( .D(cor_maj_97_port_o), .CK(clk), .Q(
        cor_port_v_0_2[6]), .QN() );
  DFF_X1 cor_m_0_1_reg_0_ ( .D(cor_maj_84_port_o), .CK(clk), .Q(
        cor_port_v_0_1[0]), .QN() );
  DFF_X1 cor_m_0_1_reg_1_ ( .D(cor_maj_85_port_o), .CK(clk), .Q(
        cor_port_v_0_1[1]), .QN() );
  DFF_X1 cor_m_0_1_reg_2_ ( .D(cor_maj_86_port_o), .CK(clk), .Q(
        cor_port_v_0_1[2]), .QN() );
  DFF_X1 cor_m_0_1_reg_3_ ( .D(cor_maj_87_port_o), .CK(clk), .Q(
        cor_port_v_0_1[3]), .QN() );
  DFF_X1 cor_m_0_1_reg_4_ ( .D(cor_maj_88_port_o), .CK(clk), .Q(
        cor_port_v_0_1[4]), .QN() );
  DFF_X1 cor_m_0_1_reg_5_ ( .D(cor_maj_89_port_o), .CK(clk), .Q(
        cor_port_v_0_1[5]), .QN() );
  DFF_X1 cor_m_0_1_reg_6_ ( .D(cor_maj_90_port_o), .CK(clk), .Q(
        cor_port_v_0_1[6]), .QN() );
  OR2_X1 cor_maj_84_U19 ( .A1(cor_maj_84_n8), .A2(cor_maj_84_n9), .ZN(
        cor_maj_84_n7) );
  NAND2_X1 cor_maj_84_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_84_n7), .ZN(
        cor_maj_84_n6) );
  NAND2_X1 cor_maj_84_U17 ( .A1(cor_maj_84_n9), .A2(cor_maj_84_n8), .ZN(
        cor_maj_84_n5) );
  NAND2_X1 cor_maj_84_U16 ( .A1(cor_maj_84_n5), .A2(cor_maj_84_n6), .ZN(
        cor_maj_84_n4) );
  NAND2_X1 cor_maj_84_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_84_n10), .ZN(
        cor_maj_84_n17) );
  NAND2_X1 cor_maj_84_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_84_n16) );
  NAND2_X1 cor_maj_84_U13 ( .A1(cor_maj_84_n16), .A2(cor_maj_84_n17), .ZN(
        cor_maj_84_n13) );
  NAND2_X1 cor_maj_84_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_84_n11), .ZN(
        cor_maj_84_n15) );
  NAND2_X1 cor_maj_84_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_84_n14) );
  NAND2_X1 cor_maj_84_U10 ( .A1(cor_maj_84_n14), .A2(cor_maj_84_n15), .ZN(
        cor_maj_84_n12) );
  XOR2_X1 cor_maj_84_U9 ( .A(v_1_0_1[2]), .B(cor_maj_84_n11), .Z(cor_maj_84_n9) );
  XOR2_X1 cor_maj_84_U8 ( .A(v_1_0_1[5]), .B(cor_maj_84_n10), .Z(cor_maj_84_n8) );
  XOR2_X1 cor_maj_84_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_84_n11)
         );
  XOR2_X1 cor_maj_84_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_84_n10)
         );
  OR2_X1 cor_maj_84_U5 ( .A1(cor_maj_84_n12), .A2(cor_maj_84_n13), .ZN(
        cor_maj_84_n3) );
  NAND2_X1 cor_maj_84_U4 ( .A1(cor_maj_84_n13), .A2(cor_maj_84_n12), .ZN(
        cor_maj_84_n1) );
  NAND2_X1 cor_maj_84_U3 ( .A1(cor_maj_84_n3), .A2(cor_maj_84_n4), .ZN(
        cor_maj_84_n2) );
  NAND2_X1 cor_maj_84_U2 ( .A1(cor_maj_84_n1), .A2(cor_maj_84_n2), .ZN(
        cor_maj_84_port_o) );
  OR2_X1 cor_maj_85_U19 ( .A1(cor_maj_85_n27), .A2(cor_maj_85_n26), .ZN(
        cor_maj_85_n28) );
  NAND2_X1 cor_maj_85_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_85_n28), .ZN(
        cor_maj_85_n29) );
  NAND2_X1 cor_maj_85_U17 ( .A1(cor_maj_85_n26), .A2(cor_maj_85_n27), .ZN(
        cor_maj_85_n30) );
  NAND2_X1 cor_maj_85_U16 ( .A1(cor_maj_85_n30), .A2(cor_maj_85_n29), .ZN(
        cor_maj_85_n31) );
  NAND2_X1 cor_maj_85_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_85_n25), .ZN(
        cor_maj_85_n18) );
  NAND2_X1 cor_maj_85_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_85_n19) );
  NAND2_X1 cor_maj_85_U13 ( .A1(cor_maj_85_n19), .A2(cor_maj_85_n18), .ZN(
        cor_maj_85_n22) );
  NAND2_X1 cor_maj_85_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_85_n24), .ZN(
        cor_maj_85_n20) );
  NAND2_X1 cor_maj_85_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_85_n21) );
  NAND2_X1 cor_maj_85_U10 ( .A1(cor_maj_85_n21), .A2(cor_maj_85_n20), .ZN(
        cor_maj_85_n23) );
  XOR2_X1 cor_maj_85_U9 ( .A(v_1_0_1[2]), .B(cor_maj_85_n24), .Z(
        cor_maj_85_n26) );
  XOR2_X1 cor_maj_85_U8 ( .A(v_1_0_1[5]), .B(cor_maj_85_n25), .Z(
        cor_maj_85_n27) );
  XOR2_X1 cor_maj_85_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_85_n24)
         );
  XOR2_X1 cor_maj_85_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_85_n25)
         );
  OR2_X1 cor_maj_85_U5 ( .A1(cor_maj_85_n23), .A2(cor_maj_85_n22), .ZN(
        cor_maj_85_n32) );
  NAND2_X1 cor_maj_85_U4 ( .A1(cor_maj_85_n22), .A2(cor_maj_85_n23), .ZN(
        cor_maj_85_n34) );
  NAND2_X1 cor_maj_85_U3 ( .A1(cor_maj_85_n32), .A2(cor_maj_85_n31), .ZN(
        cor_maj_85_n33) );
  NAND2_X1 cor_maj_85_U2 ( .A1(cor_maj_85_n34), .A2(cor_maj_85_n33), .ZN(
        cor_maj_85_port_o) );
  OR2_X1 cor_maj_86_U19 ( .A1(cor_maj_86_n27), .A2(cor_maj_86_n26), .ZN(
        cor_maj_86_n28) );
  NAND2_X1 cor_maj_86_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_86_n28), .ZN(
        cor_maj_86_n29) );
  NAND2_X1 cor_maj_86_U17 ( .A1(cor_maj_86_n26), .A2(cor_maj_86_n27), .ZN(
        cor_maj_86_n30) );
  NAND2_X1 cor_maj_86_U16 ( .A1(cor_maj_86_n30), .A2(cor_maj_86_n29), .ZN(
        cor_maj_86_n31) );
  NAND2_X1 cor_maj_86_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_86_n25), .ZN(
        cor_maj_86_n18) );
  NAND2_X1 cor_maj_86_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_86_n19) );
  NAND2_X1 cor_maj_86_U13 ( .A1(cor_maj_86_n19), .A2(cor_maj_86_n18), .ZN(
        cor_maj_86_n22) );
  NAND2_X1 cor_maj_86_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_86_n24), .ZN(
        cor_maj_86_n20) );
  NAND2_X1 cor_maj_86_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_86_n21) );
  NAND2_X1 cor_maj_86_U10 ( .A1(cor_maj_86_n21), .A2(cor_maj_86_n20), .ZN(
        cor_maj_86_n23) );
  XOR2_X1 cor_maj_86_U9 ( .A(v_1_0_1[2]), .B(cor_maj_86_n24), .Z(
        cor_maj_86_n26) );
  XOR2_X1 cor_maj_86_U8 ( .A(v_1_0_1[5]), .B(cor_maj_86_n25), .Z(
        cor_maj_86_n27) );
  XOR2_X1 cor_maj_86_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_86_n24)
         );
  XOR2_X1 cor_maj_86_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_86_n25)
         );
  OR2_X1 cor_maj_86_U5 ( .A1(cor_maj_86_n23), .A2(cor_maj_86_n22), .ZN(
        cor_maj_86_n32) );
  NAND2_X1 cor_maj_86_U4 ( .A1(cor_maj_86_n22), .A2(cor_maj_86_n23), .ZN(
        cor_maj_86_n34) );
  NAND2_X1 cor_maj_86_U3 ( .A1(cor_maj_86_n32), .A2(cor_maj_86_n31), .ZN(
        cor_maj_86_n33) );
  NAND2_X1 cor_maj_86_U2 ( .A1(cor_maj_86_n34), .A2(cor_maj_86_n33), .ZN(
        cor_maj_86_port_o) );
  OR2_X1 cor_maj_87_U19 ( .A1(cor_maj_87_n27), .A2(cor_maj_87_n26), .ZN(
        cor_maj_87_n28) );
  NAND2_X1 cor_maj_87_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_87_n28), .ZN(
        cor_maj_87_n29) );
  NAND2_X1 cor_maj_87_U17 ( .A1(cor_maj_87_n26), .A2(cor_maj_87_n27), .ZN(
        cor_maj_87_n30) );
  NAND2_X1 cor_maj_87_U16 ( .A1(cor_maj_87_n30), .A2(cor_maj_87_n29), .ZN(
        cor_maj_87_n31) );
  NAND2_X1 cor_maj_87_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_87_n25), .ZN(
        cor_maj_87_n18) );
  NAND2_X1 cor_maj_87_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_87_n19) );
  NAND2_X1 cor_maj_87_U13 ( .A1(cor_maj_87_n19), .A2(cor_maj_87_n18), .ZN(
        cor_maj_87_n22) );
  NAND2_X1 cor_maj_87_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_87_n24), .ZN(
        cor_maj_87_n20) );
  NAND2_X1 cor_maj_87_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_87_n21) );
  NAND2_X1 cor_maj_87_U10 ( .A1(cor_maj_87_n21), .A2(cor_maj_87_n20), .ZN(
        cor_maj_87_n23) );
  XOR2_X1 cor_maj_87_U9 ( .A(v_1_0_1[2]), .B(cor_maj_87_n24), .Z(
        cor_maj_87_n26) );
  XOR2_X1 cor_maj_87_U8 ( .A(v_1_0_1[5]), .B(cor_maj_87_n25), .Z(
        cor_maj_87_n27) );
  XOR2_X1 cor_maj_87_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_87_n24)
         );
  XOR2_X1 cor_maj_87_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_87_n25)
         );
  OR2_X1 cor_maj_87_U5 ( .A1(cor_maj_87_n23), .A2(cor_maj_87_n22), .ZN(
        cor_maj_87_n32) );
  NAND2_X1 cor_maj_87_U4 ( .A1(cor_maj_87_n22), .A2(cor_maj_87_n23), .ZN(
        cor_maj_87_n34) );
  NAND2_X1 cor_maj_87_U3 ( .A1(cor_maj_87_n32), .A2(cor_maj_87_n31), .ZN(
        cor_maj_87_n33) );
  NAND2_X1 cor_maj_87_U2 ( .A1(cor_maj_87_n34), .A2(cor_maj_87_n33), .ZN(
        cor_maj_87_port_o) );
  OR2_X1 cor_maj_88_U19 ( .A1(cor_maj_88_n27), .A2(cor_maj_88_n26), .ZN(
        cor_maj_88_n28) );
  NAND2_X1 cor_maj_88_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_88_n28), .ZN(
        cor_maj_88_n29) );
  NAND2_X1 cor_maj_88_U17 ( .A1(cor_maj_88_n26), .A2(cor_maj_88_n27), .ZN(
        cor_maj_88_n30) );
  NAND2_X1 cor_maj_88_U16 ( .A1(cor_maj_88_n30), .A2(cor_maj_88_n29), .ZN(
        cor_maj_88_n31) );
  NAND2_X1 cor_maj_88_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_88_n25), .ZN(
        cor_maj_88_n18) );
  NAND2_X1 cor_maj_88_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_88_n19) );
  NAND2_X1 cor_maj_88_U13 ( .A1(cor_maj_88_n19), .A2(cor_maj_88_n18), .ZN(
        cor_maj_88_n22) );
  NAND2_X1 cor_maj_88_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_88_n24), .ZN(
        cor_maj_88_n20) );
  NAND2_X1 cor_maj_88_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_88_n21) );
  NAND2_X1 cor_maj_88_U10 ( .A1(cor_maj_88_n21), .A2(cor_maj_88_n20), .ZN(
        cor_maj_88_n23) );
  XOR2_X1 cor_maj_88_U9 ( .A(v_1_0_1[2]), .B(cor_maj_88_n24), .Z(
        cor_maj_88_n26) );
  XOR2_X1 cor_maj_88_U8 ( .A(v_1_0_1[5]), .B(cor_maj_88_n25), .Z(
        cor_maj_88_n27) );
  XOR2_X1 cor_maj_88_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_88_n24)
         );
  XOR2_X1 cor_maj_88_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_88_n25)
         );
  OR2_X1 cor_maj_88_U5 ( .A1(cor_maj_88_n23), .A2(cor_maj_88_n22), .ZN(
        cor_maj_88_n32) );
  NAND2_X1 cor_maj_88_U4 ( .A1(cor_maj_88_n22), .A2(cor_maj_88_n23), .ZN(
        cor_maj_88_n34) );
  NAND2_X1 cor_maj_88_U3 ( .A1(cor_maj_88_n32), .A2(cor_maj_88_n31), .ZN(
        cor_maj_88_n33) );
  NAND2_X1 cor_maj_88_U2 ( .A1(cor_maj_88_n34), .A2(cor_maj_88_n33), .ZN(
        cor_maj_88_port_o) );
  OR2_X1 cor_maj_89_U19 ( .A1(cor_maj_89_n27), .A2(cor_maj_89_n26), .ZN(
        cor_maj_89_n28) );
  NAND2_X1 cor_maj_89_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_89_n28), .ZN(
        cor_maj_89_n29) );
  NAND2_X1 cor_maj_89_U17 ( .A1(cor_maj_89_n26), .A2(cor_maj_89_n27), .ZN(
        cor_maj_89_n30) );
  NAND2_X1 cor_maj_89_U16 ( .A1(cor_maj_89_n30), .A2(cor_maj_89_n29), .ZN(
        cor_maj_89_n31) );
  NAND2_X1 cor_maj_89_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_89_n25), .ZN(
        cor_maj_89_n18) );
  NAND2_X1 cor_maj_89_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_89_n19) );
  NAND2_X1 cor_maj_89_U13 ( .A1(cor_maj_89_n19), .A2(cor_maj_89_n18), .ZN(
        cor_maj_89_n22) );
  NAND2_X1 cor_maj_89_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_89_n24), .ZN(
        cor_maj_89_n20) );
  NAND2_X1 cor_maj_89_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_89_n21) );
  NAND2_X1 cor_maj_89_U10 ( .A1(cor_maj_89_n21), .A2(cor_maj_89_n20), .ZN(
        cor_maj_89_n23) );
  XOR2_X1 cor_maj_89_U9 ( .A(v_1_0_1[2]), .B(cor_maj_89_n24), .Z(
        cor_maj_89_n26) );
  XOR2_X1 cor_maj_89_U8 ( .A(v_1_0_1[5]), .B(cor_maj_89_n25), .Z(
        cor_maj_89_n27) );
  XOR2_X1 cor_maj_89_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_89_n24)
         );
  XOR2_X1 cor_maj_89_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_89_n25)
         );
  OR2_X1 cor_maj_89_U5 ( .A1(cor_maj_89_n23), .A2(cor_maj_89_n22), .ZN(
        cor_maj_89_n32) );
  NAND2_X1 cor_maj_89_U4 ( .A1(cor_maj_89_n22), .A2(cor_maj_89_n23), .ZN(
        cor_maj_89_n34) );
  NAND2_X1 cor_maj_89_U3 ( .A1(cor_maj_89_n32), .A2(cor_maj_89_n31), .ZN(
        cor_maj_89_n33) );
  NAND2_X1 cor_maj_89_U2 ( .A1(cor_maj_89_n34), .A2(cor_maj_89_n33), .ZN(
        cor_maj_89_port_o) );
  OR2_X1 cor_maj_90_U19 ( .A1(cor_maj_90_n27), .A2(cor_maj_90_n26), .ZN(
        cor_maj_90_n28) );
  NAND2_X1 cor_maj_90_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_90_n28), .ZN(
        cor_maj_90_n29) );
  NAND2_X1 cor_maj_90_U17 ( .A1(cor_maj_90_n26), .A2(cor_maj_90_n27), .ZN(
        cor_maj_90_n30) );
  NAND2_X1 cor_maj_90_U16 ( .A1(cor_maj_90_n30), .A2(cor_maj_90_n29), .ZN(
        cor_maj_90_n31) );
  NAND2_X1 cor_maj_90_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_90_n25), .ZN(
        cor_maj_90_n18) );
  NAND2_X1 cor_maj_90_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_90_n19) );
  NAND2_X1 cor_maj_90_U13 ( .A1(cor_maj_90_n19), .A2(cor_maj_90_n18), .ZN(
        cor_maj_90_n22) );
  NAND2_X1 cor_maj_90_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_90_n24), .ZN(
        cor_maj_90_n20) );
  NAND2_X1 cor_maj_90_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_90_n21) );
  NAND2_X1 cor_maj_90_U10 ( .A1(cor_maj_90_n21), .A2(cor_maj_90_n20), .ZN(
        cor_maj_90_n23) );
  XOR2_X1 cor_maj_90_U9 ( .A(v_1_0_1[2]), .B(cor_maj_90_n24), .Z(
        cor_maj_90_n26) );
  XOR2_X1 cor_maj_90_U8 ( .A(v_1_0_1[5]), .B(cor_maj_90_n25), .Z(
        cor_maj_90_n27) );
  XOR2_X1 cor_maj_90_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_90_n24)
         );
  XOR2_X1 cor_maj_90_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_90_n25)
         );
  OR2_X1 cor_maj_90_U5 ( .A1(cor_maj_90_n23), .A2(cor_maj_90_n22), .ZN(
        cor_maj_90_n32) );
  NAND2_X1 cor_maj_90_U4 ( .A1(cor_maj_90_n22), .A2(cor_maj_90_n23), .ZN(
        cor_maj_90_n34) );
  NAND2_X1 cor_maj_90_U3 ( .A1(cor_maj_90_n32), .A2(cor_maj_90_n31), .ZN(
        cor_maj_90_n33) );
  NAND2_X1 cor_maj_90_U2 ( .A1(cor_maj_90_n34), .A2(cor_maj_90_n33), .ZN(
        cor_maj_90_port_o) );
  OR2_X1 cor_maj_91_U19 ( .A1(cor_maj_91_n27), .A2(cor_maj_91_n26), .ZN(
        cor_maj_91_n28) );
  NAND2_X1 cor_maj_91_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_91_n28), .ZN(
        cor_maj_91_n29) );
  NAND2_X1 cor_maj_91_U17 ( .A1(cor_maj_91_n26), .A2(cor_maj_91_n27), .ZN(
        cor_maj_91_n30) );
  NAND2_X1 cor_maj_91_U16 ( .A1(cor_maj_91_n30), .A2(cor_maj_91_n29), .ZN(
        cor_maj_91_n31) );
  NAND2_X1 cor_maj_91_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_91_n25), .ZN(
        cor_maj_91_n18) );
  NAND2_X1 cor_maj_91_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_91_n19) );
  NAND2_X1 cor_maj_91_U13 ( .A1(cor_maj_91_n19), .A2(cor_maj_91_n18), .ZN(
        cor_maj_91_n22) );
  NAND2_X1 cor_maj_91_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_91_n24), .ZN(
        cor_maj_91_n20) );
  NAND2_X1 cor_maj_91_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_91_n21) );
  NAND2_X1 cor_maj_91_U10 ( .A1(cor_maj_91_n21), .A2(cor_maj_91_n20), .ZN(
        cor_maj_91_n23) );
  XOR2_X1 cor_maj_91_U9 ( .A(v_1_0_2[2]), .B(cor_maj_91_n24), .Z(
        cor_maj_91_n26) );
  XOR2_X1 cor_maj_91_U8 ( .A(v_1_0_2[5]), .B(cor_maj_91_n25), .Z(
        cor_maj_91_n27) );
  XOR2_X1 cor_maj_91_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_91_n24)
         );
  XOR2_X1 cor_maj_91_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_91_n25)
         );
  OR2_X1 cor_maj_91_U5 ( .A1(cor_maj_91_n23), .A2(cor_maj_91_n22), .ZN(
        cor_maj_91_n32) );
  NAND2_X1 cor_maj_91_U4 ( .A1(cor_maj_91_n22), .A2(cor_maj_91_n23), .ZN(
        cor_maj_91_n34) );
  NAND2_X1 cor_maj_91_U3 ( .A1(cor_maj_91_n32), .A2(cor_maj_91_n31), .ZN(
        cor_maj_91_n33) );
  NAND2_X1 cor_maj_91_U2 ( .A1(cor_maj_91_n34), .A2(cor_maj_91_n33), .ZN(
        cor_maj_91_port_o) );
  OR2_X1 cor_maj_92_U19 ( .A1(cor_maj_92_n27), .A2(cor_maj_92_n26), .ZN(
        cor_maj_92_n28) );
  NAND2_X1 cor_maj_92_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_92_n28), .ZN(
        cor_maj_92_n29) );
  NAND2_X1 cor_maj_92_U17 ( .A1(cor_maj_92_n26), .A2(cor_maj_92_n27), .ZN(
        cor_maj_92_n30) );
  NAND2_X1 cor_maj_92_U16 ( .A1(cor_maj_92_n30), .A2(cor_maj_92_n29), .ZN(
        cor_maj_92_n31) );
  NAND2_X1 cor_maj_92_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_92_n25), .ZN(
        cor_maj_92_n18) );
  NAND2_X1 cor_maj_92_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_92_n19) );
  NAND2_X1 cor_maj_92_U13 ( .A1(cor_maj_92_n19), .A2(cor_maj_92_n18), .ZN(
        cor_maj_92_n22) );
  NAND2_X1 cor_maj_92_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_92_n24), .ZN(
        cor_maj_92_n20) );
  NAND2_X1 cor_maj_92_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_92_n21) );
  NAND2_X1 cor_maj_92_U10 ( .A1(cor_maj_92_n21), .A2(cor_maj_92_n20), .ZN(
        cor_maj_92_n23) );
  XOR2_X1 cor_maj_92_U9 ( .A(v_1_0_2[2]), .B(cor_maj_92_n24), .Z(
        cor_maj_92_n26) );
  XOR2_X1 cor_maj_92_U8 ( .A(v_1_0_2[5]), .B(cor_maj_92_n25), .Z(
        cor_maj_92_n27) );
  XOR2_X1 cor_maj_92_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_92_n24)
         );
  XOR2_X1 cor_maj_92_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_92_n25)
         );
  OR2_X1 cor_maj_92_U5 ( .A1(cor_maj_92_n23), .A2(cor_maj_92_n22), .ZN(
        cor_maj_92_n32) );
  NAND2_X1 cor_maj_92_U4 ( .A1(cor_maj_92_n22), .A2(cor_maj_92_n23), .ZN(
        cor_maj_92_n34) );
  NAND2_X1 cor_maj_92_U3 ( .A1(cor_maj_92_n32), .A2(cor_maj_92_n31), .ZN(
        cor_maj_92_n33) );
  NAND2_X1 cor_maj_92_U2 ( .A1(cor_maj_92_n34), .A2(cor_maj_92_n33), .ZN(
        cor_maj_92_port_o) );
  OR2_X1 cor_maj_93_U19 ( .A1(cor_maj_93_n27), .A2(cor_maj_93_n26), .ZN(
        cor_maj_93_n28) );
  NAND2_X1 cor_maj_93_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_93_n28), .ZN(
        cor_maj_93_n29) );
  NAND2_X1 cor_maj_93_U17 ( .A1(cor_maj_93_n26), .A2(cor_maj_93_n27), .ZN(
        cor_maj_93_n30) );
  NAND2_X1 cor_maj_93_U16 ( .A1(cor_maj_93_n30), .A2(cor_maj_93_n29), .ZN(
        cor_maj_93_n31) );
  NAND2_X1 cor_maj_93_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_93_n25), .ZN(
        cor_maj_93_n18) );
  NAND2_X1 cor_maj_93_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_93_n19) );
  NAND2_X1 cor_maj_93_U13 ( .A1(cor_maj_93_n19), .A2(cor_maj_93_n18), .ZN(
        cor_maj_93_n22) );
  NAND2_X1 cor_maj_93_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_93_n24), .ZN(
        cor_maj_93_n20) );
  NAND2_X1 cor_maj_93_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_93_n21) );
  NAND2_X1 cor_maj_93_U10 ( .A1(cor_maj_93_n21), .A2(cor_maj_93_n20), .ZN(
        cor_maj_93_n23) );
  XOR2_X1 cor_maj_93_U9 ( .A(v_1_0_2[2]), .B(cor_maj_93_n24), .Z(
        cor_maj_93_n26) );
  XOR2_X1 cor_maj_93_U8 ( .A(v_1_0_2[5]), .B(cor_maj_93_n25), .Z(
        cor_maj_93_n27) );
  XOR2_X1 cor_maj_93_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_93_n24)
         );
  XOR2_X1 cor_maj_93_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_93_n25)
         );
  OR2_X1 cor_maj_93_U5 ( .A1(cor_maj_93_n23), .A2(cor_maj_93_n22), .ZN(
        cor_maj_93_n32) );
  NAND2_X1 cor_maj_93_U4 ( .A1(cor_maj_93_n22), .A2(cor_maj_93_n23), .ZN(
        cor_maj_93_n34) );
  NAND2_X1 cor_maj_93_U3 ( .A1(cor_maj_93_n32), .A2(cor_maj_93_n31), .ZN(
        cor_maj_93_n33) );
  NAND2_X1 cor_maj_93_U2 ( .A1(cor_maj_93_n34), .A2(cor_maj_93_n33), .ZN(
        cor_maj_93_port_o) );
  OR2_X1 cor_maj_94_U19 ( .A1(cor_maj_94_n27), .A2(cor_maj_94_n26), .ZN(
        cor_maj_94_n28) );
  NAND2_X1 cor_maj_94_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_94_n28), .ZN(
        cor_maj_94_n29) );
  NAND2_X1 cor_maj_94_U17 ( .A1(cor_maj_94_n26), .A2(cor_maj_94_n27), .ZN(
        cor_maj_94_n30) );
  NAND2_X1 cor_maj_94_U16 ( .A1(cor_maj_94_n30), .A2(cor_maj_94_n29), .ZN(
        cor_maj_94_n31) );
  NAND2_X1 cor_maj_94_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_94_n25), .ZN(
        cor_maj_94_n18) );
  NAND2_X1 cor_maj_94_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_94_n19) );
  NAND2_X1 cor_maj_94_U13 ( .A1(cor_maj_94_n19), .A2(cor_maj_94_n18), .ZN(
        cor_maj_94_n22) );
  NAND2_X1 cor_maj_94_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_94_n24), .ZN(
        cor_maj_94_n20) );
  NAND2_X1 cor_maj_94_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_94_n21) );
  NAND2_X1 cor_maj_94_U10 ( .A1(cor_maj_94_n21), .A2(cor_maj_94_n20), .ZN(
        cor_maj_94_n23) );
  XOR2_X1 cor_maj_94_U9 ( .A(v_1_0_2[2]), .B(cor_maj_94_n24), .Z(
        cor_maj_94_n26) );
  XOR2_X1 cor_maj_94_U8 ( .A(v_1_0_2[5]), .B(cor_maj_94_n25), .Z(
        cor_maj_94_n27) );
  XOR2_X1 cor_maj_94_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_94_n24)
         );
  XOR2_X1 cor_maj_94_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_94_n25)
         );
  OR2_X1 cor_maj_94_U5 ( .A1(cor_maj_94_n23), .A2(cor_maj_94_n22), .ZN(
        cor_maj_94_n32) );
  NAND2_X1 cor_maj_94_U4 ( .A1(cor_maj_94_n22), .A2(cor_maj_94_n23), .ZN(
        cor_maj_94_n34) );
  NAND2_X1 cor_maj_94_U3 ( .A1(cor_maj_94_n32), .A2(cor_maj_94_n31), .ZN(
        cor_maj_94_n33) );
  NAND2_X1 cor_maj_94_U2 ( .A1(cor_maj_94_n34), .A2(cor_maj_94_n33), .ZN(
        cor_maj_94_port_o) );
  OR2_X1 cor_maj_95_U19 ( .A1(cor_maj_95_n27), .A2(cor_maj_95_n26), .ZN(
        cor_maj_95_n28) );
  NAND2_X1 cor_maj_95_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_95_n28), .ZN(
        cor_maj_95_n29) );
  NAND2_X1 cor_maj_95_U17 ( .A1(cor_maj_95_n26), .A2(cor_maj_95_n27), .ZN(
        cor_maj_95_n30) );
  NAND2_X1 cor_maj_95_U16 ( .A1(cor_maj_95_n30), .A2(cor_maj_95_n29), .ZN(
        cor_maj_95_n31) );
  NAND2_X1 cor_maj_95_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_95_n25), .ZN(
        cor_maj_95_n18) );
  NAND2_X1 cor_maj_95_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_95_n19) );
  NAND2_X1 cor_maj_95_U13 ( .A1(cor_maj_95_n19), .A2(cor_maj_95_n18), .ZN(
        cor_maj_95_n22) );
  NAND2_X1 cor_maj_95_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_95_n24), .ZN(
        cor_maj_95_n20) );
  NAND2_X1 cor_maj_95_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_95_n21) );
  NAND2_X1 cor_maj_95_U10 ( .A1(cor_maj_95_n21), .A2(cor_maj_95_n20), .ZN(
        cor_maj_95_n23) );
  XOR2_X1 cor_maj_95_U9 ( .A(v_1_0_2[2]), .B(cor_maj_95_n24), .Z(
        cor_maj_95_n26) );
  XOR2_X1 cor_maj_95_U8 ( .A(v_1_0_2[5]), .B(cor_maj_95_n25), .Z(
        cor_maj_95_n27) );
  XOR2_X1 cor_maj_95_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_95_n24)
         );
  XOR2_X1 cor_maj_95_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_95_n25)
         );
  OR2_X1 cor_maj_95_U5 ( .A1(cor_maj_95_n23), .A2(cor_maj_95_n22), .ZN(
        cor_maj_95_n32) );
  NAND2_X1 cor_maj_95_U4 ( .A1(cor_maj_95_n22), .A2(cor_maj_95_n23), .ZN(
        cor_maj_95_n34) );
  NAND2_X1 cor_maj_95_U3 ( .A1(cor_maj_95_n32), .A2(cor_maj_95_n31), .ZN(
        cor_maj_95_n33) );
  NAND2_X1 cor_maj_95_U2 ( .A1(cor_maj_95_n34), .A2(cor_maj_95_n33), .ZN(
        cor_maj_95_port_o) );
  OR2_X1 cor_maj_96_U19 ( .A1(cor_maj_96_n27), .A2(cor_maj_96_n26), .ZN(
        cor_maj_96_n28) );
  NAND2_X1 cor_maj_96_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_96_n28), .ZN(
        cor_maj_96_n29) );
  NAND2_X1 cor_maj_96_U17 ( .A1(cor_maj_96_n26), .A2(cor_maj_96_n27), .ZN(
        cor_maj_96_n30) );
  NAND2_X1 cor_maj_96_U16 ( .A1(cor_maj_96_n30), .A2(cor_maj_96_n29), .ZN(
        cor_maj_96_n31) );
  NAND2_X1 cor_maj_96_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_96_n25), .ZN(
        cor_maj_96_n18) );
  NAND2_X1 cor_maj_96_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_96_n19) );
  NAND2_X1 cor_maj_96_U13 ( .A1(cor_maj_96_n19), .A2(cor_maj_96_n18), .ZN(
        cor_maj_96_n22) );
  NAND2_X1 cor_maj_96_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_96_n24), .ZN(
        cor_maj_96_n20) );
  NAND2_X1 cor_maj_96_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_96_n21) );
  NAND2_X1 cor_maj_96_U10 ( .A1(cor_maj_96_n21), .A2(cor_maj_96_n20), .ZN(
        cor_maj_96_n23) );
  XOR2_X1 cor_maj_96_U9 ( .A(v_1_0_2[2]), .B(cor_maj_96_n24), .Z(
        cor_maj_96_n26) );
  XOR2_X1 cor_maj_96_U8 ( .A(v_1_0_2[5]), .B(cor_maj_96_n25), .Z(
        cor_maj_96_n27) );
  XOR2_X1 cor_maj_96_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_96_n24)
         );
  XOR2_X1 cor_maj_96_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_96_n25)
         );
  OR2_X1 cor_maj_96_U5 ( .A1(cor_maj_96_n23), .A2(cor_maj_96_n22), .ZN(
        cor_maj_96_n32) );
  NAND2_X1 cor_maj_96_U4 ( .A1(cor_maj_96_n22), .A2(cor_maj_96_n23), .ZN(
        cor_maj_96_n34) );
  NAND2_X1 cor_maj_96_U3 ( .A1(cor_maj_96_n32), .A2(cor_maj_96_n31), .ZN(
        cor_maj_96_n33) );
  NAND2_X1 cor_maj_96_U2 ( .A1(cor_maj_96_n34), .A2(cor_maj_96_n33), .ZN(
        cor_maj_96_port_o) );
  OR2_X1 cor_maj_97_U19 ( .A1(cor_maj_97_n27), .A2(cor_maj_97_n26), .ZN(
        cor_maj_97_n28) );
  NAND2_X1 cor_maj_97_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_97_n28), .ZN(
        cor_maj_97_n29) );
  NAND2_X1 cor_maj_97_U17 ( .A1(cor_maj_97_n26), .A2(cor_maj_97_n27), .ZN(
        cor_maj_97_n30) );
  NAND2_X1 cor_maj_97_U16 ( .A1(cor_maj_97_n30), .A2(cor_maj_97_n29), .ZN(
        cor_maj_97_n31) );
  NAND2_X1 cor_maj_97_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_97_n25), .ZN(
        cor_maj_97_n18) );
  NAND2_X1 cor_maj_97_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_97_n19) );
  NAND2_X1 cor_maj_97_U13 ( .A1(cor_maj_97_n19), .A2(cor_maj_97_n18), .ZN(
        cor_maj_97_n22) );
  NAND2_X1 cor_maj_97_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_97_n24), .ZN(
        cor_maj_97_n20) );
  NAND2_X1 cor_maj_97_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_97_n21) );
  NAND2_X1 cor_maj_97_U10 ( .A1(cor_maj_97_n21), .A2(cor_maj_97_n20), .ZN(
        cor_maj_97_n23) );
  XOR2_X1 cor_maj_97_U9 ( .A(v_1_0_2[2]), .B(cor_maj_97_n24), .Z(
        cor_maj_97_n26) );
  XOR2_X1 cor_maj_97_U8 ( .A(v_1_0_2[5]), .B(cor_maj_97_n25), .Z(
        cor_maj_97_n27) );
  XOR2_X1 cor_maj_97_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_97_n24)
         );
  XOR2_X1 cor_maj_97_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_97_n25)
         );
  OR2_X1 cor_maj_97_U5 ( .A1(cor_maj_97_n23), .A2(cor_maj_97_n22), .ZN(
        cor_maj_97_n32) );
  NAND2_X1 cor_maj_97_U4 ( .A1(cor_maj_97_n22), .A2(cor_maj_97_n23), .ZN(
        cor_maj_97_n34) );
  NAND2_X1 cor_maj_97_U3 ( .A1(cor_maj_97_n32), .A2(cor_maj_97_n31), .ZN(
        cor_maj_97_n33) );
  NAND2_X1 cor_maj_97_U2 ( .A1(cor_maj_97_n34), .A2(cor_maj_97_n33), .ZN(
        cor_maj_97_port_o) );
  OR2_X1 cor_maj_98_U19 ( .A1(cor_maj_98_n27), .A2(cor_maj_98_n26), .ZN(
        cor_maj_98_n28) );
  NAND2_X1 cor_maj_98_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_98_n28), .ZN(
        cor_maj_98_n29) );
  NAND2_X1 cor_maj_98_U17 ( .A1(cor_maj_98_n26), .A2(cor_maj_98_n27), .ZN(
        cor_maj_98_n30) );
  NAND2_X1 cor_maj_98_U16 ( .A1(cor_maj_98_n30), .A2(cor_maj_98_n29), .ZN(
        cor_maj_98_n31) );
  NAND2_X1 cor_maj_98_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_98_n25), .ZN(
        cor_maj_98_n18) );
  NAND2_X1 cor_maj_98_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_98_n19) );
  NAND2_X1 cor_maj_98_U13 ( .A1(cor_maj_98_n19), .A2(cor_maj_98_n18), .ZN(
        cor_maj_98_n22) );
  NAND2_X1 cor_maj_98_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_98_n24), .ZN(
        cor_maj_98_n20) );
  NAND2_X1 cor_maj_98_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_98_n21) );
  NAND2_X1 cor_maj_98_U10 ( .A1(cor_maj_98_n21), .A2(cor_maj_98_n20), .ZN(
        cor_maj_98_n23) );
  XOR2_X1 cor_maj_98_U9 ( .A(v_1_0_3[2]), .B(cor_maj_98_n24), .Z(
        cor_maj_98_n26) );
  XOR2_X1 cor_maj_98_U8 ( .A(v_1_0_3[5]), .B(cor_maj_98_n25), .Z(
        cor_maj_98_n27) );
  XOR2_X1 cor_maj_98_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_98_n24)
         );
  XOR2_X1 cor_maj_98_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_98_n25)
         );
  OR2_X1 cor_maj_98_U5 ( .A1(cor_maj_98_n23), .A2(cor_maj_98_n22), .ZN(
        cor_maj_98_n32) );
  NAND2_X1 cor_maj_98_U4 ( .A1(cor_maj_98_n22), .A2(cor_maj_98_n23), .ZN(
        cor_maj_98_n34) );
  NAND2_X1 cor_maj_98_U3 ( .A1(cor_maj_98_n32), .A2(cor_maj_98_n31), .ZN(
        cor_maj_98_n33) );
  NAND2_X1 cor_maj_98_U2 ( .A1(cor_maj_98_n34), .A2(cor_maj_98_n33), .ZN(
        cor_maj_98_port_o) );
  OR2_X1 cor_maj_99_U19 ( .A1(cor_maj_99_n27), .A2(cor_maj_99_n26), .ZN(
        cor_maj_99_n28) );
  NAND2_X1 cor_maj_99_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_99_n28), .ZN(
        cor_maj_99_n29) );
  NAND2_X1 cor_maj_99_U17 ( .A1(cor_maj_99_n26), .A2(cor_maj_99_n27), .ZN(
        cor_maj_99_n30) );
  NAND2_X1 cor_maj_99_U16 ( .A1(cor_maj_99_n30), .A2(cor_maj_99_n29), .ZN(
        cor_maj_99_n31) );
  NAND2_X1 cor_maj_99_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_99_n25), .ZN(
        cor_maj_99_n18) );
  NAND2_X1 cor_maj_99_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_99_n19) );
  NAND2_X1 cor_maj_99_U13 ( .A1(cor_maj_99_n19), .A2(cor_maj_99_n18), .ZN(
        cor_maj_99_n22) );
  NAND2_X1 cor_maj_99_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_99_n24), .ZN(
        cor_maj_99_n20) );
  NAND2_X1 cor_maj_99_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_99_n21) );
  NAND2_X1 cor_maj_99_U10 ( .A1(cor_maj_99_n21), .A2(cor_maj_99_n20), .ZN(
        cor_maj_99_n23) );
  XOR2_X1 cor_maj_99_U9 ( .A(v_1_0_3[2]), .B(cor_maj_99_n24), .Z(
        cor_maj_99_n26) );
  XOR2_X1 cor_maj_99_U8 ( .A(v_1_0_3[5]), .B(cor_maj_99_n25), .Z(
        cor_maj_99_n27) );
  XOR2_X1 cor_maj_99_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_99_n24)
         );
  XOR2_X1 cor_maj_99_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_99_n25)
         );
  OR2_X1 cor_maj_99_U5 ( .A1(cor_maj_99_n23), .A2(cor_maj_99_n22), .ZN(
        cor_maj_99_n32) );
  NAND2_X1 cor_maj_99_U4 ( .A1(cor_maj_99_n22), .A2(cor_maj_99_n23), .ZN(
        cor_maj_99_n34) );
  NAND2_X1 cor_maj_99_U3 ( .A1(cor_maj_99_n32), .A2(cor_maj_99_n31), .ZN(
        cor_maj_99_n33) );
  NAND2_X1 cor_maj_99_U2 ( .A1(cor_maj_99_n34), .A2(cor_maj_99_n33), .ZN(
        cor_maj_99_port_o) );
  OR2_X1 cor_maj_100_U19 ( .A1(cor_maj_100_n27), .A2(cor_maj_100_n26), .ZN(
        cor_maj_100_n28) );
  NAND2_X1 cor_maj_100_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_100_n28), .ZN(
        cor_maj_100_n29) );
  NAND2_X1 cor_maj_100_U17 ( .A1(cor_maj_100_n26), .A2(cor_maj_100_n27), .ZN(
        cor_maj_100_n30) );
  NAND2_X1 cor_maj_100_U16 ( .A1(cor_maj_100_n30), .A2(cor_maj_100_n29), .ZN(
        cor_maj_100_n31) );
  NAND2_X1 cor_maj_100_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_100_n25), .ZN(
        cor_maj_100_n18) );
  NAND2_X1 cor_maj_100_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_100_n19) );
  NAND2_X1 cor_maj_100_U13 ( .A1(cor_maj_100_n19), .A2(cor_maj_100_n18), .ZN(
        cor_maj_100_n22) );
  NAND2_X1 cor_maj_100_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_100_n24), .ZN(
        cor_maj_100_n20) );
  NAND2_X1 cor_maj_100_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_100_n21) );
  NAND2_X1 cor_maj_100_U10 ( .A1(cor_maj_100_n21), .A2(cor_maj_100_n20), .ZN(
        cor_maj_100_n23) );
  XOR2_X1 cor_maj_100_U9 ( .A(v_1_0_3[2]), .B(cor_maj_100_n24), .Z(
        cor_maj_100_n26) );
  XOR2_X1 cor_maj_100_U8 ( .A(v_1_0_3[5]), .B(cor_maj_100_n25), .Z(
        cor_maj_100_n27) );
  XOR2_X1 cor_maj_100_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_100_n24)
         );
  XOR2_X1 cor_maj_100_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_100_n25)
         );
  OR2_X1 cor_maj_100_U5 ( .A1(cor_maj_100_n23), .A2(cor_maj_100_n22), .ZN(
        cor_maj_100_n32) );
  NAND2_X1 cor_maj_100_U4 ( .A1(cor_maj_100_n22), .A2(cor_maj_100_n23), .ZN(
        cor_maj_100_n34) );
  NAND2_X1 cor_maj_100_U3 ( .A1(cor_maj_100_n32), .A2(cor_maj_100_n31), .ZN(
        cor_maj_100_n33) );
  NAND2_X1 cor_maj_100_U2 ( .A1(cor_maj_100_n34), .A2(cor_maj_100_n33), .ZN(
        cor_maj_100_port_o) );
  OR2_X1 cor_maj_101_U19 ( .A1(cor_maj_101_n27), .A2(cor_maj_101_n26), .ZN(
        cor_maj_101_n28) );
  NAND2_X1 cor_maj_101_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_101_n28), .ZN(
        cor_maj_101_n29) );
  NAND2_X1 cor_maj_101_U17 ( .A1(cor_maj_101_n26), .A2(cor_maj_101_n27), .ZN(
        cor_maj_101_n30) );
  NAND2_X1 cor_maj_101_U16 ( .A1(cor_maj_101_n30), .A2(cor_maj_101_n29), .ZN(
        cor_maj_101_n31) );
  NAND2_X1 cor_maj_101_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_101_n25), .ZN(
        cor_maj_101_n18) );
  NAND2_X1 cor_maj_101_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_101_n19) );
  NAND2_X1 cor_maj_101_U13 ( .A1(cor_maj_101_n19), .A2(cor_maj_101_n18), .ZN(
        cor_maj_101_n22) );
  NAND2_X1 cor_maj_101_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_101_n24), .ZN(
        cor_maj_101_n20) );
  NAND2_X1 cor_maj_101_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_101_n21) );
  NAND2_X1 cor_maj_101_U10 ( .A1(cor_maj_101_n21), .A2(cor_maj_101_n20), .ZN(
        cor_maj_101_n23) );
  XOR2_X1 cor_maj_101_U9 ( .A(v_1_0_3[2]), .B(cor_maj_101_n24), .Z(
        cor_maj_101_n26) );
  XOR2_X1 cor_maj_101_U8 ( .A(v_1_0_3[5]), .B(cor_maj_101_n25), .Z(
        cor_maj_101_n27) );
  XOR2_X1 cor_maj_101_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_101_n24)
         );
  XOR2_X1 cor_maj_101_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_101_n25)
         );
  OR2_X1 cor_maj_101_U5 ( .A1(cor_maj_101_n23), .A2(cor_maj_101_n22), .ZN(
        cor_maj_101_n32) );
  NAND2_X1 cor_maj_101_U4 ( .A1(cor_maj_101_n22), .A2(cor_maj_101_n23), .ZN(
        cor_maj_101_n34) );
  NAND2_X1 cor_maj_101_U3 ( .A1(cor_maj_101_n32), .A2(cor_maj_101_n31), .ZN(
        cor_maj_101_n33) );
  NAND2_X1 cor_maj_101_U2 ( .A1(cor_maj_101_n34), .A2(cor_maj_101_n33), .ZN(
        cor_maj_101_port_o) );
  OR2_X1 cor_maj_102_U19 ( .A1(cor_maj_102_n27), .A2(cor_maj_102_n26), .ZN(
        cor_maj_102_n28) );
  NAND2_X1 cor_maj_102_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_102_n28), .ZN(
        cor_maj_102_n29) );
  NAND2_X1 cor_maj_102_U17 ( .A1(cor_maj_102_n26), .A2(cor_maj_102_n27), .ZN(
        cor_maj_102_n30) );
  NAND2_X1 cor_maj_102_U16 ( .A1(cor_maj_102_n30), .A2(cor_maj_102_n29), .ZN(
        cor_maj_102_n31) );
  NAND2_X1 cor_maj_102_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_102_n25), .ZN(
        cor_maj_102_n18) );
  NAND2_X1 cor_maj_102_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_102_n19) );
  NAND2_X1 cor_maj_102_U13 ( .A1(cor_maj_102_n19), .A2(cor_maj_102_n18), .ZN(
        cor_maj_102_n22) );
  NAND2_X1 cor_maj_102_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_102_n24), .ZN(
        cor_maj_102_n20) );
  NAND2_X1 cor_maj_102_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_102_n21) );
  NAND2_X1 cor_maj_102_U10 ( .A1(cor_maj_102_n21), .A2(cor_maj_102_n20), .ZN(
        cor_maj_102_n23) );
  XOR2_X1 cor_maj_102_U9 ( .A(v_1_0_3[2]), .B(cor_maj_102_n24), .Z(
        cor_maj_102_n26) );
  XOR2_X1 cor_maj_102_U8 ( .A(v_1_0_3[5]), .B(cor_maj_102_n25), .Z(
        cor_maj_102_n27) );
  XOR2_X1 cor_maj_102_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_102_n24)
         );
  XOR2_X1 cor_maj_102_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_102_n25)
         );
  OR2_X1 cor_maj_102_U5 ( .A1(cor_maj_102_n23), .A2(cor_maj_102_n22), .ZN(
        cor_maj_102_n32) );
  NAND2_X1 cor_maj_102_U4 ( .A1(cor_maj_102_n22), .A2(cor_maj_102_n23), .ZN(
        cor_maj_102_n34) );
  NAND2_X1 cor_maj_102_U3 ( .A1(cor_maj_102_n32), .A2(cor_maj_102_n31), .ZN(
        cor_maj_102_n33) );
  NAND2_X1 cor_maj_102_U2 ( .A1(cor_maj_102_n34), .A2(cor_maj_102_n33), .ZN(
        cor_maj_102_port_o) );
  OR2_X1 cor_maj_103_U19 ( .A1(cor_maj_103_n27), .A2(cor_maj_103_n26), .ZN(
        cor_maj_103_n28) );
  NAND2_X1 cor_maj_103_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_103_n28), .ZN(
        cor_maj_103_n29) );
  NAND2_X1 cor_maj_103_U17 ( .A1(cor_maj_103_n26), .A2(cor_maj_103_n27), .ZN(
        cor_maj_103_n30) );
  NAND2_X1 cor_maj_103_U16 ( .A1(cor_maj_103_n30), .A2(cor_maj_103_n29), .ZN(
        cor_maj_103_n31) );
  NAND2_X1 cor_maj_103_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_103_n25), .ZN(
        cor_maj_103_n18) );
  NAND2_X1 cor_maj_103_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_103_n19) );
  NAND2_X1 cor_maj_103_U13 ( .A1(cor_maj_103_n19), .A2(cor_maj_103_n18), .ZN(
        cor_maj_103_n22) );
  NAND2_X1 cor_maj_103_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_103_n24), .ZN(
        cor_maj_103_n20) );
  NAND2_X1 cor_maj_103_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_103_n21) );
  NAND2_X1 cor_maj_103_U10 ( .A1(cor_maj_103_n21), .A2(cor_maj_103_n20), .ZN(
        cor_maj_103_n23) );
  XOR2_X1 cor_maj_103_U9 ( .A(v_1_0_3[2]), .B(cor_maj_103_n24), .Z(
        cor_maj_103_n26) );
  XOR2_X1 cor_maj_103_U8 ( .A(v_1_0_3[5]), .B(cor_maj_103_n25), .Z(
        cor_maj_103_n27) );
  XOR2_X1 cor_maj_103_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_103_n24)
         );
  XOR2_X1 cor_maj_103_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_103_n25)
         );
  OR2_X1 cor_maj_103_U5 ( .A1(cor_maj_103_n23), .A2(cor_maj_103_n22), .ZN(
        cor_maj_103_n32) );
  NAND2_X1 cor_maj_103_U4 ( .A1(cor_maj_103_n22), .A2(cor_maj_103_n23), .ZN(
        cor_maj_103_n34) );
  NAND2_X1 cor_maj_103_U3 ( .A1(cor_maj_103_n32), .A2(cor_maj_103_n31), .ZN(
        cor_maj_103_n33) );
  NAND2_X1 cor_maj_103_U2 ( .A1(cor_maj_103_n34), .A2(cor_maj_103_n33), .ZN(
        cor_maj_103_port_o) );
  OR2_X1 cor_maj_104_U19 ( .A1(cor_maj_104_n27), .A2(cor_maj_104_n26), .ZN(
        cor_maj_104_n28) );
  NAND2_X1 cor_maj_104_U18 ( .A1(v_1_0_3[6]), .A2(cor_maj_104_n28), .ZN(
        cor_maj_104_n29) );
  NAND2_X1 cor_maj_104_U17 ( .A1(cor_maj_104_n26), .A2(cor_maj_104_n27), .ZN(
        cor_maj_104_n30) );
  NAND2_X1 cor_maj_104_U16 ( .A1(cor_maj_104_n30), .A2(cor_maj_104_n29), .ZN(
        cor_maj_104_n31) );
  NAND2_X1 cor_maj_104_U15 ( .A1(v_1_0_3[5]), .A2(cor_maj_104_n25), .ZN(
        cor_maj_104_n18) );
  NAND2_X1 cor_maj_104_U14 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_104_n19) );
  NAND2_X1 cor_maj_104_U13 ( .A1(cor_maj_104_n19), .A2(cor_maj_104_n18), .ZN(
        cor_maj_104_n22) );
  NAND2_X1 cor_maj_104_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_104_n24), .ZN(
        cor_maj_104_n20) );
  NAND2_X1 cor_maj_104_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_104_n21) );
  NAND2_X1 cor_maj_104_U10 ( .A1(cor_maj_104_n21), .A2(cor_maj_104_n20), .ZN(
        cor_maj_104_n23) );
  XOR2_X1 cor_maj_104_U9 ( .A(v_1_0_3[2]), .B(cor_maj_104_n24), .Z(
        cor_maj_104_n26) );
  XOR2_X1 cor_maj_104_U8 ( .A(v_1_0_3[5]), .B(cor_maj_104_n25), .Z(
        cor_maj_104_n27) );
  XOR2_X1 cor_maj_104_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_104_n24)
         );
  XOR2_X1 cor_maj_104_U6 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_104_n25)
         );
  OR2_X1 cor_maj_104_U5 ( .A1(cor_maj_104_n23), .A2(cor_maj_104_n22), .ZN(
        cor_maj_104_n32) );
  NAND2_X1 cor_maj_104_U4 ( .A1(cor_maj_104_n22), .A2(cor_maj_104_n23), .ZN(
        cor_maj_104_n34) );
  NAND2_X1 cor_maj_104_U3 ( .A1(cor_maj_104_n32), .A2(cor_maj_104_n31), .ZN(
        cor_maj_104_n33) );
  NAND2_X1 cor_maj_104_U2 ( .A1(cor_maj_104_n34), .A2(cor_maj_104_n33), .ZN(
        cor_maj_104_port_o) );
  OR2_X1 cor_maj_105_U19 ( .A1(cor_maj_105_n27), .A2(cor_maj_105_n26), .ZN(
        cor_maj_105_n28) );
  NAND2_X1 cor_maj_105_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_105_n28), .ZN(
        cor_maj_105_n29) );
  NAND2_X1 cor_maj_105_U17 ( .A1(cor_maj_105_n26), .A2(cor_maj_105_n27), .ZN(
        cor_maj_105_n30) );
  NAND2_X1 cor_maj_105_U16 ( .A1(cor_maj_105_n30), .A2(cor_maj_105_n29), .ZN(
        cor_maj_105_n31) );
  NAND2_X1 cor_maj_105_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_105_n25), .ZN(
        cor_maj_105_n18) );
  NAND2_X1 cor_maj_105_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_105_n19) );
  NAND2_X1 cor_maj_105_U13 ( .A1(cor_maj_105_n19), .A2(cor_maj_105_n18), .ZN(
        cor_maj_105_n22) );
  NAND2_X1 cor_maj_105_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_105_n24), .ZN(
        cor_maj_105_n20) );
  NAND2_X1 cor_maj_105_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_105_n21) );
  NAND2_X1 cor_maj_105_U10 ( .A1(cor_maj_105_n21), .A2(cor_maj_105_n20), .ZN(
        cor_maj_105_n23) );
  XOR2_X1 cor_maj_105_U9 ( .A(v_1_1_0[2]), .B(cor_maj_105_n24), .Z(
        cor_maj_105_n26) );
  XOR2_X1 cor_maj_105_U8 ( .A(v_1_1_0[5]), .B(cor_maj_105_n25), .Z(
        cor_maj_105_n27) );
  XOR2_X1 cor_maj_105_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_105_n24)
         );
  XOR2_X1 cor_maj_105_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_105_n25)
         );
  OR2_X1 cor_maj_105_U5 ( .A1(cor_maj_105_n23), .A2(cor_maj_105_n22), .ZN(
        cor_maj_105_n32) );
  NAND2_X1 cor_maj_105_U4 ( .A1(cor_maj_105_n22), .A2(cor_maj_105_n23), .ZN(
        cor_maj_105_n34) );
  NAND2_X1 cor_maj_105_U3 ( .A1(cor_maj_105_n32), .A2(cor_maj_105_n31), .ZN(
        cor_maj_105_n33) );
  NAND2_X1 cor_maj_105_U2 ( .A1(cor_maj_105_n34), .A2(cor_maj_105_n33), .ZN(
        cor_maj_105_port_o) );
  OR2_X1 cor_maj_106_U19 ( .A1(cor_maj_106_n27), .A2(cor_maj_106_n26), .ZN(
        cor_maj_106_n28) );
  NAND2_X1 cor_maj_106_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_106_n28), .ZN(
        cor_maj_106_n29) );
  NAND2_X1 cor_maj_106_U17 ( .A1(cor_maj_106_n26), .A2(cor_maj_106_n27), .ZN(
        cor_maj_106_n30) );
  NAND2_X1 cor_maj_106_U16 ( .A1(cor_maj_106_n30), .A2(cor_maj_106_n29), .ZN(
        cor_maj_106_n31) );
  NAND2_X1 cor_maj_106_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_106_n25), .ZN(
        cor_maj_106_n18) );
  NAND2_X1 cor_maj_106_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_106_n19) );
  NAND2_X1 cor_maj_106_U13 ( .A1(cor_maj_106_n19), .A2(cor_maj_106_n18), .ZN(
        cor_maj_106_n22) );
  NAND2_X1 cor_maj_106_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_106_n24), .ZN(
        cor_maj_106_n20) );
  NAND2_X1 cor_maj_106_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_106_n21) );
  NAND2_X1 cor_maj_106_U10 ( .A1(cor_maj_106_n21), .A2(cor_maj_106_n20), .ZN(
        cor_maj_106_n23) );
  XOR2_X1 cor_maj_106_U9 ( .A(v_1_1_0[2]), .B(cor_maj_106_n24), .Z(
        cor_maj_106_n26) );
  XOR2_X1 cor_maj_106_U8 ( .A(v_1_1_0[5]), .B(cor_maj_106_n25), .Z(
        cor_maj_106_n27) );
  XOR2_X1 cor_maj_106_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_106_n24)
         );
  XOR2_X1 cor_maj_106_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_106_n25)
         );
  OR2_X1 cor_maj_106_U5 ( .A1(cor_maj_106_n23), .A2(cor_maj_106_n22), .ZN(
        cor_maj_106_n32) );
  NAND2_X1 cor_maj_106_U4 ( .A1(cor_maj_106_n22), .A2(cor_maj_106_n23), .ZN(
        cor_maj_106_n34) );
  NAND2_X1 cor_maj_106_U3 ( .A1(cor_maj_106_n32), .A2(cor_maj_106_n31), .ZN(
        cor_maj_106_n33) );
  NAND2_X1 cor_maj_106_U2 ( .A1(cor_maj_106_n34), .A2(cor_maj_106_n33), .ZN(
        cor_maj_106_port_o) );
  OR2_X1 cor_maj_107_U19 ( .A1(cor_maj_107_n27), .A2(cor_maj_107_n26), .ZN(
        cor_maj_107_n28) );
  NAND2_X1 cor_maj_107_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_107_n28), .ZN(
        cor_maj_107_n29) );
  NAND2_X1 cor_maj_107_U17 ( .A1(cor_maj_107_n26), .A2(cor_maj_107_n27), .ZN(
        cor_maj_107_n30) );
  NAND2_X1 cor_maj_107_U16 ( .A1(cor_maj_107_n30), .A2(cor_maj_107_n29), .ZN(
        cor_maj_107_n31) );
  NAND2_X1 cor_maj_107_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_107_n25), .ZN(
        cor_maj_107_n18) );
  NAND2_X1 cor_maj_107_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_107_n19) );
  NAND2_X1 cor_maj_107_U13 ( .A1(cor_maj_107_n19), .A2(cor_maj_107_n18), .ZN(
        cor_maj_107_n22) );
  NAND2_X1 cor_maj_107_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_107_n24), .ZN(
        cor_maj_107_n20) );
  NAND2_X1 cor_maj_107_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_107_n21) );
  NAND2_X1 cor_maj_107_U10 ( .A1(cor_maj_107_n21), .A2(cor_maj_107_n20), .ZN(
        cor_maj_107_n23) );
  XOR2_X1 cor_maj_107_U9 ( .A(v_1_1_0[2]), .B(cor_maj_107_n24), .Z(
        cor_maj_107_n26) );
  XOR2_X1 cor_maj_107_U8 ( .A(v_1_1_0[5]), .B(cor_maj_107_n25), .Z(
        cor_maj_107_n27) );
  XOR2_X1 cor_maj_107_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_107_n24)
         );
  XOR2_X1 cor_maj_107_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_107_n25)
         );
  OR2_X1 cor_maj_107_U5 ( .A1(cor_maj_107_n23), .A2(cor_maj_107_n22), .ZN(
        cor_maj_107_n32) );
  NAND2_X1 cor_maj_107_U4 ( .A1(cor_maj_107_n22), .A2(cor_maj_107_n23), .ZN(
        cor_maj_107_n34) );
  NAND2_X1 cor_maj_107_U3 ( .A1(cor_maj_107_n32), .A2(cor_maj_107_n31), .ZN(
        cor_maj_107_n33) );
  NAND2_X1 cor_maj_107_U2 ( .A1(cor_maj_107_n34), .A2(cor_maj_107_n33), .ZN(
        cor_maj_107_port_o) );
  OR2_X1 cor_maj_108_U19 ( .A1(cor_maj_108_n27), .A2(cor_maj_108_n26), .ZN(
        cor_maj_108_n28) );
  NAND2_X1 cor_maj_108_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_108_n28), .ZN(
        cor_maj_108_n29) );
  NAND2_X1 cor_maj_108_U17 ( .A1(cor_maj_108_n26), .A2(cor_maj_108_n27), .ZN(
        cor_maj_108_n30) );
  NAND2_X1 cor_maj_108_U16 ( .A1(cor_maj_108_n30), .A2(cor_maj_108_n29), .ZN(
        cor_maj_108_n31) );
  NAND2_X1 cor_maj_108_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_108_n25), .ZN(
        cor_maj_108_n18) );
  NAND2_X1 cor_maj_108_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_108_n19) );
  NAND2_X1 cor_maj_108_U13 ( .A1(cor_maj_108_n19), .A2(cor_maj_108_n18), .ZN(
        cor_maj_108_n22) );
  NAND2_X1 cor_maj_108_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_108_n24), .ZN(
        cor_maj_108_n20) );
  NAND2_X1 cor_maj_108_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_108_n21) );
  NAND2_X1 cor_maj_108_U10 ( .A1(cor_maj_108_n21), .A2(cor_maj_108_n20), .ZN(
        cor_maj_108_n23) );
  XOR2_X1 cor_maj_108_U9 ( .A(v_1_1_0[2]), .B(cor_maj_108_n24), .Z(
        cor_maj_108_n26) );
  XOR2_X1 cor_maj_108_U8 ( .A(v_1_1_0[5]), .B(cor_maj_108_n25), .Z(
        cor_maj_108_n27) );
  XOR2_X1 cor_maj_108_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_108_n24)
         );
  XOR2_X1 cor_maj_108_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_108_n25)
         );
  OR2_X1 cor_maj_108_U5 ( .A1(cor_maj_108_n23), .A2(cor_maj_108_n22), .ZN(
        cor_maj_108_n32) );
  NAND2_X1 cor_maj_108_U4 ( .A1(cor_maj_108_n22), .A2(cor_maj_108_n23), .ZN(
        cor_maj_108_n34) );
  NAND2_X1 cor_maj_108_U3 ( .A1(cor_maj_108_n32), .A2(cor_maj_108_n31), .ZN(
        cor_maj_108_n33) );
  NAND2_X1 cor_maj_108_U2 ( .A1(cor_maj_108_n34), .A2(cor_maj_108_n33), .ZN(
        cor_maj_108_port_o) );
  OR2_X1 cor_maj_109_U19 ( .A1(cor_maj_109_n27), .A2(cor_maj_109_n26), .ZN(
        cor_maj_109_n28) );
  NAND2_X1 cor_maj_109_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_109_n28), .ZN(
        cor_maj_109_n29) );
  NAND2_X1 cor_maj_109_U17 ( .A1(cor_maj_109_n26), .A2(cor_maj_109_n27), .ZN(
        cor_maj_109_n30) );
  NAND2_X1 cor_maj_109_U16 ( .A1(cor_maj_109_n30), .A2(cor_maj_109_n29), .ZN(
        cor_maj_109_n31) );
  NAND2_X1 cor_maj_109_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_109_n25), .ZN(
        cor_maj_109_n18) );
  NAND2_X1 cor_maj_109_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_109_n19) );
  NAND2_X1 cor_maj_109_U13 ( .A1(cor_maj_109_n19), .A2(cor_maj_109_n18), .ZN(
        cor_maj_109_n22) );
  NAND2_X1 cor_maj_109_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_109_n24), .ZN(
        cor_maj_109_n20) );
  NAND2_X1 cor_maj_109_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_109_n21) );
  NAND2_X1 cor_maj_109_U10 ( .A1(cor_maj_109_n21), .A2(cor_maj_109_n20), .ZN(
        cor_maj_109_n23) );
  XOR2_X1 cor_maj_109_U9 ( .A(v_1_1_0[2]), .B(cor_maj_109_n24), .Z(
        cor_maj_109_n26) );
  XOR2_X1 cor_maj_109_U8 ( .A(v_1_1_0[5]), .B(cor_maj_109_n25), .Z(
        cor_maj_109_n27) );
  XOR2_X1 cor_maj_109_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_109_n24)
         );
  XOR2_X1 cor_maj_109_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_109_n25)
         );
  OR2_X1 cor_maj_109_U5 ( .A1(cor_maj_109_n23), .A2(cor_maj_109_n22), .ZN(
        cor_maj_109_n32) );
  NAND2_X1 cor_maj_109_U4 ( .A1(cor_maj_109_n22), .A2(cor_maj_109_n23), .ZN(
        cor_maj_109_n34) );
  NAND2_X1 cor_maj_109_U3 ( .A1(cor_maj_109_n32), .A2(cor_maj_109_n31), .ZN(
        cor_maj_109_n33) );
  NAND2_X1 cor_maj_109_U2 ( .A1(cor_maj_109_n34), .A2(cor_maj_109_n33), .ZN(
        cor_maj_109_port_o) );
  OR2_X1 cor_maj_110_U19 ( .A1(cor_maj_110_n27), .A2(cor_maj_110_n26), .ZN(
        cor_maj_110_n28) );
  NAND2_X1 cor_maj_110_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_110_n28), .ZN(
        cor_maj_110_n29) );
  NAND2_X1 cor_maj_110_U17 ( .A1(cor_maj_110_n26), .A2(cor_maj_110_n27), .ZN(
        cor_maj_110_n30) );
  NAND2_X1 cor_maj_110_U16 ( .A1(cor_maj_110_n30), .A2(cor_maj_110_n29), .ZN(
        cor_maj_110_n31) );
  NAND2_X1 cor_maj_110_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_110_n25), .ZN(
        cor_maj_110_n18) );
  NAND2_X1 cor_maj_110_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_110_n19) );
  NAND2_X1 cor_maj_110_U13 ( .A1(cor_maj_110_n19), .A2(cor_maj_110_n18), .ZN(
        cor_maj_110_n22) );
  NAND2_X1 cor_maj_110_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_110_n24), .ZN(
        cor_maj_110_n20) );
  NAND2_X1 cor_maj_110_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_110_n21) );
  NAND2_X1 cor_maj_110_U10 ( .A1(cor_maj_110_n21), .A2(cor_maj_110_n20), .ZN(
        cor_maj_110_n23) );
  XOR2_X1 cor_maj_110_U9 ( .A(v_1_1_0[2]), .B(cor_maj_110_n24), .Z(
        cor_maj_110_n26) );
  XOR2_X1 cor_maj_110_U8 ( .A(v_1_1_0[5]), .B(cor_maj_110_n25), .Z(
        cor_maj_110_n27) );
  XOR2_X1 cor_maj_110_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_110_n24)
         );
  XOR2_X1 cor_maj_110_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_110_n25)
         );
  OR2_X1 cor_maj_110_U5 ( .A1(cor_maj_110_n23), .A2(cor_maj_110_n22), .ZN(
        cor_maj_110_n32) );
  NAND2_X1 cor_maj_110_U4 ( .A1(cor_maj_110_n22), .A2(cor_maj_110_n23), .ZN(
        cor_maj_110_n34) );
  NAND2_X1 cor_maj_110_U3 ( .A1(cor_maj_110_n32), .A2(cor_maj_110_n31), .ZN(
        cor_maj_110_n33) );
  NAND2_X1 cor_maj_110_U2 ( .A1(cor_maj_110_n34), .A2(cor_maj_110_n33), .ZN(
        cor_maj_110_port_o) );
  OR2_X1 cor_maj_111_U19 ( .A1(cor_maj_111_n27), .A2(cor_maj_111_n26), .ZN(
        cor_maj_111_n28) );
  NAND2_X1 cor_maj_111_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_111_n28), .ZN(
        cor_maj_111_n29) );
  NAND2_X1 cor_maj_111_U17 ( .A1(cor_maj_111_n26), .A2(cor_maj_111_n27), .ZN(
        cor_maj_111_n30) );
  NAND2_X1 cor_maj_111_U16 ( .A1(cor_maj_111_n30), .A2(cor_maj_111_n29), .ZN(
        cor_maj_111_n31) );
  NAND2_X1 cor_maj_111_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_111_n25), .ZN(
        cor_maj_111_n18) );
  NAND2_X1 cor_maj_111_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_111_n19) );
  NAND2_X1 cor_maj_111_U13 ( .A1(cor_maj_111_n19), .A2(cor_maj_111_n18), .ZN(
        cor_maj_111_n22) );
  NAND2_X1 cor_maj_111_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_111_n24), .ZN(
        cor_maj_111_n20) );
  NAND2_X1 cor_maj_111_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_111_n21) );
  NAND2_X1 cor_maj_111_U10 ( .A1(cor_maj_111_n21), .A2(cor_maj_111_n20), .ZN(
        cor_maj_111_n23) );
  XOR2_X1 cor_maj_111_U9 ( .A(v_1_1_0[2]), .B(cor_maj_111_n24), .Z(
        cor_maj_111_n26) );
  XOR2_X1 cor_maj_111_U8 ( .A(v_1_1_0[5]), .B(cor_maj_111_n25), .Z(
        cor_maj_111_n27) );
  XOR2_X1 cor_maj_111_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_111_n24)
         );
  XOR2_X1 cor_maj_111_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_111_n25)
         );
  OR2_X1 cor_maj_111_U5 ( .A1(cor_maj_111_n23), .A2(cor_maj_111_n22), .ZN(
        cor_maj_111_n32) );
  NAND2_X1 cor_maj_111_U4 ( .A1(cor_maj_111_n22), .A2(cor_maj_111_n23), .ZN(
        cor_maj_111_n34) );
  NAND2_X1 cor_maj_111_U3 ( .A1(cor_maj_111_n32), .A2(cor_maj_111_n31), .ZN(
        cor_maj_111_n33) );
  NAND2_X1 cor_maj_111_U2 ( .A1(cor_maj_111_n34), .A2(cor_maj_111_n33), .ZN(
        cor_maj_111_port_o) );
  OR2_X1 cor_maj_112_U19 ( .A1(cor_maj_112_n27), .A2(cor_maj_112_n26), .ZN(
        cor_maj_112_n28) );
  NAND2_X1 cor_maj_112_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_112_n28), .ZN(
        cor_maj_112_n29) );
  NAND2_X1 cor_maj_112_U17 ( .A1(cor_maj_112_n26), .A2(cor_maj_112_n27), .ZN(
        cor_maj_112_n30) );
  NAND2_X1 cor_maj_112_U16 ( .A1(cor_maj_112_n30), .A2(cor_maj_112_n29), .ZN(
        cor_maj_112_n31) );
  NAND2_X1 cor_maj_112_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_112_n25), .ZN(
        cor_maj_112_n18) );
  NAND2_X1 cor_maj_112_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_112_n19) );
  NAND2_X1 cor_maj_112_U13 ( .A1(cor_maj_112_n19), .A2(cor_maj_112_n18), .ZN(
        cor_maj_112_n22) );
  NAND2_X1 cor_maj_112_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_112_n24), .ZN(
        cor_maj_112_n20) );
  NAND2_X1 cor_maj_112_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_112_n21) );
  NAND2_X1 cor_maj_112_U10 ( .A1(cor_maj_112_n21), .A2(cor_maj_112_n20), .ZN(
        cor_maj_112_n23) );
  XOR2_X1 cor_maj_112_U9 ( .A(v_1_1_2[2]), .B(cor_maj_112_n24), .Z(
        cor_maj_112_n26) );
  XOR2_X1 cor_maj_112_U8 ( .A(v_1_1_2[5]), .B(cor_maj_112_n25), .Z(
        cor_maj_112_n27) );
  XOR2_X1 cor_maj_112_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_112_n24)
         );
  XOR2_X1 cor_maj_112_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_112_n25)
         );
  OR2_X1 cor_maj_112_U5 ( .A1(cor_maj_112_n23), .A2(cor_maj_112_n22), .ZN(
        cor_maj_112_n32) );
  NAND2_X1 cor_maj_112_U4 ( .A1(cor_maj_112_n22), .A2(cor_maj_112_n23), .ZN(
        cor_maj_112_n34) );
  NAND2_X1 cor_maj_112_U3 ( .A1(cor_maj_112_n32), .A2(cor_maj_112_n31), .ZN(
        cor_maj_112_n33) );
  NAND2_X1 cor_maj_112_U2 ( .A1(cor_maj_112_n34), .A2(cor_maj_112_n33), .ZN(
        cor_maj_112_port_o) );
  OR2_X1 cor_maj_113_U19 ( .A1(cor_maj_113_n27), .A2(cor_maj_113_n26), .ZN(
        cor_maj_113_n28) );
  NAND2_X1 cor_maj_113_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_113_n28), .ZN(
        cor_maj_113_n29) );
  NAND2_X1 cor_maj_113_U17 ( .A1(cor_maj_113_n26), .A2(cor_maj_113_n27), .ZN(
        cor_maj_113_n30) );
  NAND2_X1 cor_maj_113_U16 ( .A1(cor_maj_113_n30), .A2(cor_maj_113_n29), .ZN(
        cor_maj_113_n31) );
  NAND2_X1 cor_maj_113_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_113_n25), .ZN(
        cor_maj_113_n18) );
  NAND2_X1 cor_maj_113_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_113_n19) );
  NAND2_X1 cor_maj_113_U13 ( .A1(cor_maj_113_n19), .A2(cor_maj_113_n18), .ZN(
        cor_maj_113_n22) );
  NAND2_X1 cor_maj_113_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_113_n24), .ZN(
        cor_maj_113_n20) );
  NAND2_X1 cor_maj_113_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_113_n21) );
  NAND2_X1 cor_maj_113_U10 ( .A1(cor_maj_113_n21), .A2(cor_maj_113_n20), .ZN(
        cor_maj_113_n23) );
  XOR2_X1 cor_maj_113_U9 ( .A(v_1_1_2[2]), .B(cor_maj_113_n24), .Z(
        cor_maj_113_n26) );
  XOR2_X1 cor_maj_113_U8 ( .A(v_1_1_2[5]), .B(cor_maj_113_n25), .Z(
        cor_maj_113_n27) );
  XOR2_X1 cor_maj_113_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_113_n24)
         );
  XOR2_X1 cor_maj_113_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_113_n25)
         );
  OR2_X1 cor_maj_113_U5 ( .A1(cor_maj_113_n23), .A2(cor_maj_113_n22), .ZN(
        cor_maj_113_n32) );
  NAND2_X1 cor_maj_113_U4 ( .A1(cor_maj_113_n22), .A2(cor_maj_113_n23), .ZN(
        cor_maj_113_n34) );
  NAND2_X1 cor_maj_113_U3 ( .A1(cor_maj_113_n32), .A2(cor_maj_113_n31), .ZN(
        cor_maj_113_n33) );
  NAND2_X1 cor_maj_113_U2 ( .A1(cor_maj_113_n34), .A2(cor_maj_113_n33), .ZN(
        cor_maj_113_port_o) );
  OR2_X1 cor_maj_114_U19 ( .A1(cor_maj_114_n27), .A2(cor_maj_114_n26), .ZN(
        cor_maj_114_n28) );
  NAND2_X1 cor_maj_114_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_114_n28), .ZN(
        cor_maj_114_n29) );
  NAND2_X1 cor_maj_114_U17 ( .A1(cor_maj_114_n26), .A2(cor_maj_114_n27), .ZN(
        cor_maj_114_n30) );
  NAND2_X1 cor_maj_114_U16 ( .A1(cor_maj_114_n30), .A2(cor_maj_114_n29), .ZN(
        cor_maj_114_n31) );
  NAND2_X1 cor_maj_114_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_114_n25), .ZN(
        cor_maj_114_n18) );
  NAND2_X1 cor_maj_114_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_114_n19) );
  NAND2_X1 cor_maj_114_U13 ( .A1(cor_maj_114_n19), .A2(cor_maj_114_n18), .ZN(
        cor_maj_114_n22) );
  NAND2_X1 cor_maj_114_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_114_n24), .ZN(
        cor_maj_114_n20) );
  NAND2_X1 cor_maj_114_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_114_n21) );
  NAND2_X1 cor_maj_114_U10 ( .A1(cor_maj_114_n21), .A2(cor_maj_114_n20), .ZN(
        cor_maj_114_n23) );
  XOR2_X1 cor_maj_114_U9 ( .A(v_1_1_2[2]), .B(cor_maj_114_n24), .Z(
        cor_maj_114_n26) );
  XOR2_X1 cor_maj_114_U8 ( .A(v_1_1_2[5]), .B(cor_maj_114_n25), .Z(
        cor_maj_114_n27) );
  XOR2_X1 cor_maj_114_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_114_n24)
         );
  XOR2_X1 cor_maj_114_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_114_n25)
         );
  OR2_X1 cor_maj_114_U5 ( .A1(cor_maj_114_n23), .A2(cor_maj_114_n22), .ZN(
        cor_maj_114_n32) );
  NAND2_X1 cor_maj_114_U4 ( .A1(cor_maj_114_n22), .A2(cor_maj_114_n23), .ZN(
        cor_maj_114_n34) );
  NAND2_X1 cor_maj_114_U3 ( .A1(cor_maj_114_n32), .A2(cor_maj_114_n31), .ZN(
        cor_maj_114_n33) );
  NAND2_X1 cor_maj_114_U2 ( .A1(cor_maj_114_n34), .A2(cor_maj_114_n33), .ZN(
        cor_maj_114_port_o) );
  OR2_X1 cor_maj_115_U19 ( .A1(cor_maj_115_n27), .A2(cor_maj_115_n26), .ZN(
        cor_maj_115_n28) );
  NAND2_X1 cor_maj_115_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_115_n28), .ZN(
        cor_maj_115_n29) );
  NAND2_X1 cor_maj_115_U17 ( .A1(cor_maj_115_n26), .A2(cor_maj_115_n27), .ZN(
        cor_maj_115_n30) );
  NAND2_X1 cor_maj_115_U16 ( .A1(cor_maj_115_n30), .A2(cor_maj_115_n29), .ZN(
        cor_maj_115_n31) );
  NAND2_X1 cor_maj_115_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_115_n25), .ZN(
        cor_maj_115_n18) );
  NAND2_X1 cor_maj_115_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_115_n19) );
  NAND2_X1 cor_maj_115_U13 ( .A1(cor_maj_115_n19), .A2(cor_maj_115_n18), .ZN(
        cor_maj_115_n22) );
  NAND2_X1 cor_maj_115_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_115_n24), .ZN(
        cor_maj_115_n20) );
  NAND2_X1 cor_maj_115_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_115_n21) );
  NAND2_X1 cor_maj_115_U10 ( .A1(cor_maj_115_n21), .A2(cor_maj_115_n20), .ZN(
        cor_maj_115_n23) );
  XOR2_X1 cor_maj_115_U9 ( .A(v_1_1_2[2]), .B(cor_maj_115_n24), .Z(
        cor_maj_115_n26) );
  XOR2_X1 cor_maj_115_U8 ( .A(v_1_1_2[5]), .B(cor_maj_115_n25), .Z(
        cor_maj_115_n27) );
  XOR2_X1 cor_maj_115_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_115_n24)
         );
  XOR2_X1 cor_maj_115_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_115_n25)
         );
  OR2_X1 cor_maj_115_U5 ( .A1(cor_maj_115_n23), .A2(cor_maj_115_n22), .ZN(
        cor_maj_115_n32) );
  NAND2_X1 cor_maj_115_U4 ( .A1(cor_maj_115_n22), .A2(cor_maj_115_n23), .ZN(
        cor_maj_115_n34) );
  NAND2_X1 cor_maj_115_U3 ( .A1(cor_maj_115_n32), .A2(cor_maj_115_n31), .ZN(
        cor_maj_115_n33) );
  NAND2_X1 cor_maj_115_U2 ( .A1(cor_maj_115_n34), .A2(cor_maj_115_n33), .ZN(
        cor_maj_115_port_o) );
  OR2_X1 cor_maj_116_U19 ( .A1(cor_maj_116_n27), .A2(cor_maj_116_n26), .ZN(
        cor_maj_116_n28) );
  NAND2_X1 cor_maj_116_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_116_n28), .ZN(
        cor_maj_116_n29) );
  NAND2_X1 cor_maj_116_U17 ( .A1(cor_maj_116_n26), .A2(cor_maj_116_n27), .ZN(
        cor_maj_116_n30) );
  NAND2_X1 cor_maj_116_U16 ( .A1(cor_maj_116_n30), .A2(cor_maj_116_n29), .ZN(
        cor_maj_116_n31) );
  NAND2_X1 cor_maj_116_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_116_n25), .ZN(
        cor_maj_116_n18) );
  NAND2_X1 cor_maj_116_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_116_n19) );
  NAND2_X1 cor_maj_116_U13 ( .A1(cor_maj_116_n19), .A2(cor_maj_116_n18), .ZN(
        cor_maj_116_n22) );
  NAND2_X1 cor_maj_116_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_116_n24), .ZN(
        cor_maj_116_n20) );
  NAND2_X1 cor_maj_116_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_116_n21) );
  NAND2_X1 cor_maj_116_U10 ( .A1(cor_maj_116_n21), .A2(cor_maj_116_n20), .ZN(
        cor_maj_116_n23) );
  XOR2_X1 cor_maj_116_U9 ( .A(v_1_1_2[2]), .B(cor_maj_116_n24), .Z(
        cor_maj_116_n26) );
  XOR2_X1 cor_maj_116_U8 ( .A(v_1_1_2[5]), .B(cor_maj_116_n25), .Z(
        cor_maj_116_n27) );
  XOR2_X1 cor_maj_116_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_116_n24)
         );
  XOR2_X1 cor_maj_116_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_116_n25)
         );
  OR2_X1 cor_maj_116_U5 ( .A1(cor_maj_116_n23), .A2(cor_maj_116_n22), .ZN(
        cor_maj_116_n32) );
  NAND2_X1 cor_maj_116_U4 ( .A1(cor_maj_116_n22), .A2(cor_maj_116_n23), .ZN(
        cor_maj_116_n34) );
  NAND2_X1 cor_maj_116_U3 ( .A1(cor_maj_116_n32), .A2(cor_maj_116_n31), .ZN(
        cor_maj_116_n33) );
  NAND2_X1 cor_maj_116_U2 ( .A1(cor_maj_116_n34), .A2(cor_maj_116_n33), .ZN(
        cor_maj_116_port_o) );
  OR2_X1 cor_maj_117_U19 ( .A1(cor_maj_117_n27), .A2(cor_maj_117_n26), .ZN(
        cor_maj_117_n28) );
  NAND2_X1 cor_maj_117_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_117_n28), .ZN(
        cor_maj_117_n29) );
  NAND2_X1 cor_maj_117_U17 ( .A1(cor_maj_117_n26), .A2(cor_maj_117_n27), .ZN(
        cor_maj_117_n30) );
  NAND2_X1 cor_maj_117_U16 ( .A1(cor_maj_117_n30), .A2(cor_maj_117_n29), .ZN(
        cor_maj_117_n31) );
  NAND2_X1 cor_maj_117_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_117_n25), .ZN(
        cor_maj_117_n18) );
  NAND2_X1 cor_maj_117_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_117_n19) );
  NAND2_X1 cor_maj_117_U13 ( .A1(cor_maj_117_n19), .A2(cor_maj_117_n18), .ZN(
        cor_maj_117_n22) );
  NAND2_X1 cor_maj_117_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_117_n24), .ZN(
        cor_maj_117_n20) );
  NAND2_X1 cor_maj_117_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_117_n21) );
  NAND2_X1 cor_maj_117_U10 ( .A1(cor_maj_117_n21), .A2(cor_maj_117_n20), .ZN(
        cor_maj_117_n23) );
  XOR2_X1 cor_maj_117_U9 ( .A(v_1_1_2[2]), .B(cor_maj_117_n24), .Z(
        cor_maj_117_n26) );
  XOR2_X1 cor_maj_117_U8 ( .A(v_1_1_2[5]), .B(cor_maj_117_n25), .Z(
        cor_maj_117_n27) );
  XOR2_X1 cor_maj_117_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_117_n24)
         );
  XOR2_X1 cor_maj_117_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_117_n25)
         );
  OR2_X1 cor_maj_117_U5 ( .A1(cor_maj_117_n23), .A2(cor_maj_117_n22), .ZN(
        cor_maj_117_n32) );
  NAND2_X1 cor_maj_117_U4 ( .A1(cor_maj_117_n22), .A2(cor_maj_117_n23), .ZN(
        cor_maj_117_n34) );
  NAND2_X1 cor_maj_117_U3 ( .A1(cor_maj_117_n32), .A2(cor_maj_117_n31), .ZN(
        cor_maj_117_n33) );
  NAND2_X1 cor_maj_117_U2 ( .A1(cor_maj_117_n34), .A2(cor_maj_117_n33), .ZN(
        cor_maj_117_port_o) );
  OR2_X1 cor_maj_118_U19 ( .A1(cor_maj_118_n27), .A2(cor_maj_118_n26), .ZN(
        cor_maj_118_n28) );
  NAND2_X1 cor_maj_118_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_118_n28), .ZN(
        cor_maj_118_n29) );
  NAND2_X1 cor_maj_118_U17 ( .A1(cor_maj_118_n26), .A2(cor_maj_118_n27), .ZN(
        cor_maj_118_n30) );
  NAND2_X1 cor_maj_118_U16 ( .A1(cor_maj_118_n30), .A2(cor_maj_118_n29), .ZN(
        cor_maj_118_n31) );
  NAND2_X1 cor_maj_118_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_118_n25), .ZN(
        cor_maj_118_n18) );
  NAND2_X1 cor_maj_118_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_118_n19) );
  NAND2_X1 cor_maj_118_U13 ( .A1(cor_maj_118_n19), .A2(cor_maj_118_n18), .ZN(
        cor_maj_118_n22) );
  NAND2_X1 cor_maj_118_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_118_n24), .ZN(
        cor_maj_118_n20) );
  NAND2_X1 cor_maj_118_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_118_n21) );
  NAND2_X1 cor_maj_118_U10 ( .A1(cor_maj_118_n21), .A2(cor_maj_118_n20), .ZN(
        cor_maj_118_n23) );
  XOR2_X1 cor_maj_118_U9 ( .A(v_1_1_2[2]), .B(cor_maj_118_n24), .Z(
        cor_maj_118_n26) );
  XOR2_X1 cor_maj_118_U8 ( .A(v_1_1_2[5]), .B(cor_maj_118_n25), .Z(
        cor_maj_118_n27) );
  XOR2_X1 cor_maj_118_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_118_n24)
         );
  XOR2_X1 cor_maj_118_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_118_n25)
         );
  OR2_X1 cor_maj_118_U5 ( .A1(cor_maj_118_n23), .A2(cor_maj_118_n22), .ZN(
        cor_maj_118_n32) );
  NAND2_X1 cor_maj_118_U4 ( .A1(cor_maj_118_n22), .A2(cor_maj_118_n23), .ZN(
        cor_maj_118_n34) );
  NAND2_X1 cor_maj_118_U3 ( .A1(cor_maj_118_n32), .A2(cor_maj_118_n31), .ZN(
        cor_maj_118_n33) );
  NAND2_X1 cor_maj_118_U2 ( .A1(cor_maj_118_n34), .A2(cor_maj_118_n33), .ZN(
        cor_maj_118_port_o) );
  OR2_X1 cor_maj_119_U19 ( .A1(cor_maj_119_n27), .A2(cor_maj_119_n26), .ZN(
        cor_maj_119_n28) );
  NAND2_X1 cor_maj_119_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_119_n28), .ZN(
        cor_maj_119_n29) );
  NAND2_X1 cor_maj_119_U17 ( .A1(cor_maj_119_n26), .A2(cor_maj_119_n27), .ZN(
        cor_maj_119_n30) );
  NAND2_X1 cor_maj_119_U16 ( .A1(cor_maj_119_n30), .A2(cor_maj_119_n29), .ZN(
        cor_maj_119_n31) );
  NAND2_X1 cor_maj_119_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_119_n25), .ZN(
        cor_maj_119_n18) );
  NAND2_X1 cor_maj_119_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_119_n19) );
  NAND2_X1 cor_maj_119_U13 ( .A1(cor_maj_119_n19), .A2(cor_maj_119_n18), .ZN(
        cor_maj_119_n22) );
  NAND2_X1 cor_maj_119_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_119_n24), .ZN(
        cor_maj_119_n20) );
  NAND2_X1 cor_maj_119_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_119_n21) );
  NAND2_X1 cor_maj_119_U10 ( .A1(cor_maj_119_n21), .A2(cor_maj_119_n20), .ZN(
        cor_maj_119_n23) );
  XOR2_X1 cor_maj_119_U9 ( .A(v_1_1_3[2]), .B(cor_maj_119_n24), .Z(
        cor_maj_119_n26) );
  XOR2_X1 cor_maj_119_U8 ( .A(v_1_1_3[5]), .B(cor_maj_119_n25), .Z(
        cor_maj_119_n27) );
  XOR2_X1 cor_maj_119_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_119_n24)
         );
  XOR2_X1 cor_maj_119_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_119_n25)
         );
  OR2_X1 cor_maj_119_U5 ( .A1(cor_maj_119_n23), .A2(cor_maj_119_n22), .ZN(
        cor_maj_119_n32) );
  NAND2_X1 cor_maj_119_U4 ( .A1(cor_maj_119_n22), .A2(cor_maj_119_n23), .ZN(
        cor_maj_119_n34) );
  NAND2_X1 cor_maj_119_U3 ( .A1(cor_maj_119_n32), .A2(cor_maj_119_n31), .ZN(
        cor_maj_119_n33) );
  NAND2_X1 cor_maj_119_U2 ( .A1(cor_maj_119_n34), .A2(cor_maj_119_n33), .ZN(
        cor_maj_119_port_o) );
  OR2_X1 cor_maj_120_U19 ( .A1(cor_maj_120_n27), .A2(cor_maj_120_n26), .ZN(
        cor_maj_120_n28) );
  NAND2_X1 cor_maj_120_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_120_n28), .ZN(
        cor_maj_120_n29) );
  NAND2_X1 cor_maj_120_U17 ( .A1(cor_maj_120_n26), .A2(cor_maj_120_n27), .ZN(
        cor_maj_120_n30) );
  NAND2_X1 cor_maj_120_U16 ( .A1(cor_maj_120_n30), .A2(cor_maj_120_n29), .ZN(
        cor_maj_120_n31) );
  NAND2_X1 cor_maj_120_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_120_n25), .ZN(
        cor_maj_120_n18) );
  NAND2_X1 cor_maj_120_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_120_n19) );
  NAND2_X1 cor_maj_120_U13 ( .A1(cor_maj_120_n19), .A2(cor_maj_120_n18), .ZN(
        cor_maj_120_n22) );
  NAND2_X1 cor_maj_120_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_120_n24), .ZN(
        cor_maj_120_n20) );
  NAND2_X1 cor_maj_120_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_120_n21) );
  NAND2_X1 cor_maj_120_U10 ( .A1(cor_maj_120_n21), .A2(cor_maj_120_n20), .ZN(
        cor_maj_120_n23) );
  XOR2_X1 cor_maj_120_U9 ( .A(v_1_1_3[2]), .B(cor_maj_120_n24), .Z(
        cor_maj_120_n26) );
  XOR2_X1 cor_maj_120_U8 ( .A(v_1_1_3[5]), .B(cor_maj_120_n25), .Z(
        cor_maj_120_n27) );
  XOR2_X1 cor_maj_120_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_120_n24)
         );
  XOR2_X1 cor_maj_120_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_120_n25)
         );
  OR2_X1 cor_maj_120_U5 ( .A1(cor_maj_120_n23), .A2(cor_maj_120_n22), .ZN(
        cor_maj_120_n32) );
  NAND2_X1 cor_maj_120_U4 ( .A1(cor_maj_120_n22), .A2(cor_maj_120_n23), .ZN(
        cor_maj_120_n34) );
  NAND2_X1 cor_maj_120_U3 ( .A1(cor_maj_120_n32), .A2(cor_maj_120_n31), .ZN(
        cor_maj_120_n33) );
  NAND2_X1 cor_maj_120_U2 ( .A1(cor_maj_120_n34), .A2(cor_maj_120_n33), .ZN(
        cor_maj_120_port_o) );
  OR2_X1 cor_maj_121_U19 ( .A1(cor_maj_121_n27), .A2(cor_maj_121_n26), .ZN(
        cor_maj_121_n28) );
  NAND2_X1 cor_maj_121_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_121_n28), .ZN(
        cor_maj_121_n29) );
  NAND2_X1 cor_maj_121_U17 ( .A1(cor_maj_121_n26), .A2(cor_maj_121_n27), .ZN(
        cor_maj_121_n30) );
  NAND2_X1 cor_maj_121_U16 ( .A1(cor_maj_121_n30), .A2(cor_maj_121_n29), .ZN(
        cor_maj_121_n31) );
  NAND2_X1 cor_maj_121_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_121_n25), .ZN(
        cor_maj_121_n18) );
  NAND2_X1 cor_maj_121_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_121_n19) );
  NAND2_X1 cor_maj_121_U13 ( .A1(cor_maj_121_n19), .A2(cor_maj_121_n18), .ZN(
        cor_maj_121_n22) );
  NAND2_X1 cor_maj_121_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_121_n24), .ZN(
        cor_maj_121_n20) );
  NAND2_X1 cor_maj_121_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_121_n21) );
  NAND2_X1 cor_maj_121_U10 ( .A1(cor_maj_121_n21), .A2(cor_maj_121_n20), .ZN(
        cor_maj_121_n23) );
  XOR2_X1 cor_maj_121_U9 ( .A(v_1_1_3[2]), .B(cor_maj_121_n24), .Z(
        cor_maj_121_n26) );
  XOR2_X1 cor_maj_121_U8 ( .A(v_1_1_3[5]), .B(cor_maj_121_n25), .Z(
        cor_maj_121_n27) );
  XOR2_X1 cor_maj_121_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_121_n24)
         );
  XOR2_X1 cor_maj_121_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_121_n25)
         );
  OR2_X1 cor_maj_121_U5 ( .A1(cor_maj_121_n23), .A2(cor_maj_121_n22), .ZN(
        cor_maj_121_n32) );
  NAND2_X1 cor_maj_121_U4 ( .A1(cor_maj_121_n22), .A2(cor_maj_121_n23), .ZN(
        cor_maj_121_n34) );
  NAND2_X1 cor_maj_121_U3 ( .A1(cor_maj_121_n32), .A2(cor_maj_121_n31), .ZN(
        cor_maj_121_n33) );
  NAND2_X1 cor_maj_121_U2 ( .A1(cor_maj_121_n34), .A2(cor_maj_121_n33), .ZN(
        cor_maj_121_port_o) );
  OR2_X1 cor_maj_122_U19 ( .A1(cor_maj_122_n27), .A2(cor_maj_122_n26), .ZN(
        cor_maj_122_n28) );
  NAND2_X1 cor_maj_122_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_122_n28), .ZN(
        cor_maj_122_n29) );
  NAND2_X1 cor_maj_122_U17 ( .A1(cor_maj_122_n26), .A2(cor_maj_122_n27), .ZN(
        cor_maj_122_n30) );
  NAND2_X1 cor_maj_122_U16 ( .A1(cor_maj_122_n30), .A2(cor_maj_122_n29), .ZN(
        cor_maj_122_n31) );
  NAND2_X1 cor_maj_122_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_122_n25), .ZN(
        cor_maj_122_n18) );
  NAND2_X1 cor_maj_122_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_122_n19) );
  NAND2_X1 cor_maj_122_U13 ( .A1(cor_maj_122_n19), .A2(cor_maj_122_n18), .ZN(
        cor_maj_122_n22) );
  NAND2_X1 cor_maj_122_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_122_n24), .ZN(
        cor_maj_122_n20) );
  NAND2_X1 cor_maj_122_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_122_n21) );
  NAND2_X1 cor_maj_122_U10 ( .A1(cor_maj_122_n21), .A2(cor_maj_122_n20), .ZN(
        cor_maj_122_n23) );
  XOR2_X1 cor_maj_122_U9 ( .A(v_1_1_3[2]), .B(cor_maj_122_n24), .Z(
        cor_maj_122_n26) );
  XOR2_X1 cor_maj_122_U8 ( .A(v_1_1_3[5]), .B(cor_maj_122_n25), .Z(
        cor_maj_122_n27) );
  XOR2_X1 cor_maj_122_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_122_n24)
         );
  XOR2_X1 cor_maj_122_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_122_n25)
         );
  OR2_X1 cor_maj_122_U5 ( .A1(cor_maj_122_n23), .A2(cor_maj_122_n22), .ZN(
        cor_maj_122_n32) );
  NAND2_X1 cor_maj_122_U4 ( .A1(cor_maj_122_n22), .A2(cor_maj_122_n23), .ZN(
        cor_maj_122_n34) );
  NAND2_X1 cor_maj_122_U3 ( .A1(cor_maj_122_n32), .A2(cor_maj_122_n31), .ZN(
        cor_maj_122_n33) );
  NAND2_X1 cor_maj_122_U2 ( .A1(cor_maj_122_n34), .A2(cor_maj_122_n33), .ZN(
        cor_maj_122_port_o) );
  OR2_X1 cor_maj_123_U19 ( .A1(cor_maj_123_n27), .A2(cor_maj_123_n26), .ZN(
        cor_maj_123_n28) );
  NAND2_X1 cor_maj_123_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_123_n28), .ZN(
        cor_maj_123_n29) );
  NAND2_X1 cor_maj_123_U17 ( .A1(cor_maj_123_n26), .A2(cor_maj_123_n27), .ZN(
        cor_maj_123_n30) );
  NAND2_X1 cor_maj_123_U16 ( .A1(cor_maj_123_n30), .A2(cor_maj_123_n29), .ZN(
        cor_maj_123_n31) );
  NAND2_X1 cor_maj_123_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_123_n25), .ZN(
        cor_maj_123_n18) );
  NAND2_X1 cor_maj_123_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_123_n19) );
  NAND2_X1 cor_maj_123_U13 ( .A1(cor_maj_123_n19), .A2(cor_maj_123_n18), .ZN(
        cor_maj_123_n22) );
  NAND2_X1 cor_maj_123_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_123_n24), .ZN(
        cor_maj_123_n20) );
  NAND2_X1 cor_maj_123_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_123_n21) );
  NAND2_X1 cor_maj_123_U10 ( .A1(cor_maj_123_n21), .A2(cor_maj_123_n20), .ZN(
        cor_maj_123_n23) );
  XOR2_X1 cor_maj_123_U9 ( .A(v_1_1_3[2]), .B(cor_maj_123_n24), .Z(
        cor_maj_123_n26) );
  XOR2_X1 cor_maj_123_U8 ( .A(v_1_1_3[5]), .B(cor_maj_123_n25), .Z(
        cor_maj_123_n27) );
  XOR2_X1 cor_maj_123_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_123_n24)
         );
  XOR2_X1 cor_maj_123_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_123_n25)
         );
  OR2_X1 cor_maj_123_U5 ( .A1(cor_maj_123_n23), .A2(cor_maj_123_n22), .ZN(
        cor_maj_123_n32) );
  NAND2_X1 cor_maj_123_U4 ( .A1(cor_maj_123_n22), .A2(cor_maj_123_n23), .ZN(
        cor_maj_123_n34) );
  NAND2_X1 cor_maj_123_U3 ( .A1(cor_maj_123_n32), .A2(cor_maj_123_n31), .ZN(
        cor_maj_123_n33) );
  NAND2_X1 cor_maj_123_U2 ( .A1(cor_maj_123_n34), .A2(cor_maj_123_n33), .ZN(
        cor_maj_123_port_o) );
  OR2_X1 cor_maj_124_U19 ( .A1(cor_maj_124_n27), .A2(cor_maj_124_n26), .ZN(
        cor_maj_124_n28) );
  NAND2_X1 cor_maj_124_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_124_n28), .ZN(
        cor_maj_124_n29) );
  NAND2_X1 cor_maj_124_U17 ( .A1(cor_maj_124_n26), .A2(cor_maj_124_n27), .ZN(
        cor_maj_124_n30) );
  NAND2_X1 cor_maj_124_U16 ( .A1(cor_maj_124_n30), .A2(cor_maj_124_n29), .ZN(
        cor_maj_124_n31) );
  NAND2_X1 cor_maj_124_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_124_n25), .ZN(
        cor_maj_124_n18) );
  NAND2_X1 cor_maj_124_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_124_n19) );
  NAND2_X1 cor_maj_124_U13 ( .A1(cor_maj_124_n19), .A2(cor_maj_124_n18), .ZN(
        cor_maj_124_n22) );
  NAND2_X1 cor_maj_124_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_124_n24), .ZN(
        cor_maj_124_n20) );
  NAND2_X1 cor_maj_124_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_124_n21) );
  NAND2_X1 cor_maj_124_U10 ( .A1(cor_maj_124_n21), .A2(cor_maj_124_n20), .ZN(
        cor_maj_124_n23) );
  XOR2_X1 cor_maj_124_U9 ( .A(v_1_1_3[2]), .B(cor_maj_124_n24), .Z(
        cor_maj_124_n26) );
  XOR2_X1 cor_maj_124_U8 ( .A(v_1_1_3[5]), .B(cor_maj_124_n25), .Z(
        cor_maj_124_n27) );
  XOR2_X1 cor_maj_124_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_124_n24)
         );
  XOR2_X1 cor_maj_124_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_124_n25)
         );
  OR2_X1 cor_maj_124_U5 ( .A1(cor_maj_124_n23), .A2(cor_maj_124_n22), .ZN(
        cor_maj_124_n32) );
  NAND2_X1 cor_maj_124_U4 ( .A1(cor_maj_124_n22), .A2(cor_maj_124_n23), .ZN(
        cor_maj_124_n34) );
  NAND2_X1 cor_maj_124_U3 ( .A1(cor_maj_124_n32), .A2(cor_maj_124_n31), .ZN(
        cor_maj_124_n33) );
  NAND2_X1 cor_maj_124_U2 ( .A1(cor_maj_124_n34), .A2(cor_maj_124_n33), .ZN(
        cor_maj_124_port_o) );
  OR2_X1 cor_maj_125_U19 ( .A1(cor_maj_125_n27), .A2(cor_maj_125_n26), .ZN(
        cor_maj_125_n28) );
  NAND2_X1 cor_maj_125_U18 ( .A1(v_1_1_3[6]), .A2(cor_maj_125_n28), .ZN(
        cor_maj_125_n29) );
  NAND2_X1 cor_maj_125_U17 ( .A1(cor_maj_125_n26), .A2(cor_maj_125_n27), .ZN(
        cor_maj_125_n30) );
  NAND2_X1 cor_maj_125_U16 ( .A1(cor_maj_125_n30), .A2(cor_maj_125_n29), .ZN(
        cor_maj_125_n31) );
  NAND2_X1 cor_maj_125_U15 ( .A1(v_1_1_3[5]), .A2(cor_maj_125_n25), .ZN(
        cor_maj_125_n18) );
  NAND2_X1 cor_maj_125_U14 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_125_n19) );
  NAND2_X1 cor_maj_125_U13 ( .A1(cor_maj_125_n19), .A2(cor_maj_125_n18), .ZN(
        cor_maj_125_n22) );
  NAND2_X1 cor_maj_125_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_125_n24), .ZN(
        cor_maj_125_n20) );
  NAND2_X1 cor_maj_125_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_125_n21) );
  NAND2_X1 cor_maj_125_U10 ( .A1(cor_maj_125_n21), .A2(cor_maj_125_n20), .ZN(
        cor_maj_125_n23) );
  XOR2_X1 cor_maj_125_U9 ( .A(v_1_1_3[2]), .B(cor_maj_125_n24), .Z(
        cor_maj_125_n26) );
  XOR2_X1 cor_maj_125_U8 ( .A(v_1_1_3[5]), .B(cor_maj_125_n25), .Z(
        cor_maj_125_n27) );
  XOR2_X1 cor_maj_125_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_125_n24)
         );
  XOR2_X1 cor_maj_125_U6 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_125_n25)
         );
  OR2_X1 cor_maj_125_U5 ( .A1(cor_maj_125_n23), .A2(cor_maj_125_n22), .ZN(
        cor_maj_125_n32) );
  NAND2_X1 cor_maj_125_U4 ( .A1(cor_maj_125_n22), .A2(cor_maj_125_n23), .ZN(
        cor_maj_125_n34) );
  NAND2_X1 cor_maj_125_U3 ( .A1(cor_maj_125_n32), .A2(cor_maj_125_n31), .ZN(
        cor_maj_125_n33) );
  NAND2_X1 cor_maj_125_U2 ( .A1(cor_maj_125_n34), .A2(cor_maj_125_n33), .ZN(
        cor_maj_125_port_o) );
  OR2_X1 cor_maj_126_U19 ( .A1(cor_maj_126_n27), .A2(cor_maj_126_n26), .ZN(
        cor_maj_126_n28) );
  NAND2_X1 cor_maj_126_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_126_n28), .ZN(
        cor_maj_126_n29) );
  NAND2_X1 cor_maj_126_U17 ( .A1(cor_maj_126_n26), .A2(cor_maj_126_n27), .ZN(
        cor_maj_126_n30) );
  NAND2_X1 cor_maj_126_U16 ( .A1(cor_maj_126_n30), .A2(cor_maj_126_n29), .ZN(
        cor_maj_126_n31) );
  NAND2_X1 cor_maj_126_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_126_n25), .ZN(
        cor_maj_126_n18) );
  NAND2_X1 cor_maj_126_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_126_n19) );
  NAND2_X1 cor_maj_126_U13 ( .A1(cor_maj_126_n19), .A2(cor_maj_126_n18), .ZN(
        cor_maj_126_n22) );
  NAND2_X1 cor_maj_126_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_126_n24), .ZN(
        cor_maj_126_n20) );
  NAND2_X1 cor_maj_126_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_126_n21) );
  NAND2_X1 cor_maj_126_U10 ( .A1(cor_maj_126_n21), .A2(cor_maj_126_n20), .ZN(
        cor_maj_126_n23) );
  XOR2_X1 cor_maj_126_U9 ( .A(v_1_2_0[2]), .B(cor_maj_126_n24), .Z(
        cor_maj_126_n26) );
  XOR2_X1 cor_maj_126_U8 ( .A(v_1_2_0[5]), .B(cor_maj_126_n25), .Z(
        cor_maj_126_n27) );
  XOR2_X1 cor_maj_126_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_126_n24)
         );
  XOR2_X1 cor_maj_126_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_126_n25)
         );
  OR2_X1 cor_maj_126_U5 ( .A1(cor_maj_126_n23), .A2(cor_maj_126_n22), .ZN(
        cor_maj_126_n32) );
  NAND2_X1 cor_maj_126_U4 ( .A1(cor_maj_126_n22), .A2(cor_maj_126_n23), .ZN(
        cor_maj_126_n34) );
  NAND2_X1 cor_maj_126_U3 ( .A1(cor_maj_126_n32), .A2(cor_maj_126_n31), .ZN(
        cor_maj_126_n33) );
  NAND2_X1 cor_maj_126_U2 ( .A1(cor_maj_126_n34), .A2(cor_maj_126_n33), .ZN(
        cor_maj_126_port_o) );
  OR2_X1 cor_maj_127_U19 ( .A1(cor_maj_127_n27), .A2(cor_maj_127_n26), .ZN(
        cor_maj_127_n28) );
  NAND2_X1 cor_maj_127_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_127_n28), .ZN(
        cor_maj_127_n29) );
  NAND2_X1 cor_maj_127_U17 ( .A1(cor_maj_127_n26), .A2(cor_maj_127_n27), .ZN(
        cor_maj_127_n30) );
  NAND2_X1 cor_maj_127_U16 ( .A1(cor_maj_127_n30), .A2(cor_maj_127_n29), .ZN(
        cor_maj_127_n31) );
  NAND2_X1 cor_maj_127_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_127_n25), .ZN(
        cor_maj_127_n18) );
  NAND2_X1 cor_maj_127_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_127_n19) );
  NAND2_X1 cor_maj_127_U13 ( .A1(cor_maj_127_n19), .A2(cor_maj_127_n18), .ZN(
        cor_maj_127_n22) );
  NAND2_X1 cor_maj_127_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_127_n24), .ZN(
        cor_maj_127_n20) );
  NAND2_X1 cor_maj_127_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_127_n21) );
  NAND2_X1 cor_maj_127_U10 ( .A1(cor_maj_127_n21), .A2(cor_maj_127_n20), .ZN(
        cor_maj_127_n23) );
  XOR2_X1 cor_maj_127_U9 ( .A(v_1_2_0[2]), .B(cor_maj_127_n24), .Z(
        cor_maj_127_n26) );
  XOR2_X1 cor_maj_127_U8 ( .A(v_1_2_0[5]), .B(cor_maj_127_n25), .Z(
        cor_maj_127_n27) );
  XOR2_X1 cor_maj_127_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_127_n24)
         );
  XOR2_X1 cor_maj_127_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_127_n25)
         );
  OR2_X1 cor_maj_127_U5 ( .A1(cor_maj_127_n23), .A2(cor_maj_127_n22), .ZN(
        cor_maj_127_n32) );
  NAND2_X1 cor_maj_127_U4 ( .A1(cor_maj_127_n22), .A2(cor_maj_127_n23), .ZN(
        cor_maj_127_n34) );
  NAND2_X1 cor_maj_127_U3 ( .A1(cor_maj_127_n32), .A2(cor_maj_127_n31), .ZN(
        cor_maj_127_n33) );
  NAND2_X1 cor_maj_127_U2 ( .A1(cor_maj_127_n34), .A2(cor_maj_127_n33), .ZN(
        cor_maj_127_port_o) );
  OR2_X1 cor_maj_128_U19 ( .A1(cor_maj_128_n27), .A2(cor_maj_128_n26), .ZN(
        cor_maj_128_n28) );
  NAND2_X1 cor_maj_128_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_128_n28), .ZN(
        cor_maj_128_n29) );
  NAND2_X1 cor_maj_128_U17 ( .A1(cor_maj_128_n26), .A2(cor_maj_128_n27), .ZN(
        cor_maj_128_n30) );
  NAND2_X1 cor_maj_128_U16 ( .A1(cor_maj_128_n30), .A2(cor_maj_128_n29), .ZN(
        cor_maj_128_n31) );
  NAND2_X1 cor_maj_128_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_128_n25), .ZN(
        cor_maj_128_n18) );
  NAND2_X1 cor_maj_128_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_128_n19) );
  NAND2_X1 cor_maj_128_U13 ( .A1(cor_maj_128_n19), .A2(cor_maj_128_n18), .ZN(
        cor_maj_128_n22) );
  NAND2_X1 cor_maj_128_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_128_n24), .ZN(
        cor_maj_128_n20) );
  NAND2_X1 cor_maj_128_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_128_n21) );
  NAND2_X1 cor_maj_128_U10 ( .A1(cor_maj_128_n21), .A2(cor_maj_128_n20), .ZN(
        cor_maj_128_n23) );
  XOR2_X1 cor_maj_128_U9 ( .A(v_1_2_0[2]), .B(cor_maj_128_n24), .Z(
        cor_maj_128_n26) );
  XOR2_X1 cor_maj_128_U8 ( .A(v_1_2_0[5]), .B(cor_maj_128_n25), .Z(
        cor_maj_128_n27) );
  XOR2_X1 cor_maj_128_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_128_n24)
         );
  XOR2_X1 cor_maj_128_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_128_n25)
         );
  OR2_X1 cor_maj_128_U5 ( .A1(cor_maj_128_n23), .A2(cor_maj_128_n22), .ZN(
        cor_maj_128_n32) );
  NAND2_X1 cor_maj_128_U4 ( .A1(cor_maj_128_n22), .A2(cor_maj_128_n23), .ZN(
        cor_maj_128_n34) );
  NAND2_X1 cor_maj_128_U3 ( .A1(cor_maj_128_n32), .A2(cor_maj_128_n31), .ZN(
        cor_maj_128_n33) );
  NAND2_X1 cor_maj_128_U2 ( .A1(cor_maj_128_n34), .A2(cor_maj_128_n33), .ZN(
        cor_maj_128_port_o) );
  OR2_X1 cor_maj_129_U19 ( .A1(cor_maj_129_n27), .A2(cor_maj_129_n26), .ZN(
        cor_maj_129_n28) );
  NAND2_X1 cor_maj_129_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_129_n28), .ZN(
        cor_maj_129_n29) );
  NAND2_X1 cor_maj_129_U17 ( .A1(cor_maj_129_n26), .A2(cor_maj_129_n27), .ZN(
        cor_maj_129_n30) );
  NAND2_X1 cor_maj_129_U16 ( .A1(cor_maj_129_n30), .A2(cor_maj_129_n29), .ZN(
        cor_maj_129_n31) );
  NAND2_X1 cor_maj_129_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_129_n25), .ZN(
        cor_maj_129_n18) );
  NAND2_X1 cor_maj_129_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_129_n19) );
  NAND2_X1 cor_maj_129_U13 ( .A1(cor_maj_129_n19), .A2(cor_maj_129_n18), .ZN(
        cor_maj_129_n22) );
  NAND2_X1 cor_maj_129_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_129_n24), .ZN(
        cor_maj_129_n20) );
  NAND2_X1 cor_maj_129_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_129_n21) );
  NAND2_X1 cor_maj_129_U10 ( .A1(cor_maj_129_n21), .A2(cor_maj_129_n20), .ZN(
        cor_maj_129_n23) );
  XOR2_X1 cor_maj_129_U9 ( .A(v_1_2_0[2]), .B(cor_maj_129_n24), .Z(
        cor_maj_129_n26) );
  XOR2_X1 cor_maj_129_U8 ( .A(v_1_2_0[5]), .B(cor_maj_129_n25), .Z(
        cor_maj_129_n27) );
  XOR2_X1 cor_maj_129_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_129_n24)
         );
  XOR2_X1 cor_maj_129_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_129_n25)
         );
  OR2_X1 cor_maj_129_U5 ( .A1(cor_maj_129_n23), .A2(cor_maj_129_n22), .ZN(
        cor_maj_129_n32) );
  NAND2_X1 cor_maj_129_U4 ( .A1(cor_maj_129_n22), .A2(cor_maj_129_n23), .ZN(
        cor_maj_129_n34) );
  NAND2_X1 cor_maj_129_U3 ( .A1(cor_maj_129_n32), .A2(cor_maj_129_n31), .ZN(
        cor_maj_129_n33) );
  NAND2_X1 cor_maj_129_U2 ( .A1(cor_maj_129_n34), .A2(cor_maj_129_n33), .ZN(
        cor_maj_129_port_o) );
  OR2_X1 cor_maj_130_U19 ( .A1(cor_maj_130_n27), .A2(cor_maj_130_n26), .ZN(
        cor_maj_130_n28) );
  NAND2_X1 cor_maj_130_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_130_n28), .ZN(
        cor_maj_130_n29) );
  NAND2_X1 cor_maj_130_U17 ( .A1(cor_maj_130_n26), .A2(cor_maj_130_n27), .ZN(
        cor_maj_130_n30) );
  NAND2_X1 cor_maj_130_U16 ( .A1(cor_maj_130_n30), .A2(cor_maj_130_n29), .ZN(
        cor_maj_130_n31) );
  NAND2_X1 cor_maj_130_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_130_n25), .ZN(
        cor_maj_130_n18) );
  NAND2_X1 cor_maj_130_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_130_n19) );
  NAND2_X1 cor_maj_130_U13 ( .A1(cor_maj_130_n19), .A2(cor_maj_130_n18), .ZN(
        cor_maj_130_n22) );
  NAND2_X1 cor_maj_130_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_130_n24), .ZN(
        cor_maj_130_n20) );
  NAND2_X1 cor_maj_130_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_130_n21) );
  NAND2_X1 cor_maj_130_U10 ( .A1(cor_maj_130_n21), .A2(cor_maj_130_n20), .ZN(
        cor_maj_130_n23) );
  XOR2_X1 cor_maj_130_U9 ( .A(v_1_2_0[2]), .B(cor_maj_130_n24), .Z(
        cor_maj_130_n26) );
  XOR2_X1 cor_maj_130_U8 ( .A(v_1_2_0[5]), .B(cor_maj_130_n25), .Z(
        cor_maj_130_n27) );
  XOR2_X1 cor_maj_130_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_130_n24)
         );
  XOR2_X1 cor_maj_130_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_130_n25)
         );
  OR2_X1 cor_maj_130_U5 ( .A1(cor_maj_130_n23), .A2(cor_maj_130_n22), .ZN(
        cor_maj_130_n32) );
  NAND2_X1 cor_maj_130_U4 ( .A1(cor_maj_130_n22), .A2(cor_maj_130_n23), .ZN(
        cor_maj_130_n34) );
  NAND2_X1 cor_maj_130_U3 ( .A1(cor_maj_130_n32), .A2(cor_maj_130_n31), .ZN(
        cor_maj_130_n33) );
  NAND2_X1 cor_maj_130_U2 ( .A1(cor_maj_130_n34), .A2(cor_maj_130_n33), .ZN(
        cor_maj_130_port_o) );
  OR2_X1 cor_maj_131_U19 ( .A1(cor_maj_131_n27), .A2(cor_maj_131_n26), .ZN(
        cor_maj_131_n28) );
  NAND2_X1 cor_maj_131_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_131_n28), .ZN(
        cor_maj_131_n29) );
  NAND2_X1 cor_maj_131_U17 ( .A1(cor_maj_131_n26), .A2(cor_maj_131_n27), .ZN(
        cor_maj_131_n30) );
  NAND2_X1 cor_maj_131_U16 ( .A1(cor_maj_131_n30), .A2(cor_maj_131_n29), .ZN(
        cor_maj_131_n31) );
  NAND2_X1 cor_maj_131_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_131_n25), .ZN(
        cor_maj_131_n18) );
  NAND2_X1 cor_maj_131_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_131_n19) );
  NAND2_X1 cor_maj_131_U13 ( .A1(cor_maj_131_n19), .A2(cor_maj_131_n18), .ZN(
        cor_maj_131_n22) );
  NAND2_X1 cor_maj_131_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_131_n24), .ZN(
        cor_maj_131_n20) );
  NAND2_X1 cor_maj_131_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_131_n21) );
  NAND2_X1 cor_maj_131_U10 ( .A1(cor_maj_131_n21), .A2(cor_maj_131_n20), .ZN(
        cor_maj_131_n23) );
  XOR2_X1 cor_maj_131_U9 ( .A(v_1_2_0[2]), .B(cor_maj_131_n24), .Z(
        cor_maj_131_n26) );
  XOR2_X1 cor_maj_131_U8 ( .A(v_1_2_0[5]), .B(cor_maj_131_n25), .Z(
        cor_maj_131_n27) );
  XOR2_X1 cor_maj_131_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_131_n24)
         );
  XOR2_X1 cor_maj_131_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_131_n25)
         );
  OR2_X1 cor_maj_131_U5 ( .A1(cor_maj_131_n23), .A2(cor_maj_131_n22), .ZN(
        cor_maj_131_n32) );
  NAND2_X1 cor_maj_131_U4 ( .A1(cor_maj_131_n22), .A2(cor_maj_131_n23), .ZN(
        cor_maj_131_n34) );
  NAND2_X1 cor_maj_131_U3 ( .A1(cor_maj_131_n32), .A2(cor_maj_131_n31), .ZN(
        cor_maj_131_n33) );
  NAND2_X1 cor_maj_131_U2 ( .A1(cor_maj_131_n34), .A2(cor_maj_131_n33), .ZN(
        cor_maj_131_port_o) );
  OR2_X1 cor_maj_132_U19 ( .A1(cor_maj_132_n27), .A2(cor_maj_132_n26), .ZN(
        cor_maj_132_n28) );
  NAND2_X1 cor_maj_132_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_132_n28), .ZN(
        cor_maj_132_n29) );
  NAND2_X1 cor_maj_132_U17 ( .A1(cor_maj_132_n26), .A2(cor_maj_132_n27), .ZN(
        cor_maj_132_n30) );
  NAND2_X1 cor_maj_132_U16 ( .A1(cor_maj_132_n30), .A2(cor_maj_132_n29), .ZN(
        cor_maj_132_n31) );
  NAND2_X1 cor_maj_132_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_132_n25), .ZN(
        cor_maj_132_n18) );
  NAND2_X1 cor_maj_132_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_132_n19) );
  NAND2_X1 cor_maj_132_U13 ( .A1(cor_maj_132_n19), .A2(cor_maj_132_n18), .ZN(
        cor_maj_132_n22) );
  NAND2_X1 cor_maj_132_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_132_n24), .ZN(
        cor_maj_132_n20) );
  NAND2_X1 cor_maj_132_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_132_n21) );
  NAND2_X1 cor_maj_132_U10 ( .A1(cor_maj_132_n21), .A2(cor_maj_132_n20), .ZN(
        cor_maj_132_n23) );
  XOR2_X1 cor_maj_132_U9 ( .A(v_1_2_0[2]), .B(cor_maj_132_n24), .Z(
        cor_maj_132_n26) );
  XOR2_X1 cor_maj_132_U8 ( .A(v_1_2_0[5]), .B(cor_maj_132_n25), .Z(
        cor_maj_132_n27) );
  XOR2_X1 cor_maj_132_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_132_n24)
         );
  XOR2_X1 cor_maj_132_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_132_n25)
         );
  OR2_X1 cor_maj_132_U5 ( .A1(cor_maj_132_n23), .A2(cor_maj_132_n22), .ZN(
        cor_maj_132_n32) );
  NAND2_X1 cor_maj_132_U4 ( .A1(cor_maj_132_n22), .A2(cor_maj_132_n23), .ZN(
        cor_maj_132_n34) );
  NAND2_X1 cor_maj_132_U3 ( .A1(cor_maj_132_n32), .A2(cor_maj_132_n31), .ZN(
        cor_maj_132_n33) );
  NAND2_X1 cor_maj_132_U2 ( .A1(cor_maj_132_n34), .A2(cor_maj_132_n33), .ZN(
        cor_maj_132_port_o) );
  OR2_X1 cor_maj_133_U19 ( .A1(cor_maj_133_n27), .A2(cor_maj_133_n26), .ZN(
        cor_maj_133_n28) );
  NAND2_X1 cor_maj_133_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_133_n28), .ZN(
        cor_maj_133_n29) );
  NAND2_X1 cor_maj_133_U17 ( .A1(cor_maj_133_n26), .A2(cor_maj_133_n27), .ZN(
        cor_maj_133_n30) );
  NAND2_X1 cor_maj_133_U16 ( .A1(cor_maj_133_n30), .A2(cor_maj_133_n29), .ZN(
        cor_maj_133_n31) );
  NAND2_X1 cor_maj_133_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_133_n25), .ZN(
        cor_maj_133_n18) );
  NAND2_X1 cor_maj_133_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_133_n19) );
  NAND2_X1 cor_maj_133_U13 ( .A1(cor_maj_133_n19), .A2(cor_maj_133_n18), .ZN(
        cor_maj_133_n22) );
  NAND2_X1 cor_maj_133_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_133_n24), .ZN(
        cor_maj_133_n20) );
  NAND2_X1 cor_maj_133_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_133_n21) );
  NAND2_X1 cor_maj_133_U10 ( .A1(cor_maj_133_n21), .A2(cor_maj_133_n20), .ZN(
        cor_maj_133_n23) );
  XOR2_X1 cor_maj_133_U9 ( .A(v_1_2_1[2]), .B(cor_maj_133_n24), .Z(
        cor_maj_133_n26) );
  XOR2_X1 cor_maj_133_U8 ( .A(v_1_2_1[5]), .B(cor_maj_133_n25), .Z(
        cor_maj_133_n27) );
  XOR2_X1 cor_maj_133_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_133_n24)
         );
  XOR2_X1 cor_maj_133_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_133_n25)
         );
  OR2_X1 cor_maj_133_U5 ( .A1(cor_maj_133_n23), .A2(cor_maj_133_n22), .ZN(
        cor_maj_133_n32) );
  NAND2_X1 cor_maj_133_U4 ( .A1(cor_maj_133_n22), .A2(cor_maj_133_n23), .ZN(
        cor_maj_133_n34) );
  NAND2_X1 cor_maj_133_U3 ( .A1(cor_maj_133_n32), .A2(cor_maj_133_n31), .ZN(
        cor_maj_133_n33) );
  NAND2_X1 cor_maj_133_U2 ( .A1(cor_maj_133_n34), .A2(cor_maj_133_n33), .ZN(
        cor_maj_133_port_o) );
  OR2_X1 cor_maj_134_U19 ( .A1(cor_maj_134_n27), .A2(cor_maj_134_n26), .ZN(
        cor_maj_134_n28) );
  NAND2_X1 cor_maj_134_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_134_n28), .ZN(
        cor_maj_134_n29) );
  NAND2_X1 cor_maj_134_U17 ( .A1(cor_maj_134_n26), .A2(cor_maj_134_n27), .ZN(
        cor_maj_134_n30) );
  NAND2_X1 cor_maj_134_U16 ( .A1(cor_maj_134_n30), .A2(cor_maj_134_n29), .ZN(
        cor_maj_134_n31) );
  NAND2_X1 cor_maj_134_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_134_n25), .ZN(
        cor_maj_134_n18) );
  NAND2_X1 cor_maj_134_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_134_n19) );
  NAND2_X1 cor_maj_134_U13 ( .A1(cor_maj_134_n19), .A2(cor_maj_134_n18), .ZN(
        cor_maj_134_n22) );
  NAND2_X1 cor_maj_134_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_134_n24), .ZN(
        cor_maj_134_n20) );
  NAND2_X1 cor_maj_134_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_134_n21) );
  NAND2_X1 cor_maj_134_U10 ( .A1(cor_maj_134_n21), .A2(cor_maj_134_n20), .ZN(
        cor_maj_134_n23) );
  XOR2_X1 cor_maj_134_U9 ( .A(v_1_2_1[2]), .B(cor_maj_134_n24), .Z(
        cor_maj_134_n26) );
  XOR2_X1 cor_maj_134_U8 ( .A(v_1_2_1[5]), .B(cor_maj_134_n25), .Z(
        cor_maj_134_n27) );
  XOR2_X1 cor_maj_134_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_134_n24)
         );
  XOR2_X1 cor_maj_134_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_134_n25)
         );
  OR2_X1 cor_maj_134_U5 ( .A1(cor_maj_134_n23), .A2(cor_maj_134_n22), .ZN(
        cor_maj_134_n32) );
  NAND2_X1 cor_maj_134_U4 ( .A1(cor_maj_134_n22), .A2(cor_maj_134_n23), .ZN(
        cor_maj_134_n34) );
  NAND2_X1 cor_maj_134_U3 ( .A1(cor_maj_134_n32), .A2(cor_maj_134_n31), .ZN(
        cor_maj_134_n33) );
  NAND2_X1 cor_maj_134_U2 ( .A1(cor_maj_134_n34), .A2(cor_maj_134_n33), .ZN(
        cor_maj_134_port_o) );
  OR2_X1 cor_maj_135_U19 ( .A1(cor_maj_135_n27), .A2(cor_maj_135_n26), .ZN(
        cor_maj_135_n28) );
  NAND2_X1 cor_maj_135_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_135_n28), .ZN(
        cor_maj_135_n29) );
  NAND2_X1 cor_maj_135_U17 ( .A1(cor_maj_135_n26), .A2(cor_maj_135_n27), .ZN(
        cor_maj_135_n30) );
  NAND2_X1 cor_maj_135_U16 ( .A1(cor_maj_135_n30), .A2(cor_maj_135_n29), .ZN(
        cor_maj_135_n31) );
  NAND2_X1 cor_maj_135_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_135_n25), .ZN(
        cor_maj_135_n18) );
  NAND2_X1 cor_maj_135_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_135_n19) );
  NAND2_X1 cor_maj_135_U13 ( .A1(cor_maj_135_n19), .A2(cor_maj_135_n18), .ZN(
        cor_maj_135_n22) );
  NAND2_X1 cor_maj_135_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_135_n24), .ZN(
        cor_maj_135_n20) );
  NAND2_X1 cor_maj_135_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_135_n21) );
  NAND2_X1 cor_maj_135_U10 ( .A1(cor_maj_135_n21), .A2(cor_maj_135_n20), .ZN(
        cor_maj_135_n23) );
  XOR2_X1 cor_maj_135_U9 ( .A(v_1_2_1[2]), .B(cor_maj_135_n24), .Z(
        cor_maj_135_n26) );
  XOR2_X1 cor_maj_135_U8 ( .A(v_1_2_1[5]), .B(cor_maj_135_n25), .Z(
        cor_maj_135_n27) );
  XOR2_X1 cor_maj_135_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_135_n24)
         );
  XOR2_X1 cor_maj_135_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_135_n25)
         );
  OR2_X1 cor_maj_135_U5 ( .A1(cor_maj_135_n23), .A2(cor_maj_135_n22), .ZN(
        cor_maj_135_n32) );
  NAND2_X1 cor_maj_135_U4 ( .A1(cor_maj_135_n22), .A2(cor_maj_135_n23), .ZN(
        cor_maj_135_n34) );
  NAND2_X1 cor_maj_135_U3 ( .A1(cor_maj_135_n32), .A2(cor_maj_135_n31), .ZN(
        cor_maj_135_n33) );
  NAND2_X1 cor_maj_135_U2 ( .A1(cor_maj_135_n34), .A2(cor_maj_135_n33), .ZN(
        cor_maj_135_port_o) );
  OR2_X1 cor_maj_136_U19 ( .A1(cor_maj_136_n27), .A2(cor_maj_136_n26), .ZN(
        cor_maj_136_n28) );
  NAND2_X1 cor_maj_136_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_136_n28), .ZN(
        cor_maj_136_n29) );
  NAND2_X1 cor_maj_136_U17 ( .A1(cor_maj_136_n26), .A2(cor_maj_136_n27), .ZN(
        cor_maj_136_n30) );
  NAND2_X1 cor_maj_136_U16 ( .A1(cor_maj_136_n30), .A2(cor_maj_136_n29), .ZN(
        cor_maj_136_n31) );
  NAND2_X1 cor_maj_136_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_136_n25), .ZN(
        cor_maj_136_n18) );
  NAND2_X1 cor_maj_136_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_136_n19) );
  NAND2_X1 cor_maj_136_U13 ( .A1(cor_maj_136_n19), .A2(cor_maj_136_n18), .ZN(
        cor_maj_136_n22) );
  NAND2_X1 cor_maj_136_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_136_n24), .ZN(
        cor_maj_136_n20) );
  NAND2_X1 cor_maj_136_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_136_n21) );
  NAND2_X1 cor_maj_136_U10 ( .A1(cor_maj_136_n21), .A2(cor_maj_136_n20), .ZN(
        cor_maj_136_n23) );
  XOR2_X1 cor_maj_136_U9 ( .A(v_1_2_1[2]), .B(cor_maj_136_n24), .Z(
        cor_maj_136_n26) );
  XOR2_X1 cor_maj_136_U8 ( .A(v_1_2_1[5]), .B(cor_maj_136_n25), .Z(
        cor_maj_136_n27) );
  XOR2_X1 cor_maj_136_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_136_n24)
         );
  XOR2_X1 cor_maj_136_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_136_n25)
         );
  OR2_X1 cor_maj_136_U5 ( .A1(cor_maj_136_n23), .A2(cor_maj_136_n22), .ZN(
        cor_maj_136_n32) );
  NAND2_X1 cor_maj_136_U4 ( .A1(cor_maj_136_n22), .A2(cor_maj_136_n23), .ZN(
        cor_maj_136_n34) );
  NAND2_X1 cor_maj_136_U3 ( .A1(cor_maj_136_n32), .A2(cor_maj_136_n31), .ZN(
        cor_maj_136_n33) );
  NAND2_X1 cor_maj_136_U2 ( .A1(cor_maj_136_n34), .A2(cor_maj_136_n33), .ZN(
        cor_maj_136_port_o) );
  OR2_X1 cor_maj_137_U19 ( .A1(cor_maj_137_n27), .A2(cor_maj_137_n26), .ZN(
        cor_maj_137_n28) );
  NAND2_X1 cor_maj_137_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_137_n28), .ZN(
        cor_maj_137_n29) );
  NAND2_X1 cor_maj_137_U17 ( .A1(cor_maj_137_n26), .A2(cor_maj_137_n27), .ZN(
        cor_maj_137_n30) );
  NAND2_X1 cor_maj_137_U16 ( .A1(cor_maj_137_n30), .A2(cor_maj_137_n29), .ZN(
        cor_maj_137_n31) );
  NAND2_X1 cor_maj_137_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_137_n25), .ZN(
        cor_maj_137_n18) );
  NAND2_X1 cor_maj_137_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_137_n19) );
  NAND2_X1 cor_maj_137_U13 ( .A1(cor_maj_137_n19), .A2(cor_maj_137_n18), .ZN(
        cor_maj_137_n22) );
  NAND2_X1 cor_maj_137_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_137_n24), .ZN(
        cor_maj_137_n20) );
  NAND2_X1 cor_maj_137_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_137_n21) );
  NAND2_X1 cor_maj_137_U10 ( .A1(cor_maj_137_n21), .A2(cor_maj_137_n20), .ZN(
        cor_maj_137_n23) );
  XOR2_X1 cor_maj_137_U9 ( .A(v_1_2_1[2]), .B(cor_maj_137_n24), .Z(
        cor_maj_137_n26) );
  XOR2_X1 cor_maj_137_U8 ( .A(v_1_2_1[5]), .B(cor_maj_137_n25), .Z(
        cor_maj_137_n27) );
  XOR2_X1 cor_maj_137_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_137_n24)
         );
  XOR2_X1 cor_maj_137_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_137_n25)
         );
  OR2_X1 cor_maj_137_U5 ( .A1(cor_maj_137_n23), .A2(cor_maj_137_n22), .ZN(
        cor_maj_137_n32) );
  NAND2_X1 cor_maj_137_U4 ( .A1(cor_maj_137_n22), .A2(cor_maj_137_n23), .ZN(
        cor_maj_137_n34) );
  NAND2_X1 cor_maj_137_U3 ( .A1(cor_maj_137_n32), .A2(cor_maj_137_n31), .ZN(
        cor_maj_137_n33) );
  NAND2_X1 cor_maj_137_U2 ( .A1(cor_maj_137_n34), .A2(cor_maj_137_n33), .ZN(
        cor_maj_137_port_o) );
  OR2_X1 cor_maj_138_U19 ( .A1(cor_maj_138_n27), .A2(cor_maj_138_n26), .ZN(
        cor_maj_138_n28) );
  NAND2_X1 cor_maj_138_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_138_n28), .ZN(
        cor_maj_138_n29) );
  NAND2_X1 cor_maj_138_U17 ( .A1(cor_maj_138_n26), .A2(cor_maj_138_n27), .ZN(
        cor_maj_138_n30) );
  NAND2_X1 cor_maj_138_U16 ( .A1(cor_maj_138_n30), .A2(cor_maj_138_n29), .ZN(
        cor_maj_138_n31) );
  NAND2_X1 cor_maj_138_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_138_n25), .ZN(
        cor_maj_138_n18) );
  NAND2_X1 cor_maj_138_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_138_n19) );
  NAND2_X1 cor_maj_138_U13 ( .A1(cor_maj_138_n19), .A2(cor_maj_138_n18), .ZN(
        cor_maj_138_n22) );
  NAND2_X1 cor_maj_138_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_138_n24), .ZN(
        cor_maj_138_n20) );
  NAND2_X1 cor_maj_138_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_138_n21) );
  NAND2_X1 cor_maj_138_U10 ( .A1(cor_maj_138_n21), .A2(cor_maj_138_n20), .ZN(
        cor_maj_138_n23) );
  XOR2_X1 cor_maj_138_U9 ( .A(v_1_2_1[2]), .B(cor_maj_138_n24), .Z(
        cor_maj_138_n26) );
  XOR2_X1 cor_maj_138_U8 ( .A(v_1_2_1[5]), .B(cor_maj_138_n25), .Z(
        cor_maj_138_n27) );
  XOR2_X1 cor_maj_138_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_138_n24)
         );
  XOR2_X1 cor_maj_138_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_138_n25)
         );
  OR2_X1 cor_maj_138_U5 ( .A1(cor_maj_138_n23), .A2(cor_maj_138_n22), .ZN(
        cor_maj_138_n32) );
  NAND2_X1 cor_maj_138_U4 ( .A1(cor_maj_138_n22), .A2(cor_maj_138_n23), .ZN(
        cor_maj_138_n34) );
  NAND2_X1 cor_maj_138_U3 ( .A1(cor_maj_138_n32), .A2(cor_maj_138_n31), .ZN(
        cor_maj_138_n33) );
  NAND2_X1 cor_maj_138_U2 ( .A1(cor_maj_138_n34), .A2(cor_maj_138_n33), .ZN(
        cor_maj_138_port_o) );
  OR2_X1 cor_maj_139_U19 ( .A1(cor_maj_139_n27), .A2(cor_maj_139_n26), .ZN(
        cor_maj_139_n28) );
  NAND2_X1 cor_maj_139_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_139_n28), .ZN(
        cor_maj_139_n29) );
  NAND2_X1 cor_maj_139_U17 ( .A1(cor_maj_139_n26), .A2(cor_maj_139_n27), .ZN(
        cor_maj_139_n30) );
  NAND2_X1 cor_maj_139_U16 ( .A1(cor_maj_139_n30), .A2(cor_maj_139_n29), .ZN(
        cor_maj_139_n31) );
  NAND2_X1 cor_maj_139_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_139_n25), .ZN(
        cor_maj_139_n18) );
  NAND2_X1 cor_maj_139_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_139_n19) );
  NAND2_X1 cor_maj_139_U13 ( .A1(cor_maj_139_n19), .A2(cor_maj_139_n18), .ZN(
        cor_maj_139_n22) );
  NAND2_X1 cor_maj_139_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_139_n24), .ZN(
        cor_maj_139_n20) );
  NAND2_X1 cor_maj_139_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_139_n21) );
  NAND2_X1 cor_maj_139_U10 ( .A1(cor_maj_139_n21), .A2(cor_maj_139_n20), .ZN(
        cor_maj_139_n23) );
  XOR2_X1 cor_maj_139_U9 ( .A(v_1_2_1[2]), .B(cor_maj_139_n24), .Z(
        cor_maj_139_n26) );
  XOR2_X1 cor_maj_139_U8 ( .A(v_1_2_1[5]), .B(cor_maj_139_n25), .Z(
        cor_maj_139_n27) );
  XOR2_X1 cor_maj_139_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_139_n24)
         );
  XOR2_X1 cor_maj_139_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_139_n25)
         );
  OR2_X1 cor_maj_139_U5 ( .A1(cor_maj_139_n23), .A2(cor_maj_139_n22), .ZN(
        cor_maj_139_n32) );
  NAND2_X1 cor_maj_139_U4 ( .A1(cor_maj_139_n22), .A2(cor_maj_139_n23), .ZN(
        cor_maj_139_n34) );
  NAND2_X1 cor_maj_139_U3 ( .A1(cor_maj_139_n32), .A2(cor_maj_139_n31), .ZN(
        cor_maj_139_n33) );
  NAND2_X1 cor_maj_139_U2 ( .A1(cor_maj_139_n34), .A2(cor_maj_139_n33), .ZN(
        cor_maj_139_port_o) );
  OR2_X1 cor_maj_140_U19 ( .A1(cor_maj_140_n27), .A2(cor_maj_140_n26), .ZN(
        cor_maj_140_n28) );
  NAND2_X1 cor_maj_140_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_140_n28), .ZN(
        cor_maj_140_n29) );
  NAND2_X1 cor_maj_140_U17 ( .A1(cor_maj_140_n26), .A2(cor_maj_140_n27), .ZN(
        cor_maj_140_n30) );
  NAND2_X1 cor_maj_140_U16 ( .A1(cor_maj_140_n30), .A2(cor_maj_140_n29), .ZN(
        cor_maj_140_n31) );
  NAND2_X1 cor_maj_140_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_140_n25), .ZN(
        cor_maj_140_n18) );
  NAND2_X1 cor_maj_140_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_140_n19) );
  NAND2_X1 cor_maj_140_U13 ( .A1(cor_maj_140_n19), .A2(cor_maj_140_n18), .ZN(
        cor_maj_140_n22) );
  NAND2_X1 cor_maj_140_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_140_n24), .ZN(
        cor_maj_140_n20) );
  NAND2_X1 cor_maj_140_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_140_n21) );
  NAND2_X1 cor_maj_140_U10 ( .A1(cor_maj_140_n21), .A2(cor_maj_140_n20), .ZN(
        cor_maj_140_n23) );
  XOR2_X1 cor_maj_140_U9 ( .A(v_1_2_3[2]), .B(cor_maj_140_n24), .Z(
        cor_maj_140_n26) );
  XOR2_X1 cor_maj_140_U8 ( .A(v_1_2_3[5]), .B(cor_maj_140_n25), .Z(
        cor_maj_140_n27) );
  XOR2_X1 cor_maj_140_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_140_n24)
         );
  XOR2_X1 cor_maj_140_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_140_n25)
         );
  OR2_X1 cor_maj_140_U5 ( .A1(cor_maj_140_n23), .A2(cor_maj_140_n22), .ZN(
        cor_maj_140_n32) );
  NAND2_X1 cor_maj_140_U4 ( .A1(cor_maj_140_n22), .A2(cor_maj_140_n23), .ZN(
        cor_maj_140_n34) );
  NAND2_X1 cor_maj_140_U3 ( .A1(cor_maj_140_n32), .A2(cor_maj_140_n31), .ZN(
        cor_maj_140_n33) );
  NAND2_X1 cor_maj_140_U2 ( .A1(cor_maj_140_n34), .A2(cor_maj_140_n33), .ZN(
        cor_maj_140_port_o) );
  OR2_X1 cor_maj_141_U19 ( .A1(cor_maj_141_n27), .A2(cor_maj_141_n26), .ZN(
        cor_maj_141_n28) );
  NAND2_X1 cor_maj_141_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_141_n28), .ZN(
        cor_maj_141_n29) );
  NAND2_X1 cor_maj_141_U17 ( .A1(cor_maj_141_n26), .A2(cor_maj_141_n27), .ZN(
        cor_maj_141_n30) );
  NAND2_X1 cor_maj_141_U16 ( .A1(cor_maj_141_n30), .A2(cor_maj_141_n29), .ZN(
        cor_maj_141_n31) );
  NAND2_X1 cor_maj_141_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_141_n25), .ZN(
        cor_maj_141_n18) );
  NAND2_X1 cor_maj_141_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_141_n19) );
  NAND2_X1 cor_maj_141_U13 ( .A1(cor_maj_141_n19), .A2(cor_maj_141_n18), .ZN(
        cor_maj_141_n22) );
  NAND2_X1 cor_maj_141_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_141_n24), .ZN(
        cor_maj_141_n20) );
  NAND2_X1 cor_maj_141_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_141_n21) );
  NAND2_X1 cor_maj_141_U10 ( .A1(cor_maj_141_n21), .A2(cor_maj_141_n20), .ZN(
        cor_maj_141_n23) );
  XOR2_X1 cor_maj_141_U9 ( .A(v_1_2_3[2]), .B(cor_maj_141_n24), .Z(
        cor_maj_141_n26) );
  XOR2_X1 cor_maj_141_U8 ( .A(v_1_2_3[5]), .B(cor_maj_141_n25), .Z(
        cor_maj_141_n27) );
  XOR2_X1 cor_maj_141_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_141_n24)
         );
  XOR2_X1 cor_maj_141_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_141_n25)
         );
  OR2_X1 cor_maj_141_U5 ( .A1(cor_maj_141_n23), .A2(cor_maj_141_n22), .ZN(
        cor_maj_141_n32) );
  NAND2_X1 cor_maj_141_U4 ( .A1(cor_maj_141_n22), .A2(cor_maj_141_n23), .ZN(
        cor_maj_141_n34) );
  NAND2_X1 cor_maj_141_U3 ( .A1(cor_maj_141_n32), .A2(cor_maj_141_n31), .ZN(
        cor_maj_141_n33) );
  NAND2_X1 cor_maj_141_U2 ( .A1(cor_maj_141_n34), .A2(cor_maj_141_n33), .ZN(
        cor_maj_141_port_o) );
  OR2_X1 cor_maj_142_U19 ( .A1(cor_maj_142_n27), .A2(cor_maj_142_n26), .ZN(
        cor_maj_142_n28) );
  NAND2_X1 cor_maj_142_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_142_n28), .ZN(
        cor_maj_142_n29) );
  NAND2_X1 cor_maj_142_U17 ( .A1(cor_maj_142_n26), .A2(cor_maj_142_n27), .ZN(
        cor_maj_142_n30) );
  NAND2_X1 cor_maj_142_U16 ( .A1(cor_maj_142_n30), .A2(cor_maj_142_n29), .ZN(
        cor_maj_142_n31) );
  NAND2_X1 cor_maj_142_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_142_n25), .ZN(
        cor_maj_142_n18) );
  NAND2_X1 cor_maj_142_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_142_n19) );
  NAND2_X1 cor_maj_142_U13 ( .A1(cor_maj_142_n19), .A2(cor_maj_142_n18), .ZN(
        cor_maj_142_n22) );
  NAND2_X1 cor_maj_142_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_142_n24), .ZN(
        cor_maj_142_n20) );
  NAND2_X1 cor_maj_142_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_142_n21) );
  NAND2_X1 cor_maj_142_U10 ( .A1(cor_maj_142_n21), .A2(cor_maj_142_n20), .ZN(
        cor_maj_142_n23) );
  XOR2_X1 cor_maj_142_U9 ( .A(v_1_2_3[2]), .B(cor_maj_142_n24), .Z(
        cor_maj_142_n26) );
  XOR2_X1 cor_maj_142_U8 ( .A(v_1_2_3[5]), .B(cor_maj_142_n25), .Z(
        cor_maj_142_n27) );
  XOR2_X1 cor_maj_142_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_142_n24)
         );
  XOR2_X1 cor_maj_142_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_142_n25)
         );
  OR2_X1 cor_maj_142_U5 ( .A1(cor_maj_142_n23), .A2(cor_maj_142_n22), .ZN(
        cor_maj_142_n32) );
  NAND2_X1 cor_maj_142_U4 ( .A1(cor_maj_142_n22), .A2(cor_maj_142_n23), .ZN(
        cor_maj_142_n34) );
  NAND2_X1 cor_maj_142_U3 ( .A1(cor_maj_142_n32), .A2(cor_maj_142_n31), .ZN(
        cor_maj_142_n33) );
  NAND2_X1 cor_maj_142_U2 ( .A1(cor_maj_142_n34), .A2(cor_maj_142_n33), .ZN(
        cor_maj_142_port_o) );
  OR2_X1 cor_maj_143_U19 ( .A1(cor_maj_143_n27), .A2(cor_maj_143_n26), .ZN(
        cor_maj_143_n28) );
  NAND2_X1 cor_maj_143_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_143_n28), .ZN(
        cor_maj_143_n29) );
  NAND2_X1 cor_maj_143_U17 ( .A1(cor_maj_143_n26), .A2(cor_maj_143_n27), .ZN(
        cor_maj_143_n30) );
  NAND2_X1 cor_maj_143_U16 ( .A1(cor_maj_143_n30), .A2(cor_maj_143_n29), .ZN(
        cor_maj_143_n31) );
  NAND2_X1 cor_maj_143_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_143_n25), .ZN(
        cor_maj_143_n18) );
  NAND2_X1 cor_maj_143_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_143_n19) );
  NAND2_X1 cor_maj_143_U13 ( .A1(cor_maj_143_n19), .A2(cor_maj_143_n18), .ZN(
        cor_maj_143_n22) );
  NAND2_X1 cor_maj_143_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_143_n24), .ZN(
        cor_maj_143_n20) );
  NAND2_X1 cor_maj_143_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_143_n21) );
  NAND2_X1 cor_maj_143_U10 ( .A1(cor_maj_143_n21), .A2(cor_maj_143_n20), .ZN(
        cor_maj_143_n23) );
  XOR2_X1 cor_maj_143_U9 ( .A(v_1_2_3[2]), .B(cor_maj_143_n24), .Z(
        cor_maj_143_n26) );
  XOR2_X1 cor_maj_143_U8 ( .A(v_1_2_3[5]), .B(cor_maj_143_n25), .Z(
        cor_maj_143_n27) );
  XOR2_X1 cor_maj_143_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_143_n24)
         );
  XOR2_X1 cor_maj_143_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_143_n25)
         );
  OR2_X1 cor_maj_143_U5 ( .A1(cor_maj_143_n23), .A2(cor_maj_143_n22), .ZN(
        cor_maj_143_n32) );
  NAND2_X1 cor_maj_143_U4 ( .A1(cor_maj_143_n22), .A2(cor_maj_143_n23), .ZN(
        cor_maj_143_n34) );
  NAND2_X1 cor_maj_143_U3 ( .A1(cor_maj_143_n32), .A2(cor_maj_143_n31), .ZN(
        cor_maj_143_n33) );
  NAND2_X1 cor_maj_143_U2 ( .A1(cor_maj_143_n34), .A2(cor_maj_143_n33), .ZN(
        cor_maj_143_port_o) );
  OR2_X1 cor_maj_144_U19 ( .A1(cor_maj_144_n27), .A2(cor_maj_144_n26), .ZN(
        cor_maj_144_n28) );
  NAND2_X1 cor_maj_144_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_144_n28), .ZN(
        cor_maj_144_n29) );
  NAND2_X1 cor_maj_144_U17 ( .A1(cor_maj_144_n26), .A2(cor_maj_144_n27), .ZN(
        cor_maj_144_n30) );
  NAND2_X1 cor_maj_144_U16 ( .A1(cor_maj_144_n30), .A2(cor_maj_144_n29), .ZN(
        cor_maj_144_n31) );
  NAND2_X1 cor_maj_144_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_144_n25), .ZN(
        cor_maj_144_n18) );
  NAND2_X1 cor_maj_144_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_144_n19) );
  NAND2_X1 cor_maj_144_U13 ( .A1(cor_maj_144_n19), .A2(cor_maj_144_n18), .ZN(
        cor_maj_144_n22) );
  NAND2_X1 cor_maj_144_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_144_n24), .ZN(
        cor_maj_144_n20) );
  NAND2_X1 cor_maj_144_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_144_n21) );
  NAND2_X1 cor_maj_144_U10 ( .A1(cor_maj_144_n21), .A2(cor_maj_144_n20), .ZN(
        cor_maj_144_n23) );
  XOR2_X1 cor_maj_144_U9 ( .A(v_1_2_3[2]), .B(cor_maj_144_n24), .Z(
        cor_maj_144_n26) );
  XOR2_X1 cor_maj_144_U8 ( .A(v_1_2_3[5]), .B(cor_maj_144_n25), .Z(
        cor_maj_144_n27) );
  XOR2_X1 cor_maj_144_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_144_n24)
         );
  XOR2_X1 cor_maj_144_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_144_n25)
         );
  OR2_X1 cor_maj_144_U5 ( .A1(cor_maj_144_n23), .A2(cor_maj_144_n22), .ZN(
        cor_maj_144_n32) );
  NAND2_X1 cor_maj_144_U4 ( .A1(cor_maj_144_n22), .A2(cor_maj_144_n23), .ZN(
        cor_maj_144_n34) );
  NAND2_X1 cor_maj_144_U3 ( .A1(cor_maj_144_n32), .A2(cor_maj_144_n31), .ZN(
        cor_maj_144_n33) );
  NAND2_X1 cor_maj_144_U2 ( .A1(cor_maj_144_n34), .A2(cor_maj_144_n33), .ZN(
        cor_maj_144_port_o) );
  OR2_X1 cor_maj_145_U19 ( .A1(cor_maj_145_n27), .A2(cor_maj_145_n26), .ZN(
        cor_maj_145_n28) );
  NAND2_X1 cor_maj_145_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_145_n28), .ZN(
        cor_maj_145_n29) );
  NAND2_X1 cor_maj_145_U17 ( .A1(cor_maj_145_n26), .A2(cor_maj_145_n27), .ZN(
        cor_maj_145_n30) );
  NAND2_X1 cor_maj_145_U16 ( .A1(cor_maj_145_n30), .A2(cor_maj_145_n29), .ZN(
        cor_maj_145_n31) );
  NAND2_X1 cor_maj_145_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_145_n25), .ZN(
        cor_maj_145_n18) );
  NAND2_X1 cor_maj_145_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_145_n19) );
  NAND2_X1 cor_maj_145_U13 ( .A1(cor_maj_145_n19), .A2(cor_maj_145_n18), .ZN(
        cor_maj_145_n22) );
  NAND2_X1 cor_maj_145_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_145_n24), .ZN(
        cor_maj_145_n20) );
  NAND2_X1 cor_maj_145_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_145_n21) );
  NAND2_X1 cor_maj_145_U10 ( .A1(cor_maj_145_n21), .A2(cor_maj_145_n20), .ZN(
        cor_maj_145_n23) );
  XOR2_X1 cor_maj_145_U9 ( .A(v_1_2_3[2]), .B(cor_maj_145_n24), .Z(
        cor_maj_145_n26) );
  XOR2_X1 cor_maj_145_U8 ( .A(v_1_2_3[5]), .B(cor_maj_145_n25), .Z(
        cor_maj_145_n27) );
  XOR2_X1 cor_maj_145_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_145_n24)
         );
  XOR2_X1 cor_maj_145_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_145_n25)
         );
  OR2_X1 cor_maj_145_U5 ( .A1(cor_maj_145_n23), .A2(cor_maj_145_n22), .ZN(
        cor_maj_145_n32) );
  NAND2_X1 cor_maj_145_U4 ( .A1(cor_maj_145_n22), .A2(cor_maj_145_n23), .ZN(
        cor_maj_145_n34) );
  NAND2_X1 cor_maj_145_U3 ( .A1(cor_maj_145_n32), .A2(cor_maj_145_n31), .ZN(
        cor_maj_145_n33) );
  NAND2_X1 cor_maj_145_U2 ( .A1(cor_maj_145_n34), .A2(cor_maj_145_n33), .ZN(
        cor_maj_145_port_o) );
  OR2_X1 cor_maj_146_U19 ( .A1(cor_maj_146_n27), .A2(cor_maj_146_n26), .ZN(
        cor_maj_146_n28) );
  NAND2_X1 cor_maj_146_U18 ( .A1(v_1_2_3[6]), .A2(cor_maj_146_n28), .ZN(
        cor_maj_146_n29) );
  NAND2_X1 cor_maj_146_U17 ( .A1(cor_maj_146_n26), .A2(cor_maj_146_n27), .ZN(
        cor_maj_146_n30) );
  NAND2_X1 cor_maj_146_U16 ( .A1(cor_maj_146_n30), .A2(cor_maj_146_n29), .ZN(
        cor_maj_146_n31) );
  NAND2_X1 cor_maj_146_U15 ( .A1(v_1_2_3[5]), .A2(cor_maj_146_n25), .ZN(
        cor_maj_146_n18) );
  NAND2_X1 cor_maj_146_U14 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_146_n19) );
  NAND2_X1 cor_maj_146_U13 ( .A1(cor_maj_146_n19), .A2(cor_maj_146_n18), .ZN(
        cor_maj_146_n22) );
  NAND2_X1 cor_maj_146_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_146_n24), .ZN(
        cor_maj_146_n20) );
  NAND2_X1 cor_maj_146_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_146_n21) );
  NAND2_X1 cor_maj_146_U10 ( .A1(cor_maj_146_n21), .A2(cor_maj_146_n20), .ZN(
        cor_maj_146_n23) );
  XOR2_X1 cor_maj_146_U9 ( .A(v_1_2_3[2]), .B(cor_maj_146_n24), .Z(
        cor_maj_146_n26) );
  XOR2_X1 cor_maj_146_U8 ( .A(v_1_2_3[5]), .B(cor_maj_146_n25), .Z(
        cor_maj_146_n27) );
  XOR2_X1 cor_maj_146_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_146_n24)
         );
  XOR2_X1 cor_maj_146_U6 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_146_n25)
         );
  OR2_X1 cor_maj_146_U5 ( .A1(cor_maj_146_n23), .A2(cor_maj_146_n22), .ZN(
        cor_maj_146_n32) );
  NAND2_X1 cor_maj_146_U4 ( .A1(cor_maj_146_n22), .A2(cor_maj_146_n23), .ZN(
        cor_maj_146_n34) );
  NAND2_X1 cor_maj_146_U3 ( .A1(cor_maj_146_n32), .A2(cor_maj_146_n31), .ZN(
        cor_maj_146_n33) );
  NAND2_X1 cor_maj_146_U2 ( .A1(cor_maj_146_n34), .A2(cor_maj_146_n33), .ZN(
        cor_maj_146_port_o) );
  OR2_X1 cor_maj_147_U19 ( .A1(cor_maj_147_n27), .A2(cor_maj_147_n26), .ZN(
        cor_maj_147_n28) );
  NAND2_X1 cor_maj_147_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_147_n28), .ZN(
        cor_maj_147_n29) );
  NAND2_X1 cor_maj_147_U17 ( .A1(cor_maj_147_n26), .A2(cor_maj_147_n27), .ZN(
        cor_maj_147_n30) );
  NAND2_X1 cor_maj_147_U16 ( .A1(cor_maj_147_n30), .A2(cor_maj_147_n29), .ZN(
        cor_maj_147_n31) );
  NAND2_X1 cor_maj_147_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_147_n25), .ZN(
        cor_maj_147_n18) );
  NAND2_X1 cor_maj_147_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_147_n19) );
  NAND2_X1 cor_maj_147_U13 ( .A1(cor_maj_147_n19), .A2(cor_maj_147_n18), .ZN(
        cor_maj_147_n22) );
  NAND2_X1 cor_maj_147_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_147_n24), .ZN(
        cor_maj_147_n20) );
  NAND2_X1 cor_maj_147_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_147_n21) );
  NAND2_X1 cor_maj_147_U10 ( .A1(cor_maj_147_n21), .A2(cor_maj_147_n20), .ZN(
        cor_maj_147_n23) );
  XOR2_X1 cor_maj_147_U9 ( .A(v_1_3_0[2]), .B(cor_maj_147_n24), .Z(
        cor_maj_147_n26) );
  XOR2_X1 cor_maj_147_U8 ( .A(v_1_3_0[5]), .B(cor_maj_147_n25), .Z(
        cor_maj_147_n27) );
  XOR2_X1 cor_maj_147_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_147_n24)
         );
  XOR2_X1 cor_maj_147_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_147_n25)
         );
  OR2_X1 cor_maj_147_U5 ( .A1(cor_maj_147_n23), .A2(cor_maj_147_n22), .ZN(
        cor_maj_147_n32) );
  NAND2_X1 cor_maj_147_U4 ( .A1(cor_maj_147_n22), .A2(cor_maj_147_n23), .ZN(
        cor_maj_147_n34) );
  NAND2_X1 cor_maj_147_U3 ( .A1(cor_maj_147_n32), .A2(cor_maj_147_n31), .ZN(
        cor_maj_147_n33) );
  NAND2_X1 cor_maj_147_U2 ( .A1(cor_maj_147_n34), .A2(cor_maj_147_n33), .ZN(
        cor_maj_147_port_o) );
  OR2_X1 cor_maj_148_U19 ( .A1(cor_maj_148_n27), .A2(cor_maj_148_n26), .ZN(
        cor_maj_148_n28) );
  NAND2_X1 cor_maj_148_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_148_n28), .ZN(
        cor_maj_148_n29) );
  NAND2_X1 cor_maj_148_U17 ( .A1(cor_maj_148_n26), .A2(cor_maj_148_n27), .ZN(
        cor_maj_148_n30) );
  NAND2_X1 cor_maj_148_U16 ( .A1(cor_maj_148_n30), .A2(cor_maj_148_n29), .ZN(
        cor_maj_148_n31) );
  NAND2_X1 cor_maj_148_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_148_n25), .ZN(
        cor_maj_148_n18) );
  NAND2_X1 cor_maj_148_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_148_n19) );
  NAND2_X1 cor_maj_148_U13 ( .A1(cor_maj_148_n19), .A2(cor_maj_148_n18), .ZN(
        cor_maj_148_n22) );
  NAND2_X1 cor_maj_148_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_148_n24), .ZN(
        cor_maj_148_n20) );
  NAND2_X1 cor_maj_148_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_148_n21) );
  NAND2_X1 cor_maj_148_U10 ( .A1(cor_maj_148_n21), .A2(cor_maj_148_n20), .ZN(
        cor_maj_148_n23) );
  XOR2_X1 cor_maj_148_U9 ( .A(v_1_3_0[2]), .B(cor_maj_148_n24), .Z(
        cor_maj_148_n26) );
  XOR2_X1 cor_maj_148_U8 ( .A(v_1_3_0[5]), .B(cor_maj_148_n25), .Z(
        cor_maj_148_n27) );
  XOR2_X1 cor_maj_148_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_148_n24)
         );
  XOR2_X1 cor_maj_148_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_148_n25)
         );
  OR2_X1 cor_maj_148_U5 ( .A1(cor_maj_148_n23), .A2(cor_maj_148_n22), .ZN(
        cor_maj_148_n32) );
  NAND2_X1 cor_maj_148_U4 ( .A1(cor_maj_148_n22), .A2(cor_maj_148_n23), .ZN(
        cor_maj_148_n34) );
  NAND2_X1 cor_maj_148_U3 ( .A1(cor_maj_148_n32), .A2(cor_maj_148_n31), .ZN(
        cor_maj_148_n33) );
  NAND2_X1 cor_maj_148_U2 ( .A1(cor_maj_148_n34), .A2(cor_maj_148_n33), .ZN(
        cor_maj_148_port_o) );
  OR2_X1 cor_maj_149_U19 ( .A1(cor_maj_149_n27), .A2(cor_maj_149_n26), .ZN(
        cor_maj_149_n28) );
  NAND2_X1 cor_maj_149_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_149_n28), .ZN(
        cor_maj_149_n29) );
  NAND2_X1 cor_maj_149_U17 ( .A1(cor_maj_149_n26), .A2(cor_maj_149_n27), .ZN(
        cor_maj_149_n30) );
  NAND2_X1 cor_maj_149_U16 ( .A1(cor_maj_149_n30), .A2(cor_maj_149_n29), .ZN(
        cor_maj_149_n31) );
  NAND2_X1 cor_maj_149_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_149_n25), .ZN(
        cor_maj_149_n18) );
  NAND2_X1 cor_maj_149_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_149_n19) );
  NAND2_X1 cor_maj_149_U13 ( .A1(cor_maj_149_n19), .A2(cor_maj_149_n18), .ZN(
        cor_maj_149_n22) );
  NAND2_X1 cor_maj_149_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_149_n24), .ZN(
        cor_maj_149_n20) );
  NAND2_X1 cor_maj_149_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_149_n21) );
  NAND2_X1 cor_maj_149_U10 ( .A1(cor_maj_149_n21), .A2(cor_maj_149_n20), .ZN(
        cor_maj_149_n23) );
  XOR2_X1 cor_maj_149_U9 ( .A(v_1_3_0[2]), .B(cor_maj_149_n24), .Z(
        cor_maj_149_n26) );
  XOR2_X1 cor_maj_149_U8 ( .A(v_1_3_0[5]), .B(cor_maj_149_n25), .Z(
        cor_maj_149_n27) );
  XOR2_X1 cor_maj_149_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_149_n24)
         );
  XOR2_X1 cor_maj_149_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_149_n25)
         );
  OR2_X1 cor_maj_149_U5 ( .A1(cor_maj_149_n23), .A2(cor_maj_149_n22), .ZN(
        cor_maj_149_n32) );
  NAND2_X1 cor_maj_149_U4 ( .A1(cor_maj_149_n22), .A2(cor_maj_149_n23), .ZN(
        cor_maj_149_n34) );
  NAND2_X1 cor_maj_149_U3 ( .A1(cor_maj_149_n32), .A2(cor_maj_149_n31), .ZN(
        cor_maj_149_n33) );
  NAND2_X1 cor_maj_149_U2 ( .A1(cor_maj_149_n34), .A2(cor_maj_149_n33), .ZN(
        cor_maj_149_port_o) );
  OR2_X1 cor_maj_150_U19 ( .A1(cor_maj_150_n27), .A2(cor_maj_150_n26), .ZN(
        cor_maj_150_n28) );
  NAND2_X1 cor_maj_150_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_150_n28), .ZN(
        cor_maj_150_n29) );
  NAND2_X1 cor_maj_150_U17 ( .A1(cor_maj_150_n26), .A2(cor_maj_150_n27), .ZN(
        cor_maj_150_n30) );
  NAND2_X1 cor_maj_150_U16 ( .A1(cor_maj_150_n30), .A2(cor_maj_150_n29), .ZN(
        cor_maj_150_n31) );
  NAND2_X1 cor_maj_150_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_150_n25), .ZN(
        cor_maj_150_n18) );
  NAND2_X1 cor_maj_150_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_150_n19) );
  NAND2_X1 cor_maj_150_U13 ( .A1(cor_maj_150_n19), .A2(cor_maj_150_n18), .ZN(
        cor_maj_150_n22) );
  NAND2_X1 cor_maj_150_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_150_n24), .ZN(
        cor_maj_150_n20) );
  NAND2_X1 cor_maj_150_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_150_n21) );
  NAND2_X1 cor_maj_150_U10 ( .A1(cor_maj_150_n21), .A2(cor_maj_150_n20), .ZN(
        cor_maj_150_n23) );
  XOR2_X1 cor_maj_150_U9 ( .A(v_1_3_0[2]), .B(cor_maj_150_n24), .Z(
        cor_maj_150_n26) );
  XOR2_X1 cor_maj_150_U8 ( .A(v_1_3_0[5]), .B(cor_maj_150_n25), .Z(
        cor_maj_150_n27) );
  XOR2_X1 cor_maj_150_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_150_n24)
         );
  XOR2_X1 cor_maj_150_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_150_n25)
         );
  OR2_X1 cor_maj_150_U5 ( .A1(cor_maj_150_n23), .A2(cor_maj_150_n22), .ZN(
        cor_maj_150_n32) );
  NAND2_X1 cor_maj_150_U4 ( .A1(cor_maj_150_n22), .A2(cor_maj_150_n23), .ZN(
        cor_maj_150_n34) );
  NAND2_X1 cor_maj_150_U3 ( .A1(cor_maj_150_n32), .A2(cor_maj_150_n31), .ZN(
        cor_maj_150_n33) );
  NAND2_X1 cor_maj_150_U2 ( .A1(cor_maj_150_n34), .A2(cor_maj_150_n33), .ZN(
        cor_maj_150_port_o) );
  OR2_X1 cor_maj_151_U19 ( .A1(cor_maj_151_n27), .A2(cor_maj_151_n26), .ZN(
        cor_maj_151_n28) );
  NAND2_X1 cor_maj_151_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_151_n28), .ZN(
        cor_maj_151_n29) );
  NAND2_X1 cor_maj_151_U17 ( .A1(cor_maj_151_n26), .A2(cor_maj_151_n27), .ZN(
        cor_maj_151_n30) );
  NAND2_X1 cor_maj_151_U16 ( .A1(cor_maj_151_n30), .A2(cor_maj_151_n29), .ZN(
        cor_maj_151_n31) );
  NAND2_X1 cor_maj_151_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_151_n25), .ZN(
        cor_maj_151_n18) );
  NAND2_X1 cor_maj_151_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_151_n19) );
  NAND2_X1 cor_maj_151_U13 ( .A1(cor_maj_151_n19), .A2(cor_maj_151_n18), .ZN(
        cor_maj_151_n22) );
  NAND2_X1 cor_maj_151_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_151_n24), .ZN(
        cor_maj_151_n20) );
  NAND2_X1 cor_maj_151_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_151_n21) );
  NAND2_X1 cor_maj_151_U10 ( .A1(cor_maj_151_n21), .A2(cor_maj_151_n20), .ZN(
        cor_maj_151_n23) );
  XOR2_X1 cor_maj_151_U9 ( .A(v_1_3_0[2]), .B(cor_maj_151_n24), .Z(
        cor_maj_151_n26) );
  XOR2_X1 cor_maj_151_U8 ( .A(v_1_3_0[5]), .B(cor_maj_151_n25), .Z(
        cor_maj_151_n27) );
  XOR2_X1 cor_maj_151_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_151_n24)
         );
  XOR2_X1 cor_maj_151_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_151_n25)
         );
  OR2_X1 cor_maj_151_U5 ( .A1(cor_maj_151_n23), .A2(cor_maj_151_n22), .ZN(
        cor_maj_151_n32) );
  NAND2_X1 cor_maj_151_U4 ( .A1(cor_maj_151_n22), .A2(cor_maj_151_n23), .ZN(
        cor_maj_151_n34) );
  NAND2_X1 cor_maj_151_U3 ( .A1(cor_maj_151_n32), .A2(cor_maj_151_n31), .ZN(
        cor_maj_151_n33) );
  NAND2_X1 cor_maj_151_U2 ( .A1(cor_maj_151_n34), .A2(cor_maj_151_n33), .ZN(
        cor_maj_151_port_o) );
  OR2_X1 cor_maj_152_U19 ( .A1(cor_maj_152_n27), .A2(cor_maj_152_n26), .ZN(
        cor_maj_152_n28) );
  NAND2_X1 cor_maj_152_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_152_n28), .ZN(
        cor_maj_152_n29) );
  NAND2_X1 cor_maj_152_U17 ( .A1(cor_maj_152_n26), .A2(cor_maj_152_n27), .ZN(
        cor_maj_152_n30) );
  NAND2_X1 cor_maj_152_U16 ( .A1(cor_maj_152_n30), .A2(cor_maj_152_n29), .ZN(
        cor_maj_152_n31) );
  NAND2_X1 cor_maj_152_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_152_n25), .ZN(
        cor_maj_152_n18) );
  NAND2_X1 cor_maj_152_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_152_n19) );
  NAND2_X1 cor_maj_152_U13 ( .A1(cor_maj_152_n19), .A2(cor_maj_152_n18), .ZN(
        cor_maj_152_n22) );
  NAND2_X1 cor_maj_152_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_152_n24), .ZN(
        cor_maj_152_n20) );
  NAND2_X1 cor_maj_152_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_152_n21) );
  NAND2_X1 cor_maj_152_U10 ( .A1(cor_maj_152_n21), .A2(cor_maj_152_n20), .ZN(
        cor_maj_152_n23) );
  XOR2_X1 cor_maj_152_U9 ( .A(v_1_3_0[2]), .B(cor_maj_152_n24), .Z(
        cor_maj_152_n26) );
  XOR2_X1 cor_maj_152_U8 ( .A(v_1_3_0[5]), .B(cor_maj_152_n25), .Z(
        cor_maj_152_n27) );
  XOR2_X1 cor_maj_152_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_152_n24)
         );
  XOR2_X1 cor_maj_152_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_152_n25)
         );
  OR2_X1 cor_maj_152_U5 ( .A1(cor_maj_152_n23), .A2(cor_maj_152_n22), .ZN(
        cor_maj_152_n32) );
  NAND2_X1 cor_maj_152_U4 ( .A1(cor_maj_152_n22), .A2(cor_maj_152_n23), .ZN(
        cor_maj_152_n34) );
  NAND2_X1 cor_maj_152_U3 ( .A1(cor_maj_152_n32), .A2(cor_maj_152_n31), .ZN(
        cor_maj_152_n33) );
  NAND2_X1 cor_maj_152_U2 ( .A1(cor_maj_152_n34), .A2(cor_maj_152_n33), .ZN(
        cor_maj_152_port_o) );
  OR2_X1 cor_maj_153_U19 ( .A1(cor_maj_153_n27), .A2(cor_maj_153_n26), .ZN(
        cor_maj_153_n28) );
  NAND2_X1 cor_maj_153_U18 ( .A1(v_1_3_0[6]), .A2(cor_maj_153_n28), .ZN(
        cor_maj_153_n29) );
  NAND2_X1 cor_maj_153_U17 ( .A1(cor_maj_153_n26), .A2(cor_maj_153_n27), .ZN(
        cor_maj_153_n30) );
  NAND2_X1 cor_maj_153_U16 ( .A1(cor_maj_153_n30), .A2(cor_maj_153_n29), .ZN(
        cor_maj_153_n31) );
  NAND2_X1 cor_maj_153_U15 ( .A1(v_1_3_0[5]), .A2(cor_maj_153_n25), .ZN(
        cor_maj_153_n18) );
  NAND2_X1 cor_maj_153_U14 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_153_n19) );
  NAND2_X1 cor_maj_153_U13 ( .A1(cor_maj_153_n19), .A2(cor_maj_153_n18), .ZN(
        cor_maj_153_n22) );
  NAND2_X1 cor_maj_153_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_153_n24), .ZN(
        cor_maj_153_n20) );
  NAND2_X1 cor_maj_153_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_153_n21) );
  NAND2_X1 cor_maj_153_U10 ( .A1(cor_maj_153_n21), .A2(cor_maj_153_n20), .ZN(
        cor_maj_153_n23) );
  XOR2_X1 cor_maj_153_U9 ( .A(v_1_3_0[2]), .B(cor_maj_153_n24), .Z(
        cor_maj_153_n26) );
  XOR2_X1 cor_maj_153_U8 ( .A(v_1_3_0[5]), .B(cor_maj_153_n25), .Z(
        cor_maj_153_n27) );
  XOR2_X1 cor_maj_153_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_153_n24)
         );
  XOR2_X1 cor_maj_153_U6 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_153_n25)
         );
  OR2_X1 cor_maj_153_U5 ( .A1(cor_maj_153_n23), .A2(cor_maj_153_n22), .ZN(
        cor_maj_153_n32) );
  NAND2_X1 cor_maj_153_U4 ( .A1(cor_maj_153_n22), .A2(cor_maj_153_n23), .ZN(
        cor_maj_153_n34) );
  NAND2_X1 cor_maj_153_U3 ( .A1(cor_maj_153_n32), .A2(cor_maj_153_n31), .ZN(
        cor_maj_153_n33) );
  NAND2_X1 cor_maj_153_U2 ( .A1(cor_maj_153_n34), .A2(cor_maj_153_n33), .ZN(
        cor_maj_153_port_o) );
  OR2_X1 cor_maj_154_U19 ( .A1(cor_maj_154_n27), .A2(cor_maj_154_n26), .ZN(
        cor_maj_154_n28) );
  NAND2_X1 cor_maj_154_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_154_n28), .ZN(
        cor_maj_154_n29) );
  NAND2_X1 cor_maj_154_U17 ( .A1(cor_maj_154_n26), .A2(cor_maj_154_n27), .ZN(
        cor_maj_154_n30) );
  NAND2_X1 cor_maj_154_U16 ( .A1(cor_maj_154_n30), .A2(cor_maj_154_n29), .ZN(
        cor_maj_154_n31) );
  NAND2_X1 cor_maj_154_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_154_n25), .ZN(
        cor_maj_154_n18) );
  NAND2_X1 cor_maj_154_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_154_n19) );
  NAND2_X1 cor_maj_154_U13 ( .A1(cor_maj_154_n19), .A2(cor_maj_154_n18), .ZN(
        cor_maj_154_n22) );
  NAND2_X1 cor_maj_154_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_154_n24), .ZN(
        cor_maj_154_n20) );
  NAND2_X1 cor_maj_154_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_154_n21) );
  NAND2_X1 cor_maj_154_U10 ( .A1(cor_maj_154_n21), .A2(cor_maj_154_n20), .ZN(
        cor_maj_154_n23) );
  XOR2_X1 cor_maj_154_U9 ( .A(v_1_3_1[2]), .B(cor_maj_154_n24), .Z(
        cor_maj_154_n26) );
  XOR2_X1 cor_maj_154_U8 ( .A(v_1_3_1[5]), .B(cor_maj_154_n25), .Z(
        cor_maj_154_n27) );
  XOR2_X1 cor_maj_154_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_154_n24)
         );
  XOR2_X1 cor_maj_154_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_154_n25)
         );
  OR2_X1 cor_maj_154_U5 ( .A1(cor_maj_154_n23), .A2(cor_maj_154_n22), .ZN(
        cor_maj_154_n32) );
  NAND2_X1 cor_maj_154_U4 ( .A1(cor_maj_154_n22), .A2(cor_maj_154_n23), .ZN(
        cor_maj_154_n34) );
  NAND2_X1 cor_maj_154_U3 ( .A1(cor_maj_154_n32), .A2(cor_maj_154_n31), .ZN(
        cor_maj_154_n33) );
  NAND2_X1 cor_maj_154_U2 ( .A1(cor_maj_154_n34), .A2(cor_maj_154_n33), .ZN(
        cor_maj_154_port_o) );
  OR2_X1 cor_maj_155_U19 ( .A1(cor_maj_155_n27), .A2(cor_maj_155_n26), .ZN(
        cor_maj_155_n28) );
  NAND2_X1 cor_maj_155_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_155_n28), .ZN(
        cor_maj_155_n29) );
  NAND2_X1 cor_maj_155_U17 ( .A1(cor_maj_155_n26), .A2(cor_maj_155_n27), .ZN(
        cor_maj_155_n30) );
  NAND2_X1 cor_maj_155_U16 ( .A1(cor_maj_155_n30), .A2(cor_maj_155_n29), .ZN(
        cor_maj_155_n31) );
  NAND2_X1 cor_maj_155_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_155_n25), .ZN(
        cor_maj_155_n18) );
  NAND2_X1 cor_maj_155_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_155_n19) );
  NAND2_X1 cor_maj_155_U13 ( .A1(cor_maj_155_n19), .A2(cor_maj_155_n18), .ZN(
        cor_maj_155_n22) );
  NAND2_X1 cor_maj_155_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_155_n24), .ZN(
        cor_maj_155_n20) );
  NAND2_X1 cor_maj_155_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_155_n21) );
  NAND2_X1 cor_maj_155_U10 ( .A1(cor_maj_155_n21), .A2(cor_maj_155_n20), .ZN(
        cor_maj_155_n23) );
  XOR2_X1 cor_maj_155_U9 ( .A(v_1_3_1[2]), .B(cor_maj_155_n24), .Z(
        cor_maj_155_n26) );
  XOR2_X1 cor_maj_155_U8 ( .A(v_1_3_1[5]), .B(cor_maj_155_n25), .Z(
        cor_maj_155_n27) );
  XOR2_X1 cor_maj_155_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_155_n24)
         );
  XOR2_X1 cor_maj_155_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_155_n25)
         );
  OR2_X1 cor_maj_155_U5 ( .A1(cor_maj_155_n23), .A2(cor_maj_155_n22), .ZN(
        cor_maj_155_n32) );
  NAND2_X1 cor_maj_155_U4 ( .A1(cor_maj_155_n22), .A2(cor_maj_155_n23), .ZN(
        cor_maj_155_n34) );
  NAND2_X1 cor_maj_155_U3 ( .A1(cor_maj_155_n32), .A2(cor_maj_155_n31), .ZN(
        cor_maj_155_n33) );
  NAND2_X1 cor_maj_155_U2 ( .A1(cor_maj_155_n34), .A2(cor_maj_155_n33), .ZN(
        cor_maj_155_port_o) );
  OR2_X1 cor_maj_156_U19 ( .A1(cor_maj_156_n27), .A2(cor_maj_156_n26), .ZN(
        cor_maj_156_n28) );
  NAND2_X1 cor_maj_156_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_156_n28), .ZN(
        cor_maj_156_n29) );
  NAND2_X1 cor_maj_156_U17 ( .A1(cor_maj_156_n26), .A2(cor_maj_156_n27), .ZN(
        cor_maj_156_n30) );
  NAND2_X1 cor_maj_156_U16 ( .A1(cor_maj_156_n30), .A2(cor_maj_156_n29), .ZN(
        cor_maj_156_n31) );
  NAND2_X1 cor_maj_156_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_156_n25), .ZN(
        cor_maj_156_n18) );
  NAND2_X1 cor_maj_156_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_156_n19) );
  NAND2_X1 cor_maj_156_U13 ( .A1(cor_maj_156_n19), .A2(cor_maj_156_n18), .ZN(
        cor_maj_156_n22) );
  NAND2_X1 cor_maj_156_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_156_n24), .ZN(
        cor_maj_156_n20) );
  NAND2_X1 cor_maj_156_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_156_n21) );
  NAND2_X1 cor_maj_156_U10 ( .A1(cor_maj_156_n21), .A2(cor_maj_156_n20), .ZN(
        cor_maj_156_n23) );
  XOR2_X1 cor_maj_156_U9 ( .A(v_1_3_1[2]), .B(cor_maj_156_n24), .Z(
        cor_maj_156_n26) );
  XOR2_X1 cor_maj_156_U8 ( .A(v_1_3_1[5]), .B(cor_maj_156_n25), .Z(
        cor_maj_156_n27) );
  XOR2_X1 cor_maj_156_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_156_n24)
         );
  XOR2_X1 cor_maj_156_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_156_n25)
         );
  OR2_X1 cor_maj_156_U5 ( .A1(cor_maj_156_n23), .A2(cor_maj_156_n22), .ZN(
        cor_maj_156_n32) );
  NAND2_X1 cor_maj_156_U4 ( .A1(cor_maj_156_n22), .A2(cor_maj_156_n23), .ZN(
        cor_maj_156_n34) );
  NAND2_X1 cor_maj_156_U3 ( .A1(cor_maj_156_n32), .A2(cor_maj_156_n31), .ZN(
        cor_maj_156_n33) );
  NAND2_X1 cor_maj_156_U2 ( .A1(cor_maj_156_n34), .A2(cor_maj_156_n33), .ZN(
        cor_maj_156_port_o) );
  OR2_X1 cor_maj_157_U19 ( .A1(cor_maj_157_n27), .A2(cor_maj_157_n26), .ZN(
        cor_maj_157_n28) );
  NAND2_X1 cor_maj_157_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_157_n28), .ZN(
        cor_maj_157_n29) );
  NAND2_X1 cor_maj_157_U17 ( .A1(cor_maj_157_n26), .A2(cor_maj_157_n27), .ZN(
        cor_maj_157_n30) );
  NAND2_X1 cor_maj_157_U16 ( .A1(cor_maj_157_n30), .A2(cor_maj_157_n29), .ZN(
        cor_maj_157_n31) );
  NAND2_X1 cor_maj_157_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_157_n25), .ZN(
        cor_maj_157_n18) );
  NAND2_X1 cor_maj_157_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_157_n19) );
  NAND2_X1 cor_maj_157_U13 ( .A1(cor_maj_157_n19), .A2(cor_maj_157_n18), .ZN(
        cor_maj_157_n22) );
  NAND2_X1 cor_maj_157_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_157_n24), .ZN(
        cor_maj_157_n20) );
  NAND2_X1 cor_maj_157_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_157_n21) );
  NAND2_X1 cor_maj_157_U10 ( .A1(cor_maj_157_n21), .A2(cor_maj_157_n20), .ZN(
        cor_maj_157_n23) );
  XOR2_X1 cor_maj_157_U9 ( .A(v_1_3_1[2]), .B(cor_maj_157_n24), .Z(
        cor_maj_157_n26) );
  XOR2_X1 cor_maj_157_U8 ( .A(v_1_3_1[5]), .B(cor_maj_157_n25), .Z(
        cor_maj_157_n27) );
  XOR2_X1 cor_maj_157_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_157_n24)
         );
  XOR2_X1 cor_maj_157_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_157_n25)
         );
  OR2_X1 cor_maj_157_U5 ( .A1(cor_maj_157_n23), .A2(cor_maj_157_n22), .ZN(
        cor_maj_157_n32) );
  NAND2_X1 cor_maj_157_U4 ( .A1(cor_maj_157_n22), .A2(cor_maj_157_n23), .ZN(
        cor_maj_157_n34) );
  NAND2_X1 cor_maj_157_U3 ( .A1(cor_maj_157_n32), .A2(cor_maj_157_n31), .ZN(
        cor_maj_157_n33) );
  NAND2_X1 cor_maj_157_U2 ( .A1(cor_maj_157_n34), .A2(cor_maj_157_n33), .ZN(
        cor_maj_157_port_o) );
  OR2_X1 cor_maj_158_U19 ( .A1(cor_maj_158_n27), .A2(cor_maj_158_n26), .ZN(
        cor_maj_158_n28) );
  NAND2_X1 cor_maj_158_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_158_n28), .ZN(
        cor_maj_158_n29) );
  NAND2_X1 cor_maj_158_U17 ( .A1(cor_maj_158_n26), .A2(cor_maj_158_n27), .ZN(
        cor_maj_158_n30) );
  NAND2_X1 cor_maj_158_U16 ( .A1(cor_maj_158_n30), .A2(cor_maj_158_n29), .ZN(
        cor_maj_158_n31) );
  NAND2_X1 cor_maj_158_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_158_n25), .ZN(
        cor_maj_158_n18) );
  NAND2_X1 cor_maj_158_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_158_n19) );
  NAND2_X1 cor_maj_158_U13 ( .A1(cor_maj_158_n19), .A2(cor_maj_158_n18), .ZN(
        cor_maj_158_n22) );
  NAND2_X1 cor_maj_158_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_158_n24), .ZN(
        cor_maj_158_n20) );
  NAND2_X1 cor_maj_158_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_158_n21) );
  NAND2_X1 cor_maj_158_U10 ( .A1(cor_maj_158_n21), .A2(cor_maj_158_n20), .ZN(
        cor_maj_158_n23) );
  XOR2_X1 cor_maj_158_U9 ( .A(v_1_3_1[2]), .B(cor_maj_158_n24), .Z(
        cor_maj_158_n26) );
  XOR2_X1 cor_maj_158_U8 ( .A(v_1_3_1[5]), .B(cor_maj_158_n25), .Z(
        cor_maj_158_n27) );
  XOR2_X1 cor_maj_158_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_158_n24)
         );
  XOR2_X1 cor_maj_158_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_158_n25)
         );
  OR2_X1 cor_maj_158_U5 ( .A1(cor_maj_158_n23), .A2(cor_maj_158_n22), .ZN(
        cor_maj_158_n32) );
  NAND2_X1 cor_maj_158_U4 ( .A1(cor_maj_158_n22), .A2(cor_maj_158_n23), .ZN(
        cor_maj_158_n34) );
  NAND2_X1 cor_maj_158_U3 ( .A1(cor_maj_158_n32), .A2(cor_maj_158_n31), .ZN(
        cor_maj_158_n33) );
  NAND2_X1 cor_maj_158_U2 ( .A1(cor_maj_158_n34), .A2(cor_maj_158_n33), .ZN(
        cor_maj_158_port_o) );
  OR2_X1 cor_maj_159_U19 ( .A1(cor_maj_159_n27), .A2(cor_maj_159_n26), .ZN(
        cor_maj_159_n28) );
  NAND2_X1 cor_maj_159_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_159_n28), .ZN(
        cor_maj_159_n29) );
  NAND2_X1 cor_maj_159_U17 ( .A1(cor_maj_159_n26), .A2(cor_maj_159_n27), .ZN(
        cor_maj_159_n30) );
  NAND2_X1 cor_maj_159_U16 ( .A1(cor_maj_159_n30), .A2(cor_maj_159_n29), .ZN(
        cor_maj_159_n31) );
  NAND2_X1 cor_maj_159_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_159_n25), .ZN(
        cor_maj_159_n18) );
  NAND2_X1 cor_maj_159_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_159_n19) );
  NAND2_X1 cor_maj_159_U13 ( .A1(cor_maj_159_n19), .A2(cor_maj_159_n18), .ZN(
        cor_maj_159_n22) );
  NAND2_X1 cor_maj_159_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_159_n24), .ZN(
        cor_maj_159_n20) );
  NAND2_X1 cor_maj_159_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_159_n21) );
  NAND2_X1 cor_maj_159_U10 ( .A1(cor_maj_159_n21), .A2(cor_maj_159_n20), .ZN(
        cor_maj_159_n23) );
  XOR2_X1 cor_maj_159_U9 ( .A(v_1_3_1[2]), .B(cor_maj_159_n24), .Z(
        cor_maj_159_n26) );
  XOR2_X1 cor_maj_159_U8 ( .A(v_1_3_1[5]), .B(cor_maj_159_n25), .Z(
        cor_maj_159_n27) );
  XOR2_X1 cor_maj_159_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_159_n24)
         );
  XOR2_X1 cor_maj_159_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_159_n25)
         );
  OR2_X1 cor_maj_159_U5 ( .A1(cor_maj_159_n23), .A2(cor_maj_159_n22), .ZN(
        cor_maj_159_n32) );
  NAND2_X1 cor_maj_159_U4 ( .A1(cor_maj_159_n22), .A2(cor_maj_159_n23), .ZN(
        cor_maj_159_n34) );
  NAND2_X1 cor_maj_159_U3 ( .A1(cor_maj_159_n32), .A2(cor_maj_159_n31), .ZN(
        cor_maj_159_n33) );
  NAND2_X1 cor_maj_159_U2 ( .A1(cor_maj_159_n34), .A2(cor_maj_159_n33), .ZN(
        cor_maj_159_port_o) );
  OR2_X1 cor_maj_160_U19 ( .A1(cor_maj_160_n27), .A2(cor_maj_160_n26), .ZN(
        cor_maj_160_n28) );
  NAND2_X1 cor_maj_160_U18 ( .A1(v_1_3_1[6]), .A2(cor_maj_160_n28), .ZN(
        cor_maj_160_n29) );
  NAND2_X1 cor_maj_160_U17 ( .A1(cor_maj_160_n26), .A2(cor_maj_160_n27), .ZN(
        cor_maj_160_n30) );
  NAND2_X1 cor_maj_160_U16 ( .A1(cor_maj_160_n30), .A2(cor_maj_160_n29), .ZN(
        cor_maj_160_n31) );
  NAND2_X1 cor_maj_160_U15 ( .A1(v_1_3_1[5]), .A2(cor_maj_160_n25), .ZN(
        cor_maj_160_n18) );
  NAND2_X1 cor_maj_160_U14 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_160_n19) );
  NAND2_X1 cor_maj_160_U13 ( .A1(cor_maj_160_n19), .A2(cor_maj_160_n18), .ZN(
        cor_maj_160_n22) );
  NAND2_X1 cor_maj_160_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_160_n24), .ZN(
        cor_maj_160_n20) );
  NAND2_X1 cor_maj_160_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_160_n21) );
  NAND2_X1 cor_maj_160_U10 ( .A1(cor_maj_160_n21), .A2(cor_maj_160_n20), .ZN(
        cor_maj_160_n23) );
  XOR2_X1 cor_maj_160_U9 ( .A(v_1_3_1[2]), .B(cor_maj_160_n24), .Z(
        cor_maj_160_n26) );
  XOR2_X1 cor_maj_160_U8 ( .A(v_1_3_1[5]), .B(cor_maj_160_n25), .Z(
        cor_maj_160_n27) );
  XOR2_X1 cor_maj_160_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_160_n24)
         );
  XOR2_X1 cor_maj_160_U6 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_160_n25)
         );
  OR2_X1 cor_maj_160_U5 ( .A1(cor_maj_160_n23), .A2(cor_maj_160_n22), .ZN(
        cor_maj_160_n32) );
  NAND2_X1 cor_maj_160_U4 ( .A1(cor_maj_160_n22), .A2(cor_maj_160_n23), .ZN(
        cor_maj_160_n34) );
  NAND2_X1 cor_maj_160_U3 ( .A1(cor_maj_160_n32), .A2(cor_maj_160_n31), .ZN(
        cor_maj_160_n33) );
  NAND2_X1 cor_maj_160_U2 ( .A1(cor_maj_160_n34), .A2(cor_maj_160_n33), .ZN(
        cor_maj_160_port_o) );
  OR2_X1 cor_maj_161_U19 ( .A1(cor_maj_161_n27), .A2(cor_maj_161_n26), .ZN(
        cor_maj_161_n28) );
  NAND2_X1 cor_maj_161_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_161_n28), .ZN(
        cor_maj_161_n29) );
  NAND2_X1 cor_maj_161_U17 ( .A1(cor_maj_161_n26), .A2(cor_maj_161_n27), .ZN(
        cor_maj_161_n30) );
  NAND2_X1 cor_maj_161_U16 ( .A1(cor_maj_161_n30), .A2(cor_maj_161_n29), .ZN(
        cor_maj_161_n31) );
  NAND2_X1 cor_maj_161_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_161_n25), .ZN(
        cor_maj_161_n18) );
  NAND2_X1 cor_maj_161_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_161_n19) );
  NAND2_X1 cor_maj_161_U13 ( .A1(cor_maj_161_n19), .A2(cor_maj_161_n18), .ZN(
        cor_maj_161_n22) );
  NAND2_X1 cor_maj_161_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_161_n24), .ZN(
        cor_maj_161_n20) );
  NAND2_X1 cor_maj_161_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_161_n21) );
  NAND2_X1 cor_maj_161_U10 ( .A1(cor_maj_161_n21), .A2(cor_maj_161_n20), .ZN(
        cor_maj_161_n23) );
  XOR2_X1 cor_maj_161_U9 ( .A(v_1_3_2[2]), .B(cor_maj_161_n24), .Z(
        cor_maj_161_n26) );
  XOR2_X1 cor_maj_161_U8 ( .A(v_1_3_2[5]), .B(cor_maj_161_n25), .Z(
        cor_maj_161_n27) );
  XOR2_X1 cor_maj_161_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_161_n24)
         );
  XOR2_X1 cor_maj_161_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_161_n25)
         );
  OR2_X1 cor_maj_161_U5 ( .A1(cor_maj_161_n23), .A2(cor_maj_161_n22), .ZN(
        cor_maj_161_n32) );
  NAND2_X1 cor_maj_161_U4 ( .A1(cor_maj_161_n22), .A2(cor_maj_161_n23), .ZN(
        cor_maj_161_n34) );
  NAND2_X1 cor_maj_161_U3 ( .A1(cor_maj_161_n32), .A2(cor_maj_161_n31), .ZN(
        cor_maj_161_n33) );
  NAND2_X1 cor_maj_161_U2 ( .A1(cor_maj_161_n34), .A2(cor_maj_161_n33), .ZN(
        cor_maj_161_port_o) );
  OR2_X1 cor_maj_162_U19 ( .A1(cor_maj_162_n27), .A2(cor_maj_162_n26), .ZN(
        cor_maj_162_n28) );
  NAND2_X1 cor_maj_162_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_162_n28), .ZN(
        cor_maj_162_n29) );
  NAND2_X1 cor_maj_162_U17 ( .A1(cor_maj_162_n26), .A2(cor_maj_162_n27), .ZN(
        cor_maj_162_n30) );
  NAND2_X1 cor_maj_162_U16 ( .A1(cor_maj_162_n30), .A2(cor_maj_162_n29), .ZN(
        cor_maj_162_n31) );
  NAND2_X1 cor_maj_162_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_162_n25), .ZN(
        cor_maj_162_n18) );
  NAND2_X1 cor_maj_162_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_162_n19) );
  NAND2_X1 cor_maj_162_U13 ( .A1(cor_maj_162_n19), .A2(cor_maj_162_n18), .ZN(
        cor_maj_162_n22) );
  NAND2_X1 cor_maj_162_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_162_n24), .ZN(
        cor_maj_162_n20) );
  NAND2_X1 cor_maj_162_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_162_n21) );
  NAND2_X1 cor_maj_162_U10 ( .A1(cor_maj_162_n21), .A2(cor_maj_162_n20), .ZN(
        cor_maj_162_n23) );
  XOR2_X1 cor_maj_162_U9 ( .A(v_1_3_2[2]), .B(cor_maj_162_n24), .Z(
        cor_maj_162_n26) );
  XOR2_X1 cor_maj_162_U8 ( .A(v_1_3_2[5]), .B(cor_maj_162_n25), .Z(
        cor_maj_162_n27) );
  XOR2_X1 cor_maj_162_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_162_n24)
         );
  XOR2_X1 cor_maj_162_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_162_n25)
         );
  OR2_X1 cor_maj_162_U5 ( .A1(cor_maj_162_n23), .A2(cor_maj_162_n22), .ZN(
        cor_maj_162_n32) );
  NAND2_X1 cor_maj_162_U4 ( .A1(cor_maj_162_n22), .A2(cor_maj_162_n23), .ZN(
        cor_maj_162_n34) );
  NAND2_X1 cor_maj_162_U3 ( .A1(cor_maj_162_n32), .A2(cor_maj_162_n31), .ZN(
        cor_maj_162_n33) );
  NAND2_X1 cor_maj_162_U2 ( .A1(cor_maj_162_n34), .A2(cor_maj_162_n33), .ZN(
        cor_maj_162_port_o) );
  OR2_X1 cor_maj_163_U19 ( .A1(cor_maj_163_n27), .A2(cor_maj_163_n26), .ZN(
        cor_maj_163_n28) );
  NAND2_X1 cor_maj_163_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_163_n28), .ZN(
        cor_maj_163_n29) );
  NAND2_X1 cor_maj_163_U17 ( .A1(cor_maj_163_n26), .A2(cor_maj_163_n27), .ZN(
        cor_maj_163_n30) );
  NAND2_X1 cor_maj_163_U16 ( .A1(cor_maj_163_n30), .A2(cor_maj_163_n29), .ZN(
        cor_maj_163_n31) );
  NAND2_X1 cor_maj_163_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_163_n25), .ZN(
        cor_maj_163_n18) );
  NAND2_X1 cor_maj_163_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_163_n19) );
  NAND2_X1 cor_maj_163_U13 ( .A1(cor_maj_163_n19), .A2(cor_maj_163_n18), .ZN(
        cor_maj_163_n22) );
  NAND2_X1 cor_maj_163_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_163_n24), .ZN(
        cor_maj_163_n20) );
  NAND2_X1 cor_maj_163_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_163_n21) );
  NAND2_X1 cor_maj_163_U10 ( .A1(cor_maj_163_n21), .A2(cor_maj_163_n20), .ZN(
        cor_maj_163_n23) );
  XOR2_X1 cor_maj_163_U9 ( .A(v_1_3_2[2]), .B(cor_maj_163_n24), .Z(
        cor_maj_163_n26) );
  XOR2_X1 cor_maj_163_U8 ( .A(v_1_3_2[5]), .B(cor_maj_163_n25), .Z(
        cor_maj_163_n27) );
  XOR2_X1 cor_maj_163_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_163_n24)
         );
  XOR2_X1 cor_maj_163_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_163_n25)
         );
  OR2_X1 cor_maj_163_U5 ( .A1(cor_maj_163_n23), .A2(cor_maj_163_n22), .ZN(
        cor_maj_163_n32) );
  NAND2_X1 cor_maj_163_U4 ( .A1(cor_maj_163_n22), .A2(cor_maj_163_n23), .ZN(
        cor_maj_163_n34) );
  NAND2_X1 cor_maj_163_U3 ( .A1(cor_maj_163_n32), .A2(cor_maj_163_n31), .ZN(
        cor_maj_163_n33) );
  NAND2_X1 cor_maj_163_U2 ( .A1(cor_maj_163_n34), .A2(cor_maj_163_n33), .ZN(
        cor_maj_163_port_o) );
  OR2_X1 cor_maj_164_U19 ( .A1(cor_maj_164_n27), .A2(cor_maj_164_n26), .ZN(
        cor_maj_164_n28) );
  NAND2_X1 cor_maj_164_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_164_n28), .ZN(
        cor_maj_164_n29) );
  NAND2_X1 cor_maj_164_U17 ( .A1(cor_maj_164_n26), .A2(cor_maj_164_n27), .ZN(
        cor_maj_164_n30) );
  NAND2_X1 cor_maj_164_U16 ( .A1(cor_maj_164_n30), .A2(cor_maj_164_n29), .ZN(
        cor_maj_164_n31) );
  NAND2_X1 cor_maj_164_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_164_n25), .ZN(
        cor_maj_164_n18) );
  NAND2_X1 cor_maj_164_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_164_n19) );
  NAND2_X1 cor_maj_164_U13 ( .A1(cor_maj_164_n19), .A2(cor_maj_164_n18), .ZN(
        cor_maj_164_n22) );
  NAND2_X1 cor_maj_164_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_164_n24), .ZN(
        cor_maj_164_n20) );
  NAND2_X1 cor_maj_164_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_164_n21) );
  NAND2_X1 cor_maj_164_U10 ( .A1(cor_maj_164_n21), .A2(cor_maj_164_n20), .ZN(
        cor_maj_164_n23) );
  XOR2_X1 cor_maj_164_U9 ( .A(v_1_3_2[2]), .B(cor_maj_164_n24), .Z(
        cor_maj_164_n26) );
  XOR2_X1 cor_maj_164_U8 ( .A(v_1_3_2[5]), .B(cor_maj_164_n25), .Z(
        cor_maj_164_n27) );
  XOR2_X1 cor_maj_164_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_164_n24)
         );
  XOR2_X1 cor_maj_164_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_164_n25)
         );
  OR2_X1 cor_maj_164_U5 ( .A1(cor_maj_164_n23), .A2(cor_maj_164_n22), .ZN(
        cor_maj_164_n32) );
  NAND2_X1 cor_maj_164_U4 ( .A1(cor_maj_164_n22), .A2(cor_maj_164_n23), .ZN(
        cor_maj_164_n34) );
  NAND2_X1 cor_maj_164_U3 ( .A1(cor_maj_164_n32), .A2(cor_maj_164_n31), .ZN(
        cor_maj_164_n33) );
  NAND2_X1 cor_maj_164_U2 ( .A1(cor_maj_164_n34), .A2(cor_maj_164_n33), .ZN(
        cor_maj_164_port_o) );
  OR2_X1 cor_maj_165_U19 ( .A1(cor_maj_165_n27), .A2(cor_maj_165_n26), .ZN(
        cor_maj_165_n28) );
  NAND2_X1 cor_maj_165_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_165_n28), .ZN(
        cor_maj_165_n29) );
  NAND2_X1 cor_maj_165_U17 ( .A1(cor_maj_165_n26), .A2(cor_maj_165_n27), .ZN(
        cor_maj_165_n30) );
  NAND2_X1 cor_maj_165_U16 ( .A1(cor_maj_165_n30), .A2(cor_maj_165_n29), .ZN(
        cor_maj_165_n31) );
  NAND2_X1 cor_maj_165_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_165_n25), .ZN(
        cor_maj_165_n18) );
  NAND2_X1 cor_maj_165_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_165_n19) );
  NAND2_X1 cor_maj_165_U13 ( .A1(cor_maj_165_n19), .A2(cor_maj_165_n18), .ZN(
        cor_maj_165_n22) );
  NAND2_X1 cor_maj_165_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_165_n24), .ZN(
        cor_maj_165_n20) );
  NAND2_X1 cor_maj_165_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_165_n21) );
  NAND2_X1 cor_maj_165_U10 ( .A1(cor_maj_165_n21), .A2(cor_maj_165_n20), .ZN(
        cor_maj_165_n23) );
  XOR2_X1 cor_maj_165_U9 ( .A(v_1_3_2[2]), .B(cor_maj_165_n24), .Z(
        cor_maj_165_n26) );
  XOR2_X1 cor_maj_165_U8 ( .A(v_1_3_2[5]), .B(cor_maj_165_n25), .Z(
        cor_maj_165_n27) );
  XOR2_X1 cor_maj_165_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_165_n24)
         );
  XOR2_X1 cor_maj_165_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_165_n25)
         );
  OR2_X1 cor_maj_165_U5 ( .A1(cor_maj_165_n23), .A2(cor_maj_165_n22), .ZN(
        cor_maj_165_n32) );
  NAND2_X1 cor_maj_165_U4 ( .A1(cor_maj_165_n22), .A2(cor_maj_165_n23), .ZN(
        cor_maj_165_n34) );
  NAND2_X1 cor_maj_165_U3 ( .A1(cor_maj_165_n32), .A2(cor_maj_165_n31), .ZN(
        cor_maj_165_n33) );
  NAND2_X1 cor_maj_165_U2 ( .A1(cor_maj_165_n34), .A2(cor_maj_165_n33), .ZN(
        cor_maj_165_port_o) );
  OR2_X1 cor_maj_166_U19 ( .A1(cor_maj_166_n27), .A2(cor_maj_166_n26), .ZN(
        cor_maj_166_n28) );
  NAND2_X1 cor_maj_166_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_166_n28), .ZN(
        cor_maj_166_n29) );
  NAND2_X1 cor_maj_166_U17 ( .A1(cor_maj_166_n26), .A2(cor_maj_166_n27), .ZN(
        cor_maj_166_n30) );
  NAND2_X1 cor_maj_166_U16 ( .A1(cor_maj_166_n30), .A2(cor_maj_166_n29), .ZN(
        cor_maj_166_n31) );
  NAND2_X1 cor_maj_166_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_166_n25), .ZN(
        cor_maj_166_n18) );
  NAND2_X1 cor_maj_166_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_166_n19) );
  NAND2_X1 cor_maj_166_U13 ( .A1(cor_maj_166_n19), .A2(cor_maj_166_n18), .ZN(
        cor_maj_166_n22) );
  NAND2_X1 cor_maj_166_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_166_n24), .ZN(
        cor_maj_166_n20) );
  NAND2_X1 cor_maj_166_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_166_n21) );
  NAND2_X1 cor_maj_166_U10 ( .A1(cor_maj_166_n21), .A2(cor_maj_166_n20), .ZN(
        cor_maj_166_n23) );
  XOR2_X1 cor_maj_166_U9 ( .A(v_1_3_2[2]), .B(cor_maj_166_n24), .Z(
        cor_maj_166_n26) );
  XOR2_X1 cor_maj_166_U8 ( .A(v_1_3_2[5]), .B(cor_maj_166_n25), .Z(
        cor_maj_166_n27) );
  XOR2_X1 cor_maj_166_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_166_n24)
         );
  XOR2_X1 cor_maj_166_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_166_n25)
         );
  OR2_X1 cor_maj_166_U5 ( .A1(cor_maj_166_n23), .A2(cor_maj_166_n22), .ZN(
        cor_maj_166_n32) );
  NAND2_X1 cor_maj_166_U4 ( .A1(cor_maj_166_n22), .A2(cor_maj_166_n23), .ZN(
        cor_maj_166_n34) );
  NAND2_X1 cor_maj_166_U3 ( .A1(cor_maj_166_n32), .A2(cor_maj_166_n31), .ZN(
        cor_maj_166_n33) );
  NAND2_X1 cor_maj_166_U2 ( .A1(cor_maj_166_n34), .A2(cor_maj_166_n33), .ZN(
        cor_maj_166_port_o) );
  OR2_X1 cor_maj_167_U19 ( .A1(cor_maj_167_n27), .A2(cor_maj_167_n26), .ZN(
        cor_maj_167_n28) );
  NAND2_X1 cor_maj_167_U18 ( .A1(v_1_3_2[6]), .A2(cor_maj_167_n28), .ZN(
        cor_maj_167_n29) );
  NAND2_X1 cor_maj_167_U17 ( .A1(cor_maj_167_n26), .A2(cor_maj_167_n27), .ZN(
        cor_maj_167_n30) );
  NAND2_X1 cor_maj_167_U16 ( .A1(cor_maj_167_n30), .A2(cor_maj_167_n29), .ZN(
        cor_maj_167_n31) );
  NAND2_X1 cor_maj_167_U15 ( .A1(v_1_3_2[5]), .A2(cor_maj_167_n25), .ZN(
        cor_maj_167_n18) );
  NAND2_X1 cor_maj_167_U14 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_167_n19) );
  NAND2_X1 cor_maj_167_U13 ( .A1(cor_maj_167_n19), .A2(cor_maj_167_n18), .ZN(
        cor_maj_167_n22) );
  NAND2_X1 cor_maj_167_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_167_n24), .ZN(
        cor_maj_167_n20) );
  NAND2_X1 cor_maj_167_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_167_n21) );
  NAND2_X1 cor_maj_167_U10 ( .A1(cor_maj_167_n21), .A2(cor_maj_167_n20), .ZN(
        cor_maj_167_n23) );
  XOR2_X1 cor_maj_167_U9 ( .A(v_1_3_2[2]), .B(cor_maj_167_n24), .Z(
        cor_maj_167_n26) );
  XOR2_X1 cor_maj_167_U8 ( .A(v_1_3_2[5]), .B(cor_maj_167_n25), .Z(
        cor_maj_167_n27) );
  XOR2_X1 cor_maj_167_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_167_n24)
         );
  XOR2_X1 cor_maj_167_U6 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_167_n25)
         );
  OR2_X1 cor_maj_167_U5 ( .A1(cor_maj_167_n23), .A2(cor_maj_167_n22), .ZN(
        cor_maj_167_n32) );
  NAND2_X1 cor_maj_167_U4 ( .A1(cor_maj_167_n22), .A2(cor_maj_167_n23), .ZN(
        cor_maj_167_n34) );
  NAND2_X1 cor_maj_167_U3 ( .A1(cor_maj_167_n32), .A2(cor_maj_167_n31), .ZN(
        cor_maj_167_n33) );
  NAND2_X1 cor_maj_167_U2 ( .A1(cor_maj_167_n34), .A2(cor_maj_167_n33), .ZN(
        cor_maj_167_port_o) );
  XOR2_X1 simpleXor_84_U1 ( .A(n_zz_io_c_0_4[1]), .B(u_0_1[0]), .Z(
        simpleXor_84_port_z) );
  XOR2_X1 simpleXor_85_U1 ( .A(n_zz_io_c_0_4[2]), .B(u_0_2[0]), .Z(
        simpleXor_85_port_z) );
  XOR2_X1 simpleXor_86_U1 ( .A(n_zz_io_c_0_4[3]), .B(u_0_3[0]), .Z(
        simpleXor_86_port_z) );
  XOR2_X1 simpleXor_87_U1 ( .A(n_zz_io_c_1_4[1]), .B(u_1_0[0]), .Z(
        simpleXor_87_port_z) );
  XOR2_X1 simpleXor_88_U1 ( .A(n_zz_io_c_1_4[2]), .B(u_1_2[0]), .Z(
        simpleXor_88_port_z) );
  XOR2_X1 simpleXor_89_U1 ( .A(n_zz_io_c_1_4[3]), .B(u_1_3[0]), .Z(
        simpleXor_89_port_z) );
  XOR2_X1 simpleXor_90_U1 ( .A(n_zz_io_c_2_4[1]), .B(u_2_0[0]), .Z(
        simpleXor_90_port_z) );
  XOR2_X1 simpleXor_91_U1 ( .A(n_zz_io_c_2_4[2]), .B(u_2_1[0]), .Z(
        simpleXor_91_port_z) );
  XOR2_X1 simpleXor_92_U1 ( .A(n_zz_io_c_2_4[3]), .B(u_2_3[0]), .Z(
        simpleXor_92_port_z) );
  XOR2_X1 simpleXor_93_U1 ( .A(n_zz_io_c_3_4[1]), .B(u_3_0[0]), .Z(
        simpleXor_93_port_z) );
  XOR2_X1 simpleXor_94_U1 ( .A(n_zz_io_c_3_4[2]), .B(u_3_1[0]), .Z(
        simpleXor_94_port_z) );
  XOR2_X1 simpleXor_95_U1 ( .A(n_zz_io_c_3_4[3]), .B(u_3_2[0]), .Z(
        simpleXor_95_port_z) );
  XOR2_X1 simpleXor_96_U1 ( .A(n_zz_io_c_0_9[1]), .B(u_0_1[1]), .Z(
        simpleXor_96_port_z) );
  XOR2_X1 simpleXor_97_U1 ( .A(n_zz_io_c_0_9[2]), .B(u_0_2[1]), .Z(
        simpleXor_97_port_z) );
  XOR2_X1 simpleXor_98_U1 ( .A(n_zz_io_c_0_9[3]), .B(u_0_3[1]), .Z(
        simpleXor_98_port_z) );
  XOR2_X1 simpleXor_99_U1 ( .A(n_zz_io_c_1_9[1]), .B(u_1_0[1]), .Z(
        simpleXor_99_port_z) );
  XOR2_X1 simpleXor_100_U1 ( .A(n_zz_io_c_1_9[2]), .B(u_1_2[1]), .Z(
        simpleXor_100_port_z) );
  XOR2_X1 simpleXor_101_U1 ( .A(n_zz_io_c_1_9[3]), .B(u_1_3[1]), .Z(
        simpleXor_101_port_z) );
  XOR2_X1 simpleXor_102_U1 ( .A(n_zz_io_c_2_9[1]), .B(u_2_0[1]), .Z(
        simpleXor_102_port_z) );
  XOR2_X1 simpleXor_103_U1 ( .A(n_zz_io_c_2_9[2]), .B(u_2_1[1]), .Z(
        simpleXor_103_port_z) );
  XOR2_X1 simpleXor_104_U1 ( .A(n_zz_io_c_2_9[3]), .B(u_2_3[1]), .Z(
        simpleXor_104_port_z) );
  XOR2_X1 simpleXor_105_U1 ( .A(n_zz_io_c_3_9[1]), .B(u_3_0[1]), .Z(
        simpleXor_105_port_z) );
  XOR2_X1 simpleXor_106_U1 ( .A(n_zz_io_c_3_9[2]), .B(u_3_1[1]), .Z(
        simpleXor_106_port_z) );
  XOR2_X1 simpleXor_107_U1 ( .A(n_zz_io_c_3_9[3]), .B(u_3_2[1]), .Z(
        simpleXor_107_port_z) );
  XOR2_X1 simpleXor_108_U1 ( .A(n_zz_io_c_0_14[1]), .B(u_0_1[2]), .Z(
        simpleXor_108_port_z) );
  XOR2_X1 simpleXor_109_U1 ( .A(n_zz_io_c_0_14[2]), .B(u_0_2[2]), .Z(
        simpleXor_109_port_z) );
  XOR2_X1 simpleXor_110_U1 ( .A(n_zz_io_c_0_14[3]), .B(u_0_3[2]), .Z(
        simpleXor_110_port_z) );
  XOR2_X1 simpleXor_111_U1 ( .A(n_zz_io_c_1_14[1]), .B(u_1_0[2]), .Z(
        simpleXor_111_port_z) );
  XOR2_X1 simpleXor_112_U1 ( .A(n_zz_io_c_1_14[2]), .B(u_1_2[2]), .Z(
        simpleXor_112_port_z) );
  XOR2_X1 simpleXor_113_U1 ( .A(n_zz_io_c_1_14[3]), .B(u_1_3[2]), .Z(
        simpleXor_113_port_z) );
  XOR2_X1 simpleXor_114_U1 ( .A(n_zz_io_c_2_14[1]), .B(u_2_0[2]), .Z(
        simpleXor_114_port_z) );
  XOR2_X1 simpleXor_115_U1 ( .A(n_zz_io_c_2_14[2]), .B(u_2_1[2]), .Z(
        simpleXor_115_port_z) );
  XOR2_X1 simpleXor_116_U1 ( .A(n_zz_io_c_2_14[3]), .B(u_2_3[2]), .Z(
        simpleXor_116_port_z) );
  XOR2_X1 simpleXor_117_U1 ( .A(n_zz_io_c_3_14[1]), .B(u_3_0[2]), .Z(
        simpleXor_117_port_z) );
  XOR2_X1 simpleXor_118_U1 ( .A(n_zz_io_c_3_14[2]), .B(u_3_1[2]), .Z(
        simpleXor_118_port_z) );
  XOR2_X1 simpleXor_119_U1 ( .A(n_zz_io_c_3_14[3]), .B(u_3_2[2]), .Z(
        simpleXor_119_port_z) );
  XOR2_X1 simpleXor_120_U1 ( .A(n_zz_io_c_0_19[1]), .B(u_0_1[3]), .Z(
        simpleXor_120_port_z) );
  XOR2_X1 simpleXor_121_U1 ( .A(n_zz_io_c_0_19[2]), .B(u_0_2[3]), .Z(
        simpleXor_121_port_z) );
  XOR2_X1 simpleXor_122_U1 ( .A(n_zz_io_c_0_19[3]), .B(u_0_3[3]), .Z(
        simpleXor_122_port_z) );
  XOR2_X1 simpleXor_123_U1 ( .A(n_zz_io_c_1_19[1]), .B(u_1_0[3]), .Z(
        simpleXor_123_port_z) );
  XOR2_X1 simpleXor_124_U1 ( .A(n_zz_io_c_1_19[2]), .B(u_1_2[3]), .Z(
        simpleXor_124_port_z) );
  XOR2_X1 simpleXor_125_U1 ( .A(n_zz_io_c_1_19[3]), .B(u_1_3[3]), .Z(
        simpleXor_125_port_z) );
  XOR2_X1 simpleXor_126_U1 ( .A(n_zz_io_c_2_19[1]), .B(u_2_0[3]), .Z(
        simpleXor_126_port_z) );
  XOR2_X1 simpleXor_127_U1 ( .A(n_zz_io_c_2_19[2]), .B(u_2_1[3]), .Z(
        simpleXor_127_port_z) );
  XOR2_X1 simpleXor_128_U1 ( .A(n_zz_io_c_2_19[3]), .B(u_2_3[3]), .Z(
        simpleXor_128_port_z) );
  XOR2_X1 simpleXor_129_U1 ( .A(n_zz_io_c_3_19[1]), .B(u_3_0[3]), .Z(
        simpleXor_129_port_z) );
  XOR2_X1 simpleXor_130_U1 ( .A(n_zz_io_c_3_19[2]), .B(u_3_1[3]), .Z(
        simpleXor_130_port_z) );
  XOR2_X1 simpleXor_131_U1 ( .A(n_zz_io_c_3_19[3]), .B(u_3_2[3]), .Z(
        simpleXor_131_port_z) );
  XOR2_X1 simpleXor_132_U1 ( .A(n_zz_io_c_0_24[1]), .B(u_0_1[4]), .Z(
        simpleXor_132_port_z) );
  XOR2_X1 simpleXor_133_U1 ( .A(n_zz_io_c_0_24[2]), .B(u_0_2[4]), .Z(
        simpleXor_133_port_z) );
  XOR2_X1 simpleXor_134_U1 ( .A(n_zz_io_c_0_24[3]), .B(u_0_3[4]), .Z(
        simpleXor_134_port_z) );
  XOR2_X1 simpleXor_135_U1 ( .A(n_zz_io_c_1_24[1]), .B(u_1_0[4]), .Z(
        simpleXor_135_port_z) );
  XOR2_X1 simpleXor_136_U1 ( .A(n_zz_io_c_1_24[2]), .B(u_1_2[4]), .Z(
        simpleXor_136_port_z) );
  XOR2_X1 simpleXor_137_U1 ( .A(n_zz_io_c_1_24[3]), .B(u_1_3[4]), .Z(
        simpleXor_137_port_z) );
  XOR2_X1 simpleXor_138_U1 ( .A(n_zz_io_c_2_24[1]), .B(u_2_0[4]), .Z(
        simpleXor_138_port_z) );
  XOR2_X1 simpleXor_139_U1 ( .A(n_zz_io_c_2_24[2]), .B(u_2_1[4]), .Z(
        simpleXor_139_port_z) );
  XOR2_X1 simpleXor_140_U1 ( .A(n_zz_io_c_2_24[3]), .B(u_2_3[4]), .Z(
        simpleXor_140_port_z) );
  XOR2_X1 simpleXor_141_U1 ( .A(n_zz_io_c_3_24[1]), .B(u_3_0[4]), .Z(
        simpleXor_141_port_z) );
  XOR2_X1 simpleXor_142_U1 ( .A(n_zz_io_c_3_24[2]), .B(u_3_1[4]), .Z(
        simpleXor_142_port_z) );
  XOR2_X1 simpleXor_143_U1 ( .A(n_zz_io_c_3_24[3]), .B(u_3_2[4]), .Z(
        simpleXor_143_port_z) );
  XOR2_X1 simpleXor_144_U1 ( .A(n_zz_io_c_0_29[1]), .B(u_0_1[5]), .Z(
        simpleXor_144_port_z) );
  XOR2_X1 simpleXor_145_U1 ( .A(n_zz_io_c_0_29[2]), .B(u_0_2[5]), .Z(
        simpleXor_145_port_z) );
  XOR2_X1 simpleXor_146_U1 ( .A(n_zz_io_c_0_29[3]), .B(u_0_3[5]), .Z(
        simpleXor_146_port_z) );
  XOR2_X1 simpleXor_147_U1 ( .A(n_zz_io_c_1_29[1]), .B(u_1_0[5]), .Z(
        simpleXor_147_port_z) );
  XOR2_X1 simpleXor_148_U1 ( .A(n_zz_io_c_1_29[2]), .B(u_1_2[5]), .Z(
        simpleXor_148_port_z) );
  XOR2_X1 simpleXor_149_U1 ( .A(n_zz_io_c_1_29[3]), .B(u_1_3[5]), .Z(
        simpleXor_149_port_z) );
  XOR2_X1 simpleXor_150_U1 ( .A(n_zz_io_c_2_29[1]), .B(u_2_0[5]), .Z(
        simpleXor_150_port_z) );
  XOR2_X1 simpleXor_151_U1 ( .A(n_zz_io_c_2_29[2]), .B(u_2_1[5]), .Z(
        simpleXor_151_port_z) );
  XOR2_X1 simpleXor_152_U1 ( .A(n_zz_io_c_2_29[3]), .B(u_2_3[5]), .Z(
        simpleXor_152_port_z) );
  XOR2_X1 simpleXor_153_U1 ( .A(n_zz_io_c_3_29[1]), .B(u_3_0[5]), .Z(
        simpleXor_153_port_z) );
  XOR2_X1 simpleXor_154_U1 ( .A(n_zz_io_c_3_29[2]), .B(u_3_1[5]), .Z(
        simpleXor_154_port_z) );
  XOR2_X1 simpleXor_155_U1 ( .A(n_zz_io_c_3_29[3]), .B(u_3_2[5]), .Z(
        simpleXor_155_port_z) );
  XOR2_X1 simpleXor_156_U1 ( .A(n_zz_io_c_0_34[1]), .B(u_0_1[6]), .Z(
        simpleXor_156_port_z) );
  XOR2_X1 simpleXor_157_U1 ( .A(n_zz_io_c_0_34[2]), .B(u_0_2[6]), .Z(
        simpleXor_157_port_z) );
  XOR2_X1 simpleXor_158_U1 ( .A(n_zz_io_c_0_34[3]), .B(u_0_3[6]), .Z(
        simpleXor_158_port_z) );
  XOR2_X1 simpleXor_159_U1 ( .A(n_zz_io_c_1_34[1]), .B(u_1_0[6]), .Z(
        simpleXor_159_port_z) );
  XOR2_X1 simpleXor_160_U1 ( .A(n_zz_io_c_1_34[2]), .B(u_1_2[6]), .Z(
        simpleXor_160_port_z) );
  XOR2_X1 simpleXor_161_U1 ( .A(n_zz_io_c_1_34[3]), .B(u_1_3[6]), .Z(
        simpleXor_161_port_z) );
  XOR2_X1 simpleXor_162_U1 ( .A(n_zz_io_c_2_34[1]), .B(u_2_0[6]), .Z(
        simpleXor_162_port_z) );
  XOR2_X1 simpleXor_163_U1 ( .A(n_zz_io_c_2_34[2]), .B(u_2_1[6]), .Z(
        simpleXor_163_port_z) );
  XOR2_X1 simpleXor_164_U1 ( .A(n_zz_io_c_2_34[3]), .B(u_2_3[6]), .Z(
        simpleXor_164_port_z) );
  XOR2_X1 simpleXor_165_U1 ( .A(n_zz_io_c_3_34[1]), .B(u_3_0[6]), .Z(
        simpleXor_165_port_z) );
  XOR2_X1 simpleXor_166_U1 ( .A(n_zz_io_c_3_34[2]), .B(u_3_1[6]), .Z(
        simpleXor_166_port_z) );
  XOR2_X1 simpleXor_167_U1 ( .A(n_zz_io_c_3_34[3]), .B(u_3_2[6]), .Z(
        simpleXor_167_port_z) );
endmodule

