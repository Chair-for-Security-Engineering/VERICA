
module ISW_SifaTest ( port_a_in, port_b_in, port_rand, port_det_out, clk, 
        reset );
  input [1:0] port_a_in;
  input [1:0] port_b_in;
  input [0:0] port_rand;
  output [1:0] port_det_out;
  input clk, reset;
  wire   isw_0_n5, isw_0_n4, isw_0_n3, isw_0_n2, isw_0_n1, isw_0_N6, isw_0_z_0,
         isw_0__zz_result_1_1, isw_0_N5, isw_0__zz_result_0_3,
         isw_0__zz_result_0_1, isw_0__zz_result_1, isw_0_N4,
         isw_0__zz_result_0_2, isw_0__zz_result_0, isw_0_N3, isw_0_N2,
         isw_0__zz_z_0_1, isw_0__zz_z_0, isw_0_N1, isw_0_N0, isw_1_n10,
         isw_1_n9, isw_1_n8, isw_1_n7, isw_1_n6, isw_1_N6, isw_1_z_0,
         isw_1__zz_result_1_1, isw_1_N5, isw_1__zz_result_0_3,
         isw_1__zz_result_0_1, isw_1__zz_result_1, isw_1_N4,
         isw_1__zz_result_0_2, isw_1__zz_result_0, isw_1_N3, isw_1_N2,
         isw_1__zz_z_0_1, isw_1__zz_z_0, isw_1_N1, isw_1_N0;
  wire   [1:0] n_zz_unequal_0;
  wire   [1:0] n_zz_unequal_0_1;

  XNOR2_X1 U3 ( .A(n_zz_unequal_0_1[0]), .B(n_zz_unequal_0[0]), .ZN(
        port_det_out[0]) );
  XNOR2_X1 U4 ( .A(n_zz_unequal_0_1[1]), .B(n_zz_unequal_0[1]), .ZN(
        port_det_out[1]) );
  INV_X1 isw_0_U14 ( .A(port_a_in[1]), .ZN(isw_0_n2) );
  INV_X1 isw_0_U13 ( .A(port_b_in[1]), .ZN(isw_0_n4) );
  INV_X1 isw_0_U12 ( .A(port_a_in[0]), .ZN(isw_0_n1) );
  INV_X1 isw_0_U11 ( .A(port_b_in[0]), .ZN(isw_0_n3) );
  NOR2_X1 isw_0_U10 ( .A1(isw_0_n4), .A2(isw_0_n1), .ZN(isw_0_n5) );
  XOR2_X1 isw_0_U9 ( .A(port_rand[0]), .B(isw_0_n5), .Z(isw_0_N0) );
  XOR2_X1 isw_0_U8 ( .A(isw_0__zz_z_0_1), .B(isw_0__zz_z_0), .Z(isw_0_N2) );
  XOR2_X1 isw_0_U7 ( .A(isw_0__zz_result_0_3), .B(isw_0__zz_result_0_1), .Z(
        isw_0_N5) );
  XOR2_X1 isw_0_U6 ( .A(isw_0_z_0), .B(isw_0__zz_result_1_1), .Z(isw_0_N6) );
  NOR2_X1 isw_0_U5 ( .A1(isw_0_n2), .A2(isw_0_n4), .ZN(isw_0_N4) );
  NOR2_X1 isw_0_U4 ( .A1(isw_0_n1), .A2(isw_0_n3), .ZN(isw_0_N3) );
  NOR2_X1 isw_0_U3 ( .A1(isw_0_n2), .A2(isw_0_n3), .ZN(isw_0_N1) );
  DFF_X1 isw_0_result_1_reg ( .D(isw_0_N6), .CK(clk), .Q(n_zz_unequal_0[1]), 
        .QN() );
  DFF_X1 isw_0_result_0_reg ( .D(isw_0_N5), .CK(clk), .Q(n_zz_unequal_0[0]), 
        .QN() );
  DFF_X1 isw_0__zz_result_0_3_reg ( .D(isw_0__zz_result_0_2), .CK(clk), .Q(
        isw_0__zz_result_0_3), .QN() );
  DFF_X1 isw_0__zz_result_0_2_reg ( .D(port_rand[0]), .CK(clk), .Q(
        isw_0__zz_result_0_2), .QN() );
  DFF_X1 isw_0__zz_result_1_1_reg ( .D(isw_0__zz_result_1), .CK(clk), .Q(
        isw_0__zz_result_1_1), .QN() );
  DFF_X1 isw_0__zz_result_1_reg ( .D(isw_0_N4), .CK(clk), .Q(
        isw_0__zz_result_1), .QN() );
  DFF_X1 isw_0_z_0_reg ( .D(isw_0_N2), .CK(clk), .Q(isw_0_z_0), .QN() );
  DFF_X1 isw_0__zz_z_0_reg ( .D(isw_0_N0), .CK(clk), .Q(isw_0__zz_z_0), .QN()
         );
  DFF_X1 isw_0__zz_result_0_1_reg ( .D(isw_0__zz_result_0), .CK(clk), .Q(
        isw_0__zz_result_0_1), .QN() );
  DFF_X1 isw_0__zz_z_0_1_reg ( .D(isw_0_N1), .CK(clk), .Q(isw_0__zz_z_0_1), 
        .QN() );
  DFF_X1 isw_0__zz_result_0_reg ( .D(isw_0_N3), .CK(clk), .Q(
        isw_0__zz_result_0), .QN() );
  INV_X1 isw_1_U14 ( .A(port_a_in[1]), .ZN(isw_1_n9) );
  INV_X1 isw_1_U13 ( .A(port_b_in[1]), .ZN(isw_1_n7) );
  INV_X1 isw_1_U12 ( .A(port_a_in[0]), .ZN(isw_1_n10) );
  INV_X1 isw_1_U11 ( .A(port_b_in[0]), .ZN(isw_1_n8) );
  NOR2_X1 isw_1_U10 ( .A1(isw_1_n7), .A2(isw_1_n10), .ZN(isw_1_n6) );
  XOR2_X1 isw_1_U9 ( .A(port_rand[0]), .B(isw_1_n6), .Z(isw_1_N0) );
  XOR2_X1 isw_1_U8 ( .A(isw_1__zz_z_0_1), .B(isw_1__zz_z_0), .Z(isw_1_N2) );
  XOR2_X1 isw_1_U7 ( .A(isw_1__zz_result_0_3), .B(isw_1__zz_result_0_1), .Z(
        isw_1_N5) );
  XOR2_X1 isw_1_U6 ( .A(isw_1_z_0), .B(isw_1__zz_result_1_1), .Z(isw_1_N6) );
  NOR2_X1 isw_1_U5 ( .A1(isw_1_n9), .A2(isw_1_n7), .ZN(isw_1_N4) );
  NOR2_X1 isw_1_U4 ( .A1(isw_1_n10), .A2(isw_1_n8), .ZN(isw_1_N3) );
  NOR2_X1 isw_1_U3 ( .A1(isw_1_n9), .A2(isw_1_n8), .ZN(isw_1_N1) );
  DFF_X1 isw_1_result_1_reg ( .D(isw_1_N6), .CK(clk), .Q(n_zz_unequal_0_1[1]), 
        .QN() );
  DFF_X1 isw_1_result_0_reg ( .D(isw_1_N5), .CK(clk), .Q(n_zz_unequal_0_1[0]), 
        .QN() );
  DFF_X1 isw_1__zz_result_0_3_reg ( .D(isw_1__zz_result_0_2), .CK(clk), .Q(
        isw_1__zz_result_0_3), .QN() );
  DFF_X1 isw_1__zz_result_0_2_reg ( .D(port_rand[0]), .CK(clk), .Q(
        isw_1__zz_result_0_2), .QN() );
  DFF_X1 isw_1__zz_result_1_1_reg ( .D(isw_1__zz_result_1), .CK(clk), .Q(
        isw_1__zz_result_1_1), .QN() );
  DFF_X1 isw_1__zz_result_1_reg ( .D(isw_1_N4), .CK(clk), .Q(
        isw_1__zz_result_1), .QN() );
  DFF_X1 isw_1_z_0_reg ( .D(isw_1_N2), .CK(clk), .Q(isw_1_z_0), .QN() );
  DFF_X1 isw_1__zz_z_0_reg ( .D(isw_1_N0), .CK(clk), .Q(isw_1__zz_z_0), .QN()
         );
  DFF_X1 isw_1__zz_result_0_1_reg ( .D(isw_1__zz_result_0), .CK(clk), .Q(
        isw_1__zz_result_0_1), .QN() );
  DFF_X1 isw_1__zz_z_0_1_reg ( .D(isw_1_N1), .CK(clk), .Q(isw_1__zz_z_0_1), 
        .QN() );
  DFF_X1 isw_1__zz_result_0_reg ( .D(isw_1_N3), .CK(clk), .Q(
        isw_1__zz_result_0), .QN() );
endmodule

