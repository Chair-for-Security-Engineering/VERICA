
module CINI ( io_a_0, io_a_1, io_a_2, io_b_0, io_b_1, io_b_2, io_c_0, io_c_1, 
        io_c_2, io_rand, clk, reset );
  input [6:0] io_a_0;
  input [6:0] io_a_1;
  input [6:0] io_a_2;
  input [6:0] io_b_0;
  input [6:0] io_b_1;
  input [6:0] io_b_2;
  output [6:0] io_c_0;
  output [6:0] io_c_1;
  output [6:0] io_c_2;
  input [2:0] io_rand;
  input clk, reset;
  wire   simpleNot_42_port_z, simpleNot_43_port_z, simpleNot_44_port_z,
         simpleNot_45_port_z, simpleNot_46_port_z, simpleNot_47_port_z,
         simpleNot_48_port_z, simpleNot_49_port_z, simpleNot_50_port_z,
         simpleNot_51_port_z, simpleNot_52_port_z, simpleNot_53_port_z,
         simpleNot_54_port_z, simpleNot_55_port_z, simpleNot_56_port_z,
         simpleNot_57_port_z, simpleNot_58_port_z, simpleNot_59_port_z,
         simpleNot_60_port_z, simpleNot_61_port_z, simpleNot_62_port_z,
         simpleNot_63_port_z, simpleNot_64_port_z, simpleNot_65_port_z,
         simpleNot_66_port_z, simpleNot_67_port_z, simpleNot_68_port_z,
         simpleNot_69_port_z, simpleNot_70_port_z, simpleNot_71_port_z,
         simpleNot_72_port_z, simpleNot_73_port_z, simpleNot_74_port_z,
         simpleNot_75_port_z, simpleNot_76_port_z, simpleNot_77_port_z,
         simpleNot_78_port_z, simpleNot_79_port_z, simpleNot_80_port_z,
         simpleNot_81_port_z, simpleNot_82_port_z, simpleNot_83_port_z,
         simpleXor_42_port_z, simpleXor_43_port_z, simpleXor_44_port_z,
         simpleXor_45_port_z, simpleXor_46_port_z, simpleXor_47_port_z,
         simpleXor_48_port_z, simpleXor_49_port_z, simpleXor_50_port_z,
         simpleXor_51_port_z, simpleXor_52_port_z, simpleXor_53_port_z,
         simpleXor_54_port_z, simpleXor_55_port_z, simpleXor_56_port_z,
         simpleXor_57_port_z, simpleXor_58_port_z, simpleXor_59_port_z,
         simpleXor_60_port_z, simpleXor_61_port_z, simpleXor_62_port_z,
         simpleXor_63_port_z, simpleXor_64_port_z, simpleXor_65_port_z,
         simpleXor_66_port_z, simpleXor_67_port_z, simpleXor_68_port_z,
         simpleXor_69_port_z, simpleXor_70_port_z, simpleXor_71_port_z,
         simpleXor_72_port_z, simpleXor_73_port_z, simpleXor_74_port_z,
         simpleXor_75_port_z, simpleXor_76_port_z, simpleXor_77_port_z,
         simpleXor_78_port_z, simpleXor_79_port_z, simpleXor_80_port_z,
         simpleXor_81_port_z, simpleXor_82_port_z, simpleXor_83_port_z,
         n_zz_io_c_0_0_, n_zz_io_c_1_0_, n_zz_io_c_2_0_, n_zz_io_c_0_4_0_,
         n_zz_io_c_1_4_0_, n_zz_io_c_2_4_0_, n_zz_io_c_0_8_0_,
         n_zz_io_c_1_8_0_, n_zz_io_c_2_8_0_, n_zz_io_c_0_12_0_,
         n_zz_io_c_1_12_0_, n_zz_io_c_2_12_0_, n_zz_io_c_0_16_0_,
         n_zz_io_c_1_16_0_, n_zz_io_c_2_16_0_, n_zz_io_c_0_20_0_,
         n_zz_io_c_1_20_0_, n_zz_io_c_2_20_0_, n_zz_io_c_0_24_0_,
         n_zz_io_c_1_24_0_, n_zz_io_c_2_24_0_, N0, N1, N2, N3, N4, N5, N6, N7,
         N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, cor_maj_83_port_o, cor_maj_82_port_o,
         cor_maj_81_port_o, cor_maj_80_port_o, cor_maj_79_port_o,
         cor_maj_78_port_o, cor_maj_77_port_o, cor_maj_76_port_o,
         cor_maj_75_port_o, cor_maj_74_port_o, cor_maj_73_port_o,
         cor_maj_72_port_o, cor_maj_71_port_o, cor_maj_70_port_o,
         cor_maj_69_port_o, cor_maj_68_port_o, cor_maj_67_port_o,
         cor_maj_66_port_o, cor_maj_65_port_o, cor_maj_64_port_o,
         cor_maj_63_port_o, cor_maj_62_port_o, cor_maj_61_port_o,
         cor_maj_60_port_o, cor_maj_59_port_o, cor_maj_58_port_o,
         cor_maj_57_port_o, cor_maj_56_port_o, cor_maj_55_port_o,
         cor_maj_54_port_o, cor_maj_53_port_o, cor_maj_52_port_o,
         cor_maj_51_port_o, cor_maj_50_port_o, cor_maj_49_port_o,
         cor_maj_48_port_o, cor_maj_47_port_o, cor_maj_46_port_o,
         cor_maj_45_port_o, cor_maj_44_port_o, cor_maj_43_port_o,
         cor_maj_42_port_o, cor_maj_42_n17, cor_maj_42_n16, cor_maj_42_n15,
         cor_maj_42_n14, cor_maj_42_n13, cor_maj_42_n12, cor_maj_42_n11,
         cor_maj_42_n10, cor_maj_42_n9, cor_maj_42_n8, cor_maj_42_n7,
         cor_maj_42_n6, cor_maj_42_n5, cor_maj_42_n4, cor_maj_42_n3,
         cor_maj_42_n2, cor_maj_42_n1, cor_maj_43_n34, cor_maj_43_n33,
         cor_maj_43_n32, cor_maj_43_n31, cor_maj_43_n30, cor_maj_43_n29,
         cor_maj_43_n28, cor_maj_43_n27, cor_maj_43_n26, cor_maj_43_n25,
         cor_maj_43_n24, cor_maj_43_n23, cor_maj_43_n22, cor_maj_43_n21,
         cor_maj_43_n20, cor_maj_43_n19, cor_maj_43_n18, cor_maj_44_n34,
         cor_maj_44_n33, cor_maj_44_n32, cor_maj_44_n31, cor_maj_44_n30,
         cor_maj_44_n29, cor_maj_44_n28, cor_maj_44_n27, cor_maj_44_n26,
         cor_maj_44_n25, cor_maj_44_n24, cor_maj_44_n23, cor_maj_44_n22,
         cor_maj_44_n21, cor_maj_44_n20, cor_maj_44_n19, cor_maj_44_n18,
         cor_maj_45_n34, cor_maj_45_n33, cor_maj_45_n32, cor_maj_45_n31,
         cor_maj_45_n30, cor_maj_45_n29, cor_maj_45_n28, cor_maj_45_n27,
         cor_maj_45_n26, cor_maj_45_n25, cor_maj_45_n24, cor_maj_45_n23,
         cor_maj_45_n22, cor_maj_45_n21, cor_maj_45_n20, cor_maj_45_n19,
         cor_maj_45_n18, cor_maj_46_n34, cor_maj_46_n33, cor_maj_46_n32,
         cor_maj_46_n31, cor_maj_46_n30, cor_maj_46_n29, cor_maj_46_n28,
         cor_maj_46_n27, cor_maj_46_n26, cor_maj_46_n25, cor_maj_46_n24,
         cor_maj_46_n23, cor_maj_46_n22, cor_maj_46_n21, cor_maj_46_n20,
         cor_maj_46_n19, cor_maj_46_n18, cor_maj_47_n34, cor_maj_47_n33,
         cor_maj_47_n32, cor_maj_47_n31, cor_maj_47_n30, cor_maj_47_n29,
         cor_maj_47_n28, cor_maj_47_n27, cor_maj_47_n26, cor_maj_47_n25,
         cor_maj_47_n24, cor_maj_47_n23, cor_maj_47_n22, cor_maj_47_n21,
         cor_maj_47_n20, cor_maj_47_n19, cor_maj_47_n18, cor_maj_48_n34,
         cor_maj_48_n33, cor_maj_48_n32, cor_maj_48_n31, cor_maj_48_n30,
         cor_maj_48_n29, cor_maj_48_n28, cor_maj_48_n27, cor_maj_48_n26,
         cor_maj_48_n25, cor_maj_48_n24, cor_maj_48_n23, cor_maj_48_n22,
         cor_maj_48_n21, cor_maj_48_n20, cor_maj_48_n19, cor_maj_48_n18,
         cor_maj_49_n34, cor_maj_49_n33, cor_maj_49_n32, cor_maj_49_n31,
         cor_maj_49_n30, cor_maj_49_n29, cor_maj_49_n28, cor_maj_49_n27,
         cor_maj_49_n26, cor_maj_49_n25, cor_maj_49_n24, cor_maj_49_n23,
         cor_maj_49_n22, cor_maj_49_n21, cor_maj_49_n20, cor_maj_49_n19,
         cor_maj_49_n18, cor_maj_50_n34, cor_maj_50_n33, cor_maj_50_n32,
         cor_maj_50_n31, cor_maj_50_n30, cor_maj_50_n29, cor_maj_50_n28,
         cor_maj_50_n27, cor_maj_50_n26, cor_maj_50_n25, cor_maj_50_n24,
         cor_maj_50_n23, cor_maj_50_n22, cor_maj_50_n21, cor_maj_50_n20,
         cor_maj_50_n19, cor_maj_50_n18, cor_maj_51_n34, cor_maj_51_n33,
         cor_maj_51_n32, cor_maj_51_n31, cor_maj_51_n30, cor_maj_51_n29,
         cor_maj_51_n28, cor_maj_51_n27, cor_maj_51_n26, cor_maj_51_n25,
         cor_maj_51_n24, cor_maj_51_n23, cor_maj_51_n22, cor_maj_51_n21,
         cor_maj_51_n20, cor_maj_51_n19, cor_maj_51_n18, cor_maj_52_n34,
         cor_maj_52_n33, cor_maj_52_n32, cor_maj_52_n31, cor_maj_52_n30,
         cor_maj_52_n29, cor_maj_52_n28, cor_maj_52_n27, cor_maj_52_n26,
         cor_maj_52_n25, cor_maj_52_n24, cor_maj_52_n23, cor_maj_52_n22,
         cor_maj_52_n21, cor_maj_52_n20, cor_maj_52_n19, cor_maj_52_n18,
         cor_maj_53_n34, cor_maj_53_n33, cor_maj_53_n32, cor_maj_53_n31,
         cor_maj_53_n30, cor_maj_53_n29, cor_maj_53_n28, cor_maj_53_n27,
         cor_maj_53_n26, cor_maj_53_n25, cor_maj_53_n24, cor_maj_53_n23,
         cor_maj_53_n22, cor_maj_53_n21, cor_maj_53_n20, cor_maj_53_n19,
         cor_maj_53_n18, cor_maj_54_n34, cor_maj_54_n33, cor_maj_54_n32,
         cor_maj_54_n31, cor_maj_54_n30, cor_maj_54_n29, cor_maj_54_n28,
         cor_maj_54_n27, cor_maj_54_n26, cor_maj_54_n25, cor_maj_54_n24,
         cor_maj_54_n23, cor_maj_54_n22, cor_maj_54_n21, cor_maj_54_n20,
         cor_maj_54_n19, cor_maj_54_n18, cor_maj_55_n34, cor_maj_55_n33,
         cor_maj_55_n32, cor_maj_55_n31, cor_maj_55_n30, cor_maj_55_n29,
         cor_maj_55_n28, cor_maj_55_n27, cor_maj_55_n26, cor_maj_55_n25,
         cor_maj_55_n24, cor_maj_55_n23, cor_maj_55_n22, cor_maj_55_n21,
         cor_maj_55_n20, cor_maj_55_n19, cor_maj_55_n18, cor_maj_56_n34,
         cor_maj_56_n33, cor_maj_56_n32, cor_maj_56_n31, cor_maj_56_n30,
         cor_maj_56_n29, cor_maj_56_n28, cor_maj_56_n27, cor_maj_56_n26,
         cor_maj_56_n25, cor_maj_56_n24, cor_maj_56_n23, cor_maj_56_n22,
         cor_maj_56_n21, cor_maj_56_n20, cor_maj_56_n19, cor_maj_56_n18,
         cor_maj_57_n34, cor_maj_57_n33, cor_maj_57_n32, cor_maj_57_n31,
         cor_maj_57_n30, cor_maj_57_n29, cor_maj_57_n28, cor_maj_57_n27,
         cor_maj_57_n26, cor_maj_57_n25, cor_maj_57_n24, cor_maj_57_n23,
         cor_maj_57_n22, cor_maj_57_n21, cor_maj_57_n20, cor_maj_57_n19,
         cor_maj_57_n18, cor_maj_58_n34, cor_maj_58_n33, cor_maj_58_n32,
         cor_maj_58_n31, cor_maj_58_n30, cor_maj_58_n29, cor_maj_58_n28,
         cor_maj_58_n27, cor_maj_58_n26, cor_maj_58_n25, cor_maj_58_n24,
         cor_maj_58_n23, cor_maj_58_n22, cor_maj_58_n21, cor_maj_58_n20,
         cor_maj_58_n19, cor_maj_58_n18, cor_maj_59_n34, cor_maj_59_n33,
         cor_maj_59_n32, cor_maj_59_n31, cor_maj_59_n30, cor_maj_59_n29,
         cor_maj_59_n28, cor_maj_59_n27, cor_maj_59_n26, cor_maj_59_n25,
         cor_maj_59_n24, cor_maj_59_n23, cor_maj_59_n22, cor_maj_59_n21,
         cor_maj_59_n20, cor_maj_59_n19, cor_maj_59_n18, cor_maj_60_n34,
         cor_maj_60_n33, cor_maj_60_n32, cor_maj_60_n31, cor_maj_60_n30,
         cor_maj_60_n29, cor_maj_60_n28, cor_maj_60_n27, cor_maj_60_n26,
         cor_maj_60_n25, cor_maj_60_n24, cor_maj_60_n23, cor_maj_60_n22,
         cor_maj_60_n21, cor_maj_60_n20, cor_maj_60_n19, cor_maj_60_n18,
         cor_maj_61_n34, cor_maj_61_n33, cor_maj_61_n32, cor_maj_61_n31,
         cor_maj_61_n30, cor_maj_61_n29, cor_maj_61_n28, cor_maj_61_n27,
         cor_maj_61_n26, cor_maj_61_n25, cor_maj_61_n24, cor_maj_61_n23,
         cor_maj_61_n22, cor_maj_61_n21, cor_maj_61_n20, cor_maj_61_n19,
         cor_maj_61_n18, cor_maj_62_n34, cor_maj_62_n33, cor_maj_62_n32,
         cor_maj_62_n31, cor_maj_62_n30, cor_maj_62_n29, cor_maj_62_n28,
         cor_maj_62_n27, cor_maj_62_n26, cor_maj_62_n25, cor_maj_62_n24,
         cor_maj_62_n23, cor_maj_62_n22, cor_maj_62_n21, cor_maj_62_n20,
         cor_maj_62_n19, cor_maj_62_n18, cor_maj_63_n34, cor_maj_63_n33,
         cor_maj_63_n32, cor_maj_63_n31, cor_maj_63_n30, cor_maj_63_n29,
         cor_maj_63_n28, cor_maj_63_n27, cor_maj_63_n26, cor_maj_63_n25,
         cor_maj_63_n24, cor_maj_63_n23, cor_maj_63_n22, cor_maj_63_n21,
         cor_maj_63_n20, cor_maj_63_n19, cor_maj_63_n18, cor_maj_64_n34,
         cor_maj_64_n33, cor_maj_64_n32, cor_maj_64_n31, cor_maj_64_n30,
         cor_maj_64_n29, cor_maj_64_n28, cor_maj_64_n27, cor_maj_64_n26,
         cor_maj_64_n25, cor_maj_64_n24, cor_maj_64_n23, cor_maj_64_n22,
         cor_maj_64_n21, cor_maj_64_n20, cor_maj_64_n19, cor_maj_64_n18,
         cor_maj_65_n34, cor_maj_65_n33, cor_maj_65_n32, cor_maj_65_n31,
         cor_maj_65_n30, cor_maj_65_n29, cor_maj_65_n28, cor_maj_65_n27,
         cor_maj_65_n26, cor_maj_65_n25, cor_maj_65_n24, cor_maj_65_n23,
         cor_maj_65_n22, cor_maj_65_n21, cor_maj_65_n20, cor_maj_65_n19,
         cor_maj_65_n18, cor_maj_66_n34, cor_maj_66_n33, cor_maj_66_n32,
         cor_maj_66_n31, cor_maj_66_n30, cor_maj_66_n29, cor_maj_66_n28,
         cor_maj_66_n27, cor_maj_66_n26, cor_maj_66_n25, cor_maj_66_n24,
         cor_maj_66_n23, cor_maj_66_n22, cor_maj_66_n21, cor_maj_66_n20,
         cor_maj_66_n19, cor_maj_66_n18, cor_maj_67_n34, cor_maj_67_n33,
         cor_maj_67_n32, cor_maj_67_n31, cor_maj_67_n30, cor_maj_67_n29,
         cor_maj_67_n28, cor_maj_67_n27, cor_maj_67_n26, cor_maj_67_n25,
         cor_maj_67_n24, cor_maj_67_n23, cor_maj_67_n22, cor_maj_67_n21,
         cor_maj_67_n20, cor_maj_67_n19, cor_maj_67_n18, cor_maj_68_n34,
         cor_maj_68_n33, cor_maj_68_n32, cor_maj_68_n31, cor_maj_68_n30,
         cor_maj_68_n29, cor_maj_68_n28, cor_maj_68_n27, cor_maj_68_n26,
         cor_maj_68_n25, cor_maj_68_n24, cor_maj_68_n23, cor_maj_68_n22,
         cor_maj_68_n21, cor_maj_68_n20, cor_maj_68_n19, cor_maj_68_n18,
         cor_maj_69_n34, cor_maj_69_n33, cor_maj_69_n32, cor_maj_69_n31,
         cor_maj_69_n30, cor_maj_69_n29, cor_maj_69_n28, cor_maj_69_n27,
         cor_maj_69_n26, cor_maj_69_n25, cor_maj_69_n24, cor_maj_69_n23,
         cor_maj_69_n22, cor_maj_69_n21, cor_maj_69_n20, cor_maj_69_n19,
         cor_maj_69_n18, cor_maj_70_n34, cor_maj_70_n33, cor_maj_70_n32,
         cor_maj_70_n31, cor_maj_70_n30, cor_maj_70_n29, cor_maj_70_n28,
         cor_maj_70_n27, cor_maj_70_n26, cor_maj_70_n25, cor_maj_70_n24,
         cor_maj_70_n23, cor_maj_70_n22, cor_maj_70_n21, cor_maj_70_n20,
         cor_maj_70_n19, cor_maj_70_n18, cor_maj_71_n34, cor_maj_71_n33,
         cor_maj_71_n32, cor_maj_71_n31, cor_maj_71_n30, cor_maj_71_n29,
         cor_maj_71_n28, cor_maj_71_n27, cor_maj_71_n26, cor_maj_71_n25,
         cor_maj_71_n24, cor_maj_71_n23, cor_maj_71_n22, cor_maj_71_n21,
         cor_maj_71_n20, cor_maj_71_n19, cor_maj_71_n18, cor_maj_72_n34,
         cor_maj_72_n33, cor_maj_72_n32, cor_maj_72_n31, cor_maj_72_n30,
         cor_maj_72_n29, cor_maj_72_n28, cor_maj_72_n27, cor_maj_72_n26,
         cor_maj_72_n25, cor_maj_72_n24, cor_maj_72_n23, cor_maj_72_n22,
         cor_maj_72_n21, cor_maj_72_n20, cor_maj_72_n19, cor_maj_72_n18,
         cor_maj_73_n34, cor_maj_73_n33, cor_maj_73_n32, cor_maj_73_n31,
         cor_maj_73_n30, cor_maj_73_n29, cor_maj_73_n28, cor_maj_73_n27,
         cor_maj_73_n26, cor_maj_73_n25, cor_maj_73_n24, cor_maj_73_n23,
         cor_maj_73_n22, cor_maj_73_n21, cor_maj_73_n20, cor_maj_73_n19,
         cor_maj_73_n18, cor_maj_74_n34, cor_maj_74_n33, cor_maj_74_n32,
         cor_maj_74_n31, cor_maj_74_n30, cor_maj_74_n29, cor_maj_74_n28,
         cor_maj_74_n27, cor_maj_74_n26, cor_maj_74_n25, cor_maj_74_n24,
         cor_maj_74_n23, cor_maj_74_n22, cor_maj_74_n21, cor_maj_74_n20,
         cor_maj_74_n19, cor_maj_74_n18, cor_maj_75_n34, cor_maj_75_n33,
         cor_maj_75_n32, cor_maj_75_n31, cor_maj_75_n30, cor_maj_75_n29,
         cor_maj_75_n28, cor_maj_75_n27, cor_maj_75_n26, cor_maj_75_n25,
         cor_maj_75_n24, cor_maj_75_n23, cor_maj_75_n22, cor_maj_75_n21,
         cor_maj_75_n20, cor_maj_75_n19, cor_maj_75_n18, cor_maj_76_n34,
         cor_maj_76_n33, cor_maj_76_n32, cor_maj_76_n31, cor_maj_76_n30,
         cor_maj_76_n29, cor_maj_76_n28, cor_maj_76_n27, cor_maj_76_n26,
         cor_maj_76_n25, cor_maj_76_n24, cor_maj_76_n23, cor_maj_76_n22,
         cor_maj_76_n21, cor_maj_76_n20, cor_maj_76_n19, cor_maj_76_n18,
         cor_maj_77_n34, cor_maj_77_n33, cor_maj_77_n32, cor_maj_77_n31,
         cor_maj_77_n30, cor_maj_77_n29, cor_maj_77_n28, cor_maj_77_n27,
         cor_maj_77_n26, cor_maj_77_n25, cor_maj_77_n24, cor_maj_77_n23,
         cor_maj_77_n22, cor_maj_77_n21, cor_maj_77_n20, cor_maj_77_n19,
         cor_maj_77_n18, cor_maj_78_n34, cor_maj_78_n33, cor_maj_78_n32,
         cor_maj_78_n31, cor_maj_78_n30, cor_maj_78_n29, cor_maj_78_n28,
         cor_maj_78_n27, cor_maj_78_n26, cor_maj_78_n25, cor_maj_78_n24,
         cor_maj_78_n23, cor_maj_78_n22, cor_maj_78_n21, cor_maj_78_n20,
         cor_maj_78_n19, cor_maj_78_n18, cor_maj_79_n34, cor_maj_79_n33,
         cor_maj_79_n32, cor_maj_79_n31, cor_maj_79_n30, cor_maj_79_n29,
         cor_maj_79_n28, cor_maj_79_n27, cor_maj_79_n26, cor_maj_79_n25,
         cor_maj_79_n24, cor_maj_79_n23, cor_maj_79_n22, cor_maj_79_n21,
         cor_maj_79_n20, cor_maj_79_n19, cor_maj_79_n18, cor_maj_80_n34,
         cor_maj_80_n33, cor_maj_80_n32, cor_maj_80_n31, cor_maj_80_n30,
         cor_maj_80_n29, cor_maj_80_n28, cor_maj_80_n27, cor_maj_80_n26,
         cor_maj_80_n25, cor_maj_80_n24, cor_maj_80_n23, cor_maj_80_n22,
         cor_maj_80_n21, cor_maj_80_n20, cor_maj_80_n19, cor_maj_80_n18,
         cor_maj_81_n34, cor_maj_81_n33, cor_maj_81_n32, cor_maj_81_n31,
         cor_maj_81_n30, cor_maj_81_n29, cor_maj_81_n28, cor_maj_81_n27,
         cor_maj_81_n26, cor_maj_81_n25, cor_maj_81_n24, cor_maj_81_n23,
         cor_maj_81_n22, cor_maj_81_n21, cor_maj_81_n20, cor_maj_81_n19,
         cor_maj_81_n18, cor_maj_82_n34, cor_maj_82_n33, cor_maj_82_n32,
         cor_maj_82_n31, cor_maj_82_n30, cor_maj_82_n29, cor_maj_82_n28,
         cor_maj_82_n27, cor_maj_82_n26, cor_maj_82_n25, cor_maj_82_n24,
         cor_maj_82_n23, cor_maj_82_n22, cor_maj_82_n21, cor_maj_82_n20,
         cor_maj_82_n19, cor_maj_82_n18, cor_maj_83_n34, cor_maj_83_n33,
         cor_maj_83_n32, cor_maj_83_n31, cor_maj_83_n30, cor_maj_83_n29,
         cor_maj_83_n28, cor_maj_83_n27, cor_maj_83_n26, cor_maj_83_n25,
         cor_maj_83_n24, cor_maj_83_n23, cor_maj_83_n22, cor_maj_83_n21,
         cor_maj_83_n20, cor_maj_83_n19, cor_maj_83_n18;
  wire   [6:0] v_1_0_1;
  wire   [6:0] v_1_0_2;
  wire   [6:0] v_1_1_0;
  wire   [6:0] v_1_1_2;
  wire   [6:0] v_1_2_0;
  wire   [6:0] v_1_2_1;
  wire   [6:0] cor_port_v_0_1;
  wire   [6:0] cor_port_v_0_2;
  wire   [6:0] cor_port_v_1_0;
  wire   [6:0] cor_port_v_1_2;
  wire   [6:0] cor_port_v_2_0;
  wire   [6:0] cor_port_v_2_1;
  wire   [2:1] n_zz_io_c_0_3;
  wire   [6:0] u_0_1;
  wire   [6:0] u_0_2;
  wire   [2:1] n_zz_io_c_1_3;
  wire   [6:0] u_1_0;
  wire   [6:0] u_1_2;
  wire   [2:1] n_zz_io_c_2_3;
  wire   [6:0] u_2_0;
  wire   [6:0] u_2_1;
  wire   [2:1] n_zz_io_c_0_7;
  wire   [2:1] n_zz_io_c_1_7;
  wire   [2:1] n_zz_io_c_2_7;
  wire   [2:1] n_zz_io_c_0_11;
  wire   [2:1] n_zz_io_c_1_11;
  wire   [2:1] n_zz_io_c_2_11;
  wire   [2:1] n_zz_io_c_0_15;
  wire   [2:1] n_zz_io_c_1_15;
  wire   [2:1] n_zz_io_c_2_15;
  wire   [2:1] n_zz_io_c_0_19;
  wire   [2:1] n_zz_io_c_1_19;
  wire   [2:1] n_zz_io_c_2_19;
  wire   [2:1] n_zz_io_c_0_23;
  wire   [2:1] n_zz_io_c_1_23;
  wire   [2:1] n_zz_io_c_2_23;
  wire   [2:1] n_zz_io_c_0_27;
  wire   [2:1] n_zz_io_c_1_27;
  wire   [2:1] n_zz_io_c_2_27;
  wire   [6:0] rand_reg_0;
  wire   [6:0] rand_reg_1;
  wire   [6:0] rand_reg_3;
  wire   [6:0] rand_reg_2;
  wire   [6:0] rand_reg_4;
  wire   [6:0] rand_reg_5;
  wire   [6:0] b_reg_0;
  wire   [6:0] b_reg_1;
  wire   [6:0] b_reg_2;

  DFF_X1 rand_reg_2_reg_6_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[6]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_5_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[5]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[4]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[3]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[2]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[1]), 
        .QN() );
  DFF_X1 rand_reg_2_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[0]), 
        .QN() );
  DFF_X1 b_reg_1_reg_6_ ( .D(io_b_1[6]), .CK(clk), .Q(b_reg_1[6]), .QN() );
  DFF_X1 b_reg_1_reg_5_ ( .D(io_b_1[5]), .CK(clk), .Q(b_reg_1[5]), .QN() );
  DFF_X1 b_reg_1_reg_4_ ( .D(io_b_1[4]), .CK(clk), .Q(b_reg_1[4]), .QN() );
  DFF_X1 b_reg_1_reg_3_ ( .D(io_b_1[3]), .CK(clk), .Q(b_reg_1[3]), .QN() );
  DFF_X1 b_reg_1_reg_2_ ( .D(io_b_1[2]), .CK(clk), .Q(b_reg_1[2]), .QN() );
  DFF_X1 b_reg_1_reg_1_ ( .D(io_b_1[1]), .CK(clk), .Q(b_reg_1[1]), .QN() );
  DFF_X1 b_reg_1_reg_0_ ( .D(io_b_1[0]), .CK(clk), .Q(b_reg_1[0]), .QN() );
  DFF_X1 b_reg_2_reg_6_ ( .D(io_b_2[6]), .CK(clk), .Q(b_reg_2[6]), .QN() );
  DFF_X1 b_reg_2_reg_5_ ( .D(io_b_2[5]), .CK(clk), .Q(b_reg_2[5]), .QN() );
  DFF_X1 b_reg_2_reg_4_ ( .D(io_b_2[4]), .CK(clk), .Q(b_reg_2[4]), .QN() );
  DFF_X1 b_reg_2_reg_3_ ( .D(io_b_2[3]), .CK(clk), .Q(b_reg_2[3]), .QN() );
  DFF_X1 b_reg_2_reg_2_ ( .D(io_b_2[2]), .CK(clk), .Q(b_reg_2[2]), .QN() );
  DFF_X1 b_reg_2_reg_1_ ( .D(io_b_2[1]), .CK(clk), .Q(b_reg_2[1]), .QN() );
  DFF_X1 b_reg_2_reg_0_ ( .D(io_b_2[0]), .CK(clk), .Q(b_reg_2[0]), .QN() );
  DFF_X1 u_zz_io_c_2_27_reg_2_ ( .D(N104), .CK(clk), .Q(n_zz_io_c_2_27[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_27_reg_1_ ( .D(N103), .CK(clk), .Q(n_zz_io_c_2_27[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_27_reg_0_ ( .D(N102), .CK(clk), .Q(n_zz_io_c_2_24_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_27_reg_2_ ( .D(N101), .CK(clk), .Q(n_zz_io_c_1_27[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_27_reg_1_ ( .D(N100), .CK(clk), .Q(n_zz_io_c_1_27[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_27_reg_0_ ( .D(N99), .CK(clk), .Q(n_zz_io_c_1_24_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_27_reg_2_ ( .D(N98), .CK(clk), .Q(n_zz_io_c_0_27[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_27_reg_1_ ( .D(N97), .CK(clk), .Q(n_zz_io_c_0_27[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_23_reg_2_ ( .D(N95), .CK(clk), .Q(n_zz_io_c_2_23[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_23_reg_1_ ( .D(N94), .CK(clk), .Q(n_zz_io_c_2_23[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_23_reg_0_ ( .D(N93), .CK(clk), .Q(n_zz_io_c_2_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_23_reg_2_ ( .D(N92), .CK(clk), .Q(n_zz_io_c_1_23[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_23_reg_1_ ( .D(N91), .CK(clk), .Q(n_zz_io_c_1_23[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_23_reg_0_ ( .D(N90), .CK(clk), .Q(n_zz_io_c_1_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_23_reg_2_ ( .D(N89), .CK(clk), .Q(n_zz_io_c_0_23[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_23_reg_1_ ( .D(N88), .CK(clk), .Q(n_zz_io_c_0_23[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_2_ ( .D(N86), .CK(clk), .Q(n_zz_io_c_2_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_1_ ( .D(N85), .CK(clk), .Q(n_zz_io_c_2_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_0_ ( .D(N84), .CK(clk), .Q(n_zz_io_c_2_16_0_), 
        .QN() );
  DFF_X1 rand_reg_5_reg_6_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[6]), 
        .QN() );
  DFF_X1 u_2_1_reg_6_ ( .D(N41), .CK(clk), .Q(u_2_1[6]), .QN() );
  DFF_X1 rand_reg_5_reg_5_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[5]), 
        .QN() );
  DFF_X1 u_2_1_reg_5_ ( .D(N35), .CK(clk), .Q(u_2_1[5]), .QN() );
  DFF_X1 rand_reg_5_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[4]), 
        .QN() );
  DFF_X1 u_2_1_reg_4_ ( .D(N29), .CK(clk), .Q(u_2_1[4]), .QN() );
  DFF_X1 rand_reg_5_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[3]), 
        .QN() );
  DFF_X1 u_2_1_reg_3_ ( .D(N23), .CK(clk), .Q(u_2_1[3]), .QN() );
  DFF_X1 rand_reg_5_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[2]), 
        .QN() );
  DFF_X1 u_2_1_reg_2_ ( .D(N17), .CK(clk), .Q(u_2_1[2]), .QN() );
  DFF_X1 rand_reg_5_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[1]), 
        .QN() );
  DFF_X1 u_2_1_reg_1_ ( .D(N11), .CK(clk), .Q(u_2_1[1]), .QN() );
  DFF_X1 rand_reg_5_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_5[0]), 
        .QN() );
  DFF_X1 u_2_1_reg_0_ ( .D(N5), .CK(clk), .Q(u_2_1[0]), .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_2_ ( .D(N83), .CK(clk), .Q(n_zz_io_c_1_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_1_ ( .D(N82), .CK(clk), .Q(n_zz_io_c_1_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_0_ ( .D(N81), .CK(clk), .Q(n_zz_io_c_1_16_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_2_ ( .D(N80), .CK(clk), .Q(n_zz_io_c_0_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_1_ ( .D(N79), .CK(clk), .Q(n_zz_io_c_0_19[1]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_6_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[6]), 
        .QN() );
  DFF_X1 u_0_1_reg_6_ ( .D(N36), .CK(clk), .Q(u_0_1[6]), .QN() );
  DFF_X1 rand_reg_0_reg_5_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[5]), 
        .QN() );
  DFF_X1 u_0_1_reg_5_ ( .D(N30), .CK(clk), .Q(u_0_1[5]), .QN() );
  DFF_X1 rand_reg_0_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[4]), 
        .QN() );
  DFF_X1 u_0_1_reg_4_ ( .D(N24), .CK(clk), .Q(u_0_1[4]), .QN() );
  DFF_X1 rand_reg_0_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[3]), 
        .QN() );
  DFF_X1 u_0_1_reg_3_ ( .D(N18), .CK(clk), .Q(u_0_1[3]), .QN() );
  DFF_X1 rand_reg_0_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[2]), 
        .QN() );
  DFF_X1 u_0_1_reg_2_ ( .D(N12), .CK(clk), .Q(u_0_1[2]), .QN() );
  DFF_X1 rand_reg_0_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[1]), 
        .QN() );
  DFF_X1 u_0_1_reg_1_ ( .D(N6), .CK(clk), .Q(u_0_1[1]), .QN() );
  DFF_X1 rand_reg_0_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[0]), 
        .QN() );
  DFF_X1 u_0_1_reg_0_ ( .D(N0), .CK(clk), .Q(u_0_1[0]), .QN() );
  DFF_X1 rand_reg_3_reg_6_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[6]), 
        .QN() );
  DFF_X1 u_1_0_reg_6_ ( .D(N38), .CK(clk), .Q(u_1_0[6]), .QN() );
  DFF_X1 rand_reg_3_reg_5_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[5]), 
        .QN() );
  DFF_X1 u_1_0_reg_5_ ( .D(N32), .CK(clk), .Q(u_1_0[5]), .QN() );
  DFF_X1 rand_reg_3_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[4]), 
        .QN() );
  DFF_X1 u_1_0_reg_4_ ( .D(N26), .CK(clk), .Q(u_1_0[4]), .QN() );
  DFF_X1 rand_reg_3_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[3]), 
        .QN() );
  DFF_X1 u_1_0_reg_3_ ( .D(N20), .CK(clk), .Q(u_1_0[3]), .QN() );
  DFF_X1 rand_reg_3_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[2]), 
        .QN() );
  DFF_X1 u_1_0_reg_2_ ( .D(N14), .CK(clk), .Q(u_1_0[2]), .QN() );
  DFF_X1 rand_reg_3_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[1]), 
        .QN() );
  DFF_X1 u_1_0_reg_1_ ( .D(N8), .CK(clk), .Q(u_1_0[1]), .QN() );
  DFF_X1 rand_reg_3_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_3[0]), 
        .QN() );
  DFF_X1 u_1_0_reg_0_ ( .D(N2), .CK(clk), .Q(u_1_0[0]), .QN() );
  DFF_X1 u_1_2_reg_6_ ( .D(N39), .CK(clk), .Q(u_1_2[6]), .QN() );
  DFF_X1 u_1_2_reg_5_ ( .D(N33), .CK(clk), .Q(u_1_2[5]), .QN() );
  DFF_X1 u_1_2_reg_4_ ( .D(N27), .CK(clk), .Q(u_1_2[4]), .QN() );
  DFF_X1 u_1_2_reg_3_ ( .D(N21), .CK(clk), .Q(u_1_2[3]), .QN() );
  DFF_X1 u_1_2_reg_2_ ( .D(N15), .CK(clk), .Q(u_1_2[2]), .QN() );
  DFF_X1 u_1_2_reg_1_ ( .D(N9), .CK(clk), .Q(u_1_2[1]), .QN() );
  DFF_X1 u_1_2_reg_0_ ( .D(N3), .CK(clk), .Q(u_1_2[0]), .QN() );
  DFF_X1 u_zz_io_c_2_15_reg_2_ ( .D(N77), .CK(clk), .Q(n_zz_io_c_2_15[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_15_reg_1_ ( .D(N76), .CK(clk), .Q(n_zz_io_c_2_15[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_15_reg_0_ ( .D(N75), .CK(clk), .Q(n_zz_io_c_2_12_0_), 
        .QN() );
  DFF_X1 rand_reg_1_reg_6_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[6]), 
        .QN() );
  DFF_X1 u_0_2_reg_6_ ( .D(N37), .CK(clk), .Q(u_0_2[6]), .QN() );
  DFF_X1 rand_reg_1_reg_5_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[5]), 
        .QN() );
  DFF_X1 u_0_2_reg_5_ ( .D(N31), .CK(clk), .Q(u_0_2[5]), .QN() );
  DFF_X1 rand_reg_1_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[4]), 
        .QN() );
  DFF_X1 u_0_2_reg_4_ ( .D(N25), .CK(clk), .Q(u_0_2[4]), .QN() );
  DFF_X1 rand_reg_1_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[3]), 
        .QN() );
  DFF_X1 u_0_2_reg_3_ ( .D(N19), .CK(clk), .Q(u_0_2[3]), .QN() );
  DFF_X1 rand_reg_1_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[2]), 
        .QN() );
  DFF_X1 u_0_2_reg_2_ ( .D(N13), .CK(clk), .Q(u_0_2[2]), .QN() );
  DFF_X1 rand_reg_1_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[1]), 
        .QN() );
  DFF_X1 u_0_2_reg_1_ ( .D(N7), .CK(clk), .Q(u_0_2[1]), .QN() );
  DFF_X1 rand_reg_1_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[0]), 
        .QN() );
  DFF_X1 u_0_2_reg_0_ ( .D(N1), .CK(clk), .Q(u_0_2[0]), .QN() );
  DFF_X1 rand_reg_4_reg_6_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[6]), 
        .QN() );
  DFF_X1 u_2_0_reg_6_ ( .D(N40), .CK(clk), .Q(u_2_0[6]), .QN() );
  DFF_X1 rand_reg_4_reg_5_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[5]), 
        .QN() );
  DFF_X1 u_2_0_reg_5_ ( .D(N34), .CK(clk), .Q(u_2_0[5]), .QN() );
  DFF_X1 rand_reg_4_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[4]), 
        .QN() );
  DFF_X1 u_2_0_reg_4_ ( .D(N28), .CK(clk), .Q(u_2_0[4]), .QN() );
  DFF_X1 rand_reg_4_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[3]), 
        .QN() );
  DFF_X1 u_2_0_reg_3_ ( .D(N22), .CK(clk), .Q(u_2_0[3]), .QN() );
  DFF_X1 rand_reg_4_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[2]), 
        .QN() );
  DFF_X1 u_2_0_reg_2_ ( .D(N16), .CK(clk), .Q(u_2_0[2]), .QN() );
  DFF_X1 rand_reg_4_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[1]), 
        .QN() );
  DFF_X1 u_2_0_reg_1_ ( .D(N10), .CK(clk), .Q(u_2_0[1]), .QN() );
  DFF_X1 rand_reg_4_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_4[0]), 
        .QN() );
  DFF_X1 u_2_0_reg_0_ ( .D(N4), .CK(clk), .Q(u_2_0[0]), .QN() );
  DFF_X1 b_reg_0_reg_6_ ( .D(io_b_0[6]), .CK(clk), .Q(b_reg_0[6]), .QN() );
  DFF_X1 u_zz_io_c_0_27_reg_0_ ( .D(N96), .CK(clk), .Q(n_zz_io_c_0_24_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_5_ ( .D(io_b_0[5]), .CK(clk), .Q(b_reg_0[5]), .QN() );
  DFF_X1 u_zz_io_c_0_23_reg_0_ ( .D(N87), .CK(clk), .Q(n_zz_io_c_0_20_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_4_ ( .D(io_b_0[4]), .CK(clk), .Q(b_reg_0[4]), .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_0_ ( .D(N78), .CK(clk), .Q(n_zz_io_c_0_16_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_3_ ( .D(io_b_0[3]), .CK(clk), .Q(b_reg_0[3]), .QN() );
  DFF_X1 b_reg_0_reg_2_ ( .D(io_b_0[2]), .CK(clk), .Q(b_reg_0[2]), .QN() );
  DFF_X1 b_reg_0_reg_1_ ( .D(io_b_0[1]), .CK(clk), .Q(b_reg_0[1]), .QN() );
  DFF_X1 b_reg_0_reg_0_ ( .D(io_b_0[0]), .CK(clk), .Q(b_reg_0[0]), .QN() );
  DFF_X1 u_zz_io_c_1_15_reg_2_ ( .D(N74), .CK(clk), .Q(n_zz_io_c_1_15[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_15_reg_1_ ( .D(N73), .CK(clk), .Q(n_zz_io_c_1_15[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_15_reg_0_ ( .D(N72), .CK(clk), .Q(n_zz_io_c_1_12_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_15_reg_2_ ( .D(N71), .CK(clk), .Q(n_zz_io_c_0_15[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_15_reg_1_ ( .D(N70), .CK(clk), .Q(n_zz_io_c_0_15[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_15_reg_0_ ( .D(N69), .CK(clk), .Q(n_zz_io_c_0_12_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_11_reg_2_ ( .D(N68), .CK(clk), .Q(n_zz_io_c_2_11[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_11_reg_1_ ( .D(N67), .CK(clk), .Q(n_zz_io_c_2_11[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_11_reg_0_ ( .D(N66), .CK(clk), .Q(n_zz_io_c_2_8_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_2_ ( .D(N65), .CK(clk), .Q(n_zz_io_c_1_11[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_1_ ( .D(N64), .CK(clk), .Q(n_zz_io_c_1_11[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_0_ ( .D(N63), .CK(clk), .Q(n_zz_io_c_1_8_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_2_ ( .D(N62), .CK(clk), .Q(n_zz_io_c_0_11[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_1_ ( .D(N61), .CK(clk), .Q(n_zz_io_c_0_11[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_0_ ( .D(N60), .CK(clk), .Q(n_zz_io_c_0_8_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_7_reg_2_ ( .D(N59), .CK(clk), .Q(n_zz_io_c_2_7[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_7_reg_1_ ( .D(N58), .CK(clk), .Q(n_zz_io_c_2_7[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_7_reg_0_ ( .D(N57), .CK(clk), .Q(n_zz_io_c_2_4_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_7_reg_2_ ( .D(N56), .CK(clk), .Q(n_zz_io_c_1_7[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_7_reg_1_ ( .D(N55), .CK(clk), .Q(n_zz_io_c_1_7[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_7_reg_0_ ( .D(N54), .CK(clk), .Q(n_zz_io_c_1_4_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_7_reg_2_ ( .D(N53), .CK(clk), .Q(n_zz_io_c_0_7[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_7_reg_1_ ( .D(N52), .CK(clk), .Q(n_zz_io_c_0_7[1]), .QN()
         );
  DFF_X1 u_zz_io_c_0_7_reg_0_ ( .D(N51), .CK(clk), .Q(n_zz_io_c_0_4_0_), .QN()
         );
  DFF_X1 u_zz_io_c_2_3_reg_2_ ( .D(N50), .CK(clk), .Q(n_zz_io_c_2_3[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_3_reg_1_ ( .D(N49), .CK(clk), .Q(n_zz_io_c_2_3[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_3_reg_0_ ( .D(N48), .CK(clk), .Q(n_zz_io_c_2_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_3_reg_2_ ( .D(N47), .CK(clk), .Q(n_zz_io_c_1_3[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_3_reg_1_ ( .D(N46), .CK(clk), .Q(n_zz_io_c_1_3[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_3_reg_0_ ( .D(N45), .CK(clk), .Q(n_zz_io_c_1_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_3_reg_2_ ( .D(N44), .CK(clk), .Q(n_zz_io_c_0_3[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_3_reg_1_ ( .D(N43), .CK(clk), .Q(n_zz_io_c_0_3[1]), .QN()
         );
  DFF_X1 u_zz_io_c_0_3_reg_0_ ( .D(N42), .CK(clk), .Q(n_zz_io_c_0_0_), .QN()
         );
  XOR2_X2 U4 ( .A(io_rand[2]), .B(io_b_1[5]), .Z(v_1_2_1[5]) );
  XOR2_X2 U5 ( .A(io_rand[2]), .B(io_b_1[4]), .Z(v_1_2_1[4]) );
  XOR2_X2 U6 ( .A(io_rand[2]), .B(io_b_1[3]), .Z(v_1_2_1[3]) );
  XOR2_X2 U7 ( .A(io_rand[2]), .B(io_b_1[2]), .Z(v_1_2_1[2]) );
  XOR2_X2 U8 ( .A(io_rand[2]), .B(io_b_1[1]), .Z(v_1_2_1[1]) );
  XOR2_X2 U9 ( .A(io_rand[2]), .B(io_b_1[0]), .Z(v_1_2_1[0]) );
  XOR2_X2 U11 ( .A(io_rand[1]), .B(io_b_0[5]), .Z(v_1_2_0[5]) );
  XOR2_X2 U12 ( .A(io_rand[1]), .B(io_b_0[4]), .Z(v_1_2_0[4]) );
  XOR2_X2 U13 ( .A(io_rand[1]), .B(io_b_0[3]), .Z(v_1_2_0[3]) );
  XOR2_X2 U14 ( .A(io_rand[1]), .B(io_b_0[2]), .Z(v_1_2_0[2]) );
  XOR2_X2 U15 ( .A(io_rand[1]), .B(io_b_0[1]), .Z(v_1_2_0[1]) );
  XOR2_X2 U16 ( .A(io_rand[1]), .B(io_b_0[0]), .Z(v_1_2_0[0]) );
  XOR2_X2 U18 ( .A(io_rand[2]), .B(io_b_2[5]), .Z(v_1_1_2[5]) );
  XOR2_X2 U19 ( .A(io_rand[2]), .B(io_b_2[4]), .Z(v_1_1_2[4]) );
  XOR2_X2 U20 ( .A(io_rand[2]), .B(io_b_2[3]), .Z(v_1_1_2[3]) );
  XOR2_X2 U21 ( .A(io_rand[2]), .B(io_b_2[2]), .Z(v_1_1_2[2]) );
  XOR2_X2 U22 ( .A(io_rand[2]), .B(io_b_2[1]), .Z(v_1_1_2[1]) );
  XOR2_X2 U23 ( .A(io_rand[2]), .B(io_b_2[0]), .Z(v_1_1_2[0]) );
  XOR2_X2 U25 ( .A(io_rand[0]), .B(io_b_0[5]), .Z(v_1_1_0[5]) );
  XOR2_X2 U26 ( .A(io_rand[0]), .B(io_b_0[4]), .Z(v_1_1_0[4]) );
  XOR2_X2 U27 ( .A(io_rand[0]), .B(io_b_0[3]), .Z(v_1_1_0[3]) );
  XOR2_X2 U28 ( .A(io_rand[0]), .B(io_b_0[2]), .Z(v_1_1_0[2]) );
  XOR2_X2 U29 ( .A(io_rand[0]), .B(io_b_0[1]), .Z(v_1_1_0[1]) );
  XOR2_X2 U30 ( .A(io_rand[0]), .B(io_b_0[0]), .Z(v_1_1_0[0]) );
  XOR2_X2 U32 ( .A(io_rand[1]), .B(io_b_2[5]), .Z(v_1_0_2[5]) );
  XOR2_X2 U33 ( .A(io_rand[1]), .B(io_b_2[4]), .Z(v_1_0_2[4]) );
  XOR2_X2 U34 ( .A(io_rand[1]), .B(io_b_2[3]), .Z(v_1_0_2[3]) );
  XOR2_X2 U35 ( .A(io_rand[1]), .B(io_b_2[2]), .Z(v_1_0_2[2]) );
  XOR2_X2 U36 ( .A(io_rand[1]), .B(io_b_2[1]), .Z(v_1_0_2[1]) );
  XOR2_X2 U37 ( .A(io_rand[1]), .B(io_b_2[0]), .Z(v_1_0_2[0]) );
  XOR2_X2 U39 ( .A(io_rand[0]), .B(io_b_1[5]), .Z(v_1_0_1[5]) );
  XOR2_X2 U40 ( .A(io_rand[0]), .B(io_b_1[4]), .Z(v_1_0_1[4]) );
  XOR2_X2 U41 ( .A(io_rand[0]), .B(io_b_1[3]), .Z(v_1_0_1[3]) );
  XOR2_X2 U42 ( .A(io_rand[0]), .B(io_b_1[2]), .Z(v_1_0_1[2]) );
  XOR2_X2 U43 ( .A(io_rand[0]), .B(io_b_1[1]), .Z(v_1_0_1[1]) );
  XOR2_X2 U44 ( .A(io_rand[0]), .B(io_b_1[0]), .Z(v_1_0_1[0]) );
  XOR2_X1 U192 ( .A(io_rand[2]), .B(io_b_1[6]), .Z(v_1_2_1[6]) );
  XOR2_X1 U193 ( .A(io_rand[1]), .B(io_b_0[6]), .Z(v_1_2_0[6]) );
  XOR2_X1 U194 ( .A(io_rand[2]), .B(io_b_2[6]), .Z(v_1_1_2[6]) );
  XOR2_X1 U195 ( .A(io_rand[0]), .B(io_b_0[6]), .Z(v_1_1_0[6]) );
  XOR2_X1 U196 ( .A(io_rand[1]), .B(io_b_2[6]), .Z(v_1_0_2[6]) );
  XOR2_X1 U197 ( .A(io_rand[0]), .B(io_b_1[6]), .Z(v_1_0_1[6]) );
  AND2_X1 U198 ( .A1(b_reg_0[0]), .A2(io_a_0[0]), .ZN(N42) );
  AND2_X1 U199 ( .A1(cor_port_v_0_1[0]), .A2(io_a_0[0]), .ZN(N43) );
  AND2_X1 U200 ( .A1(b_reg_1[0]), .A2(io_a_1[0]), .ZN(N45) );
  AND2_X1 U201 ( .A1(cor_port_v_1_0[0]), .A2(io_a_1[0]), .ZN(N46) );
  AND2_X1 U202 ( .A1(b_reg_2[0]), .A2(io_a_2[0]), .ZN(N48) );
  AND2_X1 U203 ( .A1(cor_port_v_2_0[0]), .A2(io_a_2[0]), .ZN(N49) );
  AND2_X1 U204 ( .A1(b_reg_0[1]), .A2(io_a_0[1]), .ZN(N51) );
  AND2_X1 U205 ( .A1(cor_port_v_0_1[1]), .A2(io_a_0[1]), .ZN(N52) );
  AND2_X1 U206 ( .A1(b_reg_1[1]), .A2(io_a_1[1]), .ZN(N54) );
  AND2_X1 U207 ( .A1(cor_port_v_1_0[1]), .A2(io_a_1[1]), .ZN(N55) );
  AND2_X1 U208 ( .A1(b_reg_2[1]), .A2(io_a_2[1]), .ZN(N57) );
  AND2_X1 U209 ( .A1(cor_port_v_2_0[1]), .A2(io_a_2[1]), .ZN(N58) );
  AND2_X1 U210 ( .A1(b_reg_0[2]), .A2(io_a_0[2]), .ZN(N60) );
  AND2_X1 U211 ( .A1(cor_port_v_0_1[2]), .A2(io_a_0[2]), .ZN(N61) );
  AND2_X1 U212 ( .A1(b_reg_1[2]), .A2(io_a_1[2]), .ZN(N63) );
  AND2_X1 U213 ( .A1(cor_port_v_1_0[2]), .A2(io_a_1[2]), .ZN(N64) );
  AND2_X1 U214 ( .A1(b_reg_2[2]), .A2(io_a_2[2]), .ZN(N66) );
  AND2_X1 U215 ( .A1(cor_port_v_2_0[2]), .A2(io_a_2[2]), .ZN(N67) );
  AND2_X1 U216 ( .A1(b_reg_0[3]), .A2(io_a_0[3]), .ZN(N69) );
  AND2_X1 U217 ( .A1(cor_port_v_0_1[3]), .A2(io_a_0[3]), .ZN(N70) );
  AND2_X1 U218 ( .A1(b_reg_1[3]), .A2(io_a_1[3]), .ZN(N72) );
  AND2_X1 U219 ( .A1(cor_port_v_1_0[3]), .A2(io_a_1[3]), .ZN(N73) );
  AND2_X1 U220 ( .A1(b_reg_0[4]), .A2(io_a_0[4]), .ZN(N78) );
  AND2_X1 U221 ( .A1(b_reg_0[5]), .A2(io_a_0[5]), .ZN(N87) );
  AND2_X1 U222 ( .A1(b_reg_0[6]), .A2(io_a_0[6]), .ZN(N96) );
  AND2_X1 U223 ( .A1(b_reg_2[3]), .A2(io_a_2[3]), .ZN(N75) );
  AND2_X1 U224 ( .A1(cor_port_v_2_0[3]), .A2(io_a_2[3]), .ZN(N76) );
  AND2_X1 U225 ( .A1(cor_port_v_0_1[4]), .A2(io_a_0[4]), .ZN(N79) );
  AND2_X1 U226 ( .A1(b_reg_1[4]), .A2(io_a_1[4]), .ZN(N81) );
  AND2_X1 U227 ( .A1(cor_port_v_1_0[4]), .A2(io_a_1[4]), .ZN(N82) );
  AND2_X1 U228 ( .A1(b_reg_2[4]), .A2(io_a_2[4]), .ZN(N84) );
  AND2_X1 U229 ( .A1(cor_port_v_2_0[4]), .A2(io_a_2[4]), .ZN(N85) );
  AND2_X1 U230 ( .A1(cor_port_v_0_1[5]), .A2(io_a_0[5]), .ZN(N88) );
  AND2_X1 U231 ( .A1(b_reg_1[5]), .A2(io_a_1[5]), .ZN(N90) );
  AND2_X1 U232 ( .A1(cor_port_v_1_0[5]), .A2(io_a_1[5]), .ZN(N91) );
  AND2_X1 U233 ( .A1(b_reg_2[5]), .A2(io_a_2[5]), .ZN(N93) );
  AND2_X1 U234 ( .A1(cor_port_v_2_0[5]), .A2(io_a_2[5]), .ZN(N94) );
  AND2_X1 U235 ( .A1(cor_port_v_0_1[6]), .A2(io_a_0[6]), .ZN(N97) );
  AND2_X1 U236 ( .A1(cor_port_v_1_0[6]), .A2(io_a_1[6]), .ZN(N100) );
  AND2_X1 U237 ( .A1(cor_port_v_1_2[6]), .A2(io_a_1[6]), .ZN(N101) );
  AND2_X1 U238 ( .A1(b_reg_2[6]), .A2(io_a_2[6]), .ZN(N102) );
  AND2_X1 U239 ( .A1(cor_port_v_2_0[6]), .A2(io_a_2[6]), .ZN(N103) );
  AND2_X1 U240 ( .A1(io_a_0[0]), .A2(cor_port_v_0_2[0]), .ZN(N44) );
  AND2_X1 U241 ( .A1(io_a_1[0]), .A2(cor_port_v_1_2[0]), .ZN(N47) );
  AND2_X1 U242 ( .A1(io_a_2[0]), .A2(cor_port_v_2_1[0]), .ZN(N50) );
  AND2_X1 U243 ( .A1(io_a_0[1]), .A2(cor_port_v_0_2[1]), .ZN(N53) );
  AND2_X1 U244 ( .A1(io_a_1[1]), .A2(cor_port_v_1_2[1]), .ZN(N56) );
  AND2_X1 U245 ( .A1(io_a_2[1]), .A2(cor_port_v_2_1[1]), .ZN(N59) );
  AND2_X1 U246 ( .A1(io_a_0[2]), .A2(cor_port_v_0_2[2]), .ZN(N62) );
  AND2_X1 U247 ( .A1(io_a_1[2]), .A2(cor_port_v_1_2[2]), .ZN(N65) );
  AND2_X1 U248 ( .A1(io_a_2[2]), .A2(cor_port_v_2_1[2]), .ZN(N68) );
  AND2_X1 U249 ( .A1(io_a_0[3]), .A2(cor_port_v_0_2[3]), .ZN(N71) );
  AND2_X1 U250 ( .A1(io_a_1[3]), .A2(cor_port_v_1_2[3]), .ZN(N74) );
  AND2_X1 U251 ( .A1(simpleNot_46_port_z), .A2(rand_reg_4[0]), .ZN(N4) );
  AND2_X1 U252 ( .A1(simpleNot_52_port_z), .A2(rand_reg_4[1]), .ZN(N10) );
  AND2_X1 U253 ( .A1(simpleNot_58_port_z), .A2(rand_reg_4[2]), .ZN(N16) );
  AND2_X1 U254 ( .A1(simpleNot_64_port_z), .A2(rand_reg_4[3]), .ZN(N22) );
  AND2_X1 U255 ( .A1(simpleNot_70_port_z), .A2(rand_reg_4[4]), .ZN(N28) );
  AND2_X1 U256 ( .A1(simpleNot_76_port_z), .A2(rand_reg_4[5]), .ZN(N34) );
  AND2_X1 U257 ( .A1(simpleNot_82_port_z), .A2(rand_reg_4[6]), .ZN(N40) );
  AND2_X1 U258 ( .A1(simpleNot_43_port_z), .A2(rand_reg_1[0]), .ZN(N1) );
  AND2_X1 U259 ( .A1(simpleNot_49_port_z), .A2(rand_reg_1[1]), .ZN(N7) );
  AND2_X1 U260 ( .A1(simpleNot_55_port_z), .A2(rand_reg_1[2]), .ZN(N13) );
  AND2_X1 U261 ( .A1(simpleNot_61_port_z), .A2(rand_reg_1[3]), .ZN(N19) );
  AND2_X1 U262 ( .A1(simpleNot_67_port_z), .A2(rand_reg_1[4]), .ZN(N25) );
  AND2_X1 U263 ( .A1(simpleNot_73_port_z), .A2(rand_reg_1[5]), .ZN(N31) );
  AND2_X1 U264 ( .A1(simpleNot_79_port_z), .A2(rand_reg_1[6]), .ZN(N37) );
  AND2_X1 U265 ( .A1(io_a_2[3]), .A2(cor_port_v_2_1[3]), .ZN(N77) );
  AND2_X1 U266 ( .A1(simpleNot_45_port_z), .A2(rand_reg_2[0]), .ZN(N3) );
  AND2_X1 U267 ( .A1(simpleNot_51_port_z), .A2(rand_reg_2[1]), .ZN(N9) );
  AND2_X1 U268 ( .A1(simpleNot_57_port_z), .A2(rand_reg_2[2]), .ZN(N15) );
  AND2_X1 U269 ( .A1(simpleNot_63_port_z), .A2(rand_reg_2[3]), .ZN(N21) );
  AND2_X1 U270 ( .A1(simpleNot_69_port_z), .A2(rand_reg_2[4]), .ZN(N27) );
  AND2_X1 U271 ( .A1(simpleNot_75_port_z), .A2(rand_reg_2[5]), .ZN(N33) );
  AND2_X1 U272 ( .A1(simpleNot_81_port_z), .A2(rand_reg_2[6]), .ZN(N39) );
  AND2_X1 U273 ( .A1(simpleNot_44_port_z), .A2(rand_reg_3[0]), .ZN(N2) );
  AND2_X1 U274 ( .A1(simpleNot_50_port_z), .A2(rand_reg_3[1]), .ZN(N8) );
  AND2_X1 U275 ( .A1(simpleNot_56_port_z), .A2(rand_reg_3[2]), .ZN(N14) );
  AND2_X1 U276 ( .A1(simpleNot_62_port_z), .A2(rand_reg_3[3]), .ZN(N20) );
  AND2_X1 U277 ( .A1(simpleNot_68_port_z), .A2(rand_reg_3[4]), .ZN(N26) );
  AND2_X1 U278 ( .A1(simpleNot_74_port_z), .A2(rand_reg_3[5]), .ZN(N32) );
  AND2_X1 U279 ( .A1(simpleNot_80_port_z), .A2(rand_reg_3[6]), .ZN(N38) );
  AND2_X1 U280 ( .A1(simpleNot_42_port_z), .A2(rand_reg_0[0]), .ZN(N0) );
  AND2_X1 U281 ( .A1(simpleNot_48_port_z), .A2(rand_reg_0[1]), .ZN(N6) );
  AND2_X1 U282 ( .A1(simpleNot_54_port_z), .A2(rand_reg_0[2]), .ZN(N12) );
  AND2_X1 U283 ( .A1(simpleNot_60_port_z), .A2(rand_reg_0[3]), .ZN(N18) );
  AND2_X1 U284 ( .A1(simpleNot_66_port_z), .A2(rand_reg_0[4]), .ZN(N24) );
  AND2_X1 U285 ( .A1(simpleNot_72_port_z), .A2(rand_reg_0[5]), .ZN(N30) );
  AND2_X1 U286 ( .A1(simpleNot_78_port_z), .A2(rand_reg_0[6]), .ZN(N36) );
  AND2_X1 U287 ( .A1(io_a_0[4]), .A2(cor_port_v_0_2[4]), .ZN(N80) );
  AND2_X1 U288 ( .A1(io_a_1[4]), .A2(cor_port_v_1_2[4]), .ZN(N83) );
  AND2_X1 U289 ( .A1(simpleNot_47_port_z), .A2(rand_reg_5[0]), .ZN(N5) );
  AND2_X1 U290 ( .A1(simpleNot_53_port_z), .A2(rand_reg_5[1]), .ZN(N11) );
  AND2_X1 U291 ( .A1(simpleNot_59_port_z), .A2(rand_reg_5[2]), .ZN(N17) );
  AND2_X1 U292 ( .A1(simpleNot_65_port_z), .A2(rand_reg_5[3]), .ZN(N23) );
  AND2_X1 U293 ( .A1(simpleNot_71_port_z), .A2(rand_reg_5[4]), .ZN(N29) );
  AND2_X1 U294 ( .A1(simpleNot_77_port_z), .A2(rand_reg_5[5]), .ZN(N35) );
  AND2_X1 U295 ( .A1(simpleNot_83_port_z), .A2(rand_reg_5[6]), .ZN(N41) );
  AND2_X1 U296 ( .A1(io_a_2[4]), .A2(cor_port_v_2_1[4]), .ZN(N86) );
  AND2_X1 U297 ( .A1(io_a_0[5]), .A2(cor_port_v_0_2[5]), .ZN(N89) );
  AND2_X1 U298 ( .A1(io_a_1[5]), .A2(cor_port_v_1_2[5]), .ZN(N92) );
  AND2_X1 U299 ( .A1(io_a_2[5]), .A2(cor_port_v_2_1[5]), .ZN(N95) );
  AND2_X1 U300 ( .A1(io_a_0[6]), .A2(cor_port_v_0_2[6]), .ZN(N98) );
  AND2_X1 U301 ( .A1(io_a_1[6]), .A2(b_reg_1[6]), .ZN(N99) );
  AND2_X1 U302 ( .A1(io_a_2[6]), .A2(cor_port_v_2_1[6]), .ZN(N104) );
  XOR2_X1 U303 ( .A(n_zz_io_c_2_0_), .B(n7), .Z(io_c_2[0]) );
  XOR2_X1 U304 ( .A(simpleXor_47_port_z), .B(simpleXor_46_port_z), .Z(n7) );
  XOR2_X1 U305 ( .A(n_zz_io_c_2_4_0_), .B(n6), .Z(io_c_2[1]) );
  XOR2_X1 U306 ( .A(simpleXor_53_port_z), .B(simpleXor_52_port_z), .Z(n6) );
  XOR2_X1 U307 ( .A(n_zz_io_c_2_8_0_), .B(n5), .Z(io_c_2[2]) );
  XOR2_X1 U308 ( .A(simpleXor_59_port_z), .B(simpleXor_58_port_z), .Z(n5) );
  XOR2_X1 U309 ( .A(n_zz_io_c_2_12_0_), .B(n4), .Z(io_c_2[3]) );
  XOR2_X1 U310 ( .A(simpleXor_65_port_z), .B(simpleXor_64_port_z), .Z(n4) );
  XOR2_X1 U311 ( .A(n_zz_io_c_2_16_0_), .B(n3), .Z(io_c_2[4]) );
  XOR2_X1 U312 ( .A(simpleXor_71_port_z), .B(simpleXor_70_port_z), .Z(n3) );
  XOR2_X1 U313 ( .A(n_zz_io_c_2_20_0_), .B(n2), .Z(io_c_2[5]) );
  XOR2_X1 U314 ( .A(simpleXor_77_port_z), .B(simpleXor_76_port_z), .Z(n2) );
  XOR2_X1 U315 ( .A(n_zz_io_c_2_24_0_), .B(n1), .Z(io_c_2[6]) );
  XOR2_X1 U316 ( .A(simpleXor_83_port_z), .B(simpleXor_82_port_z), .Z(n1) );
  XOR2_X1 U317 ( .A(n_zz_io_c_1_0_), .B(n14), .Z(io_c_1[0]) );
  XOR2_X1 U318 ( .A(simpleXor_45_port_z), .B(simpleXor_44_port_z), .Z(n14) );
  XOR2_X1 U319 ( .A(n_zz_io_c_1_4_0_), .B(n13), .Z(io_c_1[1]) );
  XOR2_X1 U320 ( .A(simpleXor_51_port_z), .B(simpleXor_50_port_z), .Z(n13) );
  XOR2_X1 U321 ( .A(n_zz_io_c_1_8_0_), .B(n12), .Z(io_c_1[2]) );
  XOR2_X1 U322 ( .A(simpleXor_57_port_z), .B(simpleXor_56_port_z), .Z(n12) );
  XOR2_X1 U323 ( .A(n_zz_io_c_1_12_0_), .B(n11), .Z(io_c_1[3]) );
  XOR2_X1 U324 ( .A(simpleXor_63_port_z), .B(simpleXor_62_port_z), .Z(n11) );
  XOR2_X1 U325 ( .A(n_zz_io_c_1_16_0_), .B(n10), .Z(io_c_1[4]) );
  XOR2_X1 U326 ( .A(simpleXor_69_port_z), .B(simpleXor_68_port_z), .Z(n10) );
  XOR2_X1 U327 ( .A(n_zz_io_c_1_20_0_), .B(n9), .Z(io_c_1[5]) );
  XOR2_X1 U328 ( .A(simpleXor_75_port_z), .B(simpleXor_74_port_z), .Z(n9) );
  XOR2_X1 U329 ( .A(n_zz_io_c_1_24_0_), .B(n8), .Z(io_c_1[6]) );
  XOR2_X1 U330 ( .A(simpleXor_81_port_z), .B(simpleXor_80_port_z), .Z(n8) );
  XOR2_X1 U331 ( .A(n_zz_io_c_0_0_), .B(n21), .Z(io_c_0[0]) );
  XOR2_X1 U332 ( .A(simpleXor_43_port_z), .B(simpleXor_42_port_z), .Z(n21) );
  XOR2_X1 U333 ( .A(n_zz_io_c_0_4_0_), .B(n20), .Z(io_c_0[1]) );
  XOR2_X1 U334 ( .A(simpleXor_49_port_z), .B(simpleXor_48_port_z), .Z(n20) );
  XOR2_X1 U335 ( .A(n_zz_io_c_0_8_0_), .B(n19), .Z(io_c_0[2]) );
  XOR2_X1 U336 ( .A(simpleXor_55_port_z), .B(simpleXor_54_port_z), .Z(n19) );
  XOR2_X1 U337 ( .A(n_zz_io_c_0_12_0_), .B(n18), .Z(io_c_0[3]) );
  XOR2_X1 U338 ( .A(simpleXor_61_port_z), .B(simpleXor_60_port_z), .Z(n18) );
  XOR2_X1 U339 ( .A(n_zz_io_c_0_16_0_), .B(n17), .Z(io_c_0[4]) );
  XOR2_X1 U340 ( .A(simpleXor_67_port_z), .B(simpleXor_66_port_z), .Z(n17) );
  XOR2_X1 U341 ( .A(n_zz_io_c_0_20_0_), .B(n16), .Z(io_c_0[5]) );
  XOR2_X1 U342 ( .A(simpleXor_73_port_z), .B(simpleXor_72_port_z), .Z(n16) );
  XOR2_X1 U343 ( .A(n_zz_io_c_0_24_0_), .B(n15), .Z(io_c_0[6]) );
  XOR2_X1 U344 ( .A(simpleXor_79_port_z), .B(simpleXor_78_port_z), .Z(n15) );
  INV_X1 simpleNot_42_U1 ( .A(io_a_0[0]), .ZN(simpleNot_42_port_z) );
  INV_X1 simpleNot_43_U1 ( .A(io_a_0[0]), .ZN(simpleNot_43_port_z) );
  INV_X1 simpleNot_44_U1 ( .A(io_a_1[0]), .ZN(simpleNot_44_port_z) );
  INV_X1 simpleNot_45_U1 ( .A(io_a_1[0]), .ZN(simpleNot_45_port_z) );
  INV_X1 simpleNot_46_U1 ( .A(io_a_2[0]), .ZN(simpleNot_46_port_z) );
  INV_X1 simpleNot_47_U1 ( .A(io_a_2[0]), .ZN(simpleNot_47_port_z) );
  INV_X1 simpleNot_48_U1 ( .A(io_a_0[1]), .ZN(simpleNot_48_port_z) );
  INV_X1 simpleNot_49_U1 ( .A(io_a_0[1]), .ZN(simpleNot_49_port_z) );
  INV_X1 simpleNot_50_U1 ( .A(io_a_1[1]), .ZN(simpleNot_50_port_z) );
  INV_X1 simpleNot_51_U1 ( .A(io_a_1[1]), .ZN(simpleNot_51_port_z) );
  INV_X1 simpleNot_52_U1 ( .A(io_a_2[1]), .ZN(simpleNot_52_port_z) );
  INV_X1 simpleNot_53_U1 ( .A(io_a_2[1]), .ZN(simpleNot_53_port_z) );
  INV_X1 simpleNot_54_U1 ( .A(io_a_0[2]), .ZN(simpleNot_54_port_z) );
  INV_X1 simpleNot_55_U1 ( .A(io_a_0[2]), .ZN(simpleNot_55_port_z) );
  INV_X1 simpleNot_56_U1 ( .A(io_a_1[2]), .ZN(simpleNot_56_port_z) );
  INV_X1 simpleNot_57_U1 ( .A(io_a_1[2]), .ZN(simpleNot_57_port_z) );
  INV_X1 simpleNot_58_U1 ( .A(io_a_2[2]), .ZN(simpleNot_58_port_z) );
  INV_X1 simpleNot_59_U1 ( .A(io_a_2[2]), .ZN(simpleNot_59_port_z) );
  INV_X1 simpleNot_60_U1 ( .A(io_a_0[3]), .ZN(simpleNot_60_port_z) );
  INV_X1 simpleNot_61_U1 ( .A(io_a_0[3]), .ZN(simpleNot_61_port_z) );
  INV_X1 simpleNot_62_U1 ( .A(io_a_1[3]), .ZN(simpleNot_62_port_z) );
  INV_X1 simpleNot_63_U1 ( .A(io_a_1[3]), .ZN(simpleNot_63_port_z) );
  INV_X1 simpleNot_64_U1 ( .A(io_a_2[3]), .ZN(simpleNot_64_port_z) );
  INV_X1 simpleNot_65_U1 ( .A(io_a_2[3]), .ZN(simpleNot_65_port_z) );
  INV_X1 simpleNot_66_U1 ( .A(io_a_0[4]), .ZN(simpleNot_66_port_z) );
  INV_X1 simpleNot_67_U1 ( .A(io_a_0[4]), .ZN(simpleNot_67_port_z) );
  INV_X1 simpleNot_68_U1 ( .A(io_a_1[4]), .ZN(simpleNot_68_port_z) );
  INV_X1 simpleNot_69_U1 ( .A(io_a_1[4]), .ZN(simpleNot_69_port_z) );
  INV_X1 simpleNot_70_U1 ( .A(io_a_2[4]), .ZN(simpleNot_70_port_z) );
  INV_X1 simpleNot_71_U1 ( .A(io_a_2[4]), .ZN(simpleNot_71_port_z) );
  INV_X1 simpleNot_72_U1 ( .A(io_a_0[5]), .ZN(simpleNot_72_port_z) );
  INV_X1 simpleNot_73_U1 ( .A(io_a_0[5]), .ZN(simpleNot_73_port_z) );
  INV_X1 simpleNot_74_U1 ( .A(io_a_1[5]), .ZN(simpleNot_74_port_z) );
  INV_X1 simpleNot_75_U1 ( .A(io_a_1[5]), .ZN(simpleNot_75_port_z) );
  INV_X1 simpleNot_76_U1 ( .A(io_a_2[5]), .ZN(simpleNot_76_port_z) );
  INV_X1 simpleNot_77_U1 ( .A(io_a_2[5]), .ZN(simpleNot_77_port_z) );
  INV_X1 simpleNot_78_U1 ( .A(io_a_0[6]), .ZN(simpleNot_78_port_z) );
  INV_X1 simpleNot_79_U1 ( .A(io_a_0[6]), .ZN(simpleNot_79_port_z) );
  INV_X1 simpleNot_80_U1 ( .A(io_a_1[6]), .ZN(simpleNot_80_port_z) );
  INV_X1 simpleNot_81_U1 ( .A(io_a_1[6]), .ZN(simpleNot_81_port_z) );
  INV_X1 simpleNot_82_U1 ( .A(io_a_2[6]), .ZN(simpleNot_82_port_z) );
  INV_X1 simpleNot_83_U1 ( .A(io_a_2[6]), .ZN(simpleNot_83_port_z) );
  DFF_X1 cor_m_2_1_reg_0_ ( .D(cor_maj_77_port_o), .CK(clk), .Q(
        cor_port_v_2_1[0]), .QN() );
  DFF_X1 cor_m_2_1_reg_1_ ( .D(cor_maj_78_port_o), .CK(clk), .Q(
        cor_port_v_2_1[1]), .QN() );
  DFF_X1 cor_m_2_1_reg_2_ ( .D(cor_maj_79_port_o), .CK(clk), .Q(
        cor_port_v_2_1[2]), .QN() );
  DFF_X1 cor_m_2_1_reg_3_ ( .D(cor_maj_80_port_o), .CK(clk), .Q(
        cor_port_v_2_1[3]), .QN() );
  DFF_X1 cor_m_2_1_reg_4_ ( .D(cor_maj_81_port_o), .CK(clk), .Q(
        cor_port_v_2_1[4]), .QN() );
  DFF_X1 cor_m_2_1_reg_5_ ( .D(cor_maj_82_port_o), .CK(clk), .Q(
        cor_port_v_2_1[5]), .QN() );
  DFF_X1 cor_m_2_1_reg_6_ ( .D(cor_maj_83_port_o), .CK(clk), .Q(
        cor_port_v_2_1[6]), .QN() );
  DFF_X1 cor_m_2_0_reg_0_ ( .D(cor_maj_70_port_o), .CK(clk), .Q(
        cor_port_v_2_0[0]), .QN() );
  DFF_X1 cor_m_2_0_reg_1_ ( .D(cor_maj_71_port_o), .CK(clk), .Q(
        cor_port_v_2_0[1]), .QN() );
  DFF_X1 cor_m_2_0_reg_2_ ( .D(cor_maj_72_port_o), .CK(clk), .Q(
        cor_port_v_2_0[2]), .QN() );
  DFF_X1 cor_m_2_0_reg_3_ ( .D(cor_maj_73_port_o), .CK(clk), .Q(
        cor_port_v_2_0[3]), .QN() );
  DFF_X1 cor_m_2_0_reg_4_ ( .D(cor_maj_74_port_o), .CK(clk), .Q(
        cor_port_v_2_0[4]), .QN() );
  DFF_X1 cor_m_2_0_reg_5_ ( .D(cor_maj_75_port_o), .CK(clk), .Q(
        cor_port_v_2_0[5]), .QN() );
  DFF_X1 cor_m_2_0_reg_6_ ( .D(cor_maj_76_port_o), .CK(clk), .Q(
        cor_port_v_2_0[6]), .QN() );
  DFF_X1 cor_m_1_2_reg_0_ ( .D(cor_maj_63_port_o), .CK(clk), .Q(
        cor_port_v_1_2[0]), .QN() );
  DFF_X1 cor_m_1_2_reg_1_ ( .D(cor_maj_64_port_o), .CK(clk), .Q(
        cor_port_v_1_2[1]), .QN() );
  DFF_X1 cor_m_1_2_reg_2_ ( .D(cor_maj_65_port_o), .CK(clk), .Q(
        cor_port_v_1_2[2]), .QN() );
  DFF_X1 cor_m_1_2_reg_3_ ( .D(cor_maj_66_port_o), .CK(clk), .Q(
        cor_port_v_1_2[3]), .QN() );
  DFF_X1 cor_m_1_2_reg_4_ ( .D(cor_maj_67_port_o), .CK(clk), .Q(
        cor_port_v_1_2[4]), .QN() );
  DFF_X1 cor_m_1_2_reg_5_ ( .D(cor_maj_68_port_o), .CK(clk), .Q(
        cor_port_v_1_2[5]), .QN() );
  DFF_X1 cor_m_1_2_reg_6_ ( .D(cor_maj_69_port_o), .CK(clk), .Q(
        cor_port_v_1_2[6]), .QN() );
  DFF_X1 cor_m_1_0_reg_0_ ( .D(cor_maj_56_port_o), .CK(clk), .Q(
        cor_port_v_1_0[0]), .QN() );
  DFF_X1 cor_m_1_0_reg_1_ ( .D(cor_maj_57_port_o), .CK(clk), .Q(
        cor_port_v_1_0[1]), .QN() );
  DFF_X1 cor_m_1_0_reg_2_ ( .D(cor_maj_58_port_o), .CK(clk), .Q(
        cor_port_v_1_0[2]), .QN() );
  DFF_X1 cor_m_1_0_reg_3_ ( .D(cor_maj_59_port_o), .CK(clk), .Q(
        cor_port_v_1_0[3]), .QN() );
  DFF_X1 cor_m_1_0_reg_4_ ( .D(cor_maj_60_port_o), .CK(clk), .Q(
        cor_port_v_1_0[4]), .QN() );
  DFF_X1 cor_m_1_0_reg_5_ ( .D(cor_maj_61_port_o), .CK(clk), .Q(
        cor_port_v_1_0[5]), .QN() );
  DFF_X1 cor_m_1_0_reg_6_ ( .D(cor_maj_62_port_o), .CK(clk), .Q(
        cor_port_v_1_0[6]), .QN() );
  DFF_X1 cor_m_0_2_reg_0_ ( .D(cor_maj_49_port_o), .CK(clk), .Q(
        cor_port_v_0_2[0]), .QN() );
  DFF_X1 cor_m_0_2_reg_1_ ( .D(cor_maj_50_port_o), .CK(clk), .Q(
        cor_port_v_0_2[1]), .QN() );
  DFF_X1 cor_m_0_2_reg_2_ ( .D(cor_maj_51_port_o), .CK(clk), .Q(
        cor_port_v_0_2[2]), .QN() );
  DFF_X1 cor_m_0_2_reg_3_ ( .D(cor_maj_52_port_o), .CK(clk), .Q(
        cor_port_v_0_2[3]), .QN() );
  DFF_X1 cor_m_0_2_reg_4_ ( .D(cor_maj_53_port_o), .CK(clk), .Q(
        cor_port_v_0_2[4]), .QN() );
  DFF_X1 cor_m_0_2_reg_5_ ( .D(cor_maj_54_port_o), .CK(clk), .Q(
        cor_port_v_0_2[5]), .QN() );
  DFF_X1 cor_m_0_2_reg_6_ ( .D(cor_maj_55_port_o), .CK(clk), .Q(
        cor_port_v_0_2[6]), .QN() );
  DFF_X1 cor_m_0_1_reg_0_ ( .D(cor_maj_42_port_o), .CK(clk), .Q(
        cor_port_v_0_1[0]), .QN() );
  DFF_X1 cor_m_0_1_reg_1_ ( .D(cor_maj_43_port_o), .CK(clk), .Q(
        cor_port_v_0_1[1]), .QN() );
  DFF_X1 cor_m_0_1_reg_2_ ( .D(cor_maj_44_port_o), .CK(clk), .Q(
        cor_port_v_0_1[2]), .QN() );
  DFF_X1 cor_m_0_1_reg_3_ ( .D(cor_maj_45_port_o), .CK(clk), .Q(
        cor_port_v_0_1[3]), .QN() );
  DFF_X1 cor_m_0_1_reg_4_ ( .D(cor_maj_46_port_o), .CK(clk), .Q(
        cor_port_v_0_1[4]), .QN() );
  DFF_X1 cor_m_0_1_reg_5_ ( .D(cor_maj_47_port_o), .CK(clk), .Q(
        cor_port_v_0_1[5]), .QN() );
  DFF_X1 cor_m_0_1_reg_6_ ( .D(cor_maj_48_port_o), .CK(clk), .Q(
        cor_port_v_0_1[6]), .QN() );
  OR2_X1 cor_maj_42_U19 ( .A1(cor_maj_42_n8), .A2(cor_maj_42_n9), .ZN(
        cor_maj_42_n7) );
  NAND2_X1 cor_maj_42_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_42_n7), .ZN(
        cor_maj_42_n6) );
  NAND2_X1 cor_maj_42_U17 ( .A1(cor_maj_42_n9), .A2(cor_maj_42_n8), .ZN(
        cor_maj_42_n5) );
  NAND2_X1 cor_maj_42_U16 ( .A1(cor_maj_42_n5), .A2(cor_maj_42_n6), .ZN(
        cor_maj_42_n4) );
  NAND2_X1 cor_maj_42_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_42_n10), .ZN(
        cor_maj_42_n17) );
  NAND2_X1 cor_maj_42_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_42_n16) );
  NAND2_X1 cor_maj_42_U13 ( .A1(cor_maj_42_n16), .A2(cor_maj_42_n17), .ZN(
        cor_maj_42_n13) );
  NAND2_X1 cor_maj_42_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_42_n11), .ZN(
        cor_maj_42_n15) );
  NAND2_X1 cor_maj_42_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_42_n14) );
  NAND2_X1 cor_maj_42_U10 ( .A1(cor_maj_42_n14), .A2(cor_maj_42_n15), .ZN(
        cor_maj_42_n12) );
  XOR2_X1 cor_maj_42_U9 ( .A(v_1_0_1[2]), .B(cor_maj_42_n11), .Z(cor_maj_42_n9) );
  XOR2_X1 cor_maj_42_U8 ( .A(v_1_0_1[5]), .B(cor_maj_42_n10), .Z(cor_maj_42_n8) );
  XOR2_X1 cor_maj_42_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_42_n11)
         );
  XOR2_X1 cor_maj_42_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_42_n10)
         );
  OR2_X1 cor_maj_42_U5 ( .A1(cor_maj_42_n12), .A2(cor_maj_42_n13), .ZN(
        cor_maj_42_n3) );
  NAND2_X1 cor_maj_42_U4 ( .A1(cor_maj_42_n13), .A2(cor_maj_42_n12), .ZN(
        cor_maj_42_n1) );
  NAND2_X1 cor_maj_42_U3 ( .A1(cor_maj_42_n3), .A2(cor_maj_42_n4), .ZN(
        cor_maj_42_n2) );
  NAND2_X1 cor_maj_42_U2 ( .A1(cor_maj_42_n1), .A2(cor_maj_42_n2), .ZN(
        cor_maj_42_port_o) );
  OR2_X1 cor_maj_43_U19 ( .A1(cor_maj_43_n27), .A2(cor_maj_43_n26), .ZN(
        cor_maj_43_n28) );
  NAND2_X1 cor_maj_43_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_43_n28), .ZN(
        cor_maj_43_n29) );
  NAND2_X1 cor_maj_43_U17 ( .A1(cor_maj_43_n26), .A2(cor_maj_43_n27), .ZN(
        cor_maj_43_n30) );
  NAND2_X1 cor_maj_43_U16 ( .A1(cor_maj_43_n30), .A2(cor_maj_43_n29), .ZN(
        cor_maj_43_n31) );
  NAND2_X1 cor_maj_43_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_43_n25), .ZN(
        cor_maj_43_n18) );
  NAND2_X1 cor_maj_43_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_43_n19) );
  NAND2_X1 cor_maj_43_U13 ( .A1(cor_maj_43_n19), .A2(cor_maj_43_n18), .ZN(
        cor_maj_43_n22) );
  NAND2_X1 cor_maj_43_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_43_n24), .ZN(
        cor_maj_43_n20) );
  NAND2_X1 cor_maj_43_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_43_n21) );
  NAND2_X1 cor_maj_43_U10 ( .A1(cor_maj_43_n21), .A2(cor_maj_43_n20), .ZN(
        cor_maj_43_n23) );
  XOR2_X1 cor_maj_43_U9 ( .A(v_1_0_1[2]), .B(cor_maj_43_n24), .Z(
        cor_maj_43_n26) );
  XOR2_X1 cor_maj_43_U8 ( .A(v_1_0_1[5]), .B(cor_maj_43_n25), .Z(
        cor_maj_43_n27) );
  XOR2_X1 cor_maj_43_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_43_n24)
         );
  XOR2_X1 cor_maj_43_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_43_n25)
         );
  OR2_X1 cor_maj_43_U5 ( .A1(cor_maj_43_n23), .A2(cor_maj_43_n22), .ZN(
        cor_maj_43_n32) );
  NAND2_X1 cor_maj_43_U4 ( .A1(cor_maj_43_n22), .A2(cor_maj_43_n23), .ZN(
        cor_maj_43_n34) );
  NAND2_X1 cor_maj_43_U3 ( .A1(cor_maj_43_n32), .A2(cor_maj_43_n31), .ZN(
        cor_maj_43_n33) );
  NAND2_X1 cor_maj_43_U2 ( .A1(cor_maj_43_n34), .A2(cor_maj_43_n33), .ZN(
        cor_maj_43_port_o) );
  OR2_X1 cor_maj_44_U19 ( .A1(cor_maj_44_n27), .A2(cor_maj_44_n26), .ZN(
        cor_maj_44_n28) );
  NAND2_X1 cor_maj_44_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_44_n28), .ZN(
        cor_maj_44_n29) );
  NAND2_X1 cor_maj_44_U17 ( .A1(cor_maj_44_n26), .A2(cor_maj_44_n27), .ZN(
        cor_maj_44_n30) );
  NAND2_X1 cor_maj_44_U16 ( .A1(cor_maj_44_n30), .A2(cor_maj_44_n29), .ZN(
        cor_maj_44_n31) );
  NAND2_X1 cor_maj_44_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_44_n25), .ZN(
        cor_maj_44_n18) );
  NAND2_X1 cor_maj_44_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_44_n19) );
  NAND2_X1 cor_maj_44_U13 ( .A1(cor_maj_44_n19), .A2(cor_maj_44_n18), .ZN(
        cor_maj_44_n22) );
  NAND2_X1 cor_maj_44_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_44_n24), .ZN(
        cor_maj_44_n20) );
  NAND2_X1 cor_maj_44_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_44_n21) );
  NAND2_X1 cor_maj_44_U10 ( .A1(cor_maj_44_n21), .A2(cor_maj_44_n20), .ZN(
        cor_maj_44_n23) );
  XOR2_X1 cor_maj_44_U9 ( .A(v_1_0_1[2]), .B(cor_maj_44_n24), .Z(
        cor_maj_44_n26) );
  XOR2_X1 cor_maj_44_U8 ( .A(v_1_0_1[5]), .B(cor_maj_44_n25), .Z(
        cor_maj_44_n27) );
  XOR2_X1 cor_maj_44_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_44_n24)
         );
  XOR2_X1 cor_maj_44_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_44_n25)
         );
  OR2_X1 cor_maj_44_U5 ( .A1(cor_maj_44_n23), .A2(cor_maj_44_n22), .ZN(
        cor_maj_44_n32) );
  NAND2_X1 cor_maj_44_U4 ( .A1(cor_maj_44_n22), .A2(cor_maj_44_n23), .ZN(
        cor_maj_44_n34) );
  NAND2_X1 cor_maj_44_U3 ( .A1(cor_maj_44_n32), .A2(cor_maj_44_n31), .ZN(
        cor_maj_44_n33) );
  NAND2_X1 cor_maj_44_U2 ( .A1(cor_maj_44_n34), .A2(cor_maj_44_n33), .ZN(
        cor_maj_44_port_o) );
  OR2_X1 cor_maj_45_U19 ( .A1(cor_maj_45_n27), .A2(cor_maj_45_n26), .ZN(
        cor_maj_45_n28) );
  NAND2_X1 cor_maj_45_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_45_n28), .ZN(
        cor_maj_45_n29) );
  NAND2_X1 cor_maj_45_U17 ( .A1(cor_maj_45_n26), .A2(cor_maj_45_n27), .ZN(
        cor_maj_45_n30) );
  NAND2_X1 cor_maj_45_U16 ( .A1(cor_maj_45_n30), .A2(cor_maj_45_n29), .ZN(
        cor_maj_45_n31) );
  NAND2_X1 cor_maj_45_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_45_n25), .ZN(
        cor_maj_45_n18) );
  NAND2_X1 cor_maj_45_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_45_n19) );
  NAND2_X1 cor_maj_45_U13 ( .A1(cor_maj_45_n19), .A2(cor_maj_45_n18), .ZN(
        cor_maj_45_n22) );
  NAND2_X1 cor_maj_45_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_45_n24), .ZN(
        cor_maj_45_n20) );
  NAND2_X1 cor_maj_45_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_45_n21) );
  NAND2_X1 cor_maj_45_U10 ( .A1(cor_maj_45_n21), .A2(cor_maj_45_n20), .ZN(
        cor_maj_45_n23) );
  XOR2_X1 cor_maj_45_U9 ( .A(v_1_0_1[2]), .B(cor_maj_45_n24), .Z(
        cor_maj_45_n26) );
  XOR2_X1 cor_maj_45_U8 ( .A(v_1_0_1[5]), .B(cor_maj_45_n25), .Z(
        cor_maj_45_n27) );
  XOR2_X1 cor_maj_45_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_45_n24)
         );
  XOR2_X1 cor_maj_45_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_45_n25)
         );
  OR2_X1 cor_maj_45_U5 ( .A1(cor_maj_45_n23), .A2(cor_maj_45_n22), .ZN(
        cor_maj_45_n32) );
  NAND2_X1 cor_maj_45_U4 ( .A1(cor_maj_45_n22), .A2(cor_maj_45_n23), .ZN(
        cor_maj_45_n34) );
  NAND2_X1 cor_maj_45_U3 ( .A1(cor_maj_45_n32), .A2(cor_maj_45_n31), .ZN(
        cor_maj_45_n33) );
  NAND2_X1 cor_maj_45_U2 ( .A1(cor_maj_45_n34), .A2(cor_maj_45_n33), .ZN(
        cor_maj_45_port_o) );
  OR2_X1 cor_maj_46_U19 ( .A1(cor_maj_46_n27), .A2(cor_maj_46_n26), .ZN(
        cor_maj_46_n28) );
  NAND2_X1 cor_maj_46_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_46_n28), .ZN(
        cor_maj_46_n29) );
  NAND2_X1 cor_maj_46_U17 ( .A1(cor_maj_46_n26), .A2(cor_maj_46_n27), .ZN(
        cor_maj_46_n30) );
  NAND2_X1 cor_maj_46_U16 ( .A1(cor_maj_46_n30), .A2(cor_maj_46_n29), .ZN(
        cor_maj_46_n31) );
  NAND2_X1 cor_maj_46_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_46_n25), .ZN(
        cor_maj_46_n18) );
  NAND2_X1 cor_maj_46_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_46_n19) );
  NAND2_X1 cor_maj_46_U13 ( .A1(cor_maj_46_n19), .A2(cor_maj_46_n18), .ZN(
        cor_maj_46_n22) );
  NAND2_X1 cor_maj_46_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_46_n24), .ZN(
        cor_maj_46_n20) );
  NAND2_X1 cor_maj_46_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_46_n21) );
  NAND2_X1 cor_maj_46_U10 ( .A1(cor_maj_46_n21), .A2(cor_maj_46_n20), .ZN(
        cor_maj_46_n23) );
  XOR2_X1 cor_maj_46_U9 ( .A(v_1_0_1[2]), .B(cor_maj_46_n24), .Z(
        cor_maj_46_n26) );
  XOR2_X1 cor_maj_46_U8 ( .A(v_1_0_1[5]), .B(cor_maj_46_n25), .Z(
        cor_maj_46_n27) );
  XOR2_X1 cor_maj_46_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_46_n24)
         );
  XOR2_X1 cor_maj_46_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_46_n25)
         );
  OR2_X1 cor_maj_46_U5 ( .A1(cor_maj_46_n23), .A2(cor_maj_46_n22), .ZN(
        cor_maj_46_n32) );
  NAND2_X1 cor_maj_46_U4 ( .A1(cor_maj_46_n22), .A2(cor_maj_46_n23), .ZN(
        cor_maj_46_n34) );
  NAND2_X1 cor_maj_46_U3 ( .A1(cor_maj_46_n32), .A2(cor_maj_46_n31), .ZN(
        cor_maj_46_n33) );
  NAND2_X1 cor_maj_46_U2 ( .A1(cor_maj_46_n34), .A2(cor_maj_46_n33), .ZN(
        cor_maj_46_port_o) );
  OR2_X1 cor_maj_47_U19 ( .A1(cor_maj_47_n27), .A2(cor_maj_47_n26), .ZN(
        cor_maj_47_n28) );
  NAND2_X1 cor_maj_47_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_47_n28), .ZN(
        cor_maj_47_n29) );
  NAND2_X1 cor_maj_47_U17 ( .A1(cor_maj_47_n26), .A2(cor_maj_47_n27), .ZN(
        cor_maj_47_n30) );
  NAND2_X1 cor_maj_47_U16 ( .A1(cor_maj_47_n30), .A2(cor_maj_47_n29), .ZN(
        cor_maj_47_n31) );
  NAND2_X1 cor_maj_47_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_47_n25), .ZN(
        cor_maj_47_n18) );
  NAND2_X1 cor_maj_47_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_47_n19) );
  NAND2_X1 cor_maj_47_U13 ( .A1(cor_maj_47_n19), .A2(cor_maj_47_n18), .ZN(
        cor_maj_47_n22) );
  NAND2_X1 cor_maj_47_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_47_n24), .ZN(
        cor_maj_47_n20) );
  NAND2_X1 cor_maj_47_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_47_n21) );
  NAND2_X1 cor_maj_47_U10 ( .A1(cor_maj_47_n21), .A2(cor_maj_47_n20), .ZN(
        cor_maj_47_n23) );
  XOR2_X1 cor_maj_47_U9 ( .A(v_1_0_1[2]), .B(cor_maj_47_n24), .Z(
        cor_maj_47_n26) );
  XOR2_X1 cor_maj_47_U8 ( .A(v_1_0_1[5]), .B(cor_maj_47_n25), .Z(
        cor_maj_47_n27) );
  XOR2_X1 cor_maj_47_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_47_n24)
         );
  XOR2_X1 cor_maj_47_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_47_n25)
         );
  OR2_X1 cor_maj_47_U5 ( .A1(cor_maj_47_n23), .A2(cor_maj_47_n22), .ZN(
        cor_maj_47_n32) );
  NAND2_X1 cor_maj_47_U4 ( .A1(cor_maj_47_n22), .A2(cor_maj_47_n23), .ZN(
        cor_maj_47_n34) );
  NAND2_X1 cor_maj_47_U3 ( .A1(cor_maj_47_n32), .A2(cor_maj_47_n31), .ZN(
        cor_maj_47_n33) );
  NAND2_X1 cor_maj_47_U2 ( .A1(cor_maj_47_n34), .A2(cor_maj_47_n33), .ZN(
        cor_maj_47_port_o) );
  OR2_X1 cor_maj_48_U19 ( .A1(cor_maj_48_n27), .A2(cor_maj_48_n26), .ZN(
        cor_maj_48_n28) );
  NAND2_X1 cor_maj_48_U18 ( .A1(v_1_0_1[6]), .A2(cor_maj_48_n28), .ZN(
        cor_maj_48_n29) );
  NAND2_X1 cor_maj_48_U17 ( .A1(cor_maj_48_n26), .A2(cor_maj_48_n27), .ZN(
        cor_maj_48_n30) );
  NAND2_X1 cor_maj_48_U16 ( .A1(cor_maj_48_n30), .A2(cor_maj_48_n29), .ZN(
        cor_maj_48_n31) );
  NAND2_X1 cor_maj_48_U15 ( .A1(v_1_0_1[5]), .A2(cor_maj_48_n25), .ZN(
        cor_maj_48_n18) );
  NAND2_X1 cor_maj_48_U14 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_48_n19) );
  NAND2_X1 cor_maj_48_U13 ( .A1(cor_maj_48_n19), .A2(cor_maj_48_n18), .ZN(
        cor_maj_48_n22) );
  NAND2_X1 cor_maj_48_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_48_n24), .ZN(
        cor_maj_48_n20) );
  NAND2_X1 cor_maj_48_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_48_n21) );
  NAND2_X1 cor_maj_48_U10 ( .A1(cor_maj_48_n21), .A2(cor_maj_48_n20), .ZN(
        cor_maj_48_n23) );
  XOR2_X1 cor_maj_48_U9 ( .A(v_1_0_1[2]), .B(cor_maj_48_n24), .Z(
        cor_maj_48_n26) );
  XOR2_X1 cor_maj_48_U8 ( .A(v_1_0_1[5]), .B(cor_maj_48_n25), .Z(
        cor_maj_48_n27) );
  XOR2_X1 cor_maj_48_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_48_n24)
         );
  XOR2_X1 cor_maj_48_U6 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_48_n25)
         );
  OR2_X1 cor_maj_48_U5 ( .A1(cor_maj_48_n23), .A2(cor_maj_48_n22), .ZN(
        cor_maj_48_n32) );
  NAND2_X1 cor_maj_48_U4 ( .A1(cor_maj_48_n22), .A2(cor_maj_48_n23), .ZN(
        cor_maj_48_n34) );
  NAND2_X1 cor_maj_48_U3 ( .A1(cor_maj_48_n32), .A2(cor_maj_48_n31), .ZN(
        cor_maj_48_n33) );
  NAND2_X1 cor_maj_48_U2 ( .A1(cor_maj_48_n34), .A2(cor_maj_48_n33), .ZN(
        cor_maj_48_port_o) );
  OR2_X1 cor_maj_49_U19 ( .A1(cor_maj_49_n27), .A2(cor_maj_49_n26), .ZN(
        cor_maj_49_n28) );
  NAND2_X1 cor_maj_49_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_49_n28), .ZN(
        cor_maj_49_n29) );
  NAND2_X1 cor_maj_49_U17 ( .A1(cor_maj_49_n26), .A2(cor_maj_49_n27), .ZN(
        cor_maj_49_n30) );
  NAND2_X1 cor_maj_49_U16 ( .A1(cor_maj_49_n30), .A2(cor_maj_49_n29), .ZN(
        cor_maj_49_n31) );
  NAND2_X1 cor_maj_49_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_49_n25), .ZN(
        cor_maj_49_n18) );
  NAND2_X1 cor_maj_49_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_49_n19) );
  NAND2_X1 cor_maj_49_U13 ( .A1(cor_maj_49_n19), .A2(cor_maj_49_n18), .ZN(
        cor_maj_49_n22) );
  NAND2_X1 cor_maj_49_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_49_n24), .ZN(
        cor_maj_49_n20) );
  NAND2_X1 cor_maj_49_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_49_n21) );
  NAND2_X1 cor_maj_49_U10 ( .A1(cor_maj_49_n21), .A2(cor_maj_49_n20), .ZN(
        cor_maj_49_n23) );
  XOR2_X1 cor_maj_49_U9 ( .A(v_1_0_2[2]), .B(cor_maj_49_n24), .Z(
        cor_maj_49_n26) );
  XOR2_X1 cor_maj_49_U8 ( .A(v_1_0_2[5]), .B(cor_maj_49_n25), .Z(
        cor_maj_49_n27) );
  XOR2_X1 cor_maj_49_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_49_n24)
         );
  XOR2_X1 cor_maj_49_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_49_n25)
         );
  OR2_X1 cor_maj_49_U5 ( .A1(cor_maj_49_n23), .A2(cor_maj_49_n22), .ZN(
        cor_maj_49_n32) );
  NAND2_X1 cor_maj_49_U4 ( .A1(cor_maj_49_n22), .A2(cor_maj_49_n23), .ZN(
        cor_maj_49_n34) );
  NAND2_X1 cor_maj_49_U3 ( .A1(cor_maj_49_n32), .A2(cor_maj_49_n31), .ZN(
        cor_maj_49_n33) );
  NAND2_X1 cor_maj_49_U2 ( .A1(cor_maj_49_n34), .A2(cor_maj_49_n33), .ZN(
        cor_maj_49_port_o) );
  OR2_X1 cor_maj_50_U19 ( .A1(cor_maj_50_n27), .A2(cor_maj_50_n26), .ZN(
        cor_maj_50_n28) );
  NAND2_X1 cor_maj_50_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_50_n28), .ZN(
        cor_maj_50_n29) );
  NAND2_X1 cor_maj_50_U17 ( .A1(cor_maj_50_n26), .A2(cor_maj_50_n27), .ZN(
        cor_maj_50_n30) );
  NAND2_X1 cor_maj_50_U16 ( .A1(cor_maj_50_n30), .A2(cor_maj_50_n29), .ZN(
        cor_maj_50_n31) );
  NAND2_X1 cor_maj_50_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_50_n25), .ZN(
        cor_maj_50_n18) );
  NAND2_X1 cor_maj_50_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_50_n19) );
  NAND2_X1 cor_maj_50_U13 ( .A1(cor_maj_50_n19), .A2(cor_maj_50_n18), .ZN(
        cor_maj_50_n22) );
  NAND2_X1 cor_maj_50_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_50_n24), .ZN(
        cor_maj_50_n20) );
  NAND2_X1 cor_maj_50_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_50_n21) );
  NAND2_X1 cor_maj_50_U10 ( .A1(cor_maj_50_n21), .A2(cor_maj_50_n20), .ZN(
        cor_maj_50_n23) );
  XOR2_X1 cor_maj_50_U9 ( .A(v_1_0_2[2]), .B(cor_maj_50_n24), .Z(
        cor_maj_50_n26) );
  XOR2_X1 cor_maj_50_U8 ( .A(v_1_0_2[5]), .B(cor_maj_50_n25), .Z(
        cor_maj_50_n27) );
  XOR2_X1 cor_maj_50_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_50_n24)
         );
  XOR2_X1 cor_maj_50_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_50_n25)
         );
  OR2_X1 cor_maj_50_U5 ( .A1(cor_maj_50_n23), .A2(cor_maj_50_n22), .ZN(
        cor_maj_50_n32) );
  NAND2_X1 cor_maj_50_U4 ( .A1(cor_maj_50_n22), .A2(cor_maj_50_n23), .ZN(
        cor_maj_50_n34) );
  NAND2_X1 cor_maj_50_U3 ( .A1(cor_maj_50_n32), .A2(cor_maj_50_n31), .ZN(
        cor_maj_50_n33) );
  NAND2_X1 cor_maj_50_U2 ( .A1(cor_maj_50_n34), .A2(cor_maj_50_n33), .ZN(
        cor_maj_50_port_o) );
  OR2_X1 cor_maj_51_U19 ( .A1(cor_maj_51_n27), .A2(cor_maj_51_n26), .ZN(
        cor_maj_51_n28) );
  NAND2_X1 cor_maj_51_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_51_n28), .ZN(
        cor_maj_51_n29) );
  NAND2_X1 cor_maj_51_U17 ( .A1(cor_maj_51_n26), .A2(cor_maj_51_n27), .ZN(
        cor_maj_51_n30) );
  NAND2_X1 cor_maj_51_U16 ( .A1(cor_maj_51_n30), .A2(cor_maj_51_n29), .ZN(
        cor_maj_51_n31) );
  NAND2_X1 cor_maj_51_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_51_n25), .ZN(
        cor_maj_51_n18) );
  NAND2_X1 cor_maj_51_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_51_n19) );
  NAND2_X1 cor_maj_51_U13 ( .A1(cor_maj_51_n19), .A2(cor_maj_51_n18), .ZN(
        cor_maj_51_n22) );
  NAND2_X1 cor_maj_51_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_51_n24), .ZN(
        cor_maj_51_n20) );
  NAND2_X1 cor_maj_51_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_51_n21) );
  NAND2_X1 cor_maj_51_U10 ( .A1(cor_maj_51_n21), .A2(cor_maj_51_n20), .ZN(
        cor_maj_51_n23) );
  XOR2_X1 cor_maj_51_U9 ( .A(v_1_0_2[2]), .B(cor_maj_51_n24), .Z(
        cor_maj_51_n26) );
  XOR2_X1 cor_maj_51_U8 ( .A(v_1_0_2[5]), .B(cor_maj_51_n25), .Z(
        cor_maj_51_n27) );
  XOR2_X1 cor_maj_51_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_51_n24)
         );
  XOR2_X1 cor_maj_51_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_51_n25)
         );
  OR2_X1 cor_maj_51_U5 ( .A1(cor_maj_51_n23), .A2(cor_maj_51_n22), .ZN(
        cor_maj_51_n32) );
  NAND2_X1 cor_maj_51_U4 ( .A1(cor_maj_51_n22), .A2(cor_maj_51_n23), .ZN(
        cor_maj_51_n34) );
  NAND2_X1 cor_maj_51_U3 ( .A1(cor_maj_51_n32), .A2(cor_maj_51_n31), .ZN(
        cor_maj_51_n33) );
  NAND2_X1 cor_maj_51_U2 ( .A1(cor_maj_51_n34), .A2(cor_maj_51_n33), .ZN(
        cor_maj_51_port_o) );
  OR2_X1 cor_maj_52_U19 ( .A1(cor_maj_52_n27), .A2(cor_maj_52_n26), .ZN(
        cor_maj_52_n28) );
  NAND2_X1 cor_maj_52_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_52_n28), .ZN(
        cor_maj_52_n29) );
  NAND2_X1 cor_maj_52_U17 ( .A1(cor_maj_52_n26), .A2(cor_maj_52_n27), .ZN(
        cor_maj_52_n30) );
  NAND2_X1 cor_maj_52_U16 ( .A1(cor_maj_52_n30), .A2(cor_maj_52_n29), .ZN(
        cor_maj_52_n31) );
  NAND2_X1 cor_maj_52_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_52_n25), .ZN(
        cor_maj_52_n18) );
  NAND2_X1 cor_maj_52_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_52_n19) );
  NAND2_X1 cor_maj_52_U13 ( .A1(cor_maj_52_n19), .A2(cor_maj_52_n18), .ZN(
        cor_maj_52_n22) );
  NAND2_X1 cor_maj_52_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_52_n24), .ZN(
        cor_maj_52_n20) );
  NAND2_X1 cor_maj_52_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_52_n21) );
  NAND2_X1 cor_maj_52_U10 ( .A1(cor_maj_52_n21), .A2(cor_maj_52_n20), .ZN(
        cor_maj_52_n23) );
  XOR2_X1 cor_maj_52_U9 ( .A(v_1_0_2[2]), .B(cor_maj_52_n24), .Z(
        cor_maj_52_n26) );
  XOR2_X1 cor_maj_52_U8 ( .A(v_1_0_2[5]), .B(cor_maj_52_n25), .Z(
        cor_maj_52_n27) );
  XOR2_X1 cor_maj_52_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_52_n24)
         );
  XOR2_X1 cor_maj_52_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_52_n25)
         );
  OR2_X1 cor_maj_52_U5 ( .A1(cor_maj_52_n23), .A2(cor_maj_52_n22), .ZN(
        cor_maj_52_n32) );
  NAND2_X1 cor_maj_52_U4 ( .A1(cor_maj_52_n22), .A2(cor_maj_52_n23), .ZN(
        cor_maj_52_n34) );
  NAND2_X1 cor_maj_52_U3 ( .A1(cor_maj_52_n32), .A2(cor_maj_52_n31), .ZN(
        cor_maj_52_n33) );
  NAND2_X1 cor_maj_52_U2 ( .A1(cor_maj_52_n34), .A2(cor_maj_52_n33), .ZN(
        cor_maj_52_port_o) );
  OR2_X1 cor_maj_53_U19 ( .A1(cor_maj_53_n27), .A2(cor_maj_53_n26), .ZN(
        cor_maj_53_n28) );
  NAND2_X1 cor_maj_53_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_53_n28), .ZN(
        cor_maj_53_n29) );
  NAND2_X1 cor_maj_53_U17 ( .A1(cor_maj_53_n26), .A2(cor_maj_53_n27), .ZN(
        cor_maj_53_n30) );
  NAND2_X1 cor_maj_53_U16 ( .A1(cor_maj_53_n30), .A2(cor_maj_53_n29), .ZN(
        cor_maj_53_n31) );
  NAND2_X1 cor_maj_53_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_53_n25), .ZN(
        cor_maj_53_n18) );
  NAND2_X1 cor_maj_53_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_53_n19) );
  NAND2_X1 cor_maj_53_U13 ( .A1(cor_maj_53_n19), .A2(cor_maj_53_n18), .ZN(
        cor_maj_53_n22) );
  NAND2_X1 cor_maj_53_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_53_n24), .ZN(
        cor_maj_53_n20) );
  NAND2_X1 cor_maj_53_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_53_n21) );
  NAND2_X1 cor_maj_53_U10 ( .A1(cor_maj_53_n21), .A2(cor_maj_53_n20), .ZN(
        cor_maj_53_n23) );
  XOR2_X1 cor_maj_53_U9 ( .A(v_1_0_2[2]), .B(cor_maj_53_n24), .Z(
        cor_maj_53_n26) );
  XOR2_X1 cor_maj_53_U8 ( .A(v_1_0_2[5]), .B(cor_maj_53_n25), .Z(
        cor_maj_53_n27) );
  XOR2_X1 cor_maj_53_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_53_n24)
         );
  XOR2_X1 cor_maj_53_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_53_n25)
         );
  OR2_X1 cor_maj_53_U5 ( .A1(cor_maj_53_n23), .A2(cor_maj_53_n22), .ZN(
        cor_maj_53_n32) );
  NAND2_X1 cor_maj_53_U4 ( .A1(cor_maj_53_n22), .A2(cor_maj_53_n23), .ZN(
        cor_maj_53_n34) );
  NAND2_X1 cor_maj_53_U3 ( .A1(cor_maj_53_n32), .A2(cor_maj_53_n31), .ZN(
        cor_maj_53_n33) );
  NAND2_X1 cor_maj_53_U2 ( .A1(cor_maj_53_n34), .A2(cor_maj_53_n33), .ZN(
        cor_maj_53_port_o) );
  OR2_X1 cor_maj_54_U19 ( .A1(cor_maj_54_n27), .A2(cor_maj_54_n26), .ZN(
        cor_maj_54_n28) );
  NAND2_X1 cor_maj_54_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_54_n28), .ZN(
        cor_maj_54_n29) );
  NAND2_X1 cor_maj_54_U17 ( .A1(cor_maj_54_n26), .A2(cor_maj_54_n27), .ZN(
        cor_maj_54_n30) );
  NAND2_X1 cor_maj_54_U16 ( .A1(cor_maj_54_n30), .A2(cor_maj_54_n29), .ZN(
        cor_maj_54_n31) );
  NAND2_X1 cor_maj_54_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_54_n25), .ZN(
        cor_maj_54_n18) );
  NAND2_X1 cor_maj_54_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_54_n19) );
  NAND2_X1 cor_maj_54_U13 ( .A1(cor_maj_54_n19), .A2(cor_maj_54_n18), .ZN(
        cor_maj_54_n22) );
  NAND2_X1 cor_maj_54_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_54_n24), .ZN(
        cor_maj_54_n20) );
  NAND2_X1 cor_maj_54_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_54_n21) );
  NAND2_X1 cor_maj_54_U10 ( .A1(cor_maj_54_n21), .A2(cor_maj_54_n20), .ZN(
        cor_maj_54_n23) );
  XOR2_X1 cor_maj_54_U9 ( .A(v_1_0_2[2]), .B(cor_maj_54_n24), .Z(
        cor_maj_54_n26) );
  XOR2_X1 cor_maj_54_U8 ( .A(v_1_0_2[5]), .B(cor_maj_54_n25), .Z(
        cor_maj_54_n27) );
  XOR2_X1 cor_maj_54_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_54_n24)
         );
  XOR2_X1 cor_maj_54_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_54_n25)
         );
  OR2_X1 cor_maj_54_U5 ( .A1(cor_maj_54_n23), .A2(cor_maj_54_n22), .ZN(
        cor_maj_54_n32) );
  NAND2_X1 cor_maj_54_U4 ( .A1(cor_maj_54_n22), .A2(cor_maj_54_n23), .ZN(
        cor_maj_54_n34) );
  NAND2_X1 cor_maj_54_U3 ( .A1(cor_maj_54_n32), .A2(cor_maj_54_n31), .ZN(
        cor_maj_54_n33) );
  NAND2_X1 cor_maj_54_U2 ( .A1(cor_maj_54_n34), .A2(cor_maj_54_n33), .ZN(
        cor_maj_54_port_o) );
  OR2_X1 cor_maj_55_U19 ( .A1(cor_maj_55_n27), .A2(cor_maj_55_n26), .ZN(
        cor_maj_55_n28) );
  NAND2_X1 cor_maj_55_U18 ( .A1(v_1_0_2[6]), .A2(cor_maj_55_n28), .ZN(
        cor_maj_55_n29) );
  NAND2_X1 cor_maj_55_U17 ( .A1(cor_maj_55_n26), .A2(cor_maj_55_n27), .ZN(
        cor_maj_55_n30) );
  NAND2_X1 cor_maj_55_U16 ( .A1(cor_maj_55_n30), .A2(cor_maj_55_n29), .ZN(
        cor_maj_55_n31) );
  NAND2_X1 cor_maj_55_U15 ( .A1(v_1_0_2[5]), .A2(cor_maj_55_n25), .ZN(
        cor_maj_55_n18) );
  NAND2_X1 cor_maj_55_U14 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_55_n19) );
  NAND2_X1 cor_maj_55_U13 ( .A1(cor_maj_55_n19), .A2(cor_maj_55_n18), .ZN(
        cor_maj_55_n22) );
  NAND2_X1 cor_maj_55_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_55_n24), .ZN(
        cor_maj_55_n20) );
  NAND2_X1 cor_maj_55_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_55_n21) );
  NAND2_X1 cor_maj_55_U10 ( .A1(cor_maj_55_n21), .A2(cor_maj_55_n20), .ZN(
        cor_maj_55_n23) );
  XOR2_X1 cor_maj_55_U9 ( .A(v_1_0_2[2]), .B(cor_maj_55_n24), .Z(
        cor_maj_55_n26) );
  XOR2_X1 cor_maj_55_U8 ( .A(v_1_0_2[5]), .B(cor_maj_55_n25), .Z(
        cor_maj_55_n27) );
  XOR2_X1 cor_maj_55_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_55_n24)
         );
  XOR2_X1 cor_maj_55_U6 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_55_n25)
         );
  OR2_X1 cor_maj_55_U5 ( .A1(cor_maj_55_n23), .A2(cor_maj_55_n22), .ZN(
        cor_maj_55_n32) );
  NAND2_X1 cor_maj_55_U4 ( .A1(cor_maj_55_n22), .A2(cor_maj_55_n23), .ZN(
        cor_maj_55_n34) );
  NAND2_X1 cor_maj_55_U3 ( .A1(cor_maj_55_n32), .A2(cor_maj_55_n31), .ZN(
        cor_maj_55_n33) );
  NAND2_X1 cor_maj_55_U2 ( .A1(cor_maj_55_n34), .A2(cor_maj_55_n33), .ZN(
        cor_maj_55_port_o) );
  OR2_X1 cor_maj_56_U19 ( .A1(cor_maj_56_n27), .A2(cor_maj_56_n26), .ZN(
        cor_maj_56_n28) );
  NAND2_X1 cor_maj_56_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_56_n28), .ZN(
        cor_maj_56_n29) );
  NAND2_X1 cor_maj_56_U17 ( .A1(cor_maj_56_n26), .A2(cor_maj_56_n27), .ZN(
        cor_maj_56_n30) );
  NAND2_X1 cor_maj_56_U16 ( .A1(cor_maj_56_n30), .A2(cor_maj_56_n29), .ZN(
        cor_maj_56_n31) );
  NAND2_X1 cor_maj_56_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_56_n25), .ZN(
        cor_maj_56_n18) );
  NAND2_X1 cor_maj_56_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_56_n19) );
  NAND2_X1 cor_maj_56_U13 ( .A1(cor_maj_56_n19), .A2(cor_maj_56_n18), .ZN(
        cor_maj_56_n22) );
  NAND2_X1 cor_maj_56_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_56_n24), .ZN(
        cor_maj_56_n20) );
  NAND2_X1 cor_maj_56_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_56_n21) );
  NAND2_X1 cor_maj_56_U10 ( .A1(cor_maj_56_n21), .A2(cor_maj_56_n20), .ZN(
        cor_maj_56_n23) );
  XOR2_X1 cor_maj_56_U9 ( .A(v_1_1_0[2]), .B(cor_maj_56_n24), .Z(
        cor_maj_56_n26) );
  XOR2_X1 cor_maj_56_U8 ( .A(v_1_1_0[5]), .B(cor_maj_56_n25), .Z(
        cor_maj_56_n27) );
  XOR2_X1 cor_maj_56_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_56_n24)
         );
  XOR2_X1 cor_maj_56_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_56_n25)
         );
  OR2_X1 cor_maj_56_U5 ( .A1(cor_maj_56_n23), .A2(cor_maj_56_n22), .ZN(
        cor_maj_56_n32) );
  NAND2_X1 cor_maj_56_U4 ( .A1(cor_maj_56_n22), .A2(cor_maj_56_n23), .ZN(
        cor_maj_56_n34) );
  NAND2_X1 cor_maj_56_U3 ( .A1(cor_maj_56_n32), .A2(cor_maj_56_n31), .ZN(
        cor_maj_56_n33) );
  NAND2_X1 cor_maj_56_U2 ( .A1(cor_maj_56_n34), .A2(cor_maj_56_n33), .ZN(
        cor_maj_56_port_o) );
  OR2_X1 cor_maj_57_U19 ( .A1(cor_maj_57_n27), .A2(cor_maj_57_n26), .ZN(
        cor_maj_57_n28) );
  NAND2_X1 cor_maj_57_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_57_n28), .ZN(
        cor_maj_57_n29) );
  NAND2_X1 cor_maj_57_U17 ( .A1(cor_maj_57_n26), .A2(cor_maj_57_n27), .ZN(
        cor_maj_57_n30) );
  NAND2_X1 cor_maj_57_U16 ( .A1(cor_maj_57_n30), .A2(cor_maj_57_n29), .ZN(
        cor_maj_57_n31) );
  NAND2_X1 cor_maj_57_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_57_n25), .ZN(
        cor_maj_57_n18) );
  NAND2_X1 cor_maj_57_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_57_n19) );
  NAND2_X1 cor_maj_57_U13 ( .A1(cor_maj_57_n19), .A2(cor_maj_57_n18), .ZN(
        cor_maj_57_n22) );
  NAND2_X1 cor_maj_57_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_57_n24), .ZN(
        cor_maj_57_n20) );
  NAND2_X1 cor_maj_57_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_57_n21) );
  NAND2_X1 cor_maj_57_U10 ( .A1(cor_maj_57_n21), .A2(cor_maj_57_n20), .ZN(
        cor_maj_57_n23) );
  XOR2_X1 cor_maj_57_U9 ( .A(v_1_1_0[2]), .B(cor_maj_57_n24), .Z(
        cor_maj_57_n26) );
  XOR2_X1 cor_maj_57_U8 ( .A(v_1_1_0[5]), .B(cor_maj_57_n25), .Z(
        cor_maj_57_n27) );
  XOR2_X1 cor_maj_57_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_57_n24)
         );
  XOR2_X1 cor_maj_57_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_57_n25)
         );
  OR2_X1 cor_maj_57_U5 ( .A1(cor_maj_57_n23), .A2(cor_maj_57_n22), .ZN(
        cor_maj_57_n32) );
  NAND2_X1 cor_maj_57_U4 ( .A1(cor_maj_57_n22), .A2(cor_maj_57_n23), .ZN(
        cor_maj_57_n34) );
  NAND2_X1 cor_maj_57_U3 ( .A1(cor_maj_57_n32), .A2(cor_maj_57_n31), .ZN(
        cor_maj_57_n33) );
  NAND2_X1 cor_maj_57_U2 ( .A1(cor_maj_57_n34), .A2(cor_maj_57_n33), .ZN(
        cor_maj_57_port_o) );
  OR2_X1 cor_maj_58_U19 ( .A1(cor_maj_58_n27), .A2(cor_maj_58_n26), .ZN(
        cor_maj_58_n28) );
  NAND2_X1 cor_maj_58_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_58_n28), .ZN(
        cor_maj_58_n29) );
  NAND2_X1 cor_maj_58_U17 ( .A1(cor_maj_58_n26), .A2(cor_maj_58_n27), .ZN(
        cor_maj_58_n30) );
  NAND2_X1 cor_maj_58_U16 ( .A1(cor_maj_58_n30), .A2(cor_maj_58_n29), .ZN(
        cor_maj_58_n31) );
  NAND2_X1 cor_maj_58_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_58_n25), .ZN(
        cor_maj_58_n18) );
  NAND2_X1 cor_maj_58_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_58_n19) );
  NAND2_X1 cor_maj_58_U13 ( .A1(cor_maj_58_n19), .A2(cor_maj_58_n18), .ZN(
        cor_maj_58_n22) );
  NAND2_X1 cor_maj_58_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_58_n24), .ZN(
        cor_maj_58_n20) );
  NAND2_X1 cor_maj_58_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_58_n21) );
  NAND2_X1 cor_maj_58_U10 ( .A1(cor_maj_58_n21), .A2(cor_maj_58_n20), .ZN(
        cor_maj_58_n23) );
  XOR2_X1 cor_maj_58_U9 ( .A(v_1_1_0[2]), .B(cor_maj_58_n24), .Z(
        cor_maj_58_n26) );
  XOR2_X1 cor_maj_58_U8 ( .A(v_1_1_0[5]), .B(cor_maj_58_n25), .Z(
        cor_maj_58_n27) );
  XOR2_X1 cor_maj_58_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_58_n24)
         );
  XOR2_X1 cor_maj_58_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_58_n25)
         );
  OR2_X1 cor_maj_58_U5 ( .A1(cor_maj_58_n23), .A2(cor_maj_58_n22), .ZN(
        cor_maj_58_n32) );
  NAND2_X1 cor_maj_58_U4 ( .A1(cor_maj_58_n22), .A2(cor_maj_58_n23), .ZN(
        cor_maj_58_n34) );
  NAND2_X1 cor_maj_58_U3 ( .A1(cor_maj_58_n32), .A2(cor_maj_58_n31), .ZN(
        cor_maj_58_n33) );
  NAND2_X1 cor_maj_58_U2 ( .A1(cor_maj_58_n34), .A2(cor_maj_58_n33), .ZN(
        cor_maj_58_port_o) );
  OR2_X1 cor_maj_59_U19 ( .A1(cor_maj_59_n27), .A2(cor_maj_59_n26), .ZN(
        cor_maj_59_n28) );
  NAND2_X1 cor_maj_59_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_59_n28), .ZN(
        cor_maj_59_n29) );
  NAND2_X1 cor_maj_59_U17 ( .A1(cor_maj_59_n26), .A2(cor_maj_59_n27), .ZN(
        cor_maj_59_n30) );
  NAND2_X1 cor_maj_59_U16 ( .A1(cor_maj_59_n30), .A2(cor_maj_59_n29), .ZN(
        cor_maj_59_n31) );
  NAND2_X1 cor_maj_59_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_59_n25), .ZN(
        cor_maj_59_n18) );
  NAND2_X1 cor_maj_59_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_59_n19) );
  NAND2_X1 cor_maj_59_U13 ( .A1(cor_maj_59_n19), .A2(cor_maj_59_n18), .ZN(
        cor_maj_59_n22) );
  NAND2_X1 cor_maj_59_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_59_n24), .ZN(
        cor_maj_59_n20) );
  NAND2_X1 cor_maj_59_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_59_n21) );
  NAND2_X1 cor_maj_59_U10 ( .A1(cor_maj_59_n21), .A2(cor_maj_59_n20), .ZN(
        cor_maj_59_n23) );
  XOR2_X1 cor_maj_59_U9 ( .A(v_1_1_0[2]), .B(cor_maj_59_n24), .Z(
        cor_maj_59_n26) );
  XOR2_X1 cor_maj_59_U8 ( .A(v_1_1_0[5]), .B(cor_maj_59_n25), .Z(
        cor_maj_59_n27) );
  XOR2_X1 cor_maj_59_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_59_n24)
         );
  XOR2_X1 cor_maj_59_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_59_n25)
         );
  OR2_X1 cor_maj_59_U5 ( .A1(cor_maj_59_n23), .A2(cor_maj_59_n22), .ZN(
        cor_maj_59_n32) );
  NAND2_X1 cor_maj_59_U4 ( .A1(cor_maj_59_n22), .A2(cor_maj_59_n23), .ZN(
        cor_maj_59_n34) );
  NAND2_X1 cor_maj_59_U3 ( .A1(cor_maj_59_n32), .A2(cor_maj_59_n31), .ZN(
        cor_maj_59_n33) );
  NAND2_X1 cor_maj_59_U2 ( .A1(cor_maj_59_n34), .A2(cor_maj_59_n33), .ZN(
        cor_maj_59_port_o) );
  OR2_X1 cor_maj_60_U19 ( .A1(cor_maj_60_n27), .A2(cor_maj_60_n26), .ZN(
        cor_maj_60_n28) );
  NAND2_X1 cor_maj_60_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_60_n28), .ZN(
        cor_maj_60_n29) );
  NAND2_X1 cor_maj_60_U17 ( .A1(cor_maj_60_n26), .A2(cor_maj_60_n27), .ZN(
        cor_maj_60_n30) );
  NAND2_X1 cor_maj_60_U16 ( .A1(cor_maj_60_n30), .A2(cor_maj_60_n29), .ZN(
        cor_maj_60_n31) );
  NAND2_X1 cor_maj_60_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_60_n25), .ZN(
        cor_maj_60_n18) );
  NAND2_X1 cor_maj_60_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_60_n19) );
  NAND2_X1 cor_maj_60_U13 ( .A1(cor_maj_60_n19), .A2(cor_maj_60_n18), .ZN(
        cor_maj_60_n22) );
  NAND2_X1 cor_maj_60_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_60_n24), .ZN(
        cor_maj_60_n20) );
  NAND2_X1 cor_maj_60_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_60_n21) );
  NAND2_X1 cor_maj_60_U10 ( .A1(cor_maj_60_n21), .A2(cor_maj_60_n20), .ZN(
        cor_maj_60_n23) );
  XOR2_X1 cor_maj_60_U9 ( .A(v_1_1_0[2]), .B(cor_maj_60_n24), .Z(
        cor_maj_60_n26) );
  XOR2_X1 cor_maj_60_U8 ( .A(v_1_1_0[5]), .B(cor_maj_60_n25), .Z(
        cor_maj_60_n27) );
  XOR2_X1 cor_maj_60_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_60_n24)
         );
  XOR2_X1 cor_maj_60_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_60_n25)
         );
  OR2_X1 cor_maj_60_U5 ( .A1(cor_maj_60_n23), .A2(cor_maj_60_n22), .ZN(
        cor_maj_60_n32) );
  NAND2_X1 cor_maj_60_U4 ( .A1(cor_maj_60_n22), .A2(cor_maj_60_n23), .ZN(
        cor_maj_60_n34) );
  NAND2_X1 cor_maj_60_U3 ( .A1(cor_maj_60_n32), .A2(cor_maj_60_n31), .ZN(
        cor_maj_60_n33) );
  NAND2_X1 cor_maj_60_U2 ( .A1(cor_maj_60_n34), .A2(cor_maj_60_n33), .ZN(
        cor_maj_60_port_o) );
  OR2_X1 cor_maj_61_U19 ( .A1(cor_maj_61_n27), .A2(cor_maj_61_n26), .ZN(
        cor_maj_61_n28) );
  NAND2_X1 cor_maj_61_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_61_n28), .ZN(
        cor_maj_61_n29) );
  NAND2_X1 cor_maj_61_U17 ( .A1(cor_maj_61_n26), .A2(cor_maj_61_n27), .ZN(
        cor_maj_61_n30) );
  NAND2_X1 cor_maj_61_U16 ( .A1(cor_maj_61_n30), .A2(cor_maj_61_n29), .ZN(
        cor_maj_61_n31) );
  NAND2_X1 cor_maj_61_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_61_n25), .ZN(
        cor_maj_61_n18) );
  NAND2_X1 cor_maj_61_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_61_n19) );
  NAND2_X1 cor_maj_61_U13 ( .A1(cor_maj_61_n19), .A2(cor_maj_61_n18), .ZN(
        cor_maj_61_n22) );
  NAND2_X1 cor_maj_61_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_61_n24), .ZN(
        cor_maj_61_n20) );
  NAND2_X1 cor_maj_61_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_61_n21) );
  NAND2_X1 cor_maj_61_U10 ( .A1(cor_maj_61_n21), .A2(cor_maj_61_n20), .ZN(
        cor_maj_61_n23) );
  XOR2_X1 cor_maj_61_U9 ( .A(v_1_1_0[2]), .B(cor_maj_61_n24), .Z(
        cor_maj_61_n26) );
  XOR2_X1 cor_maj_61_U8 ( .A(v_1_1_0[5]), .B(cor_maj_61_n25), .Z(
        cor_maj_61_n27) );
  XOR2_X1 cor_maj_61_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_61_n24)
         );
  XOR2_X1 cor_maj_61_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_61_n25)
         );
  OR2_X1 cor_maj_61_U5 ( .A1(cor_maj_61_n23), .A2(cor_maj_61_n22), .ZN(
        cor_maj_61_n32) );
  NAND2_X1 cor_maj_61_U4 ( .A1(cor_maj_61_n22), .A2(cor_maj_61_n23), .ZN(
        cor_maj_61_n34) );
  NAND2_X1 cor_maj_61_U3 ( .A1(cor_maj_61_n32), .A2(cor_maj_61_n31), .ZN(
        cor_maj_61_n33) );
  NAND2_X1 cor_maj_61_U2 ( .A1(cor_maj_61_n34), .A2(cor_maj_61_n33), .ZN(
        cor_maj_61_port_o) );
  OR2_X1 cor_maj_62_U19 ( .A1(cor_maj_62_n27), .A2(cor_maj_62_n26), .ZN(
        cor_maj_62_n28) );
  NAND2_X1 cor_maj_62_U18 ( .A1(v_1_1_0[6]), .A2(cor_maj_62_n28), .ZN(
        cor_maj_62_n29) );
  NAND2_X1 cor_maj_62_U17 ( .A1(cor_maj_62_n26), .A2(cor_maj_62_n27), .ZN(
        cor_maj_62_n30) );
  NAND2_X1 cor_maj_62_U16 ( .A1(cor_maj_62_n30), .A2(cor_maj_62_n29), .ZN(
        cor_maj_62_n31) );
  NAND2_X1 cor_maj_62_U15 ( .A1(v_1_1_0[5]), .A2(cor_maj_62_n25), .ZN(
        cor_maj_62_n18) );
  NAND2_X1 cor_maj_62_U14 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_62_n19) );
  NAND2_X1 cor_maj_62_U13 ( .A1(cor_maj_62_n19), .A2(cor_maj_62_n18), .ZN(
        cor_maj_62_n22) );
  NAND2_X1 cor_maj_62_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_62_n24), .ZN(
        cor_maj_62_n20) );
  NAND2_X1 cor_maj_62_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_62_n21) );
  NAND2_X1 cor_maj_62_U10 ( .A1(cor_maj_62_n21), .A2(cor_maj_62_n20), .ZN(
        cor_maj_62_n23) );
  XOR2_X1 cor_maj_62_U9 ( .A(v_1_1_0[2]), .B(cor_maj_62_n24), .Z(
        cor_maj_62_n26) );
  XOR2_X1 cor_maj_62_U8 ( .A(v_1_1_0[5]), .B(cor_maj_62_n25), .Z(
        cor_maj_62_n27) );
  XOR2_X1 cor_maj_62_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_62_n24)
         );
  XOR2_X1 cor_maj_62_U6 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_62_n25)
         );
  OR2_X1 cor_maj_62_U5 ( .A1(cor_maj_62_n23), .A2(cor_maj_62_n22), .ZN(
        cor_maj_62_n32) );
  NAND2_X1 cor_maj_62_U4 ( .A1(cor_maj_62_n22), .A2(cor_maj_62_n23), .ZN(
        cor_maj_62_n34) );
  NAND2_X1 cor_maj_62_U3 ( .A1(cor_maj_62_n32), .A2(cor_maj_62_n31), .ZN(
        cor_maj_62_n33) );
  NAND2_X1 cor_maj_62_U2 ( .A1(cor_maj_62_n34), .A2(cor_maj_62_n33), .ZN(
        cor_maj_62_port_o) );
  OR2_X1 cor_maj_63_U19 ( .A1(cor_maj_63_n27), .A2(cor_maj_63_n26), .ZN(
        cor_maj_63_n28) );
  NAND2_X1 cor_maj_63_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_63_n28), .ZN(
        cor_maj_63_n29) );
  NAND2_X1 cor_maj_63_U17 ( .A1(cor_maj_63_n26), .A2(cor_maj_63_n27), .ZN(
        cor_maj_63_n30) );
  NAND2_X1 cor_maj_63_U16 ( .A1(cor_maj_63_n30), .A2(cor_maj_63_n29), .ZN(
        cor_maj_63_n31) );
  NAND2_X1 cor_maj_63_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_63_n25), .ZN(
        cor_maj_63_n18) );
  NAND2_X1 cor_maj_63_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_63_n19) );
  NAND2_X1 cor_maj_63_U13 ( .A1(cor_maj_63_n19), .A2(cor_maj_63_n18), .ZN(
        cor_maj_63_n22) );
  NAND2_X1 cor_maj_63_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_63_n24), .ZN(
        cor_maj_63_n20) );
  NAND2_X1 cor_maj_63_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_63_n21) );
  NAND2_X1 cor_maj_63_U10 ( .A1(cor_maj_63_n21), .A2(cor_maj_63_n20), .ZN(
        cor_maj_63_n23) );
  XOR2_X1 cor_maj_63_U9 ( .A(v_1_1_2[2]), .B(cor_maj_63_n24), .Z(
        cor_maj_63_n26) );
  XOR2_X1 cor_maj_63_U8 ( .A(v_1_1_2[5]), .B(cor_maj_63_n25), .Z(
        cor_maj_63_n27) );
  XOR2_X1 cor_maj_63_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_63_n24)
         );
  XOR2_X1 cor_maj_63_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_63_n25)
         );
  OR2_X1 cor_maj_63_U5 ( .A1(cor_maj_63_n23), .A2(cor_maj_63_n22), .ZN(
        cor_maj_63_n32) );
  NAND2_X1 cor_maj_63_U4 ( .A1(cor_maj_63_n22), .A2(cor_maj_63_n23), .ZN(
        cor_maj_63_n34) );
  NAND2_X1 cor_maj_63_U3 ( .A1(cor_maj_63_n32), .A2(cor_maj_63_n31), .ZN(
        cor_maj_63_n33) );
  NAND2_X1 cor_maj_63_U2 ( .A1(cor_maj_63_n34), .A2(cor_maj_63_n33), .ZN(
        cor_maj_63_port_o) );
  OR2_X1 cor_maj_64_U19 ( .A1(cor_maj_64_n27), .A2(cor_maj_64_n26), .ZN(
        cor_maj_64_n28) );
  NAND2_X1 cor_maj_64_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_64_n28), .ZN(
        cor_maj_64_n29) );
  NAND2_X1 cor_maj_64_U17 ( .A1(cor_maj_64_n26), .A2(cor_maj_64_n27), .ZN(
        cor_maj_64_n30) );
  NAND2_X1 cor_maj_64_U16 ( .A1(cor_maj_64_n30), .A2(cor_maj_64_n29), .ZN(
        cor_maj_64_n31) );
  NAND2_X1 cor_maj_64_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_64_n25), .ZN(
        cor_maj_64_n18) );
  NAND2_X1 cor_maj_64_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_64_n19) );
  NAND2_X1 cor_maj_64_U13 ( .A1(cor_maj_64_n19), .A2(cor_maj_64_n18), .ZN(
        cor_maj_64_n22) );
  NAND2_X1 cor_maj_64_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_64_n24), .ZN(
        cor_maj_64_n20) );
  NAND2_X1 cor_maj_64_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_64_n21) );
  NAND2_X1 cor_maj_64_U10 ( .A1(cor_maj_64_n21), .A2(cor_maj_64_n20), .ZN(
        cor_maj_64_n23) );
  XOR2_X1 cor_maj_64_U9 ( .A(v_1_1_2[2]), .B(cor_maj_64_n24), .Z(
        cor_maj_64_n26) );
  XOR2_X1 cor_maj_64_U8 ( .A(v_1_1_2[5]), .B(cor_maj_64_n25), .Z(
        cor_maj_64_n27) );
  XOR2_X1 cor_maj_64_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_64_n24)
         );
  XOR2_X1 cor_maj_64_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_64_n25)
         );
  OR2_X1 cor_maj_64_U5 ( .A1(cor_maj_64_n23), .A2(cor_maj_64_n22), .ZN(
        cor_maj_64_n32) );
  NAND2_X1 cor_maj_64_U4 ( .A1(cor_maj_64_n22), .A2(cor_maj_64_n23), .ZN(
        cor_maj_64_n34) );
  NAND2_X1 cor_maj_64_U3 ( .A1(cor_maj_64_n32), .A2(cor_maj_64_n31), .ZN(
        cor_maj_64_n33) );
  NAND2_X1 cor_maj_64_U2 ( .A1(cor_maj_64_n34), .A2(cor_maj_64_n33), .ZN(
        cor_maj_64_port_o) );
  OR2_X1 cor_maj_65_U19 ( .A1(cor_maj_65_n27), .A2(cor_maj_65_n26), .ZN(
        cor_maj_65_n28) );
  NAND2_X1 cor_maj_65_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_65_n28), .ZN(
        cor_maj_65_n29) );
  NAND2_X1 cor_maj_65_U17 ( .A1(cor_maj_65_n26), .A2(cor_maj_65_n27), .ZN(
        cor_maj_65_n30) );
  NAND2_X1 cor_maj_65_U16 ( .A1(cor_maj_65_n30), .A2(cor_maj_65_n29), .ZN(
        cor_maj_65_n31) );
  NAND2_X1 cor_maj_65_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_65_n25), .ZN(
        cor_maj_65_n18) );
  NAND2_X1 cor_maj_65_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_65_n19) );
  NAND2_X1 cor_maj_65_U13 ( .A1(cor_maj_65_n19), .A2(cor_maj_65_n18), .ZN(
        cor_maj_65_n22) );
  NAND2_X1 cor_maj_65_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_65_n24), .ZN(
        cor_maj_65_n20) );
  NAND2_X1 cor_maj_65_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_65_n21) );
  NAND2_X1 cor_maj_65_U10 ( .A1(cor_maj_65_n21), .A2(cor_maj_65_n20), .ZN(
        cor_maj_65_n23) );
  XOR2_X1 cor_maj_65_U9 ( .A(v_1_1_2[2]), .B(cor_maj_65_n24), .Z(
        cor_maj_65_n26) );
  XOR2_X1 cor_maj_65_U8 ( .A(v_1_1_2[5]), .B(cor_maj_65_n25), .Z(
        cor_maj_65_n27) );
  XOR2_X1 cor_maj_65_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_65_n24)
         );
  XOR2_X1 cor_maj_65_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_65_n25)
         );
  OR2_X1 cor_maj_65_U5 ( .A1(cor_maj_65_n23), .A2(cor_maj_65_n22), .ZN(
        cor_maj_65_n32) );
  NAND2_X1 cor_maj_65_U4 ( .A1(cor_maj_65_n22), .A2(cor_maj_65_n23), .ZN(
        cor_maj_65_n34) );
  NAND2_X1 cor_maj_65_U3 ( .A1(cor_maj_65_n32), .A2(cor_maj_65_n31), .ZN(
        cor_maj_65_n33) );
  NAND2_X1 cor_maj_65_U2 ( .A1(cor_maj_65_n34), .A2(cor_maj_65_n33), .ZN(
        cor_maj_65_port_o) );
  OR2_X1 cor_maj_66_U19 ( .A1(cor_maj_66_n27), .A2(cor_maj_66_n26), .ZN(
        cor_maj_66_n28) );
  NAND2_X1 cor_maj_66_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_66_n28), .ZN(
        cor_maj_66_n29) );
  NAND2_X1 cor_maj_66_U17 ( .A1(cor_maj_66_n26), .A2(cor_maj_66_n27), .ZN(
        cor_maj_66_n30) );
  NAND2_X1 cor_maj_66_U16 ( .A1(cor_maj_66_n30), .A2(cor_maj_66_n29), .ZN(
        cor_maj_66_n31) );
  NAND2_X1 cor_maj_66_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_66_n25), .ZN(
        cor_maj_66_n18) );
  NAND2_X1 cor_maj_66_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_66_n19) );
  NAND2_X1 cor_maj_66_U13 ( .A1(cor_maj_66_n19), .A2(cor_maj_66_n18), .ZN(
        cor_maj_66_n22) );
  NAND2_X1 cor_maj_66_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_66_n24), .ZN(
        cor_maj_66_n20) );
  NAND2_X1 cor_maj_66_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_66_n21) );
  NAND2_X1 cor_maj_66_U10 ( .A1(cor_maj_66_n21), .A2(cor_maj_66_n20), .ZN(
        cor_maj_66_n23) );
  XOR2_X1 cor_maj_66_U9 ( .A(v_1_1_2[2]), .B(cor_maj_66_n24), .Z(
        cor_maj_66_n26) );
  XOR2_X1 cor_maj_66_U8 ( .A(v_1_1_2[5]), .B(cor_maj_66_n25), .Z(
        cor_maj_66_n27) );
  XOR2_X1 cor_maj_66_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_66_n24)
         );
  XOR2_X1 cor_maj_66_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_66_n25)
         );
  OR2_X1 cor_maj_66_U5 ( .A1(cor_maj_66_n23), .A2(cor_maj_66_n22), .ZN(
        cor_maj_66_n32) );
  NAND2_X1 cor_maj_66_U4 ( .A1(cor_maj_66_n22), .A2(cor_maj_66_n23), .ZN(
        cor_maj_66_n34) );
  NAND2_X1 cor_maj_66_U3 ( .A1(cor_maj_66_n32), .A2(cor_maj_66_n31), .ZN(
        cor_maj_66_n33) );
  NAND2_X1 cor_maj_66_U2 ( .A1(cor_maj_66_n34), .A2(cor_maj_66_n33), .ZN(
        cor_maj_66_port_o) );
  OR2_X1 cor_maj_67_U19 ( .A1(cor_maj_67_n27), .A2(cor_maj_67_n26), .ZN(
        cor_maj_67_n28) );
  NAND2_X1 cor_maj_67_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_67_n28), .ZN(
        cor_maj_67_n29) );
  NAND2_X1 cor_maj_67_U17 ( .A1(cor_maj_67_n26), .A2(cor_maj_67_n27), .ZN(
        cor_maj_67_n30) );
  NAND2_X1 cor_maj_67_U16 ( .A1(cor_maj_67_n30), .A2(cor_maj_67_n29), .ZN(
        cor_maj_67_n31) );
  NAND2_X1 cor_maj_67_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_67_n25), .ZN(
        cor_maj_67_n18) );
  NAND2_X1 cor_maj_67_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_67_n19) );
  NAND2_X1 cor_maj_67_U13 ( .A1(cor_maj_67_n19), .A2(cor_maj_67_n18), .ZN(
        cor_maj_67_n22) );
  NAND2_X1 cor_maj_67_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_67_n24), .ZN(
        cor_maj_67_n20) );
  NAND2_X1 cor_maj_67_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_67_n21) );
  NAND2_X1 cor_maj_67_U10 ( .A1(cor_maj_67_n21), .A2(cor_maj_67_n20), .ZN(
        cor_maj_67_n23) );
  XOR2_X1 cor_maj_67_U9 ( .A(v_1_1_2[2]), .B(cor_maj_67_n24), .Z(
        cor_maj_67_n26) );
  XOR2_X1 cor_maj_67_U8 ( .A(v_1_1_2[5]), .B(cor_maj_67_n25), .Z(
        cor_maj_67_n27) );
  XOR2_X1 cor_maj_67_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_67_n24)
         );
  XOR2_X1 cor_maj_67_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_67_n25)
         );
  OR2_X1 cor_maj_67_U5 ( .A1(cor_maj_67_n23), .A2(cor_maj_67_n22), .ZN(
        cor_maj_67_n32) );
  NAND2_X1 cor_maj_67_U4 ( .A1(cor_maj_67_n22), .A2(cor_maj_67_n23), .ZN(
        cor_maj_67_n34) );
  NAND2_X1 cor_maj_67_U3 ( .A1(cor_maj_67_n32), .A2(cor_maj_67_n31), .ZN(
        cor_maj_67_n33) );
  NAND2_X1 cor_maj_67_U2 ( .A1(cor_maj_67_n34), .A2(cor_maj_67_n33), .ZN(
        cor_maj_67_port_o) );
  OR2_X1 cor_maj_68_U19 ( .A1(cor_maj_68_n27), .A2(cor_maj_68_n26), .ZN(
        cor_maj_68_n28) );
  NAND2_X1 cor_maj_68_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_68_n28), .ZN(
        cor_maj_68_n29) );
  NAND2_X1 cor_maj_68_U17 ( .A1(cor_maj_68_n26), .A2(cor_maj_68_n27), .ZN(
        cor_maj_68_n30) );
  NAND2_X1 cor_maj_68_U16 ( .A1(cor_maj_68_n30), .A2(cor_maj_68_n29), .ZN(
        cor_maj_68_n31) );
  NAND2_X1 cor_maj_68_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_68_n25), .ZN(
        cor_maj_68_n18) );
  NAND2_X1 cor_maj_68_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_68_n19) );
  NAND2_X1 cor_maj_68_U13 ( .A1(cor_maj_68_n19), .A2(cor_maj_68_n18), .ZN(
        cor_maj_68_n22) );
  NAND2_X1 cor_maj_68_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_68_n24), .ZN(
        cor_maj_68_n20) );
  NAND2_X1 cor_maj_68_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_68_n21) );
  NAND2_X1 cor_maj_68_U10 ( .A1(cor_maj_68_n21), .A2(cor_maj_68_n20), .ZN(
        cor_maj_68_n23) );
  XOR2_X1 cor_maj_68_U9 ( .A(v_1_1_2[2]), .B(cor_maj_68_n24), .Z(
        cor_maj_68_n26) );
  XOR2_X1 cor_maj_68_U8 ( .A(v_1_1_2[5]), .B(cor_maj_68_n25), .Z(
        cor_maj_68_n27) );
  XOR2_X1 cor_maj_68_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_68_n24)
         );
  XOR2_X1 cor_maj_68_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_68_n25)
         );
  OR2_X1 cor_maj_68_U5 ( .A1(cor_maj_68_n23), .A2(cor_maj_68_n22), .ZN(
        cor_maj_68_n32) );
  NAND2_X1 cor_maj_68_U4 ( .A1(cor_maj_68_n22), .A2(cor_maj_68_n23), .ZN(
        cor_maj_68_n34) );
  NAND2_X1 cor_maj_68_U3 ( .A1(cor_maj_68_n32), .A2(cor_maj_68_n31), .ZN(
        cor_maj_68_n33) );
  NAND2_X1 cor_maj_68_U2 ( .A1(cor_maj_68_n34), .A2(cor_maj_68_n33), .ZN(
        cor_maj_68_port_o) );
  OR2_X1 cor_maj_69_U19 ( .A1(cor_maj_69_n27), .A2(cor_maj_69_n26), .ZN(
        cor_maj_69_n28) );
  NAND2_X1 cor_maj_69_U18 ( .A1(v_1_1_2[6]), .A2(cor_maj_69_n28), .ZN(
        cor_maj_69_n29) );
  NAND2_X1 cor_maj_69_U17 ( .A1(cor_maj_69_n26), .A2(cor_maj_69_n27), .ZN(
        cor_maj_69_n30) );
  NAND2_X1 cor_maj_69_U16 ( .A1(cor_maj_69_n30), .A2(cor_maj_69_n29), .ZN(
        cor_maj_69_n31) );
  NAND2_X1 cor_maj_69_U15 ( .A1(v_1_1_2[5]), .A2(cor_maj_69_n25), .ZN(
        cor_maj_69_n18) );
  NAND2_X1 cor_maj_69_U14 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_69_n19) );
  NAND2_X1 cor_maj_69_U13 ( .A1(cor_maj_69_n19), .A2(cor_maj_69_n18), .ZN(
        cor_maj_69_n22) );
  NAND2_X1 cor_maj_69_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_69_n24), .ZN(
        cor_maj_69_n20) );
  NAND2_X1 cor_maj_69_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_69_n21) );
  NAND2_X1 cor_maj_69_U10 ( .A1(cor_maj_69_n21), .A2(cor_maj_69_n20), .ZN(
        cor_maj_69_n23) );
  XOR2_X1 cor_maj_69_U9 ( .A(v_1_1_2[2]), .B(cor_maj_69_n24), .Z(
        cor_maj_69_n26) );
  XOR2_X1 cor_maj_69_U8 ( .A(v_1_1_2[5]), .B(cor_maj_69_n25), .Z(
        cor_maj_69_n27) );
  XOR2_X1 cor_maj_69_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_69_n24)
         );
  XOR2_X1 cor_maj_69_U6 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_69_n25)
         );
  OR2_X1 cor_maj_69_U5 ( .A1(cor_maj_69_n23), .A2(cor_maj_69_n22), .ZN(
        cor_maj_69_n32) );
  NAND2_X1 cor_maj_69_U4 ( .A1(cor_maj_69_n22), .A2(cor_maj_69_n23), .ZN(
        cor_maj_69_n34) );
  NAND2_X1 cor_maj_69_U3 ( .A1(cor_maj_69_n32), .A2(cor_maj_69_n31), .ZN(
        cor_maj_69_n33) );
  NAND2_X1 cor_maj_69_U2 ( .A1(cor_maj_69_n34), .A2(cor_maj_69_n33), .ZN(
        cor_maj_69_port_o) );
  OR2_X1 cor_maj_70_U19 ( .A1(cor_maj_70_n27), .A2(cor_maj_70_n26), .ZN(
        cor_maj_70_n28) );
  NAND2_X1 cor_maj_70_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_70_n28), .ZN(
        cor_maj_70_n29) );
  NAND2_X1 cor_maj_70_U17 ( .A1(cor_maj_70_n26), .A2(cor_maj_70_n27), .ZN(
        cor_maj_70_n30) );
  NAND2_X1 cor_maj_70_U16 ( .A1(cor_maj_70_n30), .A2(cor_maj_70_n29), .ZN(
        cor_maj_70_n31) );
  NAND2_X1 cor_maj_70_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_70_n25), .ZN(
        cor_maj_70_n18) );
  NAND2_X1 cor_maj_70_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_70_n19) );
  NAND2_X1 cor_maj_70_U13 ( .A1(cor_maj_70_n19), .A2(cor_maj_70_n18), .ZN(
        cor_maj_70_n22) );
  NAND2_X1 cor_maj_70_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_70_n24), .ZN(
        cor_maj_70_n20) );
  NAND2_X1 cor_maj_70_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_70_n21) );
  NAND2_X1 cor_maj_70_U10 ( .A1(cor_maj_70_n21), .A2(cor_maj_70_n20), .ZN(
        cor_maj_70_n23) );
  XOR2_X1 cor_maj_70_U9 ( .A(v_1_2_0[2]), .B(cor_maj_70_n24), .Z(
        cor_maj_70_n26) );
  XOR2_X1 cor_maj_70_U8 ( .A(v_1_2_0[5]), .B(cor_maj_70_n25), .Z(
        cor_maj_70_n27) );
  XOR2_X1 cor_maj_70_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_70_n24)
         );
  XOR2_X1 cor_maj_70_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_70_n25)
         );
  OR2_X1 cor_maj_70_U5 ( .A1(cor_maj_70_n23), .A2(cor_maj_70_n22), .ZN(
        cor_maj_70_n32) );
  NAND2_X1 cor_maj_70_U4 ( .A1(cor_maj_70_n22), .A2(cor_maj_70_n23), .ZN(
        cor_maj_70_n34) );
  NAND2_X1 cor_maj_70_U3 ( .A1(cor_maj_70_n32), .A2(cor_maj_70_n31), .ZN(
        cor_maj_70_n33) );
  NAND2_X1 cor_maj_70_U2 ( .A1(cor_maj_70_n34), .A2(cor_maj_70_n33), .ZN(
        cor_maj_70_port_o) );
  OR2_X1 cor_maj_71_U19 ( .A1(cor_maj_71_n27), .A2(cor_maj_71_n26), .ZN(
        cor_maj_71_n28) );
  NAND2_X1 cor_maj_71_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_71_n28), .ZN(
        cor_maj_71_n29) );
  NAND2_X1 cor_maj_71_U17 ( .A1(cor_maj_71_n26), .A2(cor_maj_71_n27), .ZN(
        cor_maj_71_n30) );
  NAND2_X1 cor_maj_71_U16 ( .A1(cor_maj_71_n30), .A2(cor_maj_71_n29), .ZN(
        cor_maj_71_n31) );
  NAND2_X1 cor_maj_71_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_71_n25), .ZN(
        cor_maj_71_n18) );
  NAND2_X1 cor_maj_71_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_71_n19) );
  NAND2_X1 cor_maj_71_U13 ( .A1(cor_maj_71_n19), .A2(cor_maj_71_n18), .ZN(
        cor_maj_71_n22) );
  NAND2_X1 cor_maj_71_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_71_n24), .ZN(
        cor_maj_71_n20) );
  NAND2_X1 cor_maj_71_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_71_n21) );
  NAND2_X1 cor_maj_71_U10 ( .A1(cor_maj_71_n21), .A2(cor_maj_71_n20), .ZN(
        cor_maj_71_n23) );
  XOR2_X1 cor_maj_71_U9 ( .A(v_1_2_0[2]), .B(cor_maj_71_n24), .Z(
        cor_maj_71_n26) );
  XOR2_X1 cor_maj_71_U8 ( .A(v_1_2_0[5]), .B(cor_maj_71_n25), .Z(
        cor_maj_71_n27) );
  XOR2_X1 cor_maj_71_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_71_n24)
         );
  XOR2_X1 cor_maj_71_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_71_n25)
         );
  OR2_X1 cor_maj_71_U5 ( .A1(cor_maj_71_n23), .A2(cor_maj_71_n22), .ZN(
        cor_maj_71_n32) );
  NAND2_X1 cor_maj_71_U4 ( .A1(cor_maj_71_n22), .A2(cor_maj_71_n23), .ZN(
        cor_maj_71_n34) );
  NAND2_X1 cor_maj_71_U3 ( .A1(cor_maj_71_n32), .A2(cor_maj_71_n31), .ZN(
        cor_maj_71_n33) );
  NAND2_X1 cor_maj_71_U2 ( .A1(cor_maj_71_n34), .A2(cor_maj_71_n33), .ZN(
        cor_maj_71_port_o) );
  OR2_X1 cor_maj_72_U19 ( .A1(cor_maj_72_n27), .A2(cor_maj_72_n26), .ZN(
        cor_maj_72_n28) );
  NAND2_X1 cor_maj_72_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_72_n28), .ZN(
        cor_maj_72_n29) );
  NAND2_X1 cor_maj_72_U17 ( .A1(cor_maj_72_n26), .A2(cor_maj_72_n27), .ZN(
        cor_maj_72_n30) );
  NAND2_X1 cor_maj_72_U16 ( .A1(cor_maj_72_n30), .A2(cor_maj_72_n29), .ZN(
        cor_maj_72_n31) );
  NAND2_X1 cor_maj_72_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_72_n25), .ZN(
        cor_maj_72_n18) );
  NAND2_X1 cor_maj_72_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_72_n19) );
  NAND2_X1 cor_maj_72_U13 ( .A1(cor_maj_72_n19), .A2(cor_maj_72_n18), .ZN(
        cor_maj_72_n22) );
  NAND2_X1 cor_maj_72_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_72_n24), .ZN(
        cor_maj_72_n20) );
  NAND2_X1 cor_maj_72_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_72_n21) );
  NAND2_X1 cor_maj_72_U10 ( .A1(cor_maj_72_n21), .A2(cor_maj_72_n20), .ZN(
        cor_maj_72_n23) );
  XOR2_X1 cor_maj_72_U9 ( .A(v_1_2_0[2]), .B(cor_maj_72_n24), .Z(
        cor_maj_72_n26) );
  XOR2_X1 cor_maj_72_U8 ( .A(v_1_2_0[5]), .B(cor_maj_72_n25), .Z(
        cor_maj_72_n27) );
  XOR2_X1 cor_maj_72_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_72_n24)
         );
  XOR2_X1 cor_maj_72_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_72_n25)
         );
  OR2_X1 cor_maj_72_U5 ( .A1(cor_maj_72_n23), .A2(cor_maj_72_n22), .ZN(
        cor_maj_72_n32) );
  NAND2_X1 cor_maj_72_U4 ( .A1(cor_maj_72_n22), .A2(cor_maj_72_n23), .ZN(
        cor_maj_72_n34) );
  NAND2_X1 cor_maj_72_U3 ( .A1(cor_maj_72_n32), .A2(cor_maj_72_n31), .ZN(
        cor_maj_72_n33) );
  NAND2_X1 cor_maj_72_U2 ( .A1(cor_maj_72_n34), .A2(cor_maj_72_n33), .ZN(
        cor_maj_72_port_o) );
  OR2_X1 cor_maj_73_U19 ( .A1(cor_maj_73_n27), .A2(cor_maj_73_n26), .ZN(
        cor_maj_73_n28) );
  NAND2_X1 cor_maj_73_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_73_n28), .ZN(
        cor_maj_73_n29) );
  NAND2_X1 cor_maj_73_U17 ( .A1(cor_maj_73_n26), .A2(cor_maj_73_n27), .ZN(
        cor_maj_73_n30) );
  NAND2_X1 cor_maj_73_U16 ( .A1(cor_maj_73_n30), .A2(cor_maj_73_n29), .ZN(
        cor_maj_73_n31) );
  NAND2_X1 cor_maj_73_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_73_n25), .ZN(
        cor_maj_73_n18) );
  NAND2_X1 cor_maj_73_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_73_n19) );
  NAND2_X1 cor_maj_73_U13 ( .A1(cor_maj_73_n19), .A2(cor_maj_73_n18), .ZN(
        cor_maj_73_n22) );
  NAND2_X1 cor_maj_73_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_73_n24), .ZN(
        cor_maj_73_n20) );
  NAND2_X1 cor_maj_73_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_73_n21) );
  NAND2_X1 cor_maj_73_U10 ( .A1(cor_maj_73_n21), .A2(cor_maj_73_n20), .ZN(
        cor_maj_73_n23) );
  XOR2_X1 cor_maj_73_U9 ( .A(v_1_2_0[2]), .B(cor_maj_73_n24), .Z(
        cor_maj_73_n26) );
  XOR2_X1 cor_maj_73_U8 ( .A(v_1_2_0[5]), .B(cor_maj_73_n25), .Z(
        cor_maj_73_n27) );
  XOR2_X1 cor_maj_73_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_73_n24)
         );
  XOR2_X1 cor_maj_73_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_73_n25)
         );
  OR2_X1 cor_maj_73_U5 ( .A1(cor_maj_73_n23), .A2(cor_maj_73_n22), .ZN(
        cor_maj_73_n32) );
  NAND2_X1 cor_maj_73_U4 ( .A1(cor_maj_73_n22), .A2(cor_maj_73_n23), .ZN(
        cor_maj_73_n34) );
  NAND2_X1 cor_maj_73_U3 ( .A1(cor_maj_73_n32), .A2(cor_maj_73_n31), .ZN(
        cor_maj_73_n33) );
  NAND2_X1 cor_maj_73_U2 ( .A1(cor_maj_73_n34), .A2(cor_maj_73_n33), .ZN(
        cor_maj_73_port_o) );
  OR2_X1 cor_maj_74_U19 ( .A1(cor_maj_74_n27), .A2(cor_maj_74_n26), .ZN(
        cor_maj_74_n28) );
  NAND2_X1 cor_maj_74_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_74_n28), .ZN(
        cor_maj_74_n29) );
  NAND2_X1 cor_maj_74_U17 ( .A1(cor_maj_74_n26), .A2(cor_maj_74_n27), .ZN(
        cor_maj_74_n30) );
  NAND2_X1 cor_maj_74_U16 ( .A1(cor_maj_74_n30), .A2(cor_maj_74_n29), .ZN(
        cor_maj_74_n31) );
  NAND2_X1 cor_maj_74_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_74_n25), .ZN(
        cor_maj_74_n18) );
  NAND2_X1 cor_maj_74_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_74_n19) );
  NAND2_X1 cor_maj_74_U13 ( .A1(cor_maj_74_n19), .A2(cor_maj_74_n18), .ZN(
        cor_maj_74_n22) );
  NAND2_X1 cor_maj_74_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_74_n24), .ZN(
        cor_maj_74_n20) );
  NAND2_X1 cor_maj_74_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_74_n21) );
  NAND2_X1 cor_maj_74_U10 ( .A1(cor_maj_74_n21), .A2(cor_maj_74_n20), .ZN(
        cor_maj_74_n23) );
  XOR2_X1 cor_maj_74_U9 ( .A(v_1_2_0[2]), .B(cor_maj_74_n24), .Z(
        cor_maj_74_n26) );
  XOR2_X1 cor_maj_74_U8 ( .A(v_1_2_0[5]), .B(cor_maj_74_n25), .Z(
        cor_maj_74_n27) );
  XOR2_X1 cor_maj_74_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_74_n24)
         );
  XOR2_X1 cor_maj_74_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_74_n25)
         );
  OR2_X1 cor_maj_74_U5 ( .A1(cor_maj_74_n23), .A2(cor_maj_74_n22), .ZN(
        cor_maj_74_n32) );
  NAND2_X1 cor_maj_74_U4 ( .A1(cor_maj_74_n22), .A2(cor_maj_74_n23), .ZN(
        cor_maj_74_n34) );
  NAND2_X1 cor_maj_74_U3 ( .A1(cor_maj_74_n32), .A2(cor_maj_74_n31), .ZN(
        cor_maj_74_n33) );
  NAND2_X1 cor_maj_74_U2 ( .A1(cor_maj_74_n34), .A2(cor_maj_74_n33), .ZN(
        cor_maj_74_port_o) );
  OR2_X1 cor_maj_75_U19 ( .A1(cor_maj_75_n27), .A2(cor_maj_75_n26), .ZN(
        cor_maj_75_n28) );
  NAND2_X1 cor_maj_75_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_75_n28), .ZN(
        cor_maj_75_n29) );
  NAND2_X1 cor_maj_75_U17 ( .A1(cor_maj_75_n26), .A2(cor_maj_75_n27), .ZN(
        cor_maj_75_n30) );
  NAND2_X1 cor_maj_75_U16 ( .A1(cor_maj_75_n30), .A2(cor_maj_75_n29), .ZN(
        cor_maj_75_n31) );
  NAND2_X1 cor_maj_75_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_75_n25), .ZN(
        cor_maj_75_n18) );
  NAND2_X1 cor_maj_75_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_75_n19) );
  NAND2_X1 cor_maj_75_U13 ( .A1(cor_maj_75_n19), .A2(cor_maj_75_n18), .ZN(
        cor_maj_75_n22) );
  NAND2_X1 cor_maj_75_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_75_n24), .ZN(
        cor_maj_75_n20) );
  NAND2_X1 cor_maj_75_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_75_n21) );
  NAND2_X1 cor_maj_75_U10 ( .A1(cor_maj_75_n21), .A2(cor_maj_75_n20), .ZN(
        cor_maj_75_n23) );
  XOR2_X1 cor_maj_75_U9 ( .A(v_1_2_0[2]), .B(cor_maj_75_n24), .Z(
        cor_maj_75_n26) );
  XOR2_X1 cor_maj_75_U8 ( .A(v_1_2_0[5]), .B(cor_maj_75_n25), .Z(
        cor_maj_75_n27) );
  XOR2_X1 cor_maj_75_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_75_n24)
         );
  XOR2_X1 cor_maj_75_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_75_n25)
         );
  OR2_X1 cor_maj_75_U5 ( .A1(cor_maj_75_n23), .A2(cor_maj_75_n22), .ZN(
        cor_maj_75_n32) );
  NAND2_X1 cor_maj_75_U4 ( .A1(cor_maj_75_n22), .A2(cor_maj_75_n23), .ZN(
        cor_maj_75_n34) );
  NAND2_X1 cor_maj_75_U3 ( .A1(cor_maj_75_n32), .A2(cor_maj_75_n31), .ZN(
        cor_maj_75_n33) );
  NAND2_X1 cor_maj_75_U2 ( .A1(cor_maj_75_n34), .A2(cor_maj_75_n33), .ZN(
        cor_maj_75_port_o) );
  OR2_X1 cor_maj_76_U19 ( .A1(cor_maj_76_n27), .A2(cor_maj_76_n26), .ZN(
        cor_maj_76_n28) );
  NAND2_X1 cor_maj_76_U18 ( .A1(v_1_2_0[6]), .A2(cor_maj_76_n28), .ZN(
        cor_maj_76_n29) );
  NAND2_X1 cor_maj_76_U17 ( .A1(cor_maj_76_n26), .A2(cor_maj_76_n27), .ZN(
        cor_maj_76_n30) );
  NAND2_X1 cor_maj_76_U16 ( .A1(cor_maj_76_n30), .A2(cor_maj_76_n29), .ZN(
        cor_maj_76_n31) );
  NAND2_X1 cor_maj_76_U15 ( .A1(v_1_2_0[5]), .A2(cor_maj_76_n25), .ZN(
        cor_maj_76_n18) );
  NAND2_X1 cor_maj_76_U14 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_76_n19) );
  NAND2_X1 cor_maj_76_U13 ( .A1(cor_maj_76_n19), .A2(cor_maj_76_n18), .ZN(
        cor_maj_76_n22) );
  NAND2_X1 cor_maj_76_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_76_n24), .ZN(
        cor_maj_76_n20) );
  NAND2_X1 cor_maj_76_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_76_n21) );
  NAND2_X1 cor_maj_76_U10 ( .A1(cor_maj_76_n21), .A2(cor_maj_76_n20), .ZN(
        cor_maj_76_n23) );
  XOR2_X1 cor_maj_76_U9 ( .A(v_1_2_0[2]), .B(cor_maj_76_n24), .Z(
        cor_maj_76_n26) );
  XOR2_X1 cor_maj_76_U8 ( .A(v_1_2_0[5]), .B(cor_maj_76_n25), .Z(
        cor_maj_76_n27) );
  XOR2_X1 cor_maj_76_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_76_n24)
         );
  XOR2_X1 cor_maj_76_U6 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_76_n25)
         );
  OR2_X1 cor_maj_76_U5 ( .A1(cor_maj_76_n23), .A2(cor_maj_76_n22), .ZN(
        cor_maj_76_n32) );
  NAND2_X1 cor_maj_76_U4 ( .A1(cor_maj_76_n22), .A2(cor_maj_76_n23), .ZN(
        cor_maj_76_n34) );
  NAND2_X1 cor_maj_76_U3 ( .A1(cor_maj_76_n32), .A2(cor_maj_76_n31), .ZN(
        cor_maj_76_n33) );
  NAND2_X1 cor_maj_76_U2 ( .A1(cor_maj_76_n34), .A2(cor_maj_76_n33), .ZN(
        cor_maj_76_port_o) );
  OR2_X1 cor_maj_77_U19 ( .A1(cor_maj_77_n27), .A2(cor_maj_77_n26), .ZN(
        cor_maj_77_n28) );
  NAND2_X1 cor_maj_77_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_77_n28), .ZN(
        cor_maj_77_n29) );
  NAND2_X1 cor_maj_77_U17 ( .A1(cor_maj_77_n26), .A2(cor_maj_77_n27), .ZN(
        cor_maj_77_n30) );
  NAND2_X1 cor_maj_77_U16 ( .A1(cor_maj_77_n30), .A2(cor_maj_77_n29), .ZN(
        cor_maj_77_n31) );
  NAND2_X1 cor_maj_77_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_77_n25), .ZN(
        cor_maj_77_n18) );
  NAND2_X1 cor_maj_77_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_77_n19) );
  NAND2_X1 cor_maj_77_U13 ( .A1(cor_maj_77_n19), .A2(cor_maj_77_n18), .ZN(
        cor_maj_77_n22) );
  NAND2_X1 cor_maj_77_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_77_n24), .ZN(
        cor_maj_77_n20) );
  NAND2_X1 cor_maj_77_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_77_n21) );
  NAND2_X1 cor_maj_77_U10 ( .A1(cor_maj_77_n21), .A2(cor_maj_77_n20), .ZN(
        cor_maj_77_n23) );
  XOR2_X1 cor_maj_77_U9 ( .A(v_1_2_1[2]), .B(cor_maj_77_n24), .Z(
        cor_maj_77_n26) );
  XOR2_X1 cor_maj_77_U8 ( .A(v_1_2_1[5]), .B(cor_maj_77_n25), .Z(
        cor_maj_77_n27) );
  XOR2_X1 cor_maj_77_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_77_n24)
         );
  XOR2_X1 cor_maj_77_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_77_n25)
         );
  OR2_X1 cor_maj_77_U5 ( .A1(cor_maj_77_n23), .A2(cor_maj_77_n22), .ZN(
        cor_maj_77_n32) );
  NAND2_X1 cor_maj_77_U4 ( .A1(cor_maj_77_n22), .A2(cor_maj_77_n23), .ZN(
        cor_maj_77_n34) );
  NAND2_X1 cor_maj_77_U3 ( .A1(cor_maj_77_n32), .A2(cor_maj_77_n31), .ZN(
        cor_maj_77_n33) );
  NAND2_X1 cor_maj_77_U2 ( .A1(cor_maj_77_n34), .A2(cor_maj_77_n33), .ZN(
        cor_maj_77_port_o) );
  OR2_X1 cor_maj_78_U19 ( .A1(cor_maj_78_n27), .A2(cor_maj_78_n26), .ZN(
        cor_maj_78_n28) );
  NAND2_X1 cor_maj_78_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_78_n28), .ZN(
        cor_maj_78_n29) );
  NAND2_X1 cor_maj_78_U17 ( .A1(cor_maj_78_n26), .A2(cor_maj_78_n27), .ZN(
        cor_maj_78_n30) );
  NAND2_X1 cor_maj_78_U16 ( .A1(cor_maj_78_n30), .A2(cor_maj_78_n29), .ZN(
        cor_maj_78_n31) );
  NAND2_X1 cor_maj_78_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_78_n25), .ZN(
        cor_maj_78_n18) );
  NAND2_X1 cor_maj_78_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_78_n19) );
  NAND2_X1 cor_maj_78_U13 ( .A1(cor_maj_78_n19), .A2(cor_maj_78_n18), .ZN(
        cor_maj_78_n22) );
  NAND2_X1 cor_maj_78_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_78_n24), .ZN(
        cor_maj_78_n20) );
  NAND2_X1 cor_maj_78_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_78_n21) );
  NAND2_X1 cor_maj_78_U10 ( .A1(cor_maj_78_n21), .A2(cor_maj_78_n20), .ZN(
        cor_maj_78_n23) );
  XOR2_X1 cor_maj_78_U9 ( .A(v_1_2_1[2]), .B(cor_maj_78_n24), .Z(
        cor_maj_78_n26) );
  XOR2_X1 cor_maj_78_U8 ( .A(v_1_2_1[5]), .B(cor_maj_78_n25), .Z(
        cor_maj_78_n27) );
  XOR2_X1 cor_maj_78_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_78_n24)
         );
  XOR2_X1 cor_maj_78_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_78_n25)
         );
  OR2_X1 cor_maj_78_U5 ( .A1(cor_maj_78_n23), .A2(cor_maj_78_n22), .ZN(
        cor_maj_78_n32) );
  NAND2_X1 cor_maj_78_U4 ( .A1(cor_maj_78_n22), .A2(cor_maj_78_n23), .ZN(
        cor_maj_78_n34) );
  NAND2_X1 cor_maj_78_U3 ( .A1(cor_maj_78_n32), .A2(cor_maj_78_n31), .ZN(
        cor_maj_78_n33) );
  NAND2_X1 cor_maj_78_U2 ( .A1(cor_maj_78_n34), .A2(cor_maj_78_n33), .ZN(
        cor_maj_78_port_o) );
  OR2_X1 cor_maj_79_U19 ( .A1(cor_maj_79_n27), .A2(cor_maj_79_n26), .ZN(
        cor_maj_79_n28) );
  NAND2_X1 cor_maj_79_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_79_n28), .ZN(
        cor_maj_79_n29) );
  NAND2_X1 cor_maj_79_U17 ( .A1(cor_maj_79_n26), .A2(cor_maj_79_n27), .ZN(
        cor_maj_79_n30) );
  NAND2_X1 cor_maj_79_U16 ( .A1(cor_maj_79_n30), .A2(cor_maj_79_n29), .ZN(
        cor_maj_79_n31) );
  NAND2_X1 cor_maj_79_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_79_n25), .ZN(
        cor_maj_79_n18) );
  NAND2_X1 cor_maj_79_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_79_n19) );
  NAND2_X1 cor_maj_79_U13 ( .A1(cor_maj_79_n19), .A2(cor_maj_79_n18), .ZN(
        cor_maj_79_n22) );
  NAND2_X1 cor_maj_79_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_79_n24), .ZN(
        cor_maj_79_n20) );
  NAND2_X1 cor_maj_79_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_79_n21) );
  NAND2_X1 cor_maj_79_U10 ( .A1(cor_maj_79_n21), .A2(cor_maj_79_n20), .ZN(
        cor_maj_79_n23) );
  XOR2_X1 cor_maj_79_U9 ( .A(v_1_2_1[2]), .B(cor_maj_79_n24), .Z(
        cor_maj_79_n26) );
  XOR2_X1 cor_maj_79_U8 ( .A(v_1_2_1[5]), .B(cor_maj_79_n25), .Z(
        cor_maj_79_n27) );
  XOR2_X1 cor_maj_79_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_79_n24)
         );
  XOR2_X1 cor_maj_79_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_79_n25)
         );
  OR2_X1 cor_maj_79_U5 ( .A1(cor_maj_79_n23), .A2(cor_maj_79_n22), .ZN(
        cor_maj_79_n32) );
  NAND2_X1 cor_maj_79_U4 ( .A1(cor_maj_79_n22), .A2(cor_maj_79_n23), .ZN(
        cor_maj_79_n34) );
  NAND2_X1 cor_maj_79_U3 ( .A1(cor_maj_79_n32), .A2(cor_maj_79_n31), .ZN(
        cor_maj_79_n33) );
  NAND2_X1 cor_maj_79_U2 ( .A1(cor_maj_79_n34), .A2(cor_maj_79_n33), .ZN(
        cor_maj_79_port_o) );
  OR2_X1 cor_maj_80_U19 ( .A1(cor_maj_80_n27), .A2(cor_maj_80_n26), .ZN(
        cor_maj_80_n28) );
  NAND2_X1 cor_maj_80_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_80_n28), .ZN(
        cor_maj_80_n29) );
  NAND2_X1 cor_maj_80_U17 ( .A1(cor_maj_80_n26), .A2(cor_maj_80_n27), .ZN(
        cor_maj_80_n30) );
  NAND2_X1 cor_maj_80_U16 ( .A1(cor_maj_80_n30), .A2(cor_maj_80_n29), .ZN(
        cor_maj_80_n31) );
  NAND2_X1 cor_maj_80_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_80_n25), .ZN(
        cor_maj_80_n18) );
  NAND2_X1 cor_maj_80_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_80_n19) );
  NAND2_X1 cor_maj_80_U13 ( .A1(cor_maj_80_n19), .A2(cor_maj_80_n18), .ZN(
        cor_maj_80_n22) );
  NAND2_X1 cor_maj_80_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_80_n24), .ZN(
        cor_maj_80_n20) );
  NAND2_X1 cor_maj_80_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_80_n21) );
  NAND2_X1 cor_maj_80_U10 ( .A1(cor_maj_80_n21), .A2(cor_maj_80_n20), .ZN(
        cor_maj_80_n23) );
  XOR2_X1 cor_maj_80_U9 ( .A(v_1_2_1[2]), .B(cor_maj_80_n24), .Z(
        cor_maj_80_n26) );
  XOR2_X1 cor_maj_80_U8 ( .A(v_1_2_1[5]), .B(cor_maj_80_n25), .Z(
        cor_maj_80_n27) );
  XOR2_X1 cor_maj_80_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_80_n24)
         );
  XOR2_X1 cor_maj_80_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_80_n25)
         );
  OR2_X1 cor_maj_80_U5 ( .A1(cor_maj_80_n23), .A2(cor_maj_80_n22), .ZN(
        cor_maj_80_n32) );
  NAND2_X1 cor_maj_80_U4 ( .A1(cor_maj_80_n22), .A2(cor_maj_80_n23), .ZN(
        cor_maj_80_n34) );
  NAND2_X1 cor_maj_80_U3 ( .A1(cor_maj_80_n32), .A2(cor_maj_80_n31), .ZN(
        cor_maj_80_n33) );
  NAND2_X1 cor_maj_80_U2 ( .A1(cor_maj_80_n34), .A2(cor_maj_80_n33), .ZN(
        cor_maj_80_port_o) );
  OR2_X1 cor_maj_81_U19 ( .A1(cor_maj_81_n27), .A2(cor_maj_81_n26), .ZN(
        cor_maj_81_n28) );
  NAND2_X1 cor_maj_81_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_81_n28), .ZN(
        cor_maj_81_n29) );
  NAND2_X1 cor_maj_81_U17 ( .A1(cor_maj_81_n26), .A2(cor_maj_81_n27), .ZN(
        cor_maj_81_n30) );
  NAND2_X1 cor_maj_81_U16 ( .A1(cor_maj_81_n30), .A2(cor_maj_81_n29), .ZN(
        cor_maj_81_n31) );
  NAND2_X1 cor_maj_81_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_81_n25), .ZN(
        cor_maj_81_n18) );
  NAND2_X1 cor_maj_81_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_81_n19) );
  NAND2_X1 cor_maj_81_U13 ( .A1(cor_maj_81_n19), .A2(cor_maj_81_n18), .ZN(
        cor_maj_81_n22) );
  NAND2_X1 cor_maj_81_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_81_n24), .ZN(
        cor_maj_81_n20) );
  NAND2_X1 cor_maj_81_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_81_n21) );
  NAND2_X1 cor_maj_81_U10 ( .A1(cor_maj_81_n21), .A2(cor_maj_81_n20), .ZN(
        cor_maj_81_n23) );
  XOR2_X1 cor_maj_81_U9 ( .A(v_1_2_1[2]), .B(cor_maj_81_n24), .Z(
        cor_maj_81_n26) );
  XOR2_X1 cor_maj_81_U8 ( .A(v_1_2_1[5]), .B(cor_maj_81_n25), .Z(
        cor_maj_81_n27) );
  XOR2_X1 cor_maj_81_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_81_n24)
         );
  XOR2_X1 cor_maj_81_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_81_n25)
         );
  OR2_X1 cor_maj_81_U5 ( .A1(cor_maj_81_n23), .A2(cor_maj_81_n22), .ZN(
        cor_maj_81_n32) );
  NAND2_X1 cor_maj_81_U4 ( .A1(cor_maj_81_n22), .A2(cor_maj_81_n23), .ZN(
        cor_maj_81_n34) );
  NAND2_X1 cor_maj_81_U3 ( .A1(cor_maj_81_n32), .A2(cor_maj_81_n31), .ZN(
        cor_maj_81_n33) );
  NAND2_X1 cor_maj_81_U2 ( .A1(cor_maj_81_n34), .A2(cor_maj_81_n33), .ZN(
        cor_maj_81_port_o) );
  OR2_X1 cor_maj_82_U19 ( .A1(cor_maj_82_n27), .A2(cor_maj_82_n26), .ZN(
        cor_maj_82_n28) );
  NAND2_X1 cor_maj_82_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_82_n28), .ZN(
        cor_maj_82_n29) );
  NAND2_X1 cor_maj_82_U17 ( .A1(cor_maj_82_n26), .A2(cor_maj_82_n27), .ZN(
        cor_maj_82_n30) );
  NAND2_X1 cor_maj_82_U16 ( .A1(cor_maj_82_n30), .A2(cor_maj_82_n29), .ZN(
        cor_maj_82_n31) );
  NAND2_X1 cor_maj_82_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_82_n25), .ZN(
        cor_maj_82_n18) );
  NAND2_X1 cor_maj_82_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_82_n19) );
  NAND2_X1 cor_maj_82_U13 ( .A1(cor_maj_82_n19), .A2(cor_maj_82_n18), .ZN(
        cor_maj_82_n22) );
  NAND2_X1 cor_maj_82_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_82_n24), .ZN(
        cor_maj_82_n20) );
  NAND2_X1 cor_maj_82_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_82_n21) );
  NAND2_X1 cor_maj_82_U10 ( .A1(cor_maj_82_n21), .A2(cor_maj_82_n20), .ZN(
        cor_maj_82_n23) );
  XOR2_X1 cor_maj_82_U9 ( .A(v_1_2_1[2]), .B(cor_maj_82_n24), .Z(
        cor_maj_82_n26) );
  XOR2_X1 cor_maj_82_U8 ( .A(v_1_2_1[5]), .B(cor_maj_82_n25), .Z(
        cor_maj_82_n27) );
  XOR2_X1 cor_maj_82_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_82_n24)
         );
  XOR2_X1 cor_maj_82_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_82_n25)
         );
  OR2_X1 cor_maj_82_U5 ( .A1(cor_maj_82_n23), .A2(cor_maj_82_n22), .ZN(
        cor_maj_82_n32) );
  NAND2_X1 cor_maj_82_U4 ( .A1(cor_maj_82_n22), .A2(cor_maj_82_n23), .ZN(
        cor_maj_82_n34) );
  NAND2_X1 cor_maj_82_U3 ( .A1(cor_maj_82_n32), .A2(cor_maj_82_n31), .ZN(
        cor_maj_82_n33) );
  NAND2_X1 cor_maj_82_U2 ( .A1(cor_maj_82_n34), .A2(cor_maj_82_n33), .ZN(
        cor_maj_82_port_o) );
  OR2_X1 cor_maj_83_U19 ( .A1(cor_maj_83_n27), .A2(cor_maj_83_n26), .ZN(
        cor_maj_83_n28) );
  NAND2_X1 cor_maj_83_U18 ( .A1(v_1_2_1[6]), .A2(cor_maj_83_n28), .ZN(
        cor_maj_83_n29) );
  NAND2_X1 cor_maj_83_U17 ( .A1(cor_maj_83_n26), .A2(cor_maj_83_n27), .ZN(
        cor_maj_83_n30) );
  NAND2_X1 cor_maj_83_U16 ( .A1(cor_maj_83_n30), .A2(cor_maj_83_n29), .ZN(
        cor_maj_83_n31) );
  NAND2_X1 cor_maj_83_U15 ( .A1(v_1_2_1[5]), .A2(cor_maj_83_n25), .ZN(
        cor_maj_83_n18) );
  NAND2_X1 cor_maj_83_U14 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_83_n19) );
  NAND2_X1 cor_maj_83_U13 ( .A1(cor_maj_83_n19), .A2(cor_maj_83_n18), .ZN(
        cor_maj_83_n22) );
  NAND2_X1 cor_maj_83_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_83_n24), .ZN(
        cor_maj_83_n20) );
  NAND2_X1 cor_maj_83_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_83_n21) );
  NAND2_X1 cor_maj_83_U10 ( .A1(cor_maj_83_n21), .A2(cor_maj_83_n20), .ZN(
        cor_maj_83_n23) );
  XOR2_X1 cor_maj_83_U9 ( .A(v_1_2_1[2]), .B(cor_maj_83_n24), .Z(
        cor_maj_83_n26) );
  XOR2_X1 cor_maj_83_U8 ( .A(v_1_2_1[5]), .B(cor_maj_83_n25), .Z(
        cor_maj_83_n27) );
  XOR2_X1 cor_maj_83_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_83_n24)
         );
  XOR2_X1 cor_maj_83_U6 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_83_n25)
         );
  OR2_X1 cor_maj_83_U5 ( .A1(cor_maj_83_n23), .A2(cor_maj_83_n22), .ZN(
        cor_maj_83_n32) );
  NAND2_X1 cor_maj_83_U4 ( .A1(cor_maj_83_n22), .A2(cor_maj_83_n23), .ZN(
        cor_maj_83_n34) );
  NAND2_X1 cor_maj_83_U3 ( .A1(cor_maj_83_n32), .A2(cor_maj_83_n31), .ZN(
        cor_maj_83_n33) );
  NAND2_X1 cor_maj_83_U2 ( .A1(cor_maj_83_n34), .A2(cor_maj_83_n33), .ZN(
        cor_maj_83_port_o) );
  XOR2_X1 simpleXor_42_U1 ( .A(n_zz_io_c_0_3[1]), .B(u_0_1[0]), .Z(
        simpleXor_42_port_z) );
  XOR2_X1 simpleXor_43_U1 ( .A(n_zz_io_c_0_3[2]), .B(u_0_2[0]), .Z(
        simpleXor_43_port_z) );
  XOR2_X1 simpleXor_44_U1 ( .A(n_zz_io_c_1_3[1]), .B(u_1_0[0]), .Z(
        simpleXor_44_port_z) );
  XOR2_X1 simpleXor_45_U1 ( .A(n_zz_io_c_1_3[2]), .B(u_1_2[0]), .Z(
        simpleXor_45_port_z) );
  XOR2_X1 simpleXor_46_U1 ( .A(n_zz_io_c_2_3[1]), .B(u_2_0[0]), .Z(
        simpleXor_46_port_z) );
  XOR2_X1 simpleXor_47_U1 ( .A(n_zz_io_c_2_3[2]), .B(u_2_1[0]), .Z(
        simpleXor_47_port_z) );
  XOR2_X1 simpleXor_48_U1 ( .A(n_zz_io_c_0_7[1]), .B(u_0_1[1]), .Z(
        simpleXor_48_port_z) );
  XOR2_X1 simpleXor_49_U1 ( .A(n_zz_io_c_0_7[2]), .B(u_0_2[1]), .Z(
        simpleXor_49_port_z) );
  XOR2_X1 simpleXor_50_U1 ( .A(n_zz_io_c_1_7[1]), .B(u_1_0[1]), .Z(
        simpleXor_50_port_z) );
  XOR2_X1 simpleXor_51_U1 ( .A(n_zz_io_c_1_7[2]), .B(u_1_2[1]), .Z(
        simpleXor_51_port_z) );
  XOR2_X1 simpleXor_52_U1 ( .A(n_zz_io_c_2_7[1]), .B(u_2_0[1]), .Z(
        simpleXor_52_port_z) );
  XOR2_X1 simpleXor_53_U1 ( .A(n_zz_io_c_2_7[2]), .B(u_2_1[1]), .Z(
        simpleXor_53_port_z) );
  XOR2_X1 simpleXor_54_U1 ( .A(n_zz_io_c_0_11[1]), .B(u_0_1[2]), .Z(
        simpleXor_54_port_z) );
  XOR2_X1 simpleXor_55_U1 ( .A(n_zz_io_c_0_11[2]), .B(u_0_2[2]), .Z(
        simpleXor_55_port_z) );
  XOR2_X1 simpleXor_56_U1 ( .A(n_zz_io_c_1_11[1]), .B(u_1_0[2]), .Z(
        simpleXor_56_port_z) );
  XOR2_X1 simpleXor_57_U1 ( .A(n_zz_io_c_1_11[2]), .B(u_1_2[2]), .Z(
        simpleXor_57_port_z) );
  XOR2_X1 simpleXor_58_U1 ( .A(n_zz_io_c_2_11[1]), .B(u_2_0[2]), .Z(
        simpleXor_58_port_z) );
  XOR2_X1 simpleXor_59_U1 ( .A(n_zz_io_c_2_11[2]), .B(u_2_1[2]), .Z(
        simpleXor_59_port_z) );
  XOR2_X1 simpleXor_60_U1 ( .A(n_zz_io_c_0_15[1]), .B(u_0_1[3]), .Z(
        simpleXor_60_port_z) );
  XOR2_X1 simpleXor_61_U1 ( .A(n_zz_io_c_0_15[2]), .B(u_0_2[3]), .Z(
        simpleXor_61_port_z) );
  XOR2_X1 simpleXor_62_U1 ( .A(n_zz_io_c_1_15[1]), .B(u_1_0[3]), .Z(
        simpleXor_62_port_z) );
  XOR2_X1 simpleXor_63_U1 ( .A(n_zz_io_c_1_15[2]), .B(u_1_2[3]), .Z(
        simpleXor_63_port_z) );
  XOR2_X1 simpleXor_64_U1 ( .A(n_zz_io_c_2_15[1]), .B(u_2_0[3]), .Z(
        simpleXor_64_port_z) );
  XOR2_X1 simpleXor_65_U1 ( .A(n_zz_io_c_2_15[2]), .B(u_2_1[3]), .Z(
        simpleXor_65_port_z) );
  XOR2_X1 simpleXor_66_U1 ( .A(n_zz_io_c_0_19[1]), .B(u_0_1[4]), .Z(
        simpleXor_66_port_z) );
  XOR2_X1 simpleXor_67_U1 ( .A(n_zz_io_c_0_19[2]), .B(u_0_2[4]), .Z(
        simpleXor_67_port_z) );
  XOR2_X1 simpleXor_68_U1 ( .A(n_zz_io_c_1_19[1]), .B(u_1_0[4]), .Z(
        simpleXor_68_port_z) );
  XOR2_X1 simpleXor_69_U1 ( .A(n_zz_io_c_1_19[2]), .B(u_1_2[4]), .Z(
        simpleXor_69_port_z) );
  XOR2_X1 simpleXor_70_U1 ( .A(n_zz_io_c_2_19[1]), .B(u_2_0[4]), .Z(
        simpleXor_70_port_z) );
  XOR2_X1 simpleXor_71_U1 ( .A(n_zz_io_c_2_19[2]), .B(u_2_1[4]), .Z(
        simpleXor_71_port_z) );
  XOR2_X1 simpleXor_72_U1 ( .A(n_zz_io_c_0_23[1]), .B(u_0_1[5]), .Z(
        simpleXor_72_port_z) );
  XOR2_X1 simpleXor_73_U1 ( .A(n_zz_io_c_0_23[2]), .B(u_0_2[5]), .Z(
        simpleXor_73_port_z) );
  XOR2_X1 simpleXor_74_U1 ( .A(n_zz_io_c_1_23[1]), .B(u_1_0[5]), .Z(
        simpleXor_74_port_z) );
  XOR2_X1 simpleXor_75_U1 ( .A(n_zz_io_c_1_23[2]), .B(u_1_2[5]), .Z(
        simpleXor_75_port_z) );
  XOR2_X1 simpleXor_76_U1 ( .A(n_zz_io_c_2_23[1]), .B(u_2_0[5]), .Z(
        simpleXor_76_port_z) );
  XOR2_X1 simpleXor_77_U1 ( .A(n_zz_io_c_2_23[2]), .B(u_2_1[5]), .Z(
        simpleXor_77_port_z) );
  XOR2_X1 simpleXor_78_U1 ( .A(n_zz_io_c_0_27[1]), .B(u_0_1[6]), .Z(
        simpleXor_78_port_z) );
  XOR2_X1 simpleXor_79_U1 ( .A(n_zz_io_c_0_27[2]), .B(u_0_2[6]), .Z(
        simpleXor_79_port_z) );
  XOR2_X1 simpleXor_80_U1 ( .A(n_zz_io_c_1_27[1]), .B(u_1_0[6]), .Z(
        simpleXor_80_port_z) );
  XOR2_X1 simpleXor_81_U1 ( .A(n_zz_io_c_1_27[2]), .B(u_1_2[6]), .Z(
        simpleXor_81_port_z) );
  XOR2_X1 simpleXor_82_U1 ( .A(n_zz_io_c_2_27[1]), .B(u_2_0[6]), .Z(
        simpleXor_82_port_z) );
  XOR2_X1 simpleXor_83_U1 ( .A(n_zz_io_c_2_27[2]), .B(u_2_1[6]), .Z(
        simpleXor_83_port_z) );
endmodule

