
module CINI ( io_a_0, io_a_1, io_a_2, io_a_3, io_b_0, io_b_1, io_b_2, io_b_3, 
        io_c_0, io_c_1, io_c_2, io_c_3, io_rand, clk, reset );
  input [4:0] io_a_0;
  input [4:0] io_a_1;
  input [4:0] io_a_2;
  input [4:0] io_a_3;
  input [4:0] io_b_0;
  input [4:0] io_b_1;
  input [4:0] io_b_2;
  input [4:0] io_b_3;
  output [4:0] io_c_0;
  output [4:0] io_c_1;
  output [4:0] io_c_2;
  output [4:0] io_c_3;
  input [5:0] io_rand;
  input clk, reset;
  wire   simpleNot_60_port_z, simpleNot_61_port_z, simpleNot_62_port_z,
         simpleNot_63_port_z, simpleNot_64_port_z, simpleNot_65_port_z,
         simpleNot_66_port_z, simpleNot_67_port_z, simpleNot_68_port_z,
         simpleNot_69_port_z, simpleNot_70_port_z, simpleNot_71_port_z,
         simpleNot_72_port_z, simpleNot_73_port_z, simpleNot_74_port_z,
         simpleNot_75_port_z, simpleNot_76_port_z, simpleNot_77_port_z,
         simpleNot_78_port_z, simpleNot_79_port_z, simpleNot_80_port_z,
         simpleNot_81_port_z, simpleNot_82_port_z, simpleNot_83_port_z,
         simpleNot_84_port_z, simpleNot_85_port_z, simpleNot_86_port_z,
         simpleNot_87_port_z, simpleNot_88_port_z, simpleNot_89_port_z,
         simpleNot_90_port_z, simpleNot_91_port_z, simpleNot_92_port_z,
         simpleNot_93_port_z, simpleNot_94_port_z, simpleNot_95_port_z,
         simpleNot_96_port_z, simpleNot_97_port_z, simpleNot_98_port_z,
         simpleNot_99_port_z, simpleNot_100_port_z, simpleNot_101_port_z,
         simpleNot_102_port_z, simpleNot_103_port_z, simpleNot_104_port_z,
         simpleNot_105_port_z, simpleNot_106_port_z, simpleNot_107_port_z,
         simpleNot_108_port_z, simpleNot_109_port_z, simpleNot_110_port_z,
         simpleNot_111_port_z, simpleNot_112_port_z, simpleNot_113_port_z,
         simpleNot_114_port_z, simpleNot_115_port_z, simpleNot_116_port_z,
         simpleNot_117_port_z, simpleNot_118_port_z, simpleNot_119_port_z,
         simpleXor_60_port_z, simpleXor_61_port_z, simpleXor_62_port_z,
         simpleXor_63_port_z, simpleXor_64_port_z, simpleXor_65_port_z,
         simpleXor_66_port_z, simpleXor_67_port_z, simpleXor_68_port_z,
         simpleXor_69_port_z, simpleXor_70_port_z, simpleXor_71_port_z,
         simpleXor_72_port_z, simpleXor_73_port_z, simpleXor_74_port_z,
         simpleXor_75_port_z, simpleXor_76_port_z, simpleXor_77_port_z,
         simpleXor_78_port_z, simpleXor_79_port_z, simpleXor_80_port_z,
         simpleXor_81_port_z, simpleXor_82_port_z, simpleXor_83_port_z,
         simpleXor_84_port_z, simpleXor_85_port_z, simpleXor_86_port_z,
         simpleXor_87_port_z, simpleXor_88_port_z, simpleXor_89_port_z,
         simpleXor_90_port_z, simpleXor_91_port_z, simpleXor_92_port_z,
         simpleXor_93_port_z, simpleXor_94_port_z, simpleXor_95_port_z,
         simpleXor_96_port_z, simpleXor_97_port_z, simpleXor_98_port_z,
         simpleXor_99_port_z, simpleXor_100_port_z, simpleXor_101_port_z,
         simpleXor_102_port_z, simpleXor_103_port_z, simpleXor_104_port_z,
         simpleXor_105_port_z, simpleXor_106_port_z, simpleXor_107_port_z,
         simpleXor_108_port_z, simpleXor_109_port_z, simpleXor_110_port_z,
         simpleXor_111_port_z, simpleXor_112_port_z, simpleXor_113_port_z,
         simpleXor_114_port_z, simpleXor_115_port_z, simpleXor_116_port_z,
         simpleXor_117_port_z, simpleXor_118_port_z, simpleXor_119_port_z,
         n_zz_io_c_0_0_, n_zz_io_c_1_0_, n_zz_io_c_2_0_, n_zz_io_c_3_0_,
         n_zz_io_c_0_5_0_, n_zz_io_c_1_5_0_, n_zz_io_c_2_5_0_,
         n_zz_io_c_3_5_0_, n_zz_io_c_0_10_0_, n_zz_io_c_1_10_0_,
         n_zz_io_c_2_10_0_, n_zz_io_c_3_10_0_, n_zz_io_c_0_15_0_,
         n_zz_io_c_1_15_0_, n_zz_io_c_2_15_0_, n_zz_io_c_3_15_0_,
         n_zz_io_c_0_20_0_, n_zz_io_c_1_20_0_, n_zz_io_c_2_20_0_,
         n_zz_io_c_3_20_0_, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11,
         N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, cor_maj_119_port_o,
         cor_maj_118_port_o, cor_maj_117_port_o, cor_maj_116_port_o,
         cor_maj_115_port_o, cor_maj_114_port_o, cor_maj_113_port_o,
         cor_maj_112_port_o, cor_maj_111_port_o, cor_maj_110_port_o,
         cor_maj_109_port_o, cor_maj_108_port_o, cor_maj_107_port_o,
         cor_maj_106_port_o, cor_maj_105_port_o, cor_maj_104_port_o,
         cor_maj_103_port_o, cor_maj_102_port_o, cor_maj_101_port_o,
         cor_maj_100_port_o, cor_maj_99_port_o, cor_maj_98_port_o,
         cor_maj_97_port_o, cor_maj_96_port_o, cor_maj_95_port_o,
         cor_maj_94_port_o, cor_maj_93_port_o, cor_maj_92_port_o,
         cor_maj_91_port_o, cor_maj_90_port_o, cor_maj_89_port_o,
         cor_maj_88_port_o, cor_maj_87_port_o, cor_maj_86_port_o,
         cor_maj_85_port_o, cor_maj_84_port_o, cor_maj_83_port_o,
         cor_maj_82_port_o, cor_maj_81_port_o, cor_maj_80_port_o,
         cor_maj_79_port_o, cor_maj_78_port_o, cor_maj_77_port_o,
         cor_maj_76_port_o, cor_maj_75_port_o, cor_maj_74_port_o,
         cor_maj_73_port_o, cor_maj_72_port_o, cor_maj_71_port_o,
         cor_maj_70_port_o, cor_maj_69_port_o, cor_maj_68_port_o,
         cor_maj_67_port_o, cor_maj_66_port_o, cor_maj_65_port_o,
         cor_maj_64_port_o, cor_maj_63_port_o, cor_maj_62_port_o,
         cor_maj_61_port_o, cor_maj_60_port_o, cor_maj_60_n13, cor_maj_60_n12,
         cor_maj_60_n11, cor_maj_60_n10, cor_maj_60_n9, cor_maj_60_n8,
         cor_maj_60_n7, cor_maj_60_n6, cor_maj_60_n5, cor_maj_60_n4,
         cor_maj_60_n3, cor_maj_60_n2, cor_maj_60_n1, cor_maj_61_n26,
         cor_maj_61_n25, cor_maj_61_n24, cor_maj_61_n23, cor_maj_61_n22,
         cor_maj_61_n21, cor_maj_61_n20, cor_maj_61_n19, cor_maj_61_n18,
         cor_maj_61_n17, cor_maj_61_n16, cor_maj_61_n15, cor_maj_61_n14,
         cor_maj_62_n26, cor_maj_62_n25, cor_maj_62_n24, cor_maj_62_n23,
         cor_maj_62_n22, cor_maj_62_n21, cor_maj_62_n20, cor_maj_62_n19,
         cor_maj_62_n18, cor_maj_62_n17, cor_maj_62_n16, cor_maj_62_n15,
         cor_maj_62_n14, cor_maj_63_n26, cor_maj_63_n25, cor_maj_63_n24,
         cor_maj_63_n23, cor_maj_63_n22, cor_maj_63_n21, cor_maj_63_n20,
         cor_maj_63_n19, cor_maj_63_n18, cor_maj_63_n17, cor_maj_63_n16,
         cor_maj_63_n15, cor_maj_63_n14, cor_maj_64_n26, cor_maj_64_n25,
         cor_maj_64_n24, cor_maj_64_n23, cor_maj_64_n22, cor_maj_64_n21,
         cor_maj_64_n20, cor_maj_64_n19, cor_maj_64_n18, cor_maj_64_n17,
         cor_maj_64_n16, cor_maj_64_n15, cor_maj_64_n14, cor_maj_65_n26,
         cor_maj_65_n25, cor_maj_65_n24, cor_maj_65_n23, cor_maj_65_n22,
         cor_maj_65_n21, cor_maj_65_n20, cor_maj_65_n19, cor_maj_65_n18,
         cor_maj_65_n17, cor_maj_65_n16, cor_maj_65_n15, cor_maj_65_n14,
         cor_maj_66_n26, cor_maj_66_n25, cor_maj_66_n24, cor_maj_66_n23,
         cor_maj_66_n22, cor_maj_66_n21, cor_maj_66_n20, cor_maj_66_n19,
         cor_maj_66_n18, cor_maj_66_n17, cor_maj_66_n16, cor_maj_66_n15,
         cor_maj_66_n14, cor_maj_67_n26, cor_maj_67_n25, cor_maj_67_n24,
         cor_maj_67_n23, cor_maj_67_n22, cor_maj_67_n21, cor_maj_67_n20,
         cor_maj_67_n19, cor_maj_67_n18, cor_maj_67_n17, cor_maj_67_n16,
         cor_maj_67_n15, cor_maj_67_n14, cor_maj_68_n26, cor_maj_68_n25,
         cor_maj_68_n24, cor_maj_68_n23, cor_maj_68_n22, cor_maj_68_n21,
         cor_maj_68_n20, cor_maj_68_n19, cor_maj_68_n18, cor_maj_68_n17,
         cor_maj_68_n16, cor_maj_68_n15, cor_maj_68_n14, cor_maj_69_n26,
         cor_maj_69_n25, cor_maj_69_n24, cor_maj_69_n23, cor_maj_69_n22,
         cor_maj_69_n21, cor_maj_69_n20, cor_maj_69_n19, cor_maj_69_n18,
         cor_maj_69_n17, cor_maj_69_n16, cor_maj_69_n15, cor_maj_69_n14,
         cor_maj_70_n26, cor_maj_70_n25, cor_maj_70_n24, cor_maj_70_n23,
         cor_maj_70_n22, cor_maj_70_n21, cor_maj_70_n20, cor_maj_70_n19,
         cor_maj_70_n18, cor_maj_70_n17, cor_maj_70_n16, cor_maj_70_n15,
         cor_maj_70_n14, cor_maj_71_n26, cor_maj_71_n25, cor_maj_71_n24,
         cor_maj_71_n23, cor_maj_71_n22, cor_maj_71_n21, cor_maj_71_n20,
         cor_maj_71_n19, cor_maj_71_n18, cor_maj_71_n17, cor_maj_71_n16,
         cor_maj_71_n15, cor_maj_71_n14, cor_maj_72_n26, cor_maj_72_n25,
         cor_maj_72_n24, cor_maj_72_n23, cor_maj_72_n22, cor_maj_72_n21,
         cor_maj_72_n20, cor_maj_72_n19, cor_maj_72_n18, cor_maj_72_n17,
         cor_maj_72_n16, cor_maj_72_n15, cor_maj_72_n14, cor_maj_73_n26,
         cor_maj_73_n25, cor_maj_73_n24, cor_maj_73_n23, cor_maj_73_n22,
         cor_maj_73_n21, cor_maj_73_n20, cor_maj_73_n19, cor_maj_73_n18,
         cor_maj_73_n17, cor_maj_73_n16, cor_maj_73_n15, cor_maj_73_n14,
         cor_maj_74_n26, cor_maj_74_n25, cor_maj_74_n24, cor_maj_74_n23,
         cor_maj_74_n22, cor_maj_74_n21, cor_maj_74_n20, cor_maj_74_n19,
         cor_maj_74_n18, cor_maj_74_n17, cor_maj_74_n16, cor_maj_74_n15,
         cor_maj_74_n14, cor_maj_75_n26, cor_maj_75_n25, cor_maj_75_n24,
         cor_maj_75_n23, cor_maj_75_n22, cor_maj_75_n21, cor_maj_75_n20,
         cor_maj_75_n19, cor_maj_75_n18, cor_maj_75_n17, cor_maj_75_n16,
         cor_maj_75_n15, cor_maj_75_n14, cor_maj_76_n26, cor_maj_76_n25,
         cor_maj_76_n24, cor_maj_76_n23, cor_maj_76_n22, cor_maj_76_n21,
         cor_maj_76_n20, cor_maj_76_n19, cor_maj_76_n18, cor_maj_76_n17,
         cor_maj_76_n16, cor_maj_76_n15, cor_maj_76_n14, cor_maj_77_n26,
         cor_maj_77_n25, cor_maj_77_n24, cor_maj_77_n23, cor_maj_77_n22,
         cor_maj_77_n21, cor_maj_77_n20, cor_maj_77_n19, cor_maj_77_n18,
         cor_maj_77_n17, cor_maj_77_n16, cor_maj_77_n15, cor_maj_77_n14,
         cor_maj_78_n26, cor_maj_78_n25, cor_maj_78_n24, cor_maj_78_n23,
         cor_maj_78_n22, cor_maj_78_n21, cor_maj_78_n20, cor_maj_78_n19,
         cor_maj_78_n18, cor_maj_78_n17, cor_maj_78_n16, cor_maj_78_n15,
         cor_maj_78_n14, cor_maj_79_n26, cor_maj_79_n25, cor_maj_79_n24,
         cor_maj_79_n23, cor_maj_79_n22, cor_maj_79_n21, cor_maj_79_n20,
         cor_maj_79_n19, cor_maj_79_n18, cor_maj_79_n17, cor_maj_79_n16,
         cor_maj_79_n15, cor_maj_79_n14, cor_maj_80_n26, cor_maj_80_n25,
         cor_maj_80_n24, cor_maj_80_n23, cor_maj_80_n22, cor_maj_80_n21,
         cor_maj_80_n20, cor_maj_80_n19, cor_maj_80_n18, cor_maj_80_n17,
         cor_maj_80_n16, cor_maj_80_n15, cor_maj_80_n14, cor_maj_81_n26,
         cor_maj_81_n25, cor_maj_81_n24, cor_maj_81_n23, cor_maj_81_n22,
         cor_maj_81_n21, cor_maj_81_n20, cor_maj_81_n19, cor_maj_81_n18,
         cor_maj_81_n17, cor_maj_81_n16, cor_maj_81_n15, cor_maj_81_n14,
         cor_maj_82_n26, cor_maj_82_n25, cor_maj_82_n24, cor_maj_82_n23,
         cor_maj_82_n22, cor_maj_82_n21, cor_maj_82_n20, cor_maj_82_n19,
         cor_maj_82_n18, cor_maj_82_n17, cor_maj_82_n16, cor_maj_82_n15,
         cor_maj_82_n14, cor_maj_83_n26, cor_maj_83_n25, cor_maj_83_n24,
         cor_maj_83_n23, cor_maj_83_n22, cor_maj_83_n21, cor_maj_83_n20,
         cor_maj_83_n19, cor_maj_83_n18, cor_maj_83_n17, cor_maj_83_n16,
         cor_maj_83_n15, cor_maj_83_n14, cor_maj_84_n26, cor_maj_84_n25,
         cor_maj_84_n24, cor_maj_84_n23, cor_maj_84_n22, cor_maj_84_n21,
         cor_maj_84_n20, cor_maj_84_n19, cor_maj_84_n18, cor_maj_84_n17,
         cor_maj_84_n16, cor_maj_84_n15, cor_maj_84_n14, cor_maj_85_n26,
         cor_maj_85_n25, cor_maj_85_n24, cor_maj_85_n23, cor_maj_85_n22,
         cor_maj_85_n21, cor_maj_85_n20, cor_maj_85_n19, cor_maj_85_n18,
         cor_maj_85_n17, cor_maj_85_n16, cor_maj_85_n15, cor_maj_85_n14,
         cor_maj_86_n26, cor_maj_86_n25, cor_maj_86_n24, cor_maj_86_n23,
         cor_maj_86_n22, cor_maj_86_n21, cor_maj_86_n20, cor_maj_86_n19,
         cor_maj_86_n18, cor_maj_86_n17, cor_maj_86_n16, cor_maj_86_n15,
         cor_maj_86_n14, cor_maj_87_n26, cor_maj_87_n25, cor_maj_87_n24,
         cor_maj_87_n23, cor_maj_87_n22, cor_maj_87_n21, cor_maj_87_n20,
         cor_maj_87_n19, cor_maj_87_n18, cor_maj_87_n17, cor_maj_87_n16,
         cor_maj_87_n15, cor_maj_87_n14, cor_maj_88_n26, cor_maj_88_n25,
         cor_maj_88_n24, cor_maj_88_n23, cor_maj_88_n22, cor_maj_88_n21,
         cor_maj_88_n20, cor_maj_88_n19, cor_maj_88_n18, cor_maj_88_n17,
         cor_maj_88_n16, cor_maj_88_n15, cor_maj_88_n14, cor_maj_89_n26,
         cor_maj_89_n25, cor_maj_89_n24, cor_maj_89_n23, cor_maj_89_n22,
         cor_maj_89_n21, cor_maj_89_n20, cor_maj_89_n19, cor_maj_89_n18,
         cor_maj_89_n17, cor_maj_89_n16, cor_maj_89_n15, cor_maj_89_n14,
         cor_maj_90_n26, cor_maj_90_n25, cor_maj_90_n24, cor_maj_90_n23,
         cor_maj_90_n22, cor_maj_90_n21, cor_maj_90_n20, cor_maj_90_n19,
         cor_maj_90_n18, cor_maj_90_n17, cor_maj_90_n16, cor_maj_90_n15,
         cor_maj_90_n14, cor_maj_91_n26, cor_maj_91_n25, cor_maj_91_n24,
         cor_maj_91_n23, cor_maj_91_n22, cor_maj_91_n21, cor_maj_91_n20,
         cor_maj_91_n19, cor_maj_91_n18, cor_maj_91_n17, cor_maj_91_n16,
         cor_maj_91_n15, cor_maj_91_n14, cor_maj_92_n26, cor_maj_92_n25,
         cor_maj_92_n24, cor_maj_92_n23, cor_maj_92_n22, cor_maj_92_n21,
         cor_maj_92_n20, cor_maj_92_n19, cor_maj_92_n18, cor_maj_92_n17,
         cor_maj_92_n16, cor_maj_92_n15, cor_maj_92_n14, cor_maj_93_n26,
         cor_maj_93_n25, cor_maj_93_n24, cor_maj_93_n23, cor_maj_93_n22,
         cor_maj_93_n21, cor_maj_93_n20, cor_maj_93_n19, cor_maj_93_n18,
         cor_maj_93_n17, cor_maj_93_n16, cor_maj_93_n15, cor_maj_93_n14,
         cor_maj_94_n26, cor_maj_94_n25, cor_maj_94_n24, cor_maj_94_n23,
         cor_maj_94_n22, cor_maj_94_n21, cor_maj_94_n20, cor_maj_94_n19,
         cor_maj_94_n18, cor_maj_94_n17, cor_maj_94_n16, cor_maj_94_n15,
         cor_maj_94_n14, cor_maj_95_n26, cor_maj_95_n25, cor_maj_95_n24,
         cor_maj_95_n23, cor_maj_95_n22, cor_maj_95_n21, cor_maj_95_n20,
         cor_maj_95_n19, cor_maj_95_n18, cor_maj_95_n17, cor_maj_95_n16,
         cor_maj_95_n15, cor_maj_95_n14, cor_maj_96_n26, cor_maj_96_n25,
         cor_maj_96_n24, cor_maj_96_n23, cor_maj_96_n22, cor_maj_96_n21,
         cor_maj_96_n20, cor_maj_96_n19, cor_maj_96_n18, cor_maj_96_n17,
         cor_maj_96_n16, cor_maj_96_n15, cor_maj_96_n14, cor_maj_97_n26,
         cor_maj_97_n25, cor_maj_97_n24, cor_maj_97_n23, cor_maj_97_n22,
         cor_maj_97_n21, cor_maj_97_n20, cor_maj_97_n19, cor_maj_97_n18,
         cor_maj_97_n17, cor_maj_97_n16, cor_maj_97_n15, cor_maj_97_n14,
         cor_maj_98_n26, cor_maj_98_n25, cor_maj_98_n24, cor_maj_98_n23,
         cor_maj_98_n22, cor_maj_98_n21, cor_maj_98_n20, cor_maj_98_n19,
         cor_maj_98_n18, cor_maj_98_n17, cor_maj_98_n16, cor_maj_98_n15,
         cor_maj_98_n14, cor_maj_99_n26, cor_maj_99_n25, cor_maj_99_n24,
         cor_maj_99_n23, cor_maj_99_n22, cor_maj_99_n21, cor_maj_99_n20,
         cor_maj_99_n19, cor_maj_99_n18, cor_maj_99_n17, cor_maj_99_n16,
         cor_maj_99_n15, cor_maj_99_n14, cor_maj_100_n26, cor_maj_100_n25,
         cor_maj_100_n24, cor_maj_100_n23, cor_maj_100_n22, cor_maj_100_n21,
         cor_maj_100_n20, cor_maj_100_n19, cor_maj_100_n18, cor_maj_100_n17,
         cor_maj_100_n16, cor_maj_100_n15, cor_maj_100_n14, cor_maj_101_n26,
         cor_maj_101_n25, cor_maj_101_n24, cor_maj_101_n23, cor_maj_101_n22,
         cor_maj_101_n21, cor_maj_101_n20, cor_maj_101_n19, cor_maj_101_n18,
         cor_maj_101_n17, cor_maj_101_n16, cor_maj_101_n15, cor_maj_101_n14,
         cor_maj_102_n26, cor_maj_102_n25, cor_maj_102_n24, cor_maj_102_n23,
         cor_maj_102_n22, cor_maj_102_n21, cor_maj_102_n20, cor_maj_102_n19,
         cor_maj_102_n18, cor_maj_102_n17, cor_maj_102_n16, cor_maj_102_n15,
         cor_maj_102_n14, cor_maj_103_n26, cor_maj_103_n25, cor_maj_103_n24,
         cor_maj_103_n23, cor_maj_103_n22, cor_maj_103_n21, cor_maj_103_n20,
         cor_maj_103_n19, cor_maj_103_n18, cor_maj_103_n17, cor_maj_103_n16,
         cor_maj_103_n15, cor_maj_103_n14, cor_maj_104_n26, cor_maj_104_n25,
         cor_maj_104_n24, cor_maj_104_n23, cor_maj_104_n22, cor_maj_104_n21,
         cor_maj_104_n20, cor_maj_104_n19, cor_maj_104_n18, cor_maj_104_n17,
         cor_maj_104_n16, cor_maj_104_n15, cor_maj_104_n14, cor_maj_105_n26,
         cor_maj_105_n25, cor_maj_105_n24, cor_maj_105_n23, cor_maj_105_n22,
         cor_maj_105_n21, cor_maj_105_n20, cor_maj_105_n19, cor_maj_105_n18,
         cor_maj_105_n17, cor_maj_105_n16, cor_maj_105_n15, cor_maj_105_n14,
         cor_maj_106_n26, cor_maj_106_n25, cor_maj_106_n24, cor_maj_106_n23,
         cor_maj_106_n22, cor_maj_106_n21, cor_maj_106_n20, cor_maj_106_n19,
         cor_maj_106_n18, cor_maj_106_n17, cor_maj_106_n16, cor_maj_106_n15,
         cor_maj_106_n14, cor_maj_107_n26, cor_maj_107_n25, cor_maj_107_n24,
         cor_maj_107_n23, cor_maj_107_n22, cor_maj_107_n21, cor_maj_107_n20,
         cor_maj_107_n19, cor_maj_107_n18, cor_maj_107_n17, cor_maj_107_n16,
         cor_maj_107_n15, cor_maj_107_n14, cor_maj_108_n26, cor_maj_108_n25,
         cor_maj_108_n24, cor_maj_108_n23, cor_maj_108_n22, cor_maj_108_n21,
         cor_maj_108_n20, cor_maj_108_n19, cor_maj_108_n18, cor_maj_108_n17,
         cor_maj_108_n16, cor_maj_108_n15, cor_maj_108_n14, cor_maj_109_n26,
         cor_maj_109_n25, cor_maj_109_n24, cor_maj_109_n23, cor_maj_109_n22,
         cor_maj_109_n21, cor_maj_109_n20, cor_maj_109_n19, cor_maj_109_n18,
         cor_maj_109_n17, cor_maj_109_n16, cor_maj_109_n15, cor_maj_109_n14,
         cor_maj_110_n26, cor_maj_110_n25, cor_maj_110_n24, cor_maj_110_n23,
         cor_maj_110_n22, cor_maj_110_n21, cor_maj_110_n20, cor_maj_110_n19,
         cor_maj_110_n18, cor_maj_110_n17, cor_maj_110_n16, cor_maj_110_n15,
         cor_maj_110_n14, cor_maj_111_n26, cor_maj_111_n25, cor_maj_111_n24,
         cor_maj_111_n23, cor_maj_111_n22, cor_maj_111_n21, cor_maj_111_n20,
         cor_maj_111_n19, cor_maj_111_n18, cor_maj_111_n17, cor_maj_111_n16,
         cor_maj_111_n15, cor_maj_111_n14, cor_maj_112_n26, cor_maj_112_n25,
         cor_maj_112_n24, cor_maj_112_n23, cor_maj_112_n22, cor_maj_112_n21,
         cor_maj_112_n20, cor_maj_112_n19, cor_maj_112_n18, cor_maj_112_n17,
         cor_maj_112_n16, cor_maj_112_n15, cor_maj_112_n14, cor_maj_113_n26,
         cor_maj_113_n25, cor_maj_113_n24, cor_maj_113_n23, cor_maj_113_n22,
         cor_maj_113_n21, cor_maj_113_n20, cor_maj_113_n19, cor_maj_113_n18,
         cor_maj_113_n17, cor_maj_113_n16, cor_maj_113_n15, cor_maj_113_n14,
         cor_maj_114_n26, cor_maj_114_n25, cor_maj_114_n24, cor_maj_114_n23,
         cor_maj_114_n22, cor_maj_114_n21, cor_maj_114_n20, cor_maj_114_n19,
         cor_maj_114_n18, cor_maj_114_n17, cor_maj_114_n16, cor_maj_114_n15,
         cor_maj_114_n14, cor_maj_115_n26, cor_maj_115_n25, cor_maj_115_n24,
         cor_maj_115_n23, cor_maj_115_n22, cor_maj_115_n21, cor_maj_115_n20,
         cor_maj_115_n19, cor_maj_115_n18, cor_maj_115_n17, cor_maj_115_n16,
         cor_maj_115_n15, cor_maj_115_n14, cor_maj_116_n26, cor_maj_116_n25,
         cor_maj_116_n24, cor_maj_116_n23, cor_maj_116_n22, cor_maj_116_n21,
         cor_maj_116_n20, cor_maj_116_n19, cor_maj_116_n18, cor_maj_116_n17,
         cor_maj_116_n16, cor_maj_116_n15, cor_maj_116_n14, cor_maj_117_n26,
         cor_maj_117_n25, cor_maj_117_n24, cor_maj_117_n23, cor_maj_117_n22,
         cor_maj_117_n21, cor_maj_117_n20, cor_maj_117_n19, cor_maj_117_n18,
         cor_maj_117_n17, cor_maj_117_n16, cor_maj_117_n15, cor_maj_117_n14,
         cor_maj_118_n26, cor_maj_118_n25, cor_maj_118_n24, cor_maj_118_n23,
         cor_maj_118_n22, cor_maj_118_n21, cor_maj_118_n20, cor_maj_118_n19,
         cor_maj_118_n18, cor_maj_118_n17, cor_maj_118_n16, cor_maj_118_n15,
         cor_maj_118_n14, cor_maj_119_n26, cor_maj_119_n25, cor_maj_119_n24,
         cor_maj_119_n23, cor_maj_119_n22, cor_maj_119_n21, cor_maj_119_n20,
         cor_maj_119_n19, cor_maj_119_n18, cor_maj_119_n17, cor_maj_119_n16,
         cor_maj_119_n15, cor_maj_119_n14;
  wire   [4:0] v_1_0_1;
  wire   [4:0] v_1_0_2;
  wire   [4:0] v_1_0_3;
  wire   [4:0] v_1_1_0;
  wire   [4:0] v_1_1_2;
  wire   [4:0] v_1_1_3;
  wire   [4:0] v_1_2_0;
  wire   [4:0] v_1_2_1;
  wire   [4:0] v_1_2_3;
  wire   [4:0] v_1_3_0;
  wire   [4:0] v_1_3_1;
  wire   [4:0] v_1_3_2;
  wire   [4:0] cor_port_v_0_1;
  wire   [4:0] cor_port_v_0_2;
  wire   [4:0] cor_port_v_0_3;
  wire   [4:0] cor_port_v_1_0;
  wire   [4:0] cor_port_v_1_2;
  wire   [4:0] cor_port_v_1_3;
  wire   [4:0] cor_port_v_2_0;
  wire   [4:0] cor_port_v_2_1;
  wire   [4:0] cor_port_v_2_3;
  wire   [4:0] cor_port_v_3_0;
  wire   [4:0] cor_port_v_3_1;
  wire   [4:0] cor_port_v_3_2;
  wire   [3:1] n_zz_io_c_0_4;
  wire   [4:0] u_0_1;
  wire   [4:0] u_0_2;
  wire   [4:0] u_0_3;
  wire   [3:1] n_zz_io_c_1_4;
  wire   [4:0] u_1_0;
  wire   [4:0] u_1_2;
  wire   [4:0] u_1_3;
  wire   [3:1] n_zz_io_c_2_4;
  wire   [4:0] u_2_0;
  wire   [4:0] u_2_1;
  wire   [4:0] u_2_3;
  wire   [3:1] n_zz_io_c_3_4;
  wire   [4:0] u_3_0;
  wire   [4:0] u_3_1;
  wire   [4:0] u_3_2;
  wire   [3:1] n_zz_io_c_0_9;
  wire   [3:1] n_zz_io_c_1_9;
  wire   [3:1] n_zz_io_c_2_9;
  wire   [3:1] n_zz_io_c_3_9;
  wire   [3:1] n_zz_io_c_0_14;
  wire   [3:1] n_zz_io_c_1_14;
  wire   [3:1] n_zz_io_c_2_14;
  wire   [3:1] n_zz_io_c_3_14;
  wire   [3:1] n_zz_io_c_0_19;
  wire   [3:1] n_zz_io_c_1_19;
  wire   [3:1] n_zz_io_c_2_19;
  wire   [3:1] n_zz_io_c_3_19;
  wire   [3:1] n_zz_io_c_0_24;
  wire   [3:1] n_zz_io_c_1_24;
  wire   [3:1] n_zz_io_c_2_24;
  wire   [3:1] n_zz_io_c_3_24;
  wire   [4:0] rand_reg_0;
  wire   [4:0] rand_reg_1;
  wire   [4:0] rand_reg_2;
  wire   [4:0] rand_reg_6;
  wire   [4:0] rand_reg_3;
  wire   [4:0] rand_reg_4;
  wire   [4:0] rand_reg_7;
  wire   [4:0] rand_reg_9;
  wire   [4:0] rand_reg_5;
  wire   [4:0] rand_reg_8;
  wire   [4:0] rand_reg_10;
  wire   [4:0] rand_reg_11;
  wire   [4:0] b_reg_0;
  wire   [4:0] b_reg_1;
  wire   [4:0] b_reg_2;
  wire   [4:0] b_reg_3;

  DFF_X1 b_reg_1_reg_4_ ( .D(io_b_1[4]), .CK(clk), .Q(b_reg_1[4]), .QN() );
  DFF_X1 b_reg_1_reg_3_ ( .D(io_b_1[3]), .CK(clk), .Q(b_reg_1[3]), .QN() );
  DFF_X1 b_reg_1_reg_2_ ( .D(io_b_1[2]), .CK(clk), .Q(b_reg_1[2]), .QN() );
  DFF_X1 b_reg_1_reg_1_ ( .D(io_b_1[1]), .CK(clk), .Q(b_reg_1[1]), .QN() );
  DFF_X1 b_reg_1_reg_0_ ( .D(io_b_1[0]), .CK(clk), .Q(b_reg_1[0]), .QN() );
  DFF_X1 b_reg_2_reg_4_ ( .D(io_b_2[4]), .CK(clk), .Q(b_reg_2[4]), .QN() );
  DFF_X1 b_reg_2_reg_3_ ( .D(io_b_2[3]), .CK(clk), .Q(b_reg_2[3]), .QN() );
  DFF_X1 b_reg_2_reg_2_ ( .D(io_b_2[2]), .CK(clk), .Q(b_reg_2[2]), .QN() );
  DFF_X1 b_reg_2_reg_1_ ( .D(io_b_2[1]), .CK(clk), .Q(b_reg_2[1]), .QN() );
  DFF_X1 b_reg_2_reg_0_ ( .D(io_b_2[0]), .CK(clk), .Q(b_reg_2[0]), .QN() );
  DFF_X1 b_reg_3_reg_4_ ( .D(io_b_3[4]), .CK(clk), .Q(b_reg_3[4]), .QN() );
  DFF_X1 b_reg_3_reg_3_ ( .D(io_b_3[3]), .CK(clk), .Q(b_reg_3[3]), .QN() );
  DFF_X1 b_reg_3_reg_2_ ( .D(io_b_3[2]), .CK(clk), .Q(b_reg_3[2]), .QN() );
  DFF_X1 b_reg_3_reg_1_ ( .D(io_b_3[1]), .CK(clk), .Q(b_reg_3[1]), .QN() );
  DFF_X1 b_reg_3_reg_0_ ( .D(io_b_3[0]), .CK(clk), .Q(b_reg_3[0]), .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_3_ ( .D(N139), .CK(clk), .Q(n_zz_io_c_3_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_2_ ( .D(N138), .CK(clk), .Q(n_zz_io_c_3_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_1_ ( .D(N137), .CK(clk), .Q(n_zz_io_c_3_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_24_reg_0_ ( .D(N136), .CK(clk), .Q(n_zz_io_c_3_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_3_ ( .D(N135), .CK(clk), .Q(n_zz_io_c_2_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_2_ ( .D(N134), .CK(clk), .Q(n_zz_io_c_2_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_1_ ( .D(N133), .CK(clk), .Q(n_zz_io_c_2_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_24_reg_0_ ( .D(N132), .CK(clk), .Q(n_zz_io_c_2_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_3_ ( .D(N131), .CK(clk), .Q(n_zz_io_c_1_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_2_ ( .D(N130), .CK(clk), .Q(n_zz_io_c_1_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_1_ ( .D(N129), .CK(clk), .Q(n_zz_io_c_1_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_24_reg_0_ ( .D(N128), .CK(clk), .Q(n_zz_io_c_1_20_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_3_ ( .D(N127), .CK(clk), .Q(n_zz_io_c_0_24[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_2_ ( .D(N126), .CK(clk), .Q(n_zz_io_c_0_24[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_1_ ( .D(N125), .CK(clk), .Q(n_zz_io_c_0_24[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_3_ ( .D(N123), .CK(clk), .Q(n_zz_io_c_3_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_2_ ( .D(N122), .CK(clk), .Q(n_zz_io_c_3_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_1_ ( .D(N121), .CK(clk), .Q(n_zz_io_c_3_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_19_reg_0_ ( .D(N120), .CK(clk), .Q(n_zz_io_c_3_15_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_3_ ( .D(N119), .CK(clk), .Q(n_zz_io_c_2_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_2_ ( .D(N118), .CK(clk), .Q(n_zz_io_c_2_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_1_ ( .D(N117), .CK(clk), .Q(n_zz_io_c_2_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_19_reg_0_ ( .D(N116), .CK(clk), .Q(n_zz_io_c_2_15_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_3_ ( .D(N115), .CK(clk), .Q(n_zz_io_c_1_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_2_ ( .D(N114), .CK(clk), .Q(n_zz_io_c_1_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_1_ ( .D(N113), .CK(clk), .Q(n_zz_io_c_1_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_19_reg_0_ ( .D(N112), .CK(clk), .Q(n_zz_io_c_1_15_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_3_ ( .D(N111), .CK(clk), .Q(n_zz_io_c_0_19[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_2_ ( .D(N110), .CK(clk), .Q(n_zz_io_c_0_19[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_1_ ( .D(N109), .CK(clk), .Q(n_zz_io_c_0_19[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_3_ ( .D(N107), .CK(clk), .Q(n_zz_io_c_3_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_2_ ( .D(N106), .CK(clk), .Q(n_zz_io_c_3_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_1_ ( .D(N105), .CK(clk), .Q(n_zz_io_c_3_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_14_reg_0_ ( .D(N104), .CK(clk), .Q(n_zz_io_c_3_10_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_3_ ( .D(N103), .CK(clk), .Q(n_zz_io_c_2_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_2_ ( .D(N102), .CK(clk), .Q(n_zz_io_c_2_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_1_ ( .D(N101), .CK(clk), .Q(n_zz_io_c_2_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_2_14_reg_0_ ( .D(N100), .CK(clk), .Q(n_zz_io_c_2_10_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_3_ ( .D(N99), .CK(clk), .Q(n_zz_io_c_1_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_2_ ( .D(N98), .CK(clk), .Q(n_zz_io_c_1_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_1_ ( .D(N97), .CK(clk), .Q(n_zz_io_c_1_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_0_ ( .D(N96), .CK(clk), .Q(n_zz_io_c_1_10_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_3_ ( .D(N95), .CK(clk), .Q(n_zz_io_c_0_14[3]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_2_ ( .D(N94), .CK(clk), .Q(n_zz_io_c_0_14[2]), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_1_ ( .D(N93), .CK(clk), .Q(n_zz_io_c_0_14[1]), 
        .QN() );
  DFF_X1 u_zz_io_c_3_9_reg_3_ ( .D(N91), .CK(clk), .Q(n_zz_io_c_3_9[3]), .QN()
         );
  DFF_X1 u_zz_io_c_3_9_reg_2_ ( .D(N90), .CK(clk), .Q(n_zz_io_c_3_9[2]), .QN()
         );
  DFF_X1 u_zz_io_c_3_9_reg_1_ ( .D(N89), .CK(clk), .Q(n_zz_io_c_3_9[1]), .QN()
         );
  DFF_X1 u_zz_io_c_3_9_reg_0_ ( .D(N88), .CK(clk), .Q(n_zz_io_c_3_5_0_), .QN()
         );
  DFF_X1 u_zz_io_c_2_9_reg_3_ ( .D(N87), .CK(clk), .Q(n_zz_io_c_2_9[3]), .QN()
         );
  DFF_X1 u_zz_io_c_2_9_reg_2_ ( .D(N86), .CK(clk), .Q(n_zz_io_c_2_9[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_9_reg_1_ ( .D(N85), .CK(clk), .Q(n_zz_io_c_2_9[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_9_reg_0_ ( .D(N84), .CK(clk), .Q(n_zz_io_c_2_5_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_9_reg_3_ ( .D(N83), .CK(clk), .Q(n_zz_io_c_1_9[3]), .QN()
         );
  DFF_X1 u_zz_io_c_1_9_reg_2_ ( .D(N82), .CK(clk), .Q(n_zz_io_c_1_9[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_9_reg_1_ ( .D(N81), .CK(clk), .Q(n_zz_io_c_1_9[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_9_reg_0_ ( .D(N80), .CK(clk), .Q(n_zz_io_c_1_5_0_), .QN()
         );
  DFF_X1 rand_reg_9_reg_4_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[4]), 
        .QN() );
  DFF_X1 u_2_1_reg_4_ ( .D(N55), .CK(clk), .Q(u_2_1[4]), .QN() );
  DFF_X1 rand_reg_9_reg_3_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[3]), 
        .QN() );
  DFF_X1 u_2_1_reg_3_ ( .D(N43), .CK(clk), .Q(u_2_1[3]), .QN() );
  DFF_X1 rand_reg_9_reg_2_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[2]), 
        .QN() );
  DFF_X1 u_2_1_reg_2_ ( .D(N31), .CK(clk), .Q(u_2_1[2]), .QN() );
  DFF_X1 rand_reg_9_reg_1_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[1]), 
        .QN() );
  DFF_X1 u_2_1_reg_1_ ( .D(N19), .CK(clk), .Q(u_2_1[1]), .QN() );
  DFF_X1 rand_reg_9_reg_0_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_9[0]), 
        .QN() );
  DFF_X1 u_2_1_reg_0_ ( .D(N7), .CK(clk), .Q(u_2_1[0]), .QN() );
  DFF_X1 u_zz_io_c_0_9_reg_3_ ( .D(N79), .CK(clk), .Q(n_zz_io_c_0_9[3]), .QN()
         );
  DFF_X1 u_zz_io_c_0_9_reg_2_ ( .D(N78), .CK(clk), .Q(n_zz_io_c_0_9[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_9_reg_1_ ( .D(N77), .CK(clk), .Q(n_zz_io_c_0_9[1]), .QN()
         );
  DFF_X1 rand_reg_1_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[4]), 
        .QN() );
  DFF_X1 u_0_2_reg_4_ ( .D(N49), .CK(clk), .Q(u_0_2[4]), .QN() );
  DFF_X1 rand_reg_1_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[3]), 
        .QN() );
  DFF_X1 u_0_2_reg_3_ ( .D(N37), .CK(clk), .Q(u_0_2[3]), .QN() );
  DFF_X1 rand_reg_1_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[2]), 
        .QN() );
  DFF_X1 u_0_2_reg_2_ ( .D(N25), .CK(clk), .Q(u_0_2[2]), .QN() );
  DFF_X1 rand_reg_1_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[1]), 
        .QN() );
  DFF_X1 u_0_2_reg_1_ ( .D(N13), .CK(clk), .Q(u_0_2[1]), .QN() );
  DFF_X1 rand_reg_1_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_1[0]), 
        .QN() );
  DFF_X1 u_0_2_reg_0_ ( .D(N1), .CK(clk), .Q(u_0_2[0]), .QN() );
  DFF_X1 u_zz_io_c_3_4_reg_3_ ( .D(N75), .CK(clk), .Q(n_zz_io_c_3_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_3_4_reg_2_ ( .D(N74), .CK(clk), .Q(n_zz_io_c_3_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_3_4_reg_1_ ( .D(N73), .CK(clk), .Q(n_zz_io_c_3_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_3_4_reg_0_ ( .D(N72), .CK(clk), .Q(n_zz_io_c_3_0_), .QN()
         );
  DFF_X1 rand_reg_0_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[4]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[3]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[2]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[1]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[0]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_4_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[4]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_3_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[3]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_2_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[2]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_1_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[1]), 
        .QN() );
  DFF_X1 rand_reg_11_reg_0_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_11[0]), 
        .QN() );
  DFF_X1 rand_reg_6_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[4]), 
        .QN() );
  DFF_X1 u_1_0_reg_4_ ( .D(N51), .CK(clk), .Q(u_1_0[4]), .QN() );
  DFF_X1 rand_reg_6_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[3]), 
        .QN() );
  DFF_X1 u_1_0_reg_3_ ( .D(N39), .CK(clk), .Q(u_1_0[3]), .QN() );
  DFF_X1 rand_reg_6_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[2]), 
        .QN() );
  DFF_X1 u_1_0_reg_2_ ( .D(N27), .CK(clk), .Q(u_1_0[2]), .QN() );
  DFF_X1 rand_reg_6_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[1]), 
        .QN() );
  DFF_X1 u_1_0_reg_1_ ( .D(N15), .CK(clk), .Q(u_1_0[1]), .QN() );
  DFF_X1 rand_reg_6_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_6[0]), 
        .QN() );
  DFF_X1 u_1_0_reg_0_ ( .D(N3), .CK(clk), .Q(u_1_0[0]), .QN() );
  DFF_X1 rand_reg_7_reg_4_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[4]), 
        .QN() );
  DFF_X1 u_2_0_reg_4_ ( .D(N54), .CK(clk), .Q(u_2_0[4]), .QN() );
  DFF_X1 rand_reg_7_reg_3_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[3]), 
        .QN() );
  DFF_X1 u_2_0_reg_3_ ( .D(N42), .CK(clk), .Q(u_2_0[3]), .QN() );
  DFF_X1 rand_reg_7_reg_2_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[2]), 
        .QN() );
  DFF_X1 u_2_0_reg_2_ ( .D(N30), .CK(clk), .Q(u_2_0[2]), .QN() );
  DFF_X1 rand_reg_7_reg_1_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[1]), 
        .QN() );
  DFF_X1 u_2_0_reg_1_ ( .D(N18), .CK(clk), .Q(u_2_0[1]), .QN() );
  DFF_X1 rand_reg_7_reg_0_ ( .D(io_rand[1]), .CK(clk), .Q(rand_reg_7[0]), 
        .QN() );
  DFF_X1 u_2_0_reg_0_ ( .D(N6), .CK(clk), .Q(u_2_0[0]), .QN() );
  DFF_X1 u_0_1_reg_4_ ( .D(N48), .CK(clk), .Q(u_0_1[4]), .QN() );
  DFF_X1 u_0_1_reg_3_ ( .D(N36), .CK(clk), .Q(u_0_1[3]), .QN() );
  DFF_X1 u_0_1_reg_2_ ( .D(N24), .CK(clk), .Q(u_0_1[2]), .QN() );
  DFF_X1 u_0_1_reg_1_ ( .D(N12), .CK(clk), .Q(u_0_1[1]), .QN() );
  DFF_X1 u_0_1_reg_0_ ( .D(N0), .CK(clk), .Q(u_0_1[0]), .QN() );
  DFF_X1 u_zz_io_c_2_4_reg_3_ ( .D(N71), .CK(clk), .Q(n_zz_io_c_2_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_2_ ( .D(N70), .CK(clk), .Q(n_zz_io_c_2_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_1_ ( .D(N69), .CK(clk), .Q(n_zz_io_c_2_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_2_4_reg_0_ ( .D(N68), .CK(clk), .Q(n_zz_io_c_2_0_), .QN()
         );
  DFF_X1 rand_reg_2_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[4]), 
        .QN() );
  DFF_X1 u_0_3_reg_4_ ( .D(N50), .CK(clk), .Q(u_0_3[4]), .QN() );
  DFF_X1 rand_reg_2_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[3]), 
        .QN() );
  DFF_X1 u_0_3_reg_3_ ( .D(N38), .CK(clk), .Q(u_0_3[3]), .QN() );
  DFF_X1 rand_reg_2_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[2]), 
        .QN() );
  DFF_X1 u_0_3_reg_2_ ( .D(N26), .CK(clk), .Q(u_0_3[2]), .QN() );
  DFF_X1 rand_reg_2_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[1]), 
        .QN() );
  DFF_X1 u_0_3_reg_1_ ( .D(N14), .CK(clk), .Q(u_0_3[1]), .QN() );
  DFF_X1 rand_reg_2_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_2[0]), 
        .QN() );
  DFF_X1 u_0_3_reg_0_ ( .D(N2), .CK(clk), .Q(u_0_3[0]), .QN() );
  DFF_X1 rand_reg_8_reg_4_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[4]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_3_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[3]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_2_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[2]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_1_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[1]), 
        .QN() );
  DFF_X1 rand_reg_8_reg_0_ ( .D(io_rand[2]), .CK(clk), .Q(rand_reg_8[0]), 
        .QN() );
  DFF_X1 rand_reg_3_reg_4_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[4]), 
        .QN() );
  DFF_X1 u_1_2_reg_4_ ( .D(N52), .CK(clk), .Q(u_1_2[4]), .QN() );
  DFF_X1 rand_reg_3_reg_3_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[3]), 
        .QN() );
  DFF_X1 u_1_2_reg_3_ ( .D(N40), .CK(clk), .Q(u_1_2[3]), .QN() );
  DFF_X1 rand_reg_3_reg_2_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[2]), 
        .QN() );
  DFF_X1 u_1_2_reg_2_ ( .D(N28), .CK(clk), .Q(u_1_2[2]), .QN() );
  DFF_X1 rand_reg_3_reg_1_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[1]), 
        .QN() );
  DFF_X1 u_1_2_reg_1_ ( .D(N16), .CK(clk), .Q(u_1_2[1]), .QN() );
  DFF_X1 rand_reg_3_reg_0_ ( .D(io_rand[3]), .CK(clk), .Q(rand_reg_3[0]), 
        .QN() );
  DFF_X1 u_1_2_reg_0_ ( .D(N4), .CK(clk), .Q(u_1_2[0]), .QN() );
  DFF_X1 rand_reg_4_reg_4_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[4]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_3_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[3]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_2_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[2]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_1_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[1]), 
        .QN() );
  DFF_X1 rand_reg_4_reg_0_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_4[0]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_4_reg_3_ ( .D(N67), .CK(clk), .Q(n_zz_io_c_1_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_2_ ( .D(N66), .CK(clk), .Q(n_zz_io_c_1_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_1_ ( .D(N65), .CK(clk), .Q(n_zz_io_c_1_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_1_4_reg_0_ ( .D(N64), .CK(clk), .Q(n_zz_io_c_1_0_), .QN()
         );
  DFF_X1 rand_reg_10_reg_4_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[4]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_3_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[3]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_2_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[2]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_1_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[1]), 
        .QN() );
  DFF_X1 rand_reg_10_reg_0_ ( .D(io_rand[4]), .CK(clk), .Q(rand_reg_10[0]), 
        .QN() );
  DFF_X1 rand_reg_5_reg_4_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[4]), 
        .QN() );
  DFF_X1 u_2_3_reg_4_ ( .D(N56), .CK(clk), .Q(u_2_3[4]), .QN() );
  DFF_X1 rand_reg_5_reg_3_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[3]), 
        .QN() );
  DFF_X1 u_2_3_reg_3_ ( .D(N44), .CK(clk), .Q(u_2_3[3]), .QN() );
  DFF_X1 rand_reg_5_reg_2_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[2]), 
        .QN() );
  DFF_X1 u_2_3_reg_2_ ( .D(N32), .CK(clk), .Q(u_2_3[2]), .QN() );
  DFF_X1 rand_reg_5_reg_1_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[1]), 
        .QN() );
  DFF_X1 u_2_3_reg_1_ ( .D(N20), .CK(clk), .Q(u_2_3[1]), .QN() );
  DFF_X1 rand_reg_5_reg_0_ ( .D(io_rand[5]), .CK(clk), .Q(rand_reg_5[0]), 
        .QN() );
  DFF_X1 u_2_3_reg_0_ ( .D(N8), .CK(clk), .Q(u_2_3[0]), .QN() );
  DFF_X1 b_reg_0_reg_4_ ( .D(io_b_0[4]), .CK(clk), .Q(b_reg_0[4]), .QN() );
  DFF_X1 u_zz_io_c_0_24_reg_0_ ( .D(N124), .CK(clk), .Q(n_zz_io_c_0_20_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_3_ ( .D(io_b_0[3]), .CK(clk), .Q(b_reg_0[3]), .QN() );
  DFF_X1 u_zz_io_c_0_19_reg_0_ ( .D(N108), .CK(clk), .Q(n_zz_io_c_0_15_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_2_ ( .D(io_b_0[2]), .CK(clk), .Q(b_reg_0[2]), .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_0_ ( .D(N92), .CK(clk), .Q(n_zz_io_c_0_10_0_), 
        .QN() );
  DFF_X1 b_reg_0_reg_1_ ( .D(io_b_0[1]), .CK(clk), .Q(b_reg_0[1]), .QN() );
  DFF_X1 u_zz_io_c_0_9_reg_0_ ( .D(N76), .CK(clk), .Q(n_zz_io_c_0_5_0_), .QN()
         );
  DFF_X1 b_reg_0_reg_0_ ( .D(io_b_0[0]), .CK(clk), .Q(b_reg_0[0]), .QN() );
  DFF_X1 u_1_3_reg_4_ ( .D(N53), .CK(clk), .Q(u_1_3[4]), .QN() );
  DFF_X1 u_1_3_reg_3_ ( .D(N41), .CK(clk), .Q(u_1_3[3]), .QN() );
  DFF_X1 u_1_3_reg_2_ ( .D(N29), .CK(clk), .Q(u_1_3[2]), .QN() );
  DFF_X1 u_1_3_reg_1_ ( .D(N17), .CK(clk), .Q(u_1_3[1]), .QN() );
  DFF_X1 u_1_3_reg_0_ ( .D(N5), .CK(clk), .Q(u_1_3[0]), .QN() );
  DFF_X1 u_zz_io_c_0_4_reg_3_ ( .D(N63), .CK(clk), .Q(n_zz_io_c_0_4[3]), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_2_ ( .D(N62), .CK(clk), .Q(n_zz_io_c_0_4[2]), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_1_ ( .D(N61), .CK(clk), .Q(n_zz_io_c_0_4[1]), .QN()
         );
  DFF_X1 u_zz_io_c_0_4_reg_0_ ( .D(N60), .CK(clk), .Q(n_zz_io_c_0_0_), .QN()
         );
  DFF_X1 u_3_2_reg_4_ ( .D(N59), .CK(clk), .Q(u_3_2[4]), .QN() );
  DFF_X1 u_3_2_reg_3_ ( .D(N47), .CK(clk), .Q(u_3_2[3]), .QN() );
  DFF_X1 u_3_2_reg_2_ ( .D(N35), .CK(clk), .Q(u_3_2[2]), .QN() );
  DFF_X1 u_3_2_reg_1_ ( .D(N23), .CK(clk), .Q(u_3_2[1]), .QN() );
  DFF_X1 u_3_2_reg_0_ ( .D(N11), .CK(clk), .Q(u_3_2[0]), .QN() );
  DFF_X1 u_3_1_reg_4_ ( .D(N58), .CK(clk), .Q(u_3_1[4]), .QN() );
  DFF_X1 u_3_1_reg_3_ ( .D(N46), .CK(clk), .Q(u_3_1[3]), .QN() );
  DFF_X1 u_3_1_reg_2_ ( .D(N34), .CK(clk), .Q(u_3_1[2]), .QN() );
  DFF_X1 u_3_1_reg_1_ ( .D(N22), .CK(clk), .Q(u_3_1[1]), .QN() );
  DFF_X1 u_3_1_reg_0_ ( .D(N10), .CK(clk), .Q(u_3_1[0]), .QN() );
  DFF_X1 u_3_0_reg_4_ ( .D(N57), .CK(clk), .Q(u_3_0[4]), .QN() );
  DFF_X1 u_3_0_reg_3_ ( .D(N45), .CK(clk), .Q(u_3_0[3]), .QN() );
  DFF_X1 u_3_0_reg_2_ ( .D(N33), .CK(clk), .Q(u_3_0[2]), .QN() );
  DFF_X1 u_3_0_reg_1_ ( .D(N21), .CK(clk), .Q(u_3_0[1]), .QN() );
  DFF_X1 u_3_0_reg_0_ ( .D(N9), .CK(clk), .Q(u_3_0[0]), .QN() );
  XOR2_X2 U3 ( .A(io_rand[5]), .B(io_b_2[4]), .Z(v_1_3_2[4]) );
  XOR2_X2 U4 ( .A(io_rand[5]), .B(io_b_2[3]), .Z(v_1_3_2[3]) );
  XOR2_X2 U5 ( .A(io_rand[5]), .B(io_b_2[2]), .Z(v_1_3_2[2]) );
  XOR2_X2 U6 ( .A(io_rand[5]), .B(io_b_2[1]), .Z(v_1_3_2[1]) );
  XOR2_X2 U7 ( .A(io_rand[5]), .B(io_b_2[0]), .Z(v_1_3_2[0]) );
  XOR2_X2 U8 ( .A(io_rand[4]), .B(io_b_1[4]), .Z(v_1_3_1[4]) );
  XOR2_X2 U9 ( .A(io_rand[4]), .B(io_b_1[3]), .Z(v_1_3_1[3]) );
  XOR2_X2 U10 ( .A(io_rand[4]), .B(io_b_1[2]), .Z(v_1_3_1[2]) );
  XOR2_X2 U11 ( .A(io_rand[4]), .B(io_b_1[1]), .Z(v_1_3_1[1]) );
  XOR2_X2 U12 ( .A(io_rand[4]), .B(io_b_1[0]), .Z(v_1_3_1[0]) );
  XOR2_X2 U13 ( .A(io_rand[2]), .B(io_b_0[4]), .Z(v_1_3_0[4]) );
  XOR2_X2 U14 ( .A(io_rand[2]), .B(io_b_0[3]), .Z(v_1_3_0[3]) );
  XOR2_X2 U15 ( .A(io_rand[2]), .B(io_b_0[2]), .Z(v_1_3_0[2]) );
  XOR2_X2 U16 ( .A(io_rand[2]), .B(io_b_0[1]), .Z(v_1_3_0[1]) );
  XOR2_X2 U17 ( .A(io_rand[2]), .B(io_b_0[0]), .Z(v_1_3_0[0]) );
  XOR2_X2 U18 ( .A(io_rand[5]), .B(io_b_3[4]), .Z(v_1_2_3[4]) );
  XOR2_X2 U19 ( .A(io_rand[5]), .B(io_b_3[3]), .Z(v_1_2_3[3]) );
  XOR2_X2 U20 ( .A(io_rand[5]), .B(io_b_3[2]), .Z(v_1_2_3[2]) );
  XOR2_X2 U21 ( .A(io_rand[5]), .B(io_b_3[1]), .Z(v_1_2_3[1]) );
  XOR2_X2 U22 ( .A(io_rand[5]), .B(io_b_3[0]), .Z(v_1_2_3[0]) );
  XOR2_X2 U23 ( .A(io_rand[3]), .B(io_b_1[4]), .Z(v_1_2_1[4]) );
  XOR2_X2 U24 ( .A(io_rand[3]), .B(io_b_1[3]), .Z(v_1_2_1[3]) );
  XOR2_X2 U25 ( .A(io_rand[3]), .B(io_b_1[2]), .Z(v_1_2_1[2]) );
  XOR2_X2 U26 ( .A(io_rand[3]), .B(io_b_1[1]), .Z(v_1_2_1[1]) );
  XOR2_X2 U27 ( .A(io_rand[3]), .B(io_b_1[0]), .Z(v_1_2_1[0]) );
  XOR2_X2 U28 ( .A(io_rand[1]), .B(io_b_0[4]), .Z(v_1_2_0[4]) );
  XOR2_X2 U29 ( .A(io_rand[1]), .B(io_b_0[3]), .Z(v_1_2_0[3]) );
  XOR2_X2 U30 ( .A(io_rand[1]), .B(io_b_0[2]), .Z(v_1_2_0[2]) );
  XOR2_X2 U31 ( .A(io_rand[1]), .B(io_b_0[1]), .Z(v_1_2_0[1]) );
  XOR2_X2 U32 ( .A(io_rand[1]), .B(io_b_0[0]), .Z(v_1_2_0[0]) );
  XOR2_X2 U33 ( .A(io_rand[4]), .B(io_b_3[4]), .Z(v_1_1_3[4]) );
  XOR2_X2 U34 ( .A(io_rand[4]), .B(io_b_3[3]), .Z(v_1_1_3[3]) );
  XOR2_X2 U35 ( .A(io_rand[4]), .B(io_b_3[2]), .Z(v_1_1_3[2]) );
  XOR2_X2 U36 ( .A(io_rand[4]), .B(io_b_3[1]), .Z(v_1_1_3[1]) );
  XOR2_X2 U37 ( .A(io_rand[4]), .B(io_b_3[0]), .Z(v_1_1_3[0]) );
  XOR2_X2 U38 ( .A(io_rand[3]), .B(io_b_2[4]), .Z(v_1_1_2[4]) );
  XOR2_X2 U39 ( .A(io_rand[3]), .B(io_b_2[3]), .Z(v_1_1_2[3]) );
  XOR2_X2 U40 ( .A(io_rand[3]), .B(io_b_2[2]), .Z(v_1_1_2[2]) );
  XOR2_X2 U41 ( .A(io_rand[3]), .B(io_b_2[1]), .Z(v_1_1_2[1]) );
  XOR2_X2 U42 ( .A(io_rand[3]), .B(io_b_2[0]), .Z(v_1_1_2[0]) );
  XOR2_X2 U43 ( .A(io_rand[0]), .B(io_b_0[4]), .Z(v_1_1_0[4]) );
  XOR2_X2 U44 ( .A(io_rand[0]), .B(io_b_0[3]), .Z(v_1_1_0[3]) );
  XOR2_X2 U45 ( .A(io_rand[0]), .B(io_b_0[2]), .Z(v_1_1_0[2]) );
  XOR2_X2 U46 ( .A(io_rand[0]), .B(io_b_0[1]), .Z(v_1_1_0[1]) );
  XOR2_X2 U47 ( .A(io_rand[0]), .B(io_b_0[0]), .Z(v_1_1_0[0]) );
  XOR2_X2 U48 ( .A(io_rand[2]), .B(io_b_3[4]), .Z(v_1_0_3[4]) );
  XOR2_X2 U49 ( .A(io_rand[2]), .B(io_b_3[3]), .Z(v_1_0_3[3]) );
  XOR2_X2 U50 ( .A(io_rand[2]), .B(io_b_3[2]), .Z(v_1_0_3[2]) );
  XOR2_X2 U51 ( .A(io_rand[2]), .B(io_b_3[1]), .Z(v_1_0_3[1]) );
  XOR2_X2 U52 ( .A(io_rand[2]), .B(io_b_3[0]), .Z(v_1_0_3[0]) );
  XOR2_X2 U53 ( .A(io_rand[1]), .B(io_b_2[4]), .Z(v_1_0_2[4]) );
  XOR2_X2 U54 ( .A(io_rand[1]), .B(io_b_2[3]), .Z(v_1_0_2[3]) );
  XOR2_X2 U55 ( .A(io_rand[1]), .B(io_b_2[2]), .Z(v_1_0_2[2]) );
  XOR2_X2 U56 ( .A(io_rand[1]), .B(io_b_2[1]), .Z(v_1_0_2[1]) );
  XOR2_X2 U57 ( .A(io_rand[1]), .B(io_b_2[0]), .Z(v_1_0_2[0]) );
  XOR2_X2 U58 ( .A(io_rand[0]), .B(io_b_1[4]), .Z(v_1_0_1[4]) );
  XOR2_X2 U59 ( .A(io_rand[0]), .B(io_b_1[3]), .Z(v_1_0_1[3]) );
  XOR2_X2 U60 ( .A(io_rand[0]), .B(io_b_1[2]), .Z(v_1_0_1[2]) );
  XOR2_X2 U61 ( .A(io_rand[0]), .B(io_b_1[1]), .Z(v_1_0_1[1]) );
  XOR2_X2 U62 ( .A(io_rand[0]), .B(io_b_1[0]), .Z(v_1_0_1[0]) );
  AND2_X1 U263 ( .A1(b_reg_0[0]), .A2(io_a_0[0]), .ZN(N60) );
  AND2_X1 U264 ( .A1(cor_port_v_0_1[0]), .A2(io_a_0[0]), .ZN(N61) );
  AND2_X1 U265 ( .A1(cor_port_v_0_2[0]), .A2(io_a_0[0]), .ZN(N62) );
  AND2_X1 U266 ( .A1(b_reg_0[1]), .A2(io_a_0[1]), .ZN(N76) );
  AND2_X1 U267 ( .A1(b_reg_0[2]), .A2(io_a_0[2]), .ZN(N92) );
  AND2_X1 U268 ( .A1(b_reg_0[3]), .A2(io_a_0[3]), .ZN(N108) );
  AND2_X1 U269 ( .A1(b_reg_0[4]), .A2(io_a_0[4]), .ZN(N124) );
  AND2_X1 U270 ( .A1(b_reg_1[0]), .A2(io_a_1[0]), .ZN(N64) );
  AND2_X1 U271 ( .A1(cor_port_v_1_0[0]), .A2(io_a_1[0]), .ZN(N65) );
  AND2_X1 U272 ( .A1(cor_port_v_1_2[0]), .A2(io_a_1[0]), .ZN(N66) );
  AND2_X1 U273 ( .A1(b_reg_2[0]), .A2(io_a_2[0]), .ZN(N68) );
  AND2_X1 U274 ( .A1(cor_port_v_2_0[0]), .A2(io_a_2[0]), .ZN(N69) );
  AND2_X1 U275 ( .A1(cor_port_v_2_1[0]), .A2(io_a_2[0]), .ZN(N70) );
  AND2_X1 U276 ( .A1(b_reg_3[0]), .A2(io_a_3[0]), .ZN(N72) );
  AND2_X1 U277 ( .A1(cor_port_v_3_0[0]), .A2(io_a_3[0]), .ZN(N73) );
  AND2_X1 U278 ( .A1(cor_port_v_3_1[0]), .A2(io_a_3[0]), .ZN(N74) );
  AND2_X1 U279 ( .A1(cor_port_v_0_1[1]), .A2(io_a_0[1]), .ZN(N77) );
  AND2_X1 U280 ( .A1(cor_port_v_0_2[1]), .A2(io_a_0[1]), .ZN(N78) );
  AND2_X1 U281 ( .A1(b_reg_1[1]), .A2(io_a_1[1]), .ZN(N80) );
  AND2_X1 U282 ( .A1(cor_port_v_1_0[1]), .A2(io_a_1[1]), .ZN(N81) );
  AND2_X1 U283 ( .A1(cor_port_v_1_2[1]), .A2(io_a_1[1]), .ZN(N82) );
  AND2_X1 U284 ( .A1(b_reg_2[1]), .A2(io_a_2[1]), .ZN(N84) );
  AND2_X1 U285 ( .A1(cor_port_v_2_0[1]), .A2(io_a_2[1]), .ZN(N85) );
  AND2_X1 U286 ( .A1(cor_port_v_2_1[1]), .A2(io_a_2[1]), .ZN(N86) );
  AND2_X1 U287 ( .A1(b_reg_3[1]), .A2(io_a_3[1]), .ZN(N88) );
  AND2_X1 U288 ( .A1(cor_port_v_3_0[1]), .A2(io_a_3[1]), .ZN(N89) );
  AND2_X1 U289 ( .A1(cor_port_v_3_1[1]), .A2(io_a_3[1]), .ZN(N90) );
  AND2_X1 U290 ( .A1(cor_port_v_0_1[2]), .A2(io_a_0[2]), .ZN(N93) );
  AND2_X1 U291 ( .A1(cor_port_v_0_2[2]), .A2(io_a_0[2]), .ZN(N94) );
  AND2_X1 U292 ( .A1(b_reg_1[2]), .A2(io_a_1[2]), .ZN(N96) );
  AND2_X1 U293 ( .A1(cor_port_v_1_0[2]), .A2(io_a_1[2]), .ZN(N97) );
  AND2_X1 U294 ( .A1(cor_port_v_1_2[2]), .A2(io_a_1[2]), .ZN(N98) );
  AND2_X1 U295 ( .A1(b_reg_2[2]), .A2(io_a_2[2]), .ZN(N100) );
  AND2_X1 U296 ( .A1(cor_port_v_2_0[2]), .A2(io_a_2[2]), .ZN(N101) );
  AND2_X1 U297 ( .A1(cor_port_v_2_1[2]), .A2(io_a_2[2]), .ZN(N102) );
  AND2_X1 U298 ( .A1(b_reg_3[2]), .A2(io_a_3[2]), .ZN(N104) );
  AND2_X1 U299 ( .A1(cor_port_v_3_0[2]), .A2(io_a_3[2]), .ZN(N105) );
  AND2_X1 U300 ( .A1(cor_port_v_3_1[2]), .A2(io_a_3[2]), .ZN(N106) );
  AND2_X1 U301 ( .A1(cor_port_v_0_1[3]), .A2(io_a_0[3]), .ZN(N109) );
  AND2_X1 U302 ( .A1(cor_port_v_0_2[3]), .A2(io_a_0[3]), .ZN(N110) );
  AND2_X1 U303 ( .A1(b_reg_1[3]), .A2(io_a_1[3]), .ZN(N112) );
  AND2_X1 U304 ( .A1(cor_port_v_1_0[3]), .A2(io_a_1[3]), .ZN(N113) );
  AND2_X1 U305 ( .A1(cor_port_v_1_2[3]), .A2(io_a_1[3]), .ZN(N114) );
  AND2_X1 U306 ( .A1(b_reg_2[3]), .A2(io_a_2[3]), .ZN(N116) );
  AND2_X1 U307 ( .A1(cor_port_v_2_0[3]), .A2(io_a_2[3]), .ZN(N117) );
  AND2_X1 U308 ( .A1(cor_port_v_2_1[3]), .A2(io_a_2[3]), .ZN(N118) );
  AND2_X1 U309 ( .A1(b_reg_3[3]), .A2(io_a_3[3]), .ZN(N120) );
  AND2_X1 U310 ( .A1(cor_port_v_3_0[3]), .A2(io_a_3[3]), .ZN(N121) );
  AND2_X1 U311 ( .A1(cor_port_v_3_1[3]), .A2(io_a_3[3]), .ZN(N122) );
  AND2_X1 U312 ( .A1(cor_port_v_0_1[4]), .A2(io_a_0[4]), .ZN(N125) );
  AND2_X1 U313 ( .A1(cor_port_v_0_2[4]), .A2(io_a_0[4]), .ZN(N126) );
  AND2_X1 U314 ( .A1(b_reg_1[4]), .A2(io_a_1[4]), .ZN(N128) );
  AND2_X1 U315 ( .A1(cor_port_v_1_0[4]), .A2(io_a_1[4]), .ZN(N129) );
  AND2_X1 U316 ( .A1(cor_port_v_1_2[4]), .A2(io_a_1[4]), .ZN(N130) );
  AND2_X1 U317 ( .A1(b_reg_2[4]), .A2(io_a_2[4]), .ZN(N132) );
  AND2_X1 U318 ( .A1(cor_port_v_2_0[4]), .A2(io_a_2[4]), .ZN(N133) );
  AND2_X1 U319 ( .A1(cor_port_v_2_1[4]), .A2(io_a_2[4]), .ZN(N134) );
  AND2_X1 U320 ( .A1(b_reg_3[4]), .A2(io_a_3[4]), .ZN(N136) );
  AND2_X1 U321 ( .A1(cor_port_v_3_0[4]), .A2(io_a_3[4]), .ZN(N137) );
  AND2_X1 U322 ( .A1(cor_port_v_3_1[4]), .A2(io_a_3[4]), .ZN(N138) );
  AND2_X1 U323 ( .A1(simpleNot_69_port_z), .A2(rand_reg_8[0]), .ZN(N9) );
  AND2_X1 U324 ( .A1(simpleNot_81_port_z), .A2(rand_reg_8[1]), .ZN(N21) );
  AND2_X1 U325 ( .A1(simpleNot_93_port_z), .A2(rand_reg_8[2]), .ZN(N33) );
  AND2_X1 U326 ( .A1(simpleNot_105_port_z), .A2(rand_reg_8[3]), .ZN(N45) );
  AND2_X1 U327 ( .A1(simpleNot_117_port_z), .A2(rand_reg_8[4]), .ZN(N57) );
  AND2_X1 U328 ( .A1(simpleNot_70_port_z), .A2(rand_reg_10[0]), .ZN(N10) );
  AND2_X1 U329 ( .A1(simpleNot_82_port_z), .A2(rand_reg_10[1]), .ZN(N22) );
  AND2_X1 U330 ( .A1(simpleNot_94_port_z), .A2(rand_reg_10[2]), .ZN(N34) );
  AND2_X1 U331 ( .A1(simpleNot_106_port_z), .A2(rand_reg_10[3]), .ZN(N46) );
  AND2_X1 U332 ( .A1(simpleNot_118_port_z), .A2(rand_reg_10[4]), .ZN(N58) );
  AND2_X1 U333 ( .A1(simpleNot_71_port_z), .A2(rand_reg_11[0]), .ZN(N11) );
  AND2_X1 U334 ( .A1(simpleNot_83_port_z), .A2(rand_reg_11[1]), .ZN(N23) );
  AND2_X1 U335 ( .A1(simpleNot_95_port_z), .A2(rand_reg_11[2]), .ZN(N35) );
  AND2_X1 U336 ( .A1(simpleNot_107_port_z), .A2(rand_reg_11[3]), .ZN(N47) );
  AND2_X1 U337 ( .A1(simpleNot_119_port_z), .A2(rand_reg_11[4]), .ZN(N59) );
  AND2_X1 U338 ( .A1(io_a_0[0]), .A2(cor_port_v_0_3[0]), .ZN(N63) );
  AND2_X1 U339 ( .A1(simpleNot_65_port_z), .A2(rand_reg_4[0]), .ZN(N5) );
  AND2_X1 U340 ( .A1(simpleNot_77_port_z), .A2(rand_reg_4[1]), .ZN(N17) );
  AND2_X1 U341 ( .A1(simpleNot_89_port_z), .A2(rand_reg_4[2]), .ZN(N29) );
  AND2_X1 U342 ( .A1(simpleNot_101_port_z), .A2(rand_reg_4[3]), .ZN(N41) );
  AND2_X1 U343 ( .A1(simpleNot_113_port_z), .A2(rand_reg_4[4]), .ZN(N53) );
  AND2_X1 U344 ( .A1(simpleNot_68_port_z), .A2(rand_reg_5[0]), .ZN(N8) );
  AND2_X1 U345 ( .A1(simpleNot_80_port_z), .A2(rand_reg_5[1]), .ZN(N20) );
  AND2_X1 U346 ( .A1(simpleNot_92_port_z), .A2(rand_reg_5[2]), .ZN(N32) );
  AND2_X1 U347 ( .A1(simpleNot_104_port_z), .A2(rand_reg_5[3]), .ZN(N44) );
  AND2_X1 U348 ( .A1(simpleNot_116_port_z), .A2(rand_reg_5[4]), .ZN(N56) );
  AND2_X1 U349 ( .A1(io_a_1[0]), .A2(cor_port_v_1_3[0]), .ZN(N67) );
  AND2_X1 U350 ( .A1(simpleNot_64_port_z), .A2(rand_reg_3[0]), .ZN(N4) );
  AND2_X1 U351 ( .A1(simpleNot_76_port_z), .A2(rand_reg_3[1]), .ZN(N16) );
  AND2_X1 U352 ( .A1(simpleNot_88_port_z), .A2(rand_reg_3[2]), .ZN(N28) );
  AND2_X1 U353 ( .A1(simpleNot_100_port_z), .A2(rand_reg_3[3]), .ZN(N40) );
  AND2_X1 U354 ( .A1(simpleNot_112_port_z), .A2(rand_reg_3[4]), .ZN(N52) );
  AND2_X1 U355 ( .A1(simpleNot_62_port_z), .A2(rand_reg_2[0]), .ZN(N2) );
  AND2_X1 U356 ( .A1(simpleNot_74_port_z), .A2(rand_reg_2[1]), .ZN(N14) );
  AND2_X1 U357 ( .A1(simpleNot_86_port_z), .A2(rand_reg_2[2]), .ZN(N26) );
  AND2_X1 U358 ( .A1(simpleNot_98_port_z), .A2(rand_reg_2[3]), .ZN(N38) );
  AND2_X1 U359 ( .A1(simpleNot_110_port_z), .A2(rand_reg_2[4]), .ZN(N50) );
  AND2_X1 U360 ( .A1(io_a_2[0]), .A2(cor_port_v_2_3[0]), .ZN(N71) );
  AND2_X1 U361 ( .A1(simpleNot_60_port_z), .A2(rand_reg_0[0]), .ZN(N0) );
  AND2_X1 U362 ( .A1(simpleNot_72_port_z), .A2(rand_reg_0[1]), .ZN(N12) );
  AND2_X1 U363 ( .A1(simpleNot_84_port_z), .A2(rand_reg_0[2]), .ZN(N24) );
  AND2_X1 U364 ( .A1(simpleNot_96_port_z), .A2(rand_reg_0[3]), .ZN(N36) );
  AND2_X1 U365 ( .A1(simpleNot_108_port_z), .A2(rand_reg_0[4]), .ZN(N48) );
  AND2_X1 U366 ( .A1(simpleNot_66_port_z), .A2(rand_reg_7[0]), .ZN(N6) );
  AND2_X1 U367 ( .A1(simpleNot_78_port_z), .A2(rand_reg_7[1]), .ZN(N18) );
  AND2_X1 U368 ( .A1(simpleNot_90_port_z), .A2(rand_reg_7[2]), .ZN(N30) );
  AND2_X1 U369 ( .A1(simpleNot_102_port_z), .A2(rand_reg_7[3]), .ZN(N42) );
  AND2_X1 U370 ( .A1(simpleNot_114_port_z), .A2(rand_reg_7[4]), .ZN(N54) );
  AND2_X1 U371 ( .A1(simpleNot_63_port_z), .A2(rand_reg_6[0]), .ZN(N3) );
  AND2_X1 U372 ( .A1(simpleNot_75_port_z), .A2(rand_reg_6[1]), .ZN(N15) );
  AND2_X1 U373 ( .A1(simpleNot_87_port_z), .A2(rand_reg_6[2]), .ZN(N27) );
  AND2_X1 U374 ( .A1(simpleNot_99_port_z), .A2(rand_reg_6[3]), .ZN(N39) );
  AND2_X1 U375 ( .A1(simpleNot_111_port_z), .A2(rand_reg_6[4]), .ZN(N51) );
  AND2_X1 U376 ( .A1(io_a_3[0]), .A2(cor_port_v_3_2[0]), .ZN(N75) );
  AND2_X1 U377 ( .A1(simpleNot_61_port_z), .A2(rand_reg_1[0]), .ZN(N1) );
  AND2_X1 U378 ( .A1(simpleNot_73_port_z), .A2(rand_reg_1[1]), .ZN(N13) );
  AND2_X1 U379 ( .A1(simpleNot_85_port_z), .A2(rand_reg_1[2]), .ZN(N25) );
  AND2_X1 U380 ( .A1(simpleNot_97_port_z), .A2(rand_reg_1[3]), .ZN(N37) );
  AND2_X1 U381 ( .A1(simpleNot_109_port_z), .A2(rand_reg_1[4]), .ZN(N49) );
  AND2_X1 U382 ( .A1(io_a_0[1]), .A2(cor_port_v_0_3[1]), .ZN(N79) );
  AND2_X1 U383 ( .A1(simpleNot_67_port_z), .A2(rand_reg_9[0]), .ZN(N7) );
  AND2_X1 U384 ( .A1(simpleNot_79_port_z), .A2(rand_reg_9[1]), .ZN(N19) );
  AND2_X1 U385 ( .A1(simpleNot_91_port_z), .A2(rand_reg_9[2]), .ZN(N31) );
  AND2_X1 U386 ( .A1(simpleNot_103_port_z), .A2(rand_reg_9[3]), .ZN(N43) );
  AND2_X1 U387 ( .A1(simpleNot_115_port_z), .A2(rand_reg_9[4]), .ZN(N55) );
  AND2_X1 U388 ( .A1(io_a_1[1]), .A2(cor_port_v_1_3[1]), .ZN(N83) );
  AND2_X1 U389 ( .A1(io_a_2[1]), .A2(cor_port_v_2_3[1]), .ZN(N87) );
  AND2_X1 U390 ( .A1(io_a_3[1]), .A2(cor_port_v_3_2[1]), .ZN(N91) );
  AND2_X1 U391 ( .A1(io_a_0[2]), .A2(cor_port_v_0_3[2]), .ZN(N95) );
  AND2_X1 U392 ( .A1(io_a_1[2]), .A2(cor_port_v_1_3[2]), .ZN(N99) );
  AND2_X1 U393 ( .A1(io_a_2[2]), .A2(cor_port_v_2_3[2]), .ZN(N103) );
  AND2_X1 U394 ( .A1(io_a_3[2]), .A2(cor_port_v_3_2[2]), .ZN(N107) );
  AND2_X1 U395 ( .A1(io_a_0[3]), .A2(cor_port_v_0_3[3]), .ZN(N111) );
  AND2_X1 U396 ( .A1(io_a_1[3]), .A2(cor_port_v_1_3[3]), .ZN(N115) );
  AND2_X1 U397 ( .A1(io_a_2[3]), .A2(cor_port_v_2_3[3]), .ZN(N119) );
  AND2_X1 U398 ( .A1(io_a_3[3]), .A2(cor_port_v_3_2[3]), .ZN(N123) );
  AND2_X1 U399 ( .A1(io_a_0[4]), .A2(cor_port_v_0_3[4]), .ZN(N127) );
  AND2_X1 U400 ( .A1(io_a_1[4]), .A2(cor_port_v_1_3[4]), .ZN(N131) );
  AND2_X1 U401 ( .A1(io_a_2[4]), .A2(cor_port_v_2_3[4]), .ZN(N135) );
  AND2_X1 U402 ( .A1(io_a_3[4]), .A2(cor_port_v_3_2[4]), .ZN(N139) );
  XOR2_X1 U403 ( .A(n9), .B(n10), .Z(io_c_3[0]) );
  XNOR2_X1 U404 ( .A(simpleXor_71_port_z), .B(simpleXor_70_port_z), .ZN(n9) );
  XNOR2_X1 U405 ( .A(simpleXor_69_port_z), .B(n_zz_io_c_3_0_), .ZN(n10) );
  XOR2_X1 U406 ( .A(n7), .B(n8), .Z(io_c_3[1]) );
  XNOR2_X1 U407 ( .A(simpleXor_83_port_z), .B(simpleXor_82_port_z), .ZN(n7) );
  XNOR2_X1 U408 ( .A(simpleXor_81_port_z), .B(n_zz_io_c_3_5_0_), .ZN(n8) );
  XOR2_X1 U409 ( .A(n5), .B(n6), .Z(io_c_3[2]) );
  XNOR2_X1 U410 ( .A(simpleXor_95_port_z), .B(simpleXor_94_port_z), .ZN(n5) );
  XNOR2_X1 U411 ( .A(simpleXor_93_port_z), .B(n_zz_io_c_3_10_0_), .ZN(n6) );
  XOR2_X1 U412 ( .A(n3), .B(n4), .Z(io_c_3[3]) );
  XNOR2_X1 U413 ( .A(simpleXor_107_port_z), .B(simpleXor_106_port_z), .ZN(n3)
         );
  XNOR2_X1 U414 ( .A(simpleXor_105_port_z), .B(n_zz_io_c_3_15_0_), .ZN(n4) );
  XOR2_X1 U415 ( .A(n1), .B(n2), .Z(io_c_3[4]) );
  XNOR2_X1 U416 ( .A(simpleXor_119_port_z), .B(simpleXor_118_port_z), .ZN(n1)
         );
  XNOR2_X1 U417 ( .A(simpleXor_117_port_z), .B(n_zz_io_c_3_20_0_), .ZN(n2) );
  XOR2_X1 U418 ( .A(n19), .B(n20), .Z(io_c_2[0]) );
  XNOR2_X1 U419 ( .A(simpleXor_68_port_z), .B(simpleXor_67_port_z), .ZN(n19)
         );
  XNOR2_X1 U420 ( .A(simpleXor_66_port_z), .B(n_zz_io_c_2_0_), .ZN(n20) );
  XOR2_X1 U421 ( .A(n17), .B(n18), .Z(io_c_2[1]) );
  XNOR2_X1 U422 ( .A(simpleXor_80_port_z), .B(simpleXor_79_port_z), .ZN(n17)
         );
  XNOR2_X1 U423 ( .A(simpleXor_78_port_z), .B(n_zz_io_c_2_5_0_), .ZN(n18) );
  XOR2_X1 U424 ( .A(n15), .B(n16), .Z(io_c_2[2]) );
  XNOR2_X1 U425 ( .A(simpleXor_92_port_z), .B(simpleXor_91_port_z), .ZN(n15)
         );
  XNOR2_X1 U426 ( .A(simpleXor_90_port_z), .B(n_zz_io_c_2_10_0_), .ZN(n16) );
  XOR2_X1 U427 ( .A(n13), .B(n14), .Z(io_c_2[3]) );
  XNOR2_X1 U428 ( .A(simpleXor_104_port_z), .B(simpleXor_103_port_z), .ZN(n13)
         );
  XNOR2_X1 U429 ( .A(simpleXor_102_port_z), .B(n_zz_io_c_2_15_0_), .ZN(n14) );
  XOR2_X1 U430 ( .A(n11), .B(n12), .Z(io_c_2[4]) );
  XNOR2_X1 U431 ( .A(simpleXor_116_port_z), .B(simpleXor_115_port_z), .ZN(n11)
         );
  XNOR2_X1 U432 ( .A(simpleXor_114_port_z), .B(n_zz_io_c_2_20_0_), .ZN(n12) );
  XOR2_X1 U433 ( .A(n29), .B(n30), .Z(io_c_1[0]) );
  XNOR2_X1 U434 ( .A(simpleXor_65_port_z), .B(simpleXor_64_port_z), .ZN(n29)
         );
  XNOR2_X1 U435 ( .A(simpleXor_63_port_z), .B(n_zz_io_c_1_0_), .ZN(n30) );
  XOR2_X1 U436 ( .A(n27), .B(n28), .Z(io_c_1[1]) );
  XNOR2_X1 U437 ( .A(simpleXor_77_port_z), .B(simpleXor_76_port_z), .ZN(n27)
         );
  XNOR2_X1 U438 ( .A(simpleXor_75_port_z), .B(n_zz_io_c_1_5_0_), .ZN(n28) );
  XOR2_X1 U439 ( .A(n25), .B(n26), .Z(io_c_1[2]) );
  XNOR2_X1 U440 ( .A(simpleXor_89_port_z), .B(simpleXor_88_port_z), .ZN(n25)
         );
  XNOR2_X1 U441 ( .A(simpleXor_87_port_z), .B(n_zz_io_c_1_10_0_), .ZN(n26) );
  XOR2_X1 U442 ( .A(n23), .B(n24), .Z(io_c_1[3]) );
  XNOR2_X1 U443 ( .A(simpleXor_99_port_z), .B(simpleXor_101_port_z), .ZN(n23)
         );
  XNOR2_X1 U444 ( .A(simpleXor_100_port_z), .B(n_zz_io_c_1_15_0_), .ZN(n24) );
  XOR2_X1 U445 ( .A(n21), .B(n22), .Z(io_c_1[4]) );
  XNOR2_X1 U446 ( .A(simpleXor_113_port_z), .B(simpleXor_112_port_z), .ZN(n21)
         );
  XNOR2_X1 U447 ( .A(simpleXor_111_port_z), .B(n_zz_io_c_1_20_0_), .ZN(n22) );
  XOR2_X1 U448 ( .A(n39), .B(n40), .Z(io_c_0[0]) );
  XNOR2_X1 U449 ( .A(simpleXor_62_port_z), .B(simpleXor_61_port_z), .ZN(n39)
         );
  XNOR2_X1 U450 ( .A(simpleXor_60_port_z), .B(n_zz_io_c_0_0_), .ZN(n40) );
  XOR2_X1 U451 ( .A(n37), .B(n38), .Z(io_c_0[1]) );
  XNOR2_X1 U452 ( .A(simpleXor_74_port_z), .B(simpleXor_73_port_z), .ZN(n37)
         );
  XNOR2_X1 U453 ( .A(simpleXor_72_port_z), .B(n_zz_io_c_0_5_0_), .ZN(n38) );
  XOR2_X1 U454 ( .A(n35), .B(n36), .Z(io_c_0[2]) );
  XNOR2_X1 U455 ( .A(simpleXor_86_port_z), .B(simpleXor_85_port_z), .ZN(n35)
         );
  XNOR2_X1 U456 ( .A(simpleXor_84_port_z), .B(n_zz_io_c_0_10_0_), .ZN(n36) );
  XOR2_X1 U457 ( .A(n33), .B(n34), .Z(io_c_0[3]) );
  XNOR2_X1 U458 ( .A(simpleXor_98_port_z), .B(simpleXor_97_port_z), .ZN(n33)
         );
  XNOR2_X1 U459 ( .A(simpleXor_96_port_z), .B(n_zz_io_c_0_15_0_), .ZN(n34) );
  XOR2_X1 U460 ( .A(n31), .B(n32), .Z(io_c_0[4]) );
  XNOR2_X1 U461 ( .A(simpleXor_110_port_z), .B(simpleXor_109_port_z), .ZN(n31)
         );
  XNOR2_X1 U462 ( .A(simpleXor_108_port_z), .B(n_zz_io_c_0_20_0_), .ZN(n32) );
  INV_X1 simpleNot_60_U1 ( .A(io_a_0[0]), .ZN(simpleNot_60_port_z) );
  INV_X1 simpleNot_61_U1 ( .A(io_a_0[0]), .ZN(simpleNot_61_port_z) );
  INV_X1 simpleNot_62_U1 ( .A(io_a_0[0]), .ZN(simpleNot_62_port_z) );
  INV_X1 simpleNot_63_U1 ( .A(io_a_1[0]), .ZN(simpleNot_63_port_z) );
  INV_X1 simpleNot_64_U1 ( .A(io_a_1[0]), .ZN(simpleNot_64_port_z) );
  INV_X1 simpleNot_65_U1 ( .A(io_a_1[0]), .ZN(simpleNot_65_port_z) );
  INV_X1 simpleNot_66_U1 ( .A(io_a_2[0]), .ZN(simpleNot_66_port_z) );
  INV_X1 simpleNot_67_U1 ( .A(io_a_2[0]), .ZN(simpleNot_67_port_z) );
  INV_X1 simpleNot_68_U1 ( .A(io_a_2[0]), .ZN(simpleNot_68_port_z) );
  INV_X1 simpleNot_69_U1 ( .A(io_a_3[0]), .ZN(simpleNot_69_port_z) );
  INV_X1 simpleNot_70_U1 ( .A(io_a_3[0]), .ZN(simpleNot_70_port_z) );
  INV_X1 simpleNot_71_U1 ( .A(io_a_3[0]), .ZN(simpleNot_71_port_z) );
  INV_X1 simpleNot_72_U1 ( .A(io_a_0[1]), .ZN(simpleNot_72_port_z) );
  INV_X1 simpleNot_73_U1 ( .A(io_a_0[1]), .ZN(simpleNot_73_port_z) );
  INV_X1 simpleNot_74_U1 ( .A(io_a_0[1]), .ZN(simpleNot_74_port_z) );
  INV_X1 simpleNot_75_U1 ( .A(io_a_1[1]), .ZN(simpleNot_75_port_z) );
  INV_X1 simpleNot_76_U1 ( .A(io_a_1[1]), .ZN(simpleNot_76_port_z) );
  INV_X1 simpleNot_77_U1 ( .A(io_a_1[1]), .ZN(simpleNot_77_port_z) );
  INV_X1 simpleNot_78_U1 ( .A(io_a_2[1]), .ZN(simpleNot_78_port_z) );
  INV_X1 simpleNot_79_U1 ( .A(io_a_2[1]), .ZN(simpleNot_79_port_z) );
  INV_X1 simpleNot_80_U1 ( .A(io_a_2[1]), .ZN(simpleNot_80_port_z) );
  INV_X1 simpleNot_81_U1 ( .A(io_a_3[1]), .ZN(simpleNot_81_port_z) );
  INV_X1 simpleNot_82_U1 ( .A(io_a_3[1]), .ZN(simpleNot_82_port_z) );
  INV_X1 simpleNot_83_U1 ( .A(io_a_3[1]), .ZN(simpleNot_83_port_z) );
  INV_X1 simpleNot_84_U1 ( .A(io_a_0[2]), .ZN(simpleNot_84_port_z) );
  INV_X1 simpleNot_85_U1 ( .A(io_a_0[2]), .ZN(simpleNot_85_port_z) );
  INV_X1 simpleNot_86_U1 ( .A(io_a_0[2]), .ZN(simpleNot_86_port_z) );
  INV_X1 simpleNot_87_U1 ( .A(io_a_1[2]), .ZN(simpleNot_87_port_z) );
  INV_X1 simpleNot_88_U1 ( .A(io_a_1[2]), .ZN(simpleNot_88_port_z) );
  INV_X1 simpleNot_89_U1 ( .A(io_a_1[2]), .ZN(simpleNot_89_port_z) );
  INV_X1 simpleNot_90_U1 ( .A(io_a_2[2]), .ZN(simpleNot_90_port_z) );
  INV_X1 simpleNot_91_U1 ( .A(io_a_2[2]), .ZN(simpleNot_91_port_z) );
  INV_X1 simpleNot_92_U1 ( .A(io_a_2[2]), .ZN(simpleNot_92_port_z) );
  INV_X1 simpleNot_93_U1 ( .A(io_a_3[2]), .ZN(simpleNot_93_port_z) );
  INV_X1 simpleNot_94_U1 ( .A(io_a_3[2]), .ZN(simpleNot_94_port_z) );
  INV_X1 simpleNot_95_U1 ( .A(io_a_3[2]), .ZN(simpleNot_95_port_z) );
  INV_X1 simpleNot_96_U1 ( .A(io_a_0[3]), .ZN(simpleNot_96_port_z) );
  INV_X1 simpleNot_97_U1 ( .A(io_a_0[3]), .ZN(simpleNot_97_port_z) );
  INV_X1 simpleNot_98_U1 ( .A(io_a_0[3]), .ZN(simpleNot_98_port_z) );
  INV_X1 simpleNot_99_U1 ( .A(io_a_1[3]), .ZN(simpleNot_99_port_z) );
  INV_X1 simpleNot_100_U1 ( .A(io_a_1[3]), .ZN(simpleNot_100_port_z) );
  INV_X1 simpleNot_101_U1 ( .A(io_a_1[3]), .ZN(simpleNot_101_port_z) );
  INV_X1 simpleNot_102_U1 ( .A(io_a_2[3]), .ZN(simpleNot_102_port_z) );
  INV_X1 simpleNot_103_U1 ( .A(io_a_2[3]), .ZN(simpleNot_103_port_z) );
  INV_X1 simpleNot_104_U1 ( .A(io_a_2[3]), .ZN(simpleNot_104_port_z) );
  INV_X1 simpleNot_105_U1 ( .A(io_a_3[3]), .ZN(simpleNot_105_port_z) );
  INV_X1 simpleNot_106_U1 ( .A(io_a_3[3]), .ZN(simpleNot_106_port_z) );
  INV_X1 simpleNot_107_U1 ( .A(io_a_3[3]), .ZN(simpleNot_107_port_z) );
  INV_X1 simpleNot_108_U1 ( .A(io_a_0[4]), .ZN(simpleNot_108_port_z) );
  INV_X1 simpleNot_109_U1 ( .A(io_a_0[4]), .ZN(simpleNot_109_port_z) );
  INV_X1 simpleNot_110_U1 ( .A(io_a_0[4]), .ZN(simpleNot_110_port_z) );
  INV_X1 simpleNot_111_U1 ( .A(io_a_1[4]), .ZN(simpleNot_111_port_z) );
  INV_X1 simpleNot_112_U1 ( .A(io_a_1[4]), .ZN(simpleNot_112_port_z) );
  INV_X1 simpleNot_113_U1 ( .A(io_a_1[4]), .ZN(simpleNot_113_port_z) );
  INV_X1 simpleNot_114_U1 ( .A(io_a_2[4]), .ZN(simpleNot_114_port_z) );
  INV_X1 simpleNot_115_U1 ( .A(io_a_2[4]), .ZN(simpleNot_115_port_z) );
  INV_X1 simpleNot_116_U1 ( .A(io_a_2[4]), .ZN(simpleNot_116_port_z) );
  INV_X1 simpleNot_117_U1 ( .A(io_a_3[4]), .ZN(simpleNot_117_port_z) );
  INV_X1 simpleNot_118_U1 ( .A(io_a_3[4]), .ZN(simpleNot_118_port_z) );
  INV_X1 simpleNot_119_U1 ( .A(io_a_3[4]), .ZN(simpleNot_119_port_z) );
  DFF_X1 cor_m_3_2_reg_0_ ( .D(cor_maj_115_port_o), .CK(clk), .Q(
        cor_port_v_3_2[0]), .QN() );
  DFF_X1 cor_m_3_2_reg_1_ ( .D(cor_maj_116_port_o), .CK(clk), .Q(
        cor_port_v_3_2[1]), .QN() );
  DFF_X1 cor_m_3_2_reg_2_ ( .D(cor_maj_117_port_o), .CK(clk), .Q(
        cor_port_v_3_2[2]), .QN() );
  DFF_X1 cor_m_3_2_reg_3_ ( .D(cor_maj_118_port_o), .CK(clk), .Q(
        cor_port_v_3_2[3]), .QN() );
  DFF_X1 cor_m_3_2_reg_4_ ( .D(cor_maj_119_port_o), .CK(clk), .Q(
        cor_port_v_3_2[4]), .QN() );
  DFF_X1 cor_m_3_1_reg_0_ ( .D(cor_maj_110_port_o), .CK(clk), .Q(
        cor_port_v_3_1[0]), .QN() );
  DFF_X1 cor_m_3_1_reg_1_ ( .D(cor_maj_111_port_o), .CK(clk), .Q(
        cor_port_v_3_1[1]), .QN() );
  DFF_X1 cor_m_3_1_reg_2_ ( .D(cor_maj_112_port_o), .CK(clk), .Q(
        cor_port_v_3_1[2]), .QN() );
  DFF_X1 cor_m_3_1_reg_3_ ( .D(cor_maj_113_port_o), .CK(clk), .Q(
        cor_port_v_3_1[3]), .QN() );
  DFF_X1 cor_m_3_1_reg_4_ ( .D(cor_maj_114_port_o), .CK(clk), .Q(
        cor_port_v_3_1[4]), .QN() );
  DFF_X1 cor_m_3_0_reg_0_ ( .D(cor_maj_105_port_o), .CK(clk), .Q(
        cor_port_v_3_0[0]), .QN() );
  DFF_X1 cor_m_3_0_reg_1_ ( .D(cor_maj_106_port_o), .CK(clk), .Q(
        cor_port_v_3_0[1]), .QN() );
  DFF_X1 cor_m_3_0_reg_2_ ( .D(cor_maj_107_port_o), .CK(clk), .Q(
        cor_port_v_3_0[2]), .QN() );
  DFF_X1 cor_m_3_0_reg_3_ ( .D(cor_maj_108_port_o), .CK(clk), .Q(
        cor_port_v_3_0[3]), .QN() );
  DFF_X1 cor_m_3_0_reg_4_ ( .D(cor_maj_109_port_o), .CK(clk), .Q(
        cor_port_v_3_0[4]), .QN() );
  DFF_X1 cor_m_2_3_reg_0_ ( .D(cor_maj_100_port_o), .CK(clk), .Q(
        cor_port_v_2_3[0]), .QN() );
  DFF_X1 cor_m_2_3_reg_1_ ( .D(cor_maj_101_port_o), .CK(clk), .Q(
        cor_port_v_2_3[1]), .QN() );
  DFF_X1 cor_m_2_3_reg_2_ ( .D(cor_maj_102_port_o), .CK(clk), .Q(
        cor_port_v_2_3[2]), .QN() );
  DFF_X1 cor_m_2_3_reg_3_ ( .D(cor_maj_103_port_o), .CK(clk), .Q(
        cor_port_v_2_3[3]), .QN() );
  DFF_X1 cor_m_2_3_reg_4_ ( .D(cor_maj_104_port_o), .CK(clk), .Q(
        cor_port_v_2_3[4]), .QN() );
  DFF_X1 cor_m_2_1_reg_0_ ( .D(cor_maj_95_port_o), .CK(clk), .Q(
        cor_port_v_2_1[0]), .QN() );
  DFF_X1 cor_m_2_1_reg_1_ ( .D(cor_maj_96_port_o), .CK(clk), .Q(
        cor_port_v_2_1[1]), .QN() );
  DFF_X1 cor_m_2_1_reg_2_ ( .D(cor_maj_97_port_o), .CK(clk), .Q(
        cor_port_v_2_1[2]), .QN() );
  DFF_X1 cor_m_2_1_reg_3_ ( .D(cor_maj_98_port_o), .CK(clk), .Q(
        cor_port_v_2_1[3]), .QN() );
  DFF_X1 cor_m_2_1_reg_4_ ( .D(cor_maj_99_port_o), .CK(clk), .Q(
        cor_port_v_2_1[4]), .QN() );
  DFF_X1 cor_m_2_0_reg_0_ ( .D(cor_maj_90_port_o), .CK(clk), .Q(
        cor_port_v_2_0[0]), .QN() );
  DFF_X1 cor_m_2_0_reg_1_ ( .D(cor_maj_91_port_o), .CK(clk), .Q(
        cor_port_v_2_0[1]), .QN() );
  DFF_X1 cor_m_2_0_reg_2_ ( .D(cor_maj_92_port_o), .CK(clk), .Q(
        cor_port_v_2_0[2]), .QN() );
  DFF_X1 cor_m_2_0_reg_3_ ( .D(cor_maj_93_port_o), .CK(clk), .Q(
        cor_port_v_2_0[3]), .QN() );
  DFF_X1 cor_m_2_0_reg_4_ ( .D(cor_maj_94_port_o), .CK(clk), .Q(
        cor_port_v_2_0[4]), .QN() );
  DFF_X1 cor_m_1_3_reg_0_ ( .D(cor_maj_85_port_o), .CK(clk), .Q(
        cor_port_v_1_3[0]), .QN() );
  DFF_X1 cor_m_1_3_reg_1_ ( .D(cor_maj_86_port_o), .CK(clk), .Q(
        cor_port_v_1_3[1]), .QN() );
  DFF_X1 cor_m_1_3_reg_2_ ( .D(cor_maj_87_port_o), .CK(clk), .Q(
        cor_port_v_1_3[2]), .QN() );
  DFF_X1 cor_m_1_3_reg_3_ ( .D(cor_maj_88_port_o), .CK(clk), .Q(
        cor_port_v_1_3[3]), .QN() );
  DFF_X1 cor_m_1_3_reg_4_ ( .D(cor_maj_89_port_o), .CK(clk), .Q(
        cor_port_v_1_3[4]), .QN() );
  DFF_X1 cor_m_1_2_reg_0_ ( .D(cor_maj_80_port_o), .CK(clk), .Q(
        cor_port_v_1_2[0]), .QN() );
  DFF_X1 cor_m_1_2_reg_1_ ( .D(cor_maj_81_port_o), .CK(clk), .Q(
        cor_port_v_1_2[1]), .QN() );
  DFF_X1 cor_m_1_2_reg_2_ ( .D(cor_maj_82_port_o), .CK(clk), .Q(
        cor_port_v_1_2[2]), .QN() );
  DFF_X1 cor_m_1_2_reg_3_ ( .D(cor_maj_83_port_o), .CK(clk), .Q(
        cor_port_v_1_2[3]), .QN() );
  DFF_X1 cor_m_1_2_reg_4_ ( .D(cor_maj_84_port_o), .CK(clk), .Q(
        cor_port_v_1_2[4]), .QN() );
  DFF_X1 cor_m_1_0_reg_0_ ( .D(cor_maj_75_port_o), .CK(clk), .Q(
        cor_port_v_1_0[0]), .QN() );
  DFF_X1 cor_m_1_0_reg_1_ ( .D(cor_maj_76_port_o), .CK(clk), .Q(
        cor_port_v_1_0[1]), .QN() );
  DFF_X1 cor_m_1_0_reg_2_ ( .D(cor_maj_77_port_o), .CK(clk), .Q(
        cor_port_v_1_0[2]), .QN() );
  DFF_X1 cor_m_1_0_reg_3_ ( .D(cor_maj_78_port_o), .CK(clk), .Q(
        cor_port_v_1_0[3]), .QN() );
  DFF_X1 cor_m_1_0_reg_4_ ( .D(cor_maj_79_port_o), .CK(clk), .Q(
        cor_port_v_1_0[4]), .QN() );
  DFF_X1 cor_m_0_3_reg_0_ ( .D(cor_maj_70_port_o), .CK(clk), .Q(
        cor_port_v_0_3[0]), .QN() );
  DFF_X1 cor_m_0_3_reg_1_ ( .D(cor_maj_71_port_o), .CK(clk), .Q(
        cor_port_v_0_3[1]), .QN() );
  DFF_X1 cor_m_0_3_reg_2_ ( .D(cor_maj_72_port_o), .CK(clk), .Q(
        cor_port_v_0_3[2]), .QN() );
  DFF_X1 cor_m_0_3_reg_3_ ( .D(cor_maj_73_port_o), .CK(clk), .Q(
        cor_port_v_0_3[3]), .QN() );
  DFF_X1 cor_m_0_3_reg_4_ ( .D(cor_maj_74_port_o), .CK(clk), .Q(
        cor_port_v_0_3[4]), .QN() );
  DFF_X1 cor_m_0_2_reg_0_ ( .D(cor_maj_65_port_o), .CK(clk), .Q(
        cor_port_v_0_2[0]), .QN() );
  DFF_X1 cor_m_0_2_reg_1_ ( .D(cor_maj_66_port_o), .CK(clk), .Q(
        cor_port_v_0_2[1]), .QN() );
  DFF_X1 cor_m_0_2_reg_2_ ( .D(cor_maj_67_port_o), .CK(clk), .Q(
        cor_port_v_0_2[2]), .QN() );
  DFF_X1 cor_m_0_2_reg_3_ ( .D(cor_maj_68_port_o), .CK(clk), .Q(
        cor_port_v_0_2[3]), .QN() );
  DFF_X1 cor_m_0_2_reg_4_ ( .D(cor_maj_69_port_o), .CK(clk), .Q(
        cor_port_v_0_2[4]), .QN() );
  DFF_X1 cor_m_0_1_reg_0_ ( .D(cor_maj_60_port_o), .CK(clk), .Q(
        cor_port_v_0_1[0]), .QN() );
  DFF_X1 cor_m_0_1_reg_1_ ( .D(cor_maj_61_port_o), .CK(clk), .Q(
        cor_port_v_0_1[1]), .QN() );
  DFF_X1 cor_m_0_1_reg_2_ ( .D(cor_maj_62_port_o), .CK(clk), .Q(
        cor_port_v_0_1[2]), .QN() );
  DFF_X1 cor_m_0_1_reg_3_ ( .D(cor_maj_63_port_o), .CK(clk), .Q(
        cor_port_v_0_1[3]), .QN() );
  DFF_X1 cor_m_0_1_reg_4_ ( .D(cor_maj_64_port_o), .CK(clk), .Q(
        cor_port_v_0_1[4]), .QN() );
  NAND2_X1 cor_maj_60_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_60_n9) );
  NAND2_X1 cor_maj_60_U14 ( .A1(cor_maj_60_n6), .A2(cor_maj_60_n5), .ZN(
        cor_maj_60_n10) );
  NAND2_X1 cor_maj_60_U13 ( .A1(cor_maj_60_n9), .A2(cor_maj_60_n10), .ZN(
        cor_maj_60_n8) );
  NAND2_X1 cor_maj_60_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_60_n11), .ZN(
        cor_maj_60_n13) );
  NAND2_X1 cor_maj_60_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_60_n12) );
  NAND2_X1 cor_maj_60_U10 ( .A1(cor_maj_60_n12), .A2(cor_maj_60_n13), .ZN(
        cor_maj_60_n7) );
  XOR2_X1 cor_maj_60_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_60_n5) );
  XOR2_X1 cor_maj_60_U8 ( .A(v_1_0_1[2]), .B(cor_maj_60_n11), .Z(cor_maj_60_n6) );
  XOR2_X1 cor_maj_60_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_60_n11)
         );
  OR2_X1 cor_maj_60_U6 ( .A1(cor_maj_60_n7), .A2(cor_maj_60_n8), .ZN(
        cor_maj_60_n3) );
  NAND2_X1 cor_maj_60_U5 ( .A1(cor_maj_60_n3), .A2(cor_maj_60_n4), .ZN(
        cor_maj_60_n2) );
  NAND2_X1 cor_maj_60_U4 ( .A1(cor_maj_60_n7), .A2(cor_maj_60_n8), .ZN(
        cor_maj_60_n1) );
  NAND2_X1 cor_maj_60_U3 ( .A1(cor_maj_60_n1), .A2(cor_maj_60_n2), .ZN(
        cor_maj_60_port_o) );
  XOR2_X1 cor_maj_60_U2 ( .A(cor_maj_60_n5), .B(cor_maj_60_n6), .Z(
        cor_maj_60_n4) );
  NAND2_X1 cor_maj_61_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_61_n18) );
  NAND2_X1 cor_maj_61_U14 ( .A1(cor_maj_61_n21), .A2(cor_maj_61_n22), .ZN(
        cor_maj_61_n17) );
  NAND2_X1 cor_maj_61_U13 ( .A1(cor_maj_61_n18), .A2(cor_maj_61_n17), .ZN(
        cor_maj_61_n19) );
  NAND2_X1 cor_maj_61_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_61_n16), .ZN(
        cor_maj_61_n14) );
  NAND2_X1 cor_maj_61_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_61_n15) );
  NAND2_X1 cor_maj_61_U10 ( .A1(cor_maj_61_n15), .A2(cor_maj_61_n14), .ZN(
        cor_maj_61_n20) );
  XOR2_X1 cor_maj_61_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_61_n22)
         );
  XOR2_X1 cor_maj_61_U8 ( .A(v_1_0_1[2]), .B(cor_maj_61_n16), .Z(
        cor_maj_61_n21) );
  XOR2_X1 cor_maj_61_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_61_n16)
         );
  OR2_X1 cor_maj_61_U6 ( .A1(cor_maj_61_n20), .A2(cor_maj_61_n19), .ZN(
        cor_maj_61_n24) );
  NAND2_X1 cor_maj_61_U5 ( .A1(cor_maj_61_n24), .A2(cor_maj_61_n23), .ZN(
        cor_maj_61_n25) );
  NAND2_X1 cor_maj_61_U4 ( .A1(cor_maj_61_n20), .A2(cor_maj_61_n19), .ZN(
        cor_maj_61_n26) );
  NAND2_X1 cor_maj_61_U3 ( .A1(cor_maj_61_n26), .A2(cor_maj_61_n25), .ZN(
        cor_maj_61_port_o) );
  XOR2_X1 cor_maj_61_U2 ( .A(cor_maj_61_n22), .B(cor_maj_61_n21), .Z(
        cor_maj_61_n23) );
  NAND2_X1 cor_maj_62_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_62_n18) );
  NAND2_X1 cor_maj_62_U14 ( .A1(cor_maj_62_n21), .A2(cor_maj_62_n22), .ZN(
        cor_maj_62_n17) );
  NAND2_X1 cor_maj_62_U13 ( .A1(cor_maj_62_n18), .A2(cor_maj_62_n17), .ZN(
        cor_maj_62_n19) );
  NAND2_X1 cor_maj_62_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_62_n16), .ZN(
        cor_maj_62_n14) );
  NAND2_X1 cor_maj_62_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_62_n15) );
  NAND2_X1 cor_maj_62_U10 ( .A1(cor_maj_62_n15), .A2(cor_maj_62_n14), .ZN(
        cor_maj_62_n20) );
  XOR2_X1 cor_maj_62_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_62_n22)
         );
  XOR2_X1 cor_maj_62_U8 ( .A(v_1_0_1[2]), .B(cor_maj_62_n16), .Z(
        cor_maj_62_n21) );
  XOR2_X1 cor_maj_62_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_62_n16)
         );
  OR2_X1 cor_maj_62_U6 ( .A1(cor_maj_62_n20), .A2(cor_maj_62_n19), .ZN(
        cor_maj_62_n24) );
  NAND2_X1 cor_maj_62_U5 ( .A1(cor_maj_62_n24), .A2(cor_maj_62_n23), .ZN(
        cor_maj_62_n25) );
  NAND2_X1 cor_maj_62_U4 ( .A1(cor_maj_62_n20), .A2(cor_maj_62_n19), .ZN(
        cor_maj_62_n26) );
  NAND2_X1 cor_maj_62_U3 ( .A1(cor_maj_62_n26), .A2(cor_maj_62_n25), .ZN(
        cor_maj_62_port_o) );
  XOR2_X1 cor_maj_62_U2 ( .A(cor_maj_62_n22), .B(cor_maj_62_n21), .Z(
        cor_maj_62_n23) );
  NAND2_X1 cor_maj_63_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_63_n18) );
  NAND2_X1 cor_maj_63_U14 ( .A1(cor_maj_63_n21), .A2(cor_maj_63_n22), .ZN(
        cor_maj_63_n17) );
  NAND2_X1 cor_maj_63_U13 ( .A1(cor_maj_63_n18), .A2(cor_maj_63_n17), .ZN(
        cor_maj_63_n19) );
  NAND2_X1 cor_maj_63_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_63_n16), .ZN(
        cor_maj_63_n14) );
  NAND2_X1 cor_maj_63_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_63_n15) );
  NAND2_X1 cor_maj_63_U10 ( .A1(cor_maj_63_n15), .A2(cor_maj_63_n14), .ZN(
        cor_maj_63_n20) );
  XOR2_X1 cor_maj_63_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_63_n22)
         );
  XOR2_X1 cor_maj_63_U8 ( .A(v_1_0_1[2]), .B(cor_maj_63_n16), .Z(
        cor_maj_63_n21) );
  XOR2_X1 cor_maj_63_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_63_n16)
         );
  OR2_X1 cor_maj_63_U6 ( .A1(cor_maj_63_n20), .A2(cor_maj_63_n19), .ZN(
        cor_maj_63_n24) );
  NAND2_X1 cor_maj_63_U5 ( .A1(cor_maj_63_n24), .A2(cor_maj_63_n23), .ZN(
        cor_maj_63_n25) );
  NAND2_X1 cor_maj_63_U4 ( .A1(cor_maj_63_n20), .A2(cor_maj_63_n19), .ZN(
        cor_maj_63_n26) );
  NAND2_X1 cor_maj_63_U3 ( .A1(cor_maj_63_n26), .A2(cor_maj_63_n25), .ZN(
        cor_maj_63_port_o) );
  XOR2_X1 cor_maj_63_U2 ( .A(cor_maj_63_n22), .B(cor_maj_63_n21), .Z(
        cor_maj_63_n23) );
  NAND2_X1 cor_maj_64_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_64_n18) );
  NAND2_X1 cor_maj_64_U14 ( .A1(cor_maj_64_n21), .A2(cor_maj_64_n22), .ZN(
        cor_maj_64_n17) );
  NAND2_X1 cor_maj_64_U13 ( .A1(cor_maj_64_n18), .A2(cor_maj_64_n17), .ZN(
        cor_maj_64_n19) );
  NAND2_X1 cor_maj_64_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_64_n16), .ZN(
        cor_maj_64_n14) );
  NAND2_X1 cor_maj_64_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_64_n15) );
  NAND2_X1 cor_maj_64_U10 ( .A1(cor_maj_64_n15), .A2(cor_maj_64_n14), .ZN(
        cor_maj_64_n20) );
  XOR2_X1 cor_maj_64_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_64_n22)
         );
  XOR2_X1 cor_maj_64_U8 ( .A(v_1_0_1[2]), .B(cor_maj_64_n16), .Z(
        cor_maj_64_n21) );
  XOR2_X1 cor_maj_64_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_64_n16)
         );
  OR2_X1 cor_maj_64_U6 ( .A1(cor_maj_64_n20), .A2(cor_maj_64_n19), .ZN(
        cor_maj_64_n24) );
  NAND2_X1 cor_maj_64_U5 ( .A1(cor_maj_64_n24), .A2(cor_maj_64_n23), .ZN(
        cor_maj_64_n25) );
  NAND2_X1 cor_maj_64_U4 ( .A1(cor_maj_64_n20), .A2(cor_maj_64_n19), .ZN(
        cor_maj_64_n26) );
  NAND2_X1 cor_maj_64_U3 ( .A1(cor_maj_64_n26), .A2(cor_maj_64_n25), .ZN(
        cor_maj_64_port_o) );
  XOR2_X1 cor_maj_64_U2 ( .A(cor_maj_64_n22), .B(cor_maj_64_n21), .Z(
        cor_maj_64_n23) );
  NAND2_X1 cor_maj_65_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_65_n18) );
  NAND2_X1 cor_maj_65_U14 ( .A1(cor_maj_65_n21), .A2(cor_maj_65_n22), .ZN(
        cor_maj_65_n17) );
  NAND2_X1 cor_maj_65_U13 ( .A1(cor_maj_65_n18), .A2(cor_maj_65_n17), .ZN(
        cor_maj_65_n19) );
  NAND2_X1 cor_maj_65_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_65_n16), .ZN(
        cor_maj_65_n14) );
  NAND2_X1 cor_maj_65_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_65_n15) );
  NAND2_X1 cor_maj_65_U10 ( .A1(cor_maj_65_n15), .A2(cor_maj_65_n14), .ZN(
        cor_maj_65_n20) );
  XOR2_X1 cor_maj_65_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_65_n22)
         );
  XOR2_X1 cor_maj_65_U8 ( .A(v_1_0_2[2]), .B(cor_maj_65_n16), .Z(
        cor_maj_65_n21) );
  XOR2_X1 cor_maj_65_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_65_n16)
         );
  OR2_X1 cor_maj_65_U6 ( .A1(cor_maj_65_n20), .A2(cor_maj_65_n19), .ZN(
        cor_maj_65_n24) );
  NAND2_X1 cor_maj_65_U5 ( .A1(cor_maj_65_n24), .A2(cor_maj_65_n23), .ZN(
        cor_maj_65_n25) );
  NAND2_X1 cor_maj_65_U4 ( .A1(cor_maj_65_n20), .A2(cor_maj_65_n19), .ZN(
        cor_maj_65_n26) );
  NAND2_X1 cor_maj_65_U3 ( .A1(cor_maj_65_n26), .A2(cor_maj_65_n25), .ZN(
        cor_maj_65_port_o) );
  XOR2_X1 cor_maj_65_U2 ( .A(cor_maj_65_n22), .B(cor_maj_65_n21), .Z(
        cor_maj_65_n23) );
  NAND2_X1 cor_maj_66_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_66_n18) );
  NAND2_X1 cor_maj_66_U14 ( .A1(cor_maj_66_n21), .A2(cor_maj_66_n22), .ZN(
        cor_maj_66_n17) );
  NAND2_X1 cor_maj_66_U13 ( .A1(cor_maj_66_n18), .A2(cor_maj_66_n17), .ZN(
        cor_maj_66_n19) );
  NAND2_X1 cor_maj_66_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_66_n16), .ZN(
        cor_maj_66_n14) );
  NAND2_X1 cor_maj_66_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_66_n15) );
  NAND2_X1 cor_maj_66_U10 ( .A1(cor_maj_66_n15), .A2(cor_maj_66_n14), .ZN(
        cor_maj_66_n20) );
  XOR2_X1 cor_maj_66_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_66_n22)
         );
  XOR2_X1 cor_maj_66_U8 ( .A(v_1_0_2[2]), .B(cor_maj_66_n16), .Z(
        cor_maj_66_n21) );
  XOR2_X1 cor_maj_66_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_66_n16)
         );
  OR2_X1 cor_maj_66_U6 ( .A1(cor_maj_66_n20), .A2(cor_maj_66_n19), .ZN(
        cor_maj_66_n24) );
  NAND2_X1 cor_maj_66_U5 ( .A1(cor_maj_66_n24), .A2(cor_maj_66_n23), .ZN(
        cor_maj_66_n25) );
  NAND2_X1 cor_maj_66_U4 ( .A1(cor_maj_66_n20), .A2(cor_maj_66_n19), .ZN(
        cor_maj_66_n26) );
  NAND2_X1 cor_maj_66_U3 ( .A1(cor_maj_66_n26), .A2(cor_maj_66_n25), .ZN(
        cor_maj_66_port_o) );
  XOR2_X1 cor_maj_66_U2 ( .A(cor_maj_66_n22), .B(cor_maj_66_n21), .Z(
        cor_maj_66_n23) );
  NAND2_X1 cor_maj_67_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_67_n18) );
  NAND2_X1 cor_maj_67_U14 ( .A1(cor_maj_67_n21), .A2(cor_maj_67_n22), .ZN(
        cor_maj_67_n17) );
  NAND2_X1 cor_maj_67_U13 ( .A1(cor_maj_67_n18), .A2(cor_maj_67_n17), .ZN(
        cor_maj_67_n19) );
  NAND2_X1 cor_maj_67_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_67_n16), .ZN(
        cor_maj_67_n14) );
  NAND2_X1 cor_maj_67_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_67_n15) );
  NAND2_X1 cor_maj_67_U10 ( .A1(cor_maj_67_n15), .A2(cor_maj_67_n14), .ZN(
        cor_maj_67_n20) );
  XOR2_X1 cor_maj_67_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_67_n22)
         );
  XOR2_X1 cor_maj_67_U8 ( .A(v_1_0_2[2]), .B(cor_maj_67_n16), .Z(
        cor_maj_67_n21) );
  XOR2_X1 cor_maj_67_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_67_n16)
         );
  OR2_X1 cor_maj_67_U6 ( .A1(cor_maj_67_n20), .A2(cor_maj_67_n19), .ZN(
        cor_maj_67_n24) );
  NAND2_X1 cor_maj_67_U5 ( .A1(cor_maj_67_n24), .A2(cor_maj_67_n23), .ZN(
        cor_maj_67_n25) );
  NAND2_X1 cor_maj_67_U4 ( .A1(cor_maj_67_n20), .A2(cor_maj_67_n19), .ZN(
        cor_maj_67_n26) );
  NAND2_X1 cor_maj_67_U3 ( .A1(cor_maj_67_n26), .A2(cor_maj_67_n25), .ZN(
        cor_maj_67_port_o) );
  XOR2_X1 cor_maj_67_U2 ( .A(cor_maj_67_n22), .B(cor_maj_67_n21), .Z(
        cor_maj_67_n23) );
  NAND2_X1 cor_maj_68_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_68_n18) );
  NAND2_X1 cor_maj_68_U14 ( .A1(cor_maj_68_n21), .A2(cor_maj_68_n22), .ZN(
        cor_maj_68_n17) );
  NAND2_X1 cor_maj_68_U13 ( .A1(cor_maj_68_n18), .A2(cor_maj_68_n17), .ZN(
        cor_maj_68_n19) );
  NAND2_X1 cor_maj_68_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_68_n16), .ZN(
        cor_maj_68_n14) );
  NAND2_X1 cor_maj_68_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_68_n15) );
  NAND2_X1 cor_maj_68_U10 ( .A1(cor_maj_68_n15), .A2(cor_maj_68_n14), .ZN(
        cor_maj_68_n20) );
  XOR2_X1 cor_maj_68_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_68_n22)
         );
  XOR2_X1 cor_maj_68_U8 ( .A(v_1_0_2[2]), .B(cor_maj_68_n16), .Z(
        cor_maj_68_n21) );
  XOR2_X1 cor_maj_68_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_68_n16)
         );
  OR2_X1 cor_maj_68_U6 ( .A1(cor_maj_68_n20), .A2(cor_maj_68_n19), .ZN(
        cor_maj_68_n24) );
  NAND2_X1 cor_maj_68_U5 ( .A1(cor_maj_68_n24), .A2(cor_maj_68_n23), .ZN(
        cor_maj_68_n25) );
  NAND2_X1 cor_maj_68_U4 ( .A1(cor_maj_68_n20), .A2(cor_maj_68_n19), .ZN(
        cor_maj_68_n26) );
  NAND2_X1 cor_maj_68_U3 ( .A1(cor_maj_68_n26), .A2(cor_maj_68_n25), .ZN(
        cor_maj_68_port_o) );
  XOR2_X1 cor_maj_68_U2 ( .A(cor_maj_68_n22), .B(cor_maj_68_n21), .Z(
        cor_maj_68_n23) );
  NAND2_X1 cor_maj_69_U15 ( .A1(v_1_0_2[3]), .A2(v_1_0_2[4]), .ZN(
        cor_maj_69_n18) );
  NAND2_X1 cor_maj_69_U14 ( .A1(cor_maj_69_n21), .A2(cor_maj_69_n22), .ZN(
        cor_maj_69_n17) );
  NAND2_X1 cor_maj_69_U13 ( .A1(cor_maj_69_n18), .A2(cor_maj_69_n17), .ZN(
        cor_maj_69_n19) );
  NAND2_X1 cor_maj_69_U12 ( .A1(v_1_0_2[2]), .A2(cor_maj_69_n16), .ZN(
        cor_maj_69_n14) );
  NAND2_X1 cor_maj_69_U11 ( .A1(v_1_0_2[0]), .A2(v_1_0_2[1]), .ZN(
        cor_maj_69_n15) );
  NAND2_X1 cor_maj_69_U10 ( .A1(cor_maj_69_n15), .A2(cor_maj_69_n14), .ZN(
        cor_maj_69_n20) );
  XOR2_X1 cor_maj_69_U9 ( .A(v_1_0_2[3]), .B(v_1_0_2[4]), .Z(cor_maj_69_n22)
         );
  XOR2_X1 cor_maj_69_U8 ( .A(v_1_0_2[2]), .B(cor_maj_69_n16), .Z(
        cor_maj_69_n21) );
  XOR2_X1 cor_maj_69_U7 ( .A(v_1_0_2[0]), .B(v_1_0_2[1]), .Z(cor_maj_69_n16)
         );
  OR2_X1 cor_maj_69_U6 ( .A1(cor_maj_69_n20), .A2(cor_maj_69_n19), .ZN(
        cor_maj_69_n24) );
  NAND2_X1 cor_maj_69_U5 ( .A1(cor_maj_69_n24), .A2(cor_maj_69_n23), .ZN(
        cor_maj_69_n25) );
  NAND2_X1 cor_maj_69_U4 ( .A1(cor_maj_69_n20), .A2(cor_maj_69_n19), .ZN(
        cor_maj_69_n26) );
  NAND2_X1 cor_maj_69_U3 ( .A1(cor_maj_69_n26), .A2(cor_maj_69_n25), .ZN(
        cor_maj_69_port_o) );
  XOR2_X1 cor_maj_69_U2 ( .A(cor_maj_69_n22), .B(cor_maj_69_n21), .Z(
        cor_maj_69_n23) );
  NAND2_X1 cor_maj_70_U15 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_70_n18) );
  NAND2_X1 cor_maj_70_U14 ( .A1(cor_maj_70_n21), .A2(cor_maj_70_n22), .ZN(
        cor_maj_70_n17) );
  NAND2_X1 cor_maj_70_U13 ( .A1(cor_maj_70_n18), .A2(cor_maj_70_n17), .ZN(
        cor_maj_70_n19) );
  NAND2_X1 cor_maj_70_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_70_n16), .ZN(
        cor_maj_70_n14) );
  NAND2_X1 cor_maj_70_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_70_n15) );
  NAND2_X1 cor_maj_70_U10 ( .A1(cor_maj_70_n15), .A2(cor_maj_70_n14), .ZN(
        cor_maj_70_n20) );
  XOR2_X1 cor_maj_70_U9 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_70_n22)
         );
  XOR2_X1 cor_maj_70_U8 ( .A(v_1_0_3[2]), .B(cor_maj_70_n16), .Z(
        cor_maj_70_n21) );
  XOR2_X1 cor_maj_70_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_70_n16)
         );
  OR2_X1 cor_maj_70_U6 ( .A1(cor_maj_70_n20), .A2(cor_maj_70_n19), .ZN(
        cor_maj_70_n24) );
  NAND2_X1 cor_maj_70_U5 ( .A1(cor_maj_70_n24), .A2(cor_maj_70_n23), .ZN(
        cor_maj_70_n25) );
  NAND2_X1 cor_maj_70_U4 ( .A1(cor_maj_70_n20), .A2(cor_maj_70_n19), .ZN(
        cor_maj_70_n26) );
  NAND2_X1 cor_maj_70_U3 ( .A1(cor_maj_70_n26), .A2(cor_maj_70_n25), .ZN(
        cor_maj_70_port_o) );
  XOR2_X1 cor_maj_70_U2 ( .A(cor_maj_70_n22), .B(cor_maj_70_n21), .Z(
        cor_maj_70_n23) );
  NAND2_X1 cor_maj_71_U15 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_71_n18) );
  NAND2_X1 cor_maj_71_U14 ( .A1(cor_maj_71_n21), .A2(cor_maj_71_n22), .ZN(
        cor_maj_71_n17) );
  NAND2_X1 cor_maj_71_U13 ( .A1(cor_maj_71_n18), .A2(cor_maj_71_n17), .ZN(
        cor_maj_71_n19) );
  NAND2_X1 cor_maj_71_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_71_n16), .ZN(
        cor_maj_71_n14) );
  NAND2_X1 cor_maj_71_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_71_n15) );
  NAND2_X1 cor_maj_71_U10 ( .A1(cor_maj_71_n15), .A2(cor_maj_71_n14), .ZN(
        cor_maj_71_n20) );
  XOR2_X1 cor_maj_71_U9 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_71_n22)
         );
  XOR2_X1 cor_maj_71_U8 ( .A(v_1_0_3[2]), .B(cor_maj_71_n16), .Z(
        cor_maj_71_n21) );
  XOR2_X1 cor_maj_71_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_71_n16)
         );
  OR2_X1 cor_maj_71_U6 ( .A1(cor_maj_71_n20), .A2(cor_maj_71_n19), .ZN(
        cor_maj_71_n24) );
  NAND2_X1 cor_maj_71_U5 ( .A1(cor_maj_71_n24), .A2(cor_maj_71_n23), .ZN(
        cor_maj_71_n25) );
  NAND2_X1 cor_maj_71_U4 ( .A1(cor_maj_71_n20), .A2(cor_maj_71_n19), .ZN(
        cor_maj_71_n26) );
  NAND2_X1 cor_maj_71_U3 ( .A1(cor_maj_71_n26), .A2(cor_maj_71_n25), .ZN(
        cor_maj_71_port_o) );
  XOR2_X1 cor_maj_71_U2 ( .A(cor_maj_71_n22), .B(cor_maj_71_n21), .Z(
        cor_maj_71_n23) );
  NAND2_X1 cor_maj_72_U15 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_72_n18) );
  NAND2_X1 cor_maj_72_U14 ( .A1(cor_maj_72_n21), .A2(cor_maj_72_n22), .ZN(
        cor_maj_72_n17) );
  NAND2_X1 cor_maj_72_U13 ( .A1(cor_maj_72_n18), .A2(cor_maj_72_n17), .ZN(
        cor_maj_72_n19) );
  NAND2_X1 cor_maj_72_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_72_n16), .ZN(
        cor_maj_72_n14) );
  NAND2_X1 cor_maj_72_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_72_n15) );
  NAND2_X1 cor_maj_72_U10 ( .A1(cor_maj_72_n15), .A2(cor_maj_72_n14), .ZN(
        cor_maj_72_n20) );
  XOR2_X1 cor_maj_72_U9 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_72_n22)
         );
  XOR2_X1 cor_maj_72_U8 ( .A(v_1_0_3[2]), .B(cor_maj_72_n16), .Z(
        cor_maj_72_n21) );
  XOR2_X1 cor_maj_72_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_72_n16)
         );
  OR2_X1 cor_maj_72_U6 ( .A1(cor_maj_72_n20), .A2(cor_maj_72_n19), .ZN(
        cor_maj_72_n24) );
  NAND2_X1 cor_maj_72_U5 ( .A1(cor_maj_72_n24), .A2(cor_maj_72_n23), .ZN(
        cor_maj_72_n25) );
  NAND2_X1 cor_maj_72_U4 ( .A1(cor_maj_72_n20), .A2(cor_maj_72_n19), .ZN(
        cor_maj_72_n26) );
  NAND2_X1 cor_maj_72_U3 ( .A1(cor_maj_72_n26), .A2(cor_maj_72_n25), .ZN(
        cor_maj_72_port_o) );
  XOR2_X1 cor_maj_72_U2 ( .A(cor_maj_72_n22), .B(cor_maj_72_n21), .Z(
        cor_maj_72_n23) );
  NAND2_X1 cor_maj_73_U15 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_73_n18) );
  NAND2_X1 cor_maj_73_U14 ( .A1(cor_maj_73_n21), .A2(cor_maj_73_n22), .ZN(
        cor_maj_73_n17) );
  NAND2_X1 cor_maj_73_U13 ( .A1(cor_maj_73_n18), .A2(cor_maj_73_n17), .ZN(
        cor_maj_73_n19) );
  NAND2_X1 cor_maj_73_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_73_n16), .ZN(
        cor_maj_73_n14) );
  NAND2_X1 cor_maj_73_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_73_n15) );
  NAND2_X1 cor_maj_73_U10 ( .A1(cor_maj_73_n15), .A2(cor_maj_73_n14), .ZN(
        cor_maj_73_n20) );
  XOR2_X1 cor_maj_73_U9 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_73_n22)
         );
  XOR2_X1 cor_maj_73_U8 ( .A(v_1_0_3[2]), .B(cor_maj_73_n16), .Z(
        cor_maj_73_n21) );
  XOR2_X1 cor_maj_73_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_73_n16)
         );
  OR2_X1 cor_maj_73_U6 ( .A1(cor_maj_73_n20), .A2(cor_maj_73_n19), .ZN(
        cor_maj_73_n24) );
  NAND2_X1 cor_maj_73_U5 ( .A1(cor_maj_73_n24), .A2(cor_maj_73_n23), .ZN(
        cor_maj_73_n25) );
  NAND2_X1 cor_maj_73_U4 ( .A1(cor_maj_73_n20), .A2(cor_maj_73_n19), .ZN(
        cor_maj_73_n26) );
  NAND2_X1 cor_maj_73_U3 ( .A1(cor_maj_73_n26), .A2(cor_maj_73_n25), .ZN(
        cor_maj_73_port_o) );
  XOR2_X1 cor_maj_73_U2 ( .A(cor_maj_73_n22), .B(cor_maj_73_n21), .Z(
        cor_maj_73_n23) );
  NAND2_X1 cor_maj_74_U15 ( .A1(v_1_0_3[3]), .A2(v_1_0_3[4]), .ZN(
        cor_maj_74_n18) );
  NAND2_X1 cor_maj_74_U14 ( .A1(cor_maj_74_n21), .A2(cor_maj_74_n22), .ZN(
        cor_maj_74_n17) );
  NAND2_X1 cor_maj_74_U13 ( .A1(cor_maj_74_n18), .A2(cor_maj_74_n17), .ZN(
        cor_maj_74_n19) );
  NAND2_X1 cor_maj_74_U12 ( .A1(v_1_0_3[2]), .A2(cor_maj_74_n16), .ZN(
        cor_maj_74_n14) );
  NAND2_X1 cor_maj_74_U11 ( .A1(v_1_0_3[0]), .A2(v_1_0_3[1]), .ZN(
        cor_maj_74_n15) );
  NAND2_X1 cor_maj_74_U10 ( .A1(cor_maj_74_n15), .A2(cor_maj_74_n14), .ZN(
        cor_maj_74_n20) );
  XOR2_X1 cor_maj_74_U9 ( .A(v_1_0_3[3]), .B(v_1_0_3[4]), .Z(cor_maj_74_n22)
         );
  XOR2_X1 cor_maj_74_U8 ( .A(v_1_0_3[2]), .B(cor_maj_74_n16), .Z(
        cor_maj_74_n21) );
  XOR2_X1 cor_maj_74_U7 ( .A(v_1_0_3[0]), .B(v_1_0_3[1]), .Z(cor_maj_74_n16)
         );
  OR2_X1 cor_maj_74_U6 ( .A1(cor_maj_74_n20), .A2(cor_maj_74_n19), .ZN(
        cor_maj_74_n24) );
  NAND2_X1 cor_maj_74_U5 ( .A1(cor_maj_74_n24), .A2(cor_maj_74_n23), .ZN(
        cor_maj_74_n25) );
  NAND2_X1 cor_maj_74_U4 ( .A1(cor_maj_74_n20), .A2(cor_maj_74_n19), .ZN(
        cor_maj_74_n26) );
  NAND2_X1 cor_maj_74_U3 ( .A1(cor_maj_74_n26), .A2(cor_maj_74_n25), .ZN(
        cor_maj_74_port_o) );
  XOR2_X1 cor_maj_74_U2 ( .A(cor_maj_74_n22), .B(cor_maj_74_n21), .Z(
        cor_maj_74_n23) );
  NAND2_X1 cor_maj_75_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_75_n18) );
  NAND2_X1 cor_maj_75_U14 ( .A1(cor_maj_75_n21), .A2(cor_maj_75_n22), .ZN(
        cor_maj_75_n17) );
  NAND2_X1 cor_maj_75_U13 ( .A1(cor_maj_75_n18), .A2(cor_maj_75_n17), .ZN(
        cor_maj_75_n19) );
  NAND2_X1 cor_maj_75_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_75_n16), .ZN(
        cor_maj_75_n14) );
  NAND2_X1 cor_maj_75_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_75_n15) );
  NAND2_X1 cor_maj_75_U10 ( .A1(cor_maj_75_n15), .A2(cor_maj_75_n14), .ZN(
        cor_maj_75_n20) );
  XOR2_X1 cor_maj_75_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_75_n22)
         );
  XOR2_X1 cor_maj_75_U8 ( .A(v_1_1_0[2]), .B(cor_maj_75_n16), .Z(
        cor_maj_75_n21) );
  XOR2_X1 cor_maj_75_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_75_n16)
         );
  OR2_X1 cor_maj_75_U6 ( .A1(cor_maj_75_n20), .A2(cor_maj_75_n19), .ZN(
        cor_maj_75_n24) );
  NAND2_X1 cor_maj_75_U5 ( .A1(cor_maj_75_n24), .A2(cor_maj_75_n23), .ZN(
        cor_maj_75_n25) );
  NAND2_X1 cor_maj_75_U4 ( .A1(cor_maj_75_n20), .A2(cor_maj_75_n19), .ZN(
        cor_maj_75_n26) );
  NAND2_X1 cor_maj_75_U3 ( .A1(cor_maj_75_n26), .A2(cor_maj_75_n25), .ZN(
        cor_maj_75_port_o) );
  XOR2_X1 cor_maj_75_U2 ( .A(cor_maj_75_n22), .B(cor_maj_75_n21), .Z(
        cor_maj_75_n23) );
  NAND2_X1 cor_maj_76_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_76_n18) );
  NAND2_X1 cor_maj_76_U14 ( .A1(cor_maj_76_n21), .A2(cor_maj_76_n22), .ZN(
        cor_maj_76_n17) );
  NAND2_X1 cor_maj_76_U13 ( .A1(cor_maj_76_n18), .A2(cor_maj_76_n17), .ZN(
        cor_maj_76_n19) );
  NAND2_X1 cor_maj_76_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_76_n16), .ZN(
        cor_maj_76_n14) );
  NAND2_X1 cor_maj_76_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_76_n15) );
  NAND2_X1 cor_maj_76_U10 ( .A1(cor_maj_76_n15), .A2(cor_maj_76_n14), .ZN(
        cor_maj_76_n20) );
  XOR2_X1 cor_maj_76_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_76_n22)
         );
  XOR2_X1 cor_maj_76_U8 ( .A(v_1_1_0[2]), .B(cor_maj_76_n16), .Z(
        cor_maj_76_n21) );
  XOR2_X1 cor_maj_76_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_76_n16)
         );
  OR2_X1 cor_maj_76_U6 ( .A1(cor_maj_76_n20), .A2(cor_maj_76_n19), .ZN(
        cor_maj_76_n24) );
  NAND2_X1 cor_maj_76_U5 ( .A1(cor_maj_76_n24), .A2(cor_maj_76_n23), .ZN(
        cor_maj_76_n25) );
  NAND2_X1 cor_maj_76_U4 ( .A1(cor_maj_76_n20), .A2(cor_maj_76_n19), .ZN(
        cor_maj_76_n26) );
  NAND2_X1 cor_maj_76_U3 ( .A1(cor_maj_76_n26), .A2(cor_maj_76_n25), .ZN(
        cor_maj_76_port_o) );
  XOR2_X1 cor_maj_76_U2 ( .A(cor_maj_76_n22), .B(cor_maj_76_n21), .Z(
        cor_maj_76_n23) );
  NAND2_X1 cor_maj_77_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_77_n18) );
  NAND2_X1 cor_maj_77_U14 ( .A1(cor_maj_77_n21), .A2(cor_maj_77_n22), .ZN(
        cor_maj_77_n17) );
  NAND2_X1 cor_maj_77_U13 ( .A1(cor_maj_77_n18), .A2(cor_maj_77_n17), .ZN(
        cor_maj_77_n19) );
  NAND2_X1 cor_maj_77_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_77_n16), .ZN(
        cor_maj_77_n14) );
  NAND2_X1 cor_maj_77_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_77_n15) );
  NAND2_X1 cor_maj_77_U10 ( .A1(cor_maj_77_n15), .A2(cor_maj_77_n14), .ZN(
        cor_maj_77_n20) );
  XOR2_X1 cor_maj_77_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_77_n22)
         );
  XOR2_X1 cor_maj_77_U8 ( .A(v_1_1_0[2]), .B(cor_maj_77_n16), .Z(
        cor_maj_77_n21) );
  XOR2_X1 cor_maj_77_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_77_n16)
         );
  OR2_X1 cor_maj_77_U6 ( .A1(cor_maj_77_n20), .A2(cor_maj_77_n19), .ZN(
        cor_maj_77_n24) );
  NAND2_X1 cor_maj_77_U5 ( .A1(cor_maj_77_n24), .A2(cor_maj_77_n23), .ZN(
        cor_maj_77_n25) );
  NAND2_X1 cor_maj_77_U4 ( .A1(cor_maj_77_n20), .A2(cor_maj_77_n19), .ZN(
        cor_maj_77_n26) );
  NAND2_X1 cor_maj_77_U3 ( .A1(cor_maj_77_n26), .A2(cor_maj_77_n25), .ZN(
        cor_maj_77_port_o) );
  XOR2_X1 cor_maj_77_U2 ( .A(cor_maj_77_n22), .B(cor_maj_77_n21), .Z(
        cor_maj_77_n23) );
  NAND2_X1 cor_maj_78_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_78_n18) );
  NAND2_X1 cor_maj_78_U14 ( .A1(cor_maj_78_n21), .A2(cor_maj_78_n22), .ZN(
        cor_maj_78_n17) );
  NAND2_X1 cor_maj_78_U13 ( .A1(cor_maj_78_n18), .A2(cor_maj_78_n17), .ZN(
        cor_maj_78_n19) );
  NAND2_X1 cor_maj_78_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_78_n16), .ZN(
        cor_maj_78_n14) );
  NAND2_X1 cor_maj_78_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_78_n15) );
  NAND2_X1 cor_maj_78_U10 ( .A1(cor_maj_78_n15), .A2(cor_maj_78_n14), .ZN(
        cor_maj_78_n20) );
  XOR2_X1 cor_maj_78_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_78_n22)
         );
  XOR2_X1 cor_maj_78_U8 ( .A(v_1_1_0[2]), .B(cor_maj_78_n16), .Z(
        cor_maj_78_n21) );
  XOR2_X1 cor_maj_78_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_78_n16)
         );
  OR2_X1 cor_maj_78_U6 ( .A1(cor_maj_78_n20), .A2(cor_maj_78_n19), .ZN(
        cor_maj_78_n24) );
  NAND2_X1 cor_maj_78_U5 ( .A1(cor_maj_78_n24), .A2(cor_maj_78_n23), .ZN(
        cor_maj_78_n25) );
  NAND2_X1 cor_maj_78_U4 ( .A1(cor_maj_78_n20), .A2(cor_maj_78_n19), .ZN(
        cor_maj_78_n26) );
  NAND2_X1 cor_maj_78_U3 ( .A1(cor_maj_78_n26), .A2(cor_maj_78_n25), .ZN(
        cor_maj_78_port_o) );
  XOR2_X1 cor_maj_78_U2 ( .A(cor_maj_78_n22), .B(cor_maj_78_n21), .Z(
        cor_maj_78_n23) );
  NAND2_X1 cor_maj_79_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_79_n18) );
  NAND2_X1 cor_maj_79_U14 ( .A1(cor_maj_79_n21), .A2(cor_maj_79_n22), .ZN(
        cor_maj_79_n17) );
  NAND2_X1 cor_maj_79_U13 ( .A1(cor_maj_79_n18), .A2(cor_maj_79_n17), .ZN(
        cor_maj_79_n19) );
  NAND2_X1 cor_maj_79_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_79_n16), .ZN(
        cor_maj_79_n14) );
  NAND2_X1 cor_maj_79_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_79_n15) );
  NAND2_X1 cor_maj_79_U10 ( .A1(cor_maj_79_n15), .A2(cor_maj_79_n14), .ZN(
        cor_maj_79_n20) );
  XOR2_X1 cor_maj_79_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_79_n22)
         );
  XOR2_X1 cor_maj_79_U8 ( .A(v_1_1_0[2]), .B(cor_maj_79_n16), .Z(
        cor_maj_79_n21) );
  XOR2_X1 cor_maj_79_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_79_n16)
         );
  OR2_X1 cor_maj_79_U6 ( .A1(cor_maj_79_n20), .A2(cor_maj_79_n19), .ZN(
        cor_maj_79_n24) );
  NAND2_X1 cor_maj_79_U5 ( .A1(cor_maj_79_n24), .A2(cor_maj_79_n23), .ZN(
        cor_maj_79_n25) );
  NAND2_X1 cor_maj_79_U4 ( .A1(cor_maj_79_n20), .A2(cor_maj_79_n19), .ZN(
        cor_maj_79_n26) );
  NAND2_X1 cor_maj_79_U3 ( .A1(cor_maj_79_n26), .A2(cor_maj_79_n25), .ZN(
        cor_maj_79_port_o) );
  XOR2_X1 cor_maj_79_U2 ( .A(cor_maj_79_n22), .B(cor_maj_79_n21), .Z(
        cor_maj_79_n23) );
  NAND2_X1 cor_maj_80_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_80_n18) );
  NAND2_X1 cor_maj_80_U14 ( .A1(cor_maj_80_n21), .A2(cor_maj_80_n22), .ZN(
        cor_maj_80_n17) );
  NAND2_X1 cor_maj_80_U13 ( .A1(cor_maj_80_n18), .A2(cor_maj_80_n17), .ZN(
        cor_maj_80_n19) );
  NAND2_X1 cor_maj_80_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_80_n16), .ZN(
        cor_maj_80_n14) );
  NAND2_X1 cor_maj_80_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_80_n15) );
  NAND2_X1 cor_maj_80_U10 ( .A1(cor_maj_80_n15), .A2(cor_maj_80_n14), .ZN(
        cor_maj_80_n20) );
  XOR2_X1 cor_maj_80_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_80_n22)
         );
  XOR2_X1 cor_maj_80_U8 ( .A(v_1_1_2[2]), .B(cor_maj_80_n16), .Z(
        cor_maj_80_n21) );
  XOR2_X1 cor_maj_80_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_80_n16)
         );
  OR2_X1 cor_maj_80_U6 ( .A1(cor_maj_80_n20), .A2(cor_maj_80_n19), .ZN(
        cor_maj_80_n24) );
  NAND2_X1 cor_maj_80_U5 ( .A1(cor_maj_80_n24), .A2(cor_maj_80_n23), .ZN(
        cor_maj_80_n25) );
  NAND2_X1 cor_maj_80_U4 ( .A1(cor_maj_80_n20), .A2(cor_maj_80_n19), .ZN(
        cor_maj_80_n26) );
  NAND2_X1 cor_maj_80_U3 ( .A1(cor_maj_80_n26), .A2(cor_maj_80_n25), .ZN(
        cor_maj_80_port_o) );
  XOR2_X1 cor_maj_80_U2 ( .A(cor_maj_80_n22), .B(cor_maj_80_n21), .Z(
        cor_maj_80_n23) );
  NAND2_X1 cor_maj_81_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_81_n18) );
  NAND2_X1 cor_maj_81_U14 ( .A1(cor_maj_81_n21), .A2(cor_maj_81_n22), .ZN(
        cor_maj_81_n17) );
  NAND2_X1 cor_maj_81_U13 ( .A1(cor_maj_81_n18), .A2(cor_maj_81_n17), .ZN(
        cor_maj_81_n19) );
  NAND2_X1 cor_maj_81_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_81_n16), .ZN(
        cor_maj_81_n14) );
  NAND2_X1 cor_maj_81_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_81_n15) );
  NAND2_X1 cor_maj_81_U10 ( .A1(cor_maj_81_n15), .A2(cor_maj_81_n14), .ZN(
        cor_maj_81_n20) );
  XOR2_X1 cor_maj_81_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_81_n22)
         );
  XOR2_X1 cor_maj_81_U8 ( .A(v_1_1_2[2]), .B(cor_maj_81_n16), .Z(
        cor_maj_81_n21) );
  XOR2_X1 cor_maj_81_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_81_n16)
         );
  OR2_X1 cor_maj_81_U6 ( .A1(cor_maj_81_n20), .A2(cor_maj_81_n19), .ZN(
        cor_maj_81_n24) );
  NAND2_X1 cor_maj_81_U5 ( .A1(cor_maj_81_n24), .A2(cor_maj_81_n23), .ZN(
        cor_maj_81_n25) );
  NAND2_X1 cor_maj_81_U4 ( .A1(cor_maj_81_n20), .A2(cor_maj_81_n19), .ZN(
        cor_maj_81_n26) );
  NAND2_X1 cor_maj_81_U3 ( .A1(cor_maj_81_n26), .A2(cor_maj_81_n25), .ZN(
        cor_maj_81_port_o) );
  XOR2_X1 cor_maj_81_U2 ( .A(cor_maj_81_n22), .B(cor_maj_81_n21), .Z(
        cor_maj_81_n23) );
  NAND2_X1 cor_maj_82_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_82_n18) );
  NAND2_X1 cor_maj_82_U14 ( .A1(cor_maj_82_n21), .A2(cor_maj_82_n22), .ZN(
        cor_maj_82_n17) );
  NAND2_X1 cor_maj_82_U13 ( .A1(cor_maj_82_n18), .A2(cor_maj_82_n17), .ZN(
        cor_maj_82_n19) );
  NAND2_X1 cor_maj_82_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_82_n16), .ZN(
        cor_maj_82_n14) );
  NAND2_X1 cor_maj_82_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_82_n15) );
  NAND2_X1 cor_maj_82_U10 ( .A1(cor_maj_82_n15), .A2(cor_maj_82_n14), .ZN(
        cor_maj_82_n20) );
  XOR2_X1 cor_maj_82_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_82_n22)
         );
  XOR2_X1 cor_maj_82_U8 ( .A(v_1_1_2[2]), .B(cor_maj_82_n16), .Z(
        cor_maj_82_n21) );
  XOR2_X1 cor_maj_82_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_82_n16)
         );
  OR2_X1 cor_maj_82_U6 ( .A1(cor_maj_82_n20), .A2(cor_maj_82_n19), .ZN(
        cor_maj_82_n24) );
  NAND2_X1 cor_maj_82_U5 ( .A1(cor_maj_82_n24), .A2(cor_maj_82_n23), .ZN(
        cor_maj_82_n25) );
  NAND2_X1 cor_maj_82_U4 ( .A1(cor_maj_82_n20), .A2(cor_maj_82_n19), .ZN(
        cor_maj_82_n26) );
  NAND2_X1 cor_maj_82_U3 ( .A1(cor_maj_82_n26), .A2(cor_maj_82_n25), .ZN(
        cor_maj_82_port_o) );
  XOR2_X1 cor_maj_82_U2 ( .A(cor_maj_82_n22), .B(cor_maj_82_n21), .Z(
        cor_maj_82_n23) );
  NAND2_X1 cor_maj_83_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_83_n18) );
  NAND2_X1 cor_maj_83_U14 ( .A1(cor_maj_83_n21), .A2(cor_maj_83_n22), .ZN(
        cor_maj_83_n17) );
  NAND2_X1 cor_maj_83_U13 ( .A1(cor_maj_83_n18), .A2(cor_maj_83_n17), .ZN(
        cor_maj_83_n19) );
  NAND2_X1 cor_maj_83_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_83_n16), .ZN(
        cor_maj_83_n14) );
  NAND2_X1 cor_maj_83_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_83_n15) );
  NAND2_X1 cor_maj_83_U10 ( .A1(cor_maj_83_n15), .A2(cor_maj_83_n14), .ZN(
        cor_maj_83_n20) );
  XOR2_X1 cor_maj_83_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_83_n22)
         );
  XOR2_X1 cor_maj_83_U8 ( .A(v_1_1_2[2]), .B(cor_maj_83_n16), .Z(
        cor_maj_83_n21) );
  XOR2_X1 cor_maj_83_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_83_n16)
         );
  OR2_X1 cor_maj_83_U6 ( .A1(cor_maj_83_n20), .A2(cor_maj_83_n19), .ZN(
        cor_maj_83_n24) );
  NAND2_X1 cor_maj_83_U5 ( .A1(cor_maj_83_n24), .A2(cor_maj_83_n23), .ZN(
        cor_maj_83_n25) );
  NAND2_X1 cor_maj_83_U4 ( .A1(cor_maj_83_n20), .A2(cor_maj_83_n19), .ZN(
        cor_maj_83_n26) );
  NAND2_X1 cor_maj_83_U3 ( .A1(cor_maj_83_n26), .A2(cor_maj_83_n25), .ZN(
        cor_maj_83_port_o) );
  XOR2_X1 cor_maj_83_U2 ( .A(cor_maj_83_n22), .B(cor_maj_83_n21), .Z(
        cor_maj_83_n23) );
  NAND2_X1 cor_maj_84_U15 ( .A1(v_1_1_2[3]), .A2(v_1_1_2[4]), .ZN(
        cor_maj_84_n18) );
  NAND2_X1 cor_maj_84_U14 ( .A1(cor_maj_84_n21), .A2(cor_maj_84_n22), .ZN(
        cor_maj_84_n17) );
  NAND2_X1 cor_maj_84_U13 ( .A1(cor_maj_84_n18), .A2(cor_maj_84_n17), .ZN(
        cor_maj_84_n19) );
  NAND2_X1 cor_maj_84_U12 ( .A1(v_1_1_2[2]), .A2(cor_maj_84_n16), .ZN(
        cor_maj_84_n14) );
  NAND2_X1 cor_maj_84_U11 ( .A1(v_1_1_2[0]), .A2(v_1_1_2[1]), .ZN(
        cor_maj_84_n15) );
  NAND2_X1 cor_maj_84_U10 ( .A1(cor_maj_84_n15), .A2(cor_maj_84_n14), .ZN(
        cor_maj_84_n20) );
  XOR2_X1 cor_maj_84_U9 ( .A(v_1_1_2[3]), .B(v_1_1_2[4]), .Z(cor_maj_84_n22)
         );
  XOR2_X1 cor_maj_84_U8 ( .A(v_1_1_2[2]), .B(cor_maj_84_n16), .Z(
        cor_maj_84_n21) );
  XOR2_X1 cor_maj_84_U7 ( .A(v_1_1_2[0]), .B(v_1_1_2[1]), .Z(cor_maj_84_n16)
         );
  OR2_X1 cor_maj_84_U6 ( .A1(cor_maj_84_n20), .A2(cor_maj_84_n19), .ZN(
        cor_maj_84_n24) );
  NAND2_X1 cor_maj_84_U5 ( .A1(cor_maj_84_n24), .A2(cor_maj_84_n23), .ZN(
        cor_maj_84_n25) );
  NAND2_X1 cor_maj_84_U4 ( .A1(cor_maj_84_n20), .A2(cor_maj_84_n19), .ZN(
        cor_maj_84_n26) );
  NAND2_X1 cor_maj_84_U3 ( .A1(cor_maj_84_n26), .A2(cor_maj_84_n25), .ZN(
        cor_maj_84_port_o) );
  XOR2_X1 cor_maj_84_U2 ( .A(cor_maj_84_n22), .B(cor_maj_84_n21), .Z(
        cor_maj_84_n23) );
  NAND2_X1 cor_maj_85_U15 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_85_n18) );
  NAND2_X1 cor_maj_85_U14 ( .A1(cor_maj_85_n21), .A2(cor_maj_85_n22), .ZN(
        cor_maj_85_n17) );
  NAND2_X1 cor_maj_85_U13 ( .A1(cor_maj_85_n18), .A2(cor_maj_85_n17), .ZN(
        cor_maj_85_n19) );
  NAND2_X1 cor_maj_85_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_85_n16), .ZN(
        cor_maj_85_n14) );
  NAND2_X1 cor_maj_85_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_85_n15) );
  NAND2_X1 cor_maj_85_U10 ( .A1(cor_maj_85_n15), .A2(cor_maj_85_n14), .ZN(
        cor_maj_85_n20) );
  XOR2_X1 cor_maj_85_U9 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_85_n22)
         );
  XOR2_X1 cor_maj_85_U8 ( .A(v_1_1_3[2]), .B(cor_maj_85_n16), .Z(
        cor_maj_85_n21) );
  XOR2_X1 cor_maj_85_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_85_n16)
         );
  OR2_X1 cor_maj_85_U6 ( .A1(cor_maj_85_n20), .A2(cor_maj_85_n19), .ZN(
        cor_maj_85_n24) );
  NAND2_X1 cor_maj_85_U5 ( .A1(cor_maj_85_n24), .A2(cor_maj_85_n23), .ZN(
        cor_maj_85_n25) );
  NAND2_X1 cor_maj_85_U4 ( .A1(cor_maj_85_n20), .A2(cor_maj_85_n19), .ZN(
        cor_maj_85_n26) );
  NAND2_X1 cor_maj_85_U3 ( .A1(cor_maj_85_n26), .A2(cor_maj_85_n25), .ZN(
        cor_maj_85_port_o) );
  XOR2_X1 cor_maj_85_U2 ( .A(cor_maj_85_n22), .B(cor_maj_85_n21), .Z(
        cor_maj_85_n23) );
  NAND2_X1 cor_maj_86_U15 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_86_n18) );
  NAND2_X1 cor_maj_86_U14 ( .A1(cor_maj_86_n21), .A2(cor_maj_86_n22), .ZN(
        cor_maj_86_n17) );
  NAND2_X1 cor_maj_86_U13 ( .A1(cor_maj_86_n18), .A2(cor_maj_86_n17), .ZN(
        cor_maj_86_n19) );
  NAND2_X1 cor_maj_86_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_86_n16), .ZN(
        cor_maj_86_n14) );
  NAND2_X1 cor_maj_86_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_86_n15) );
  NAND2_X1 cor_maj_86_U10 ( .A1(cor_maj_86_n15), .A2(cor_maj_86_n14), .ZN(
        cor_maj_86_n20) );
  XOR2_X1 cor_maj_86_U9 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_86_n22)
         );
  XOR2_X1 cor_maj_86_U8 ( .A(v_1_1_3[2]), .B(cor_maj_86_n16), .Z(
        cor_maj_86_n21) );
  XOR2_X1 cor_maj_86_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_86_n16)
         );
  OR2_X1 cor_maj_86_U6 ( .A1(cor_maj_86_n20), .A2(cor_maj_86_n19), .ZN(
        cor_maj_86_n24) );
  NAND2_X1 cor_maj_86_U5 ( .A1(cor_maj_86_n24), .A2(cor_maj_86_n23), .ZN(
        cor_maj_86_n25) );
  NAND2_X1 cor_maj_86_U4 ( .A1(cor_maj_86_n20), .A2(cor_maj_86_n19), .ZN(
        cor_maj_86_n26) );
  NAND2_X1 cor_maj_86_U3 ( .A1(cor_maj_86_n26), .A2(cor_maj_86_n25), .ZN(
        cor_maj_86_port_o) );
  XOR2_X1 cor_maj_86_U2 ( .A(cor_maj_86_n22), .B(cor_maj_86_n21), .Z(
        cor_maj_86_n23) );
  NAND2_X1 cor_maj_87_U15 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_87_n18) );
  NAND2_X1 cor_maj_87_U14 ( .A1(cor_maj_87_n21), .A2(cor_maj_87_n22), .ZN(
        cor_maj_87_n17) );
  NAND2_X1 cor_maj_87_U13 ( .A1(cor_maj_87_n18), .A2(cor_maj_87_n17), .ZN(
        cor_maj_87_n19) );
  NAND2_X1 cor_maj_87_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_87_n16), .ZN(
        cor_maj_87_n14) );
  NAND2_X1 cor_maj_87_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_87_n15) );
  NAND2_X1 cor_maj_87_U10 ( .A1(cor_maj_87_n15), .A2(cor_maj_87_n14), .ZN(
        cor_maj_87_n20) );
  XOR2_X1 cor_maj_87_U9 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_87_n22)
         );
  XOR2_X1 cor_maj_87_U8 ( .A(v_1_1_3[2]), .B(cor_maj_87_n16), .Z(
        cor_maj_87_n21) );
  XOR2_X1 cor_maj_87_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_87_n16)
         );
  OR2_X1 cor_maj_87_U6 ( .A1(cor_maj_87_n20), .A2(cor_maj_87_n19), .ZN(
        cor_maj_87_n24) );
  NAND2_X1 cor_maj_87_U5 ( .A1(cor_maj_87_n24), .A2(cor_maj_87_n23), .ZN(
        cor_maj_87_n25) );
  NAND2_X1 cor_maj_87_U4 ( .A1(cor_maj_87_n20), .A2(cor_maj_87_n19), .ZN(
        cor_maj_87_n26) );
  NAND2_X1 cor_maj_87_U3 ( .A1(cor_maj_87_n26), .A2(cor_maj_87_n25), .ZN(
        cor_maj_87_port_o) );
  XOR2_X1 cor_maj_87_U2 ( .A(cor_maj_87_n22), .B(cor_maj_87_n21), .Z(
        cor_maj_87_n23) );
  NAND2_X1 cor_maj_88_U15 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_88_n18) );
  NAND2_X1 cor_maj_88_U14 ( .A1(cor_maj_88_n21), .A2(cor_maj_88_n22), .ZN(
        cor_maj_88_n17) );
  NAND2_X1 cor_maj_88_U13 ( .A1(cor_maj_88_n18), .A2(cor_maj_88_n17), .ZN(
        cor_maj_88_n19) );
  NAND2_X1 cor_maj_88_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_88_n16), .ZN(
        cor_maj_88_n14) );
  NAND2_X1 cor_maj_88_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_88_n15) );
  NAND2_X1 cor_maj_88_U10 ( .A1(cor_maj_88_n15), .A2(cor_maj_88_n14), .ZN(
        cor_maj_88_n20) );
  XOR2_X1 cor_maj_88_U9 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_88_n22)
         );
  XOR2_X1 cor_maj_88_U8 ( .A(v_1_1_3[2]), .B(cor_maj_88_n16), .Z(
        cor_maj_88_n21) );
  XOR2_X1 cor_maj_88_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_88_n16)
         );
  OR2_X1 cor_maj_88_U6 ( .A1(cor_maj_88_n20), .A2(cor_maj_88_n19), .ZN(
        cor_maj_88_n24) );
  NAND2_X1 cor_maj_88_U5 ( .A1(cor_maj_88_n24), .A2(cor_maj_88_n23), .ZN(
        cor_maj_88_n25) );
  NAND2_X1 cor_maj_88_U4 ( .A1(cor_maj_88_n20), .A2(cor_maj_88_n19), .ZN(
        cor_maj_88_n26) );
  NAND2_X1 cor_maj_88_U3 ( .A1(cor_maj_88_n26), .A2(cor_maj_88_n25), .ZN(
        cor_maj_88_port_o) );
  XOR2_X1 cor_maj_88_U2 ( .A(cor_maj_88_n22), .B(cor_maj_88_n21), .Z(
        cor_maj_88_n23) );
  NAND2_X1 cor_maj_89_U15 ( .A1(v_1_1_3[3]), .A2(v_1_1_3[4]), .ZN(
        cor_maj_89_n18) );
  NAND2_X1 cor_maj_89_U14 ( .A1(cor_maj_89_n21), .A2(cor_maj_89_n22), .ZN(
        cor_maj_89_n17) );
  NAND2_X1 cor_maj_89_U13 ( .A1(cor_maj_89_n18), .A2(cor_maj_89_n17), .ZN(
        cor_maj_89_n19) );
  NAND2_X1 cor_maj_89_U12 ( .A1(v_1_1_3[2]), .A2(cor_maj_89_n16), .ZN(
        cor_maj_89_n14) );
  NAND2_X1 cor_maj_89_U11 ( .A1(v_1_1_3[0]), .A2(v_1_1_3[1]), .ZN(
        cor_maj_89_n15) );
  NAND2_X1 cor_maj_89_U10 ( .A1(cor_maj_89_n15), .A2(cor_maj_89_n14), .ZN(
        cor_maj_89_n20) );
  XOR2_X1 cor_maj_89_U9 ( .A(v_1_1_3[3]), .B(v_1_1_3[4]), .Z(cor_maj_89_n22)
         );
  XOR2_X1 cor_maj_89_U8 ( .A(v_1_1_3[2]), .B(cor_maj_89_n16), .Z(
        cor_maj_89_n21) );
  XOR2_X1 cor_maj_89_U7 ( .A(v_1_1_3[0]), .B(v_1_1_3[1]), .Z(cor_maj_89_n16)
         );
  OR2_X1 cor_maj_89_U6 ( .A1(cor_maj_89_n20), .A2(cor_maj_89_n19), .ZN(
        cor_maj_89_n24) );
  NAND2_X1 cor_maj_89_U5 ( .A1(cor_maj_89_n24), .A2(cor_maj_89_n23), .ZN(
        cor_maj_89_n25) );
  NAND2_X1 cor_maj_89_U4 ( .A1(cor_maj_89_n20), .A2(cor_maj_89_n19), .ZN(
        cor_maj_89_n26) );
  NAND2_X1 cor_maj_89_U3 ( .A1(cor_maj_89_n26), .A2(cor_maj_89_n25), .ZN(
        cor_maj_89_port_o) );
  XOR2_X1 cor_maj_89_U2 ( .A(cor_maj_89_n22), .B(cor_maj_89_n21), .Z(
        cor_maj_89_n23) );
  NAND2_X1 cor_maj_90_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_90_n18) );
  NAND2_X1 cor_maj_90_U14 ( .A1(cor_maj_90_n21), .A2(cor_maj_90_n22), .ZN(
        cor_maj_90_n17) );
  NAND2_X1 cor_maj_90_U13 ( .A1(cor_maj_90_n18), .A2(cor_maj_90_n17), .ZN(
        cor_maj_90_n19) );
  NAND2_X1 cor_maj_90_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_90_n16), .ZN(
        cor_maj_90_n14) );
  NAND2_X1 cor_maj_90_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_90_n15) );
  NAND2_X1 cor_maj_90_U10 ( .A1(cor_maj_90_n15), .A2(cor_maj_90_n14), .ZN(
        cor_maj_90_n20) );
  XOR2_X1 cor_maj_90_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_90_n22)
         );
  XOR2_X1 cor_maj_90_U8 ( .A(v_1_2_0[2]), .B(cor_maj_90_n16), .Z(
        cor_maj_90_n21) );
  XOR2_X1 cor_maj_90_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_90_n16)
         );
  OR2_X1 cor_maj_90_U6 ( .A1(cor_maj_90_n20), .A2(cor_maj_90_n19), .ZN(
        cor_maj_90_n24) );
  NAND2_X1 cor_maj_90_U5 ( .A1(cor_maj_90_n24), .A2(cor_maj_90_n23), .ZN(
        cor_maj_90_n25) );
  NAND2_X1 cor_maj_90_U4 ( .A1(cor_maj_90_n20), .A2(cor_maj_90_n19), .ZN(
        cor_maj_90_n26) );
  NAND2_X1 cor_maj_90_U3 ( .A1(cor_maj_90_n26), .A2(cor_maj_90_n25), .ZN(
        cor_maj_90_port_o) );
  XOR2_X1 cor_maj_90_U2 ( .A(cor_maj_90_n22), .B(cor_maj_90_n21), .Z(
        cor_maj_90_n23) );
  NAND2_X1 cor_maj_91_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_91_n18) );
  NAND2_X1 cor_maj_91_U14 ( .A1(cor_maj_91_n21), .A2(cor_maj_91_n22), .ZN(
        cor_maj_91_n17) );
  NAND2_X1 cor_maj_91_U13 ( .A1(cor_maj_91_n18), .A2(cor_maj_91_n17), .ZN(
        cor_maj_91_n19) );
  NAND2_X1 cor_maj_91_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_91_n16), .ZN(
        cor_maj_91_n14) );
  NAND2_X1 cor_maj_91_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_91_n15) );
  NAND2_X1 cor_maj_91_U10 ( .A1(cor_maj_91_n15), .A2(cor_maj_91_n14), .ZN(
        cor_maj_91_n20) );
  XOR2_X1 cor_maj_91_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_91_n22)
         );
  XOR2_X1 cor_maj_91_U8 ( .A(v_1_2_0[2]), .B(cor_maj_91_n16), .Z(
        cor_maj_91_n21) );
  XOR2_X1 cor_maj_91_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_91_n16)
         );
  OR2_X1 cor_maj_91_U6 ( .A1(cor_maj_91_n20), .A2(cor_maj_91_n19), .ZN(
        cor_maj_91_n24) );
  NAND2_X1 cor_maj_91_U5 ( .A1(cor_maj_91_n24), .A2(cor_maj_91_n23), .ZN(
        cor_maj_91_n25) );
  NAND2_X1 cor_maj_91_U4 ( .A1(cor_maj_91_n20), .A2(cor_maj_91_n19), .ZN(
        cor_maj_91_n26) );
  NAND2_X1 cor_maj_91_U3 ( .A1(cor_maj_91_n26), .A2(cor_maj_91_n25), .ZN(
        cor_maj_91_port_o) );
  XOR2_X1 cor_maj_91_U2 ( .A(cor_maj_91_n22), .B(cor_maj_91_n21), .Z(
        cor_maj_91_n23) );
  NAND2_X1 cor_maj_92_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_92_n18) );
  NAND2_X1 cor_maj_92_U14 ( .A1(cor_maj_92_n21), .A2(cor_maj_92_n22), .ZN(
        cor_maj_92_n17) );
  NAND2_X1 cor_maj_92_U13 ( .A1(cor_maj_92_n18), .A2(cor_maj_92_n17), .ZN(
        cor_maj_92_n19) );
  NAND2_X1 cor_maj_92_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_92_n16), .ZN(
        cor_maj_92_n14) );
  NAND2_X1 cor_maj_92_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_92_n15) );
  NAND2_X1 cor_maj_92_U10 ( .A1(cor_maj_92_n15), .A2(cor_maj_92_n14), .ZN(
        cor_maj_92_n20) );
  XOR2_X1 cor_maj_92_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_92_n22)
         );
  XOR2_X1 cor_maj_92_U8 ( .A(v_1_2_0[2]), .B(cor_maj_92_n16), .Z(
        cor_maj_92_n21) );
  XOR2_X1 cor_maj_92_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_92_n16)
         );
  OR2_X1 cor_maj_92_U6 ( .A1(cor_maj_92_n20), .A2(cor_maj_92_n19), .ZN(
        cor_maj_92_n24) );
  NAND2_X1 cor_maj_92_U5 ( .A1(cor_maj_92_n24), .A2(cor_maj_92_n23), .ZN(
        cor_maj_92_n25) );
  NAND2_X1 cor_maj_92_U4 ( .A1(cor_maj_92_n20), .A2(cor_maj_92_n19), .ZN(
        cor_maj_92_n26) );
  NAND2_X1 cor_maj_92_U3 ( .A1(cor_maj_92_n26), .A2(cor_maj_92_n25), .ZN(
        cor_maj_92_port_o) );
  XOR2_X1 cor_maj_92_U2 ( .A(cor_maj_92_n22), .B(cor_maj_92_n21), .Z(
        cor_maj_92_n23) );
  NAND2_X1 cor_maj_93_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_93_n18) );
  NAND2_X1 cor_maj_93_U14 ( .A1(cor_maj_93_n21), .A2(cor_maj_93_n22), .ZN(
        cor_maj_93_n17) );
  NAND2_X1 cor_maj_93_U13 ( .A1(cor_maj_93_n18), .A2(cor_maj_93_n17), .ZN(
        cor_maj_93_n19) );
  NAND2_X1 cor_maj_93_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_93_n16), .ZN(
        cor_maj_93_n14) );
  NAND2_X1 cor_maj_93_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_93_n15) );
  NAND2_X1 cor_maj_93_U10 ( .A1(cor_maj_93_n15), .A2(cor_maj_93_n14), .ZN(
        cor_maj_93_n20) );
  XOR2_X1 cor_maj_93_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_93_n22)
         );
  XOR2_X1 cor_maj_93_U8 ( .A(v_1_2_0[2]), .B(cor_maj_93_n16), .Z(
        cor_maj_93_n21) );
  XOR2_X1 cor_maj_93_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_93_n16)
         );
  OR2_X1 cor_maj_93_U6 ( .A1(cor_maj_93_n20), .A2(cor_maj_93_n19), .ZN(
        cor_maj_93_n24) );
  NAND2_X1 cor_maj_93_U5 ( .A1(cor_maj_93_n24), .A2(cor_maj_93_n23), .ZN(
        cor_maj_93_n25) );
  NAND2_X1 cor_maj_93_U4 ( .A1(cor_maj_93_n20), .A2(cor_maj_93_n19), .ZN(
        cor_maj_93_n26) );
  NAND2_X1 cor_maj_93_U3 ( .A1(cor_maj_93_n26), .A2(cor_maj_93_n25), .ZN(
        cor_maj_93_port_o) );
  XOR2_X1 cor_maj_93_U2 ( .A(cor_maj_93_n22), .B(cor_maj_93_n21), .Z(
        cor_maj_93_n23) );
  NAND2_X1 cor_maj_94_U15 ( .A1(v_1_2_0[3]), .A2(v_1_2_0[4]), .ZN(
        cor_maj_94_n18) );
  NAND2_X1 cor_maj_94_U14 ( .A1(cor_maj_94_n21), .A2(cor_maj_94_n22), .ZN(
        cor_maj_94_n17) );
  NAND2_X1 cor_maj_94_U13 ( .A1(cor_maj_94_n18), .A2(cor_maj_94_n17), .ZN(
        cor_maj_94_n19) );
  NAND2_X1 cor_maj_94_U12 ( .A1(v_1_2_0[2]), .A2(cor_maj_94_n16), .ZN(
        cor_maj_94_n14) );
  NAND2_X1 cor_maj_94_U11 ( .A1(v_1_2_0[0]), .A2(v_1_2_0[1]), .ZN(
        cor_maj_94_n15) );
  NAND2_X1 cor_maj_94_U10 ( .A1(cor_maj_94_n15), .A2(cor_maj_94_n14), .ZN(
        cor_maj_94_n20) );
  XOR2_X1 cor_maj_94_U9 ( .A(v_1_2_0[3]), .B(v_1_2_0[4]), .Z(cor_maj_94_n22)
         );
  XOR2_X1 cor_maj_94_U8 ( .A(v_1_2_0[2]), .B(cor_maj_94_n16), .Z(
        cor_maj_94_n21) );
  XOR2_X1 cor_maj_94_U7 ( .A(v_1_2_0[0]), .B(v_1_2_0[1]), .Z(cor_maj_94_n16)
         );
  OR2_X1 cor_maj_94_U6 ( .A1(cor_maj_94_n20), .A2(cor_maj_94_n19), .ZN(
        cor_maj_94_n24) );
  NAND2_X1 cor_maj_94_U5 ( .A1(cor_maj_94_n24), .A2(cor_maj_94_n23), .ZN(
        cor_maj_94_n25) );
  NAND2_X1 cor_maj_94_U4 ( .A1(cor_maj_94_n20), .A2(cor_maj_94_n19), .ZN(
        cor_maj_94_n26) );
  NAND2_X1 cor_maj_94_U3 ( .A1(cor_maj_94_n26), .A2(cor_maj_94_n25), .ZN(
        cor_maj_94_port_o) );
  XOR2_X1 cor_maj_94_U2 ( .A(cor_maj_94_n22), .B(cor_maj_94_n21), .Z(
        cor_maj_94_n23) );
  NAND2_X1 cor_maj_95_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_95_n18) );
  NAND2_X1 cor_maj_95_U14 ( .A1(cor_maj_95_n21), .A2(cor_maj_95_n22), .ZN(
        cor_maj_95_n17) );
  NAND2_X1 cor_maj_95_U13 ( .A1(cor_maj_95_n18), .A2(cor_maj_95_n17), .ZN(
        cor_maj_95_n19) );
  NAND2_X1 cor_maj_95_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_95_n16), .ZN(
        cor_maj_95_n14) );
  NAND2_X1 cor_maj_95_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_95_n15) );
  NAND2_X1 cor_maj_95_U10 ( .A1(cor_maj_95_n15), .A2(cor_maj_95_n14), .ZN(
        cor_maj_95_n20) );
  XOR2_X1 cor_maj_95_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_95_n22)
         );
  XOR2_X1 cor_maj_95_U8 ( .A(v_1_2_1[2]), .B(cor_maj_95_n16), .Z(
        cor_maj_95_n21) );
  XOR2_X1 cor_maj_95_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_95_n16)
         );
  OR2_X1 cor_maj_95_U6 ( .A1(cor_maj_95_n20), .A2(cor_maj_95_n19), .ZN(
        cor_maj_95_n24) );
  NAND2_X1 cor_maj_95_U5 ( .A1(cor_maj_95_n24), .A2(cor_maj_95_n23), .ZN(
        cor_maj_95_n25) );
  NAND2_X1 cor_maj_95_U4 ( .A1(cor_maj_95_n20), .A2(cor_maj_95_n19), .ZN(
        cor_maj_95_n26) );
  NAND2_X1 cor_maj_95_U3 ( .A1(cor_maj_95_n26), .A2(cor_maj_95_n25), .ZN(
        cor_maj_95_port_o) );
  XOR2_X1 cor_maj_95_U2 ( .A(cor_maj_95_n22), .B(cor_maj_95_n21), .Z(
        cor_maj_95_n23) );
  NAND2_X1 cor_maj_96_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_96_n18) );
  NAND2_X1 cor_maj_96_U14 ( .A1(cor_maj_96_n21), .A2(cor_maj_96_n22), .ZN(
        cor_maj_96_n17) );
  NAND2_X1 cor_maj_96_U13 ( .A1(cor_maj_96_n18), .A2(cor_maj_96_n17), .ZN(
        cor_maj_96_n19) );
  NAND2_X1 cor_maj_96_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_96_n16), .ZN(
        cor_maj_96_n14) );
  NAND2_X1 cor_maj_96_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_96_n15) );
  NAND2_X1 cor_maj_96_U10 ( .A1(cor_maj_96_n15), .A2(cor_maj_96_n14), .ZN(
        cor_maj_96_n20) );
  XOR2_X1 cor_maj_96_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_96_n22)
         );
  XOR2_X1 cor_maj_96_U8 ( .A(v_1_2_1[2]), .B(cor_maj_96_n16), .Z(
        cor_maj_96_n21) );
  XOR2_X1 cor_maj_96_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_96_n16)
         );
  OR2_X1 cor_maj_96_U6 ( .A1(cor_maj_96_n20), .A2(cor_maj_96_n19), .ZN(
        cor_maj_96_n24) );
  NAND2_X1 cor_maj_96_U5 ( .A1(cor_maj_96_n24), .A2(cor_maj_96_n23), .ZN(
        cor_maj_96_n25) );
  NAND2_X1 cor_maj_96_U4 ( .A1(cor_maj_96_n20), .A2(cor_maj_96_n19), .ZN(
        cor_maj_96_n26) );
  NAND2_X1 cor_maj_96_U3 ( .A1(cor_maj_96_n26), .A2(cor_maj_96_n25), .ZN(
        cor_maj_96_port_o) );
  XOR2_X1 cor_maj_96_U2 ( .A(cor_maj_96_n22), .B(cor_maj_96_n21), .Z(
        cor_maj_96_n23) );
  NAND2_X1 cor_maj_97_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_97_n18) );
  NAND2_X1 cor_maj_97_U14 ( .A1(cor_maj_97_n21), .A2(cor_maj_97_n22), .ZN(
        cor_maj_97_n17) );
  NAND2_X1 cor_maj_97_U13 ( .A1(cor_maj_97_n18), .A2(cor_maj_97_n17), .ZN(
        cor_maj_97_n19) );
  NAND2_X1 cor_maj_97_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_97_n16), .ZN(
        cor_maj_97_n14) );
  NAND2_X1 cor_maj_97_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_97_n15) );
  NAND2_X1 cor_maj_97_U10 ( .A1(cor_maj_97_n15), .A2(cor_maj_97_n14), .ZN(
        cor_maj_97_n20) );
  XOR2_X1 cor_maj_97_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_97_n22)
         );
  XOR2_X1 cor_maj_97_U8 ( .A(v_1_2_1[2]), .B(cor_maj_97_n16), .Z(
        cor_maj_97_n21) );
  XOR2_X1 cor_maj_97_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_97_n16)
         );
  OR2_X1 cor_maj_97_U6 ( .A1(cor_maj_97_n20), .A2(cor_maj_97_n19), .ZN(
        cor_maj_97_n24) );
  NAND2_X1 cor_maj_97_U5 ( .A1(cor_maj_97_n24), .A2(cor_maj_97_n23), .ZN(
        cor_maj_97_n25) );
  NAND2_X1 cor_maj_97_U4 ( .A1(cor_maj_97_n20), .A2(cor_maj_97_n19), .ZN(
        cor_maj_97_n26) );
  NAND2_X1 cor_maj_97_U3 ( .A1(cor_maj_97_n26), .A2(cor_maj_97_n25), .ZN(
        cor_maj_97_port_o) );
  XOR2_X1 cor_maj_97_U2 ( .A(cor_maj_97_n22), .B(cor_maj_97_n21), .Z(
        cor_maj_97_n23) );
  NAND2_X1 cor_maj_98_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_98_n18) );
  NAND2_X1 cor_maj_98_U14 ( .A1(cor_maj_98_n21), .A2(cor_maj_98_n22), .ZN(
        cor_maj_98_n17) );
  NAND2_X1 cor_maj_98_U13 ( .A1(cor_maj_98_n18), .A2(cor_maj_98_n17), .ZN(
        cor_maj_98_n19) );
  NAND2_X1 cor_maj_98_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_98_n16), .ZN(
        cor_maj_98_n14) );
  NAND2_X1 cor_maj_98_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_98_n15) );
  NAND2_X1 cor_maj_98_U10 ( .A1(cor_maj_98_n15), .A2(cor_maj_98_n14), .ZN(
        cor_maj_98_n20) );
  XOR2_X1 cor_maj_98_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_98_n22)
         );
  XOR2_X1 cor_maj_98_U8 ( .A(v_1_2_1[2]), .B(cor_maj_98_n16), .Z(
        cor_maj_98_n21) );
  XOR2_X1 cor_maj_98_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_98_n16)
         );
  OR2_X1 cor_maj_98_U6 ( .A1(cor_maj_98_n20), .A2(cor_maj_98_n19), .ZN(
        cor_maj_98_n24) );
  NAND2_X1 cor_maj_98_U5 ( .A1(cor_maj_98_n24), .A2(cor_maj_98_n23), .ZN(
        cor_maj_98_n25) );
  NAND2_X1 cor_maj_98_U4 ( .A1(cor_maj_98_n20), .A2(cor_maj_98_n19), .ZN(
        cor_maj_98_n26) );
  NAND2_X1 cor_maj_98_U3 ( .A1(cor_maj_98_n26), .A2(cor_maj_98_n25), .ZN(
        cor_maj_98_port_o) );
  XOR2_X1 cor_maj_98_U2 ( .A(cor_maj_98_n22), .B(cor_maj_98_n21), .Z(
        cor_maj_98_n23) );
  NAND2_X1 cor_maj_99_U15 ( .A1(v_1_2_1[3]), .A2(v_1_2_1[4]), .ZN(
        cor_maj_99_n18) );
  NAND2_X1 cor_maj_99_U14 ( .A1(cor_maj_99_n21), .A2(cor_maj_99_n22), .ZN(
        cor_maj_99_n17) );
  NAND2_X1 cor_maj_99_U13 ( .A1(cor_maj_99_n18), .A2(cor_maj_99_n17), .ZN(
        cor_maj_99_n19) );
  NAND2_X1 cor_maj_99_U12 ( .A1(v_1_2_1[2]), .A2(cor_maj_99_n16), .ZN(
        cor_maj_99_n14) );
  NAND2_X1 cor_maj_99_U11 ( .A1(v_1_2_1[0]), .A2(v_1_2_1[1]), .ZN(
        cor_maj_99_n15) );
  NAND2_X1 cor_maj_99_U10 ( .A1(cor_maj_99_n15), .A2(cor_maj_99_n14), .ZN(
        cor_maj_99_n20) );
  XOR2_X1 cor_maj_99_U9 ( .A(v_1_2_1[3]), .B(v_1_2_1[4]), .Z(cor_maj_99_n22)
         );
  XOR2_X1 cor_maj_99_U8 ( .A(v_1_2_1[2]), .B(cor_maj_99_n16), .Z(
        cor_maj_99_n21) );
  XOR2_X1 cor_maj_99_U7 ( .A(v_1_2_1[0]), .B(v_1_2_1[1]), .Z(cor_maj_99_n16)
         );
  OR2_X1 cor_maj_99_U6 ( .A1(cor_maj_99_n20), .A2(cor_maj_99_n19), .ZN(
        cor_maj_99_n24) );
  NAND2_X1 cor_maj_99_U5 ( .A1(cor_maj_99_n24), .A2(cor_maj_99_n23), .ZN(
        cor_maj_99_n25) );
  NAND2_X1 cor_maj_99_U4 ( .A1(cor_maj_99_n20), .A2(cor_maj_99_n19), .ZN(
        cor_maj_99_n26) );
  NAND2_X1 cor_maj_99_U3 ( .A1(cor_maj_99_n26), .A2(cor_maj_99_n25), .ZN(
        cor_maj_99_port_o) );
  XOR2_X1 cor_maj_99_U2 ( .A(cor_maj_99_n22), .B(cor_maj_99_n21), .Z(
        cor_maj_99_n23) );
  NAND2_X1 cor_maj_100_U15 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_100_n18) );
  NAND2_X1 cor_maj_100_U14 ( .A1(cor_maj_100_n21), .A2(cor_maj_100_n22), .ZN(
        cor_maj_100_n17) );
  NAND2_X1 cor_maj_100_U13 ( .A1(cor_maj_100_n18), .A2(cor_maj_100_n17), .ZN(
        cor_maj_100_n19) );
  NAND2_X1 cor_maj_100_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_100_n16), .ZN(
        cor_maj_100_n14) );
  NAND2_X1 cor_maj_100_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_100_n15) );
  NAND2_X1 cor_maj_100_U10 ( .A1(cor_maj_100_n15), .A2(cor_maj_100_n14), .ZN(
        cor_maj_100_n20) );
  XOR2_X1 cor_maj_100_U9 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_100_n22)
         );
  XOR2_X1 cor_maj_100_U8 ( .A(v_1_2_3[2]), .B(cor_maj_100_n16), .Z(
        cor_maj_100_n21) );
  XOR2_X1 cor_maj_100_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_100_n16)
         );
  OR2_X1 cor_maj_100_U6 ( .A1(cor_maj_100_n20), .A2(cor_maj_100_n19), .ZN(
        cor_maj_100_n24) );
  NAND2_X1 cor_maj_100_U5 ( .A1(cor_maj_100_n24), .A2(cor_maj_100_n23), .ZN(
        cor_maj_100_n25) );
  NAND2_X1 cor_maj_100_U4 ( .A1(cor_maj_100_n20), .A2(cor_maj_100_n19), .ZN(
        cor_maj_100_n26) );
  NAND2_X1 cor_maj_100_U3 ( .A1(cor_maj_100_n26), .A2(cor_maj_100_n25), .ZN(
        cor_maj_100_port_o) );
  XOR2_X1 cor_maj_100_U2 ( .A(cor_maj_100_n22), .B(cor_maj_100_n21), .Z(
        cor_maj_100_n23) );
  NAND2_X1 cor_maj_101_U15 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_101_n18) );
  NAND2_X1 cor_maj_101_U14 ( .A1(cor_maj_101_n21), .A2(cor_maj_101_n22), .ZN(
        cor_maj_101_n17) );
  NAND2_X1 cor_maj_101_U13 ( .A1(cor_maj_101_n18), .A2(cor_maj_101_n17), .ZN(
        cor_maj_101_n19) );
  NAND2_X1 cor_maj_101_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_101_n16), .ZN(
        cor_maj_101_n14) );
  NAND2_X1 cor_maj_101_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_101_n15) );
  NAND2_X1 cor_maj_101_U10 ( .A1(cor_maj_101_n15), .A2(cor_maj_101_n14), .ZN(
        cor_maj_101_n20) );
  XOR2_X1 cor_maj_101_U9 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_101_n22)
         );
  XOR2_X1 cor_maj_101_U8 ( .A(v_1_2_3[2]), .B(cor_maj_101_n16), .Z(
        cor_maj_101_n21) );
  XOR2_X1 cor_maj_101_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_101_n16)
         );
  OR2_X1 cor_maj_101_U6 ( .A1(cor_maj_101_n20), .A2(cor_maj_101_n19), .ZN(
        cor_maj_101_n24) );
  NAND2_X1 cor_maj_101_U5 ( .A1(cor_maj_101_n24), .A2(cor_maj_101_n23), .ZN(
        cor_maj_101_n25) );
  NAND2_X1 cor_maj_101_U4 ( .A1(cor_maj_101_n20), .A2(cor_maj_101_n19), .ZN(
        cor_maj_101_n26) );
  NAND2_X1 cor_maj_101_U3 ( .A1(cor_maj_101_n26), .A2(cor_maj_101_n25), .ZN(
        cor_maj_101_port_o) );
  XOR2_X1 cor_maj_101_U2 ( .A(cor_maj_101_n22), .B(cor_maj_101_n21), .Z(
        cor_maj_101_n23) );
  NAND2_X1 cor_maj_102_U15 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_102_n18) );
  NAND2_X1 cor_maj_102_U14 ( .A1(cor_maj_102_n21), .A2(cor_maj_102_n22), .ZN(
        cor_maj_102_n17) );
  NAND2_X1 cor_maj_102_U13 ( .A1(cor_maj_102_n18), .A2(cor_maj_102_n17), .ZN(
        cor_maj_102_n19) );
  NAND2_X1 cor_maj_102_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_102_n16), .ZN(
        cor_maj_102_n14) );
  NAND2_X1 cor_maj_102_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_102_n15) );
  NAND2_X1 cor_maj_102_U10 ( .A1(cor_maj_102_n15), .A2(cor_maj_102_n14), .ZN(
        cor_maj_102_n20) );
  XOR2_X1 cor_maj_102_U9 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_102_n22)
         );
  XOR2_X1 cor_maj_102_U8 ( .A(v_1_2_3[2]), .B(cor_maj_102_n16), .Z(
        cor_maj_102_n21) );
  XOR2_X1 cor_maj_102_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_102_n16)
         );
  OR2_X1 cor_maj_102_U6 ( .A1(cor_maj_102_n20), .A2(cor_maj_102_n19), .ZN(
        cor_maj_102_n24) );
  NAND2_X1 cor_maj_102_U5 ( .A1(cor_maj_102_n24), .A2(cor_maj_102_n23), .ZN(
        cor_maj_102_n25) );
  NAND2_X1 cor_maj_102_U4 ( .A1(cor_maj_102_n20), .A2(cor_maj_102_n19), .ZN(
        cor_maj_102_n26) );
  NAND2_X1 cor_maj_102_U3 ( .A1(cor_maj_102_n26), .A2(cor_maj_102_n25), .ZN(
        cor_maj_102_port_o) );
  XOR2_X1 cor_maj_102_U2 ( .A(cor_maj_102_n22), .B(cor_maj_102_n21), .Z(
        cor_maj_102_n23) );
  NAND2_X1 cor_maj_103_U15 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_103_n18) );
  NAND2_X1 cor_maj_103_U14 ( .A1(cor_maj_103_n21), .A2(cor_maj_103_n22), .ZN(
        cor_maj_103_n17) );
  NAND2_X1 cor_maj_103_U13 ( .A1(cor_maj_103_n18), .A2(cor_maj_103_n17), .ZN(
        cor_maj_103_n19) );
  NAND2_X1 cor_maj_103_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_103_n16), .ZN(
        cor_maj_103_n14) );
  NAND2_X1 cor_maj_103_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_103_n15) );
  NAND2_X1 cor_maj_103_U10 ( .A1(cor_maj_103_n15), .A2(cor_maj_103_n14), .ZN(
        cor_maj_103_n20) );
  XOR2_X1 cor_maj_103_U9 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_103_n22)
         );
  XOR2_X1 cor_maj_103_U8 ( .A(v_1_2_3[2]), .B(cor_maj_103_n16), .Z(
        cor_maj_103_n21) );
  XOR2_X1 cor_maj_103_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_103_n16)
         );
  OR2_X1 cor_maj_103_U6 ( .A1(cor_maj_103_n20), .A2(cor_maj_103_n19), .ZN(
        cor_maj_103_n24) );
  NAND2_X1 cor_maj_103_U5 ( .A1(cor_maj_103_n24), .A2(cor_maj_103_n23), .ZN(
        cor_maj_103_n25) );
  NAND2_X1 cor_maj_103_U4 ( .A1(cor_maj_103_n20), .A2(cor_maj_103_n19), .ZN(
        cor_maj_103_n26) );
  NAND2_X1 cor_maj_103_U3 ( .A1(cor_maj_103_n26), .A2(cor_maj_103_n25), .ZN(
        cor_maj_103_port_o) );
  XOR2_X1 cor_maj_103_U2 ( .A(cor_maj_103_n22), .B(cor_maj_103_n21), .Z(
        cor_maj_103_n23) );
  NAND2_X1 cor_maj_104_U15 ( .A1(v_1_2_3[3]), .A2(v_1_2_3[4]), .ZN(
        cor_maj_104_n18) );
  NAND2_X1 cor_maj_104_U14 ( .A1(cor_maj_104_n21), .A2(cor_maj_104_n22), .ZN(
        cor_maj_104_n17) );
  NAND2_X1 cor_maj_104_U13 ( .A1(cor_maj_104_n18), .A2(cor_maj_104_n17), .ZN(
        cor_maj_104_n19) );
  NAND2_X1 cor_maj_104_U12 ( .A1(v_1_2_3[2]), .A2(cor_maj_104_n16), .ZN(
        cor_maj_104_n14) );
  NAND2_X1 cor_maj_104_U11 ( .A1(v_1_2_3[0]), .A2(v_1_2_3[1]), .ZN(
        cor_maj_104_n15) );
  NAND2_X1 cor_maj_104_U10 ( .A1(cor_maj_104_n15), .A2(cor_maj_104_n14), .ZN(
        cor_maj_104_n20) );
  XOR2_X1 cor_maj_104_U9 ( .A(v_1_2_3[3]), .B(v_1_2_3[4]), .Z(cor_maj_104_n22)
         );
  XOR2_X1 cor_maj_104_U8 ( .A(v_1_2_3[2]), .B(cor_maj_104_n16), .Z(
        cor_maj_104_n21) );
  XOR2_X1 cor_maj_104_U7 ( .A(v_1_2_3[0]), .B(v_1_2_3[1]), .Z(cor_maj_104_n16)
         );
  OR2_X1 cor_maj_104_U6 ( .A1(cor_maj_104_n20), .A2(cor_maj_104_n19), .ZN(
        cor_maj_104_n24) );
  NAND2_X1 cor_maj_104_U5 ( .A1(cor_maj_104_n24), .A2(cor_maj_104_n23), .ZN(
        cor_maj_104_n25) );
  NAND2_X1 cor_maj_104_U4 ( .A1(cor_maj_104_n20), .A2(cor_maj_104_n19), .ZN(
        cor_maj_104_n26) );
  NAND2_X1 cor_maj_104_U3 ( .A1(cor_maj_104_n26), .A2(cor_maj_104_n25), .ZN(
        cor_maj_104_port_o) );
  XOR2_X1 cor_maj_104_U2 ( .A(cor_maj_104_n22), .B(cor_maj_104_n21), .Z(
        cor_maj_104_n23) );
  NAND2_X1 cor_maj_105_U15 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_105_n18) );
  NAND2_X1 cor_maj_105_U14 ( .A1(cor_maj_105_n21), .A2(cor_maj_105_n22), .ZN(
        cor_maj_105_n17) );
  NAND2_X1 cor_maj_105_U13 ( .A1(cor_maj_105_n18), .A2(cor_maj_105_n17), .ZN(
        cor_maj_105_n19) );
  NAND2_X1 cor_maj_105_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_105_n16), .ZN(
        cor_maj_105_n14) );
  NAND2_X1 cor_maj_105_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_105_n15) );
  NAND2_X1 cor_maj_105_U10 ( .A1(cor_maj_105_n15), .A2(cor_maj_105_n14), .ZN(
        cor_maj_105_n20) );
  XOR2_X1 cor_maj_105_U9 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_105_n22)
         );
  XOR2_X1 cor_maj_105_U8 ( .A(v_1_3_0[2]), .B(cor_maj_105_n16), .Z(
        cor_maj_105_n21) );
  XOR2_X1 cor_maj_105_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_105_n16)
         );
  OR2_X1 cor_maj_105_U6 ( .A1(cor_maj_105_n20), .A2(cor_maj_105_n19), .ZN(
        cor_maj_105_n24) );
  NAND2_X1 cor_maj_105_U5 ( .A1(cor_maj_105_n24), .A2(cor_maj_105_n23), .ZN(
        cor_maj_105_n25) );
  NAND2_X1 cor_maj_105_U4 ( .A1(cor_maj_105_n20), .A2(cor_maj_105_n19), .ZN(
        cor_maj_105_n26) );
  NAND2_X1 cor_maj_105_U3 ( .A1(cor_maj_105_n26), .A2(cor_maj_105_n25), .ZN(
        cor_maj_105_port_o) );
  XOR2_X1 cor_maj_105_U2 ( .A(cor_maj_105_n22), .B(cor_maj_105_n21), .Z(
        cor_maj_105_n23) );
  NAND2_X1 cor_maj_106_U15 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_106_n18) );
  NAND2_X1 cor_maj_106_U14 ( .A1(cor_maj_106_n21), .A2(cor_maj_106_n22), .ZN(
        cor_maj_106_n17) );
  NAND2_X1 cor_maj_106_U13 ( .A1(cor_maj_106_n18), .A2(cor_maj_106_n17), .ZN(
        cor_maj_106_n19) );
  NAND2_X1 cor_maj_106_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_106_n16), .ZN(
        cor_maj_106_n14) );
  NAND2_X1 cor_maj_106_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_106_n15) );
  NAND2_X1 cor_maj_106_U10 ( .A1(cor_maj_106_n15), .A2(cor_maj_106_n14), .ZN(
        cor_maj_106_n20) );
  XOR2_X1 cor_maj_106_U9 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_106_n22)
         );
  XOR2_X1 cor_maj_106_U8 ( .A(v_1_3_0[2]), .B(cor_maj_106_n16), .Z(
        cor_maj_106_n21) );
  XOR2_X1 cor_maj_106_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_106_n16)
         );
  OR2_X1 cor_maj_106_U6 ( .A1(cor_maj_106_n20), .A2(cor_maj_106_n19), .ZN(
        cor_maj_106_n24) );
  NAND2_X1 cor_maj_106_U5 ( .A1(cor_maj_106_n24), .A2(cor_maj_106_n23), .ZN(
        cor_maj_106_n25) );
  NAND2_X1 cor_maj_106_U4 ( .A1(cor_maj_106_n20), .A2(cor_maj_106_n19), .ZN(
        cor_maj_106_n26) );
  NAND2_X1 cor_maj_106_U3 ( .A1(cor_maj_106_n26), .A2(cor_maj_106_n25), .ZN(
        cor_maj_106_port_o) );
  XOR2_X1 cor_maj_106_U2 ( .A(cor_maj_106_n22), .B(cor_maj_106_n21), .Z(
        cor_maj_106_n23) );
  NAND2_X1 cor_maj_107_U15 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_107_n18) );
  NAND2_X1 cor_maj_107_U14 ( .A1(cor_maj_107_n21), .A2(cor_maj_107_n22), .ZN(
        cor_maj_107_n17) );
  NAND2_X1 cor_maj_107_U13 ( .A1(cor_maj_107_n18), .A2(cor_maj_107_n17), .ZN(
        cor_maj_107_n19) );
  NAND2_X1 cor_maj_107_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_107_n16), .ZN(
        cor_maj_107_n14) );
  NAND2_X1 cor_maj_107_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_107_n15) );
  NAND2_X1 cor_maj_107_U10 ( .A1(cor_maj_107_n15), .A2(cor_maj_107_n14), .ZN(
        cor_maj_107_n20) );
  XOR2_X1 cor_maj_107_U9 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_107_n22)
         );
  XOR2_X1 cor_maj_107_U8 ( .A(v_1_3_0[2]), .B(cor_maj_107_n16), .Z(
        cor_maj_107_n21) );
  XOR2_X1 cor_maj_107_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_107_n16)
         );
  OR2_X1 cor_maj_107_U6 ( .A1(cor_maj_107_n20), .A2(cor_maj_107_n19), .ZN(
        cor_maj_107_n24) );
  NAND2_X1 cor_maj_107_U5 ( .A1(cor_maj_107_n24), .A2(cor_maj_107_n23), .ZN(
        cor_maj_107_n25) );
  NAND2_X1 cor_maj_107_U4 ( .A1(cor_maj_107_n20), .A2(cor_maj_107_n19), .ZN(
        cor_maj_107_n26) );
  NAND2_X1 cor_maj_107_U3 ( .A1(cor_maj_107_n26), .A2(cor_maj_107_n25), .ZN(
        cor_maj_107_port_o) );
  XOR2_X1 cor_maj_107_U2 ( .A(cor_maj_107_n22), .B(cor_maj_107_n21), .Z(
        cor_maj_107_n23) );
  NAND2_X1 cor_maj_108_U15 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_108_n18) );
  NAND2_X1 cor_maj_108_U14 ( .A1(cor_maj_108_n21), .A2(cor_maj_108_n22), .ZN(
        cor_maj_108_n17) );
  NAND2_X1 cor_maj_108_U13 ( .A1(cor_maj_108_n18), .A2(cor_maj_108_n17), .ZN(
        cor_maj_108_n19) );
  NAND2_X1 cor_maj_108_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_108_n16), .ZN(
        cor_maj_108_n14) );
  NAND2_X1 cor_maj_108_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_108_n15) );
  NAND2_X1 cor_maj_108_U10 ( .A1(cor_maj_108_n15), .A2(cor_maj_108_n14), .ZN(
        cor_maj_108_n20) );
  XOR2_X1 cor_maj_108_U9 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_108_n22)
         );
  XOR2_X1 cor_maj_108_U8 ( .A(v_1_3_0[2]), .B(cor_maj_108_n16), .Z(
        cor_maj_108_n21) );
  XOR2_X1 cor_maj_108_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_108_n16)
         );
  OR2_X1 cor_maj_108_U6 ( .A1(cor_maj_108_n20), .A2(cor_maj_108_n19), .ZN(
        cor_maj_108_n24) );
  NAND2_X1 cor_maj_108_U5 ( .A1(cor_maj_108_n24), .A2(cor_maj_108_n23), .ZN(
        cor_maj_108_n25) );
  NAND2_X1 cor_maj_108_U4 ( .A1(cor_maj_108_n20), .A2(cor_maj_108_n19), .ZN(
        cor_maj_108_n26) );
  NAND2_X1 cor_maj_108_U3 ( .A1(cor_maj_108_n26), .A2(cor_maj_108_n25), .ZN(
        cor_maj_108_port_o) );
  XOR2_X1 cor_maj_108_U2 ( .A(cor_maj_108_n22), .B(cor_maj_108_n21), .Z(
        cor_maj_108_n23) );
  NAND2_X1 cor_maj_109_U15 ( .A1(v_1_3_0[3]), .A2(v_1_3_0[4]), .ZN(
        cor_maj_109_n18) );
  NAND2_X1 cor_maj_109_U14 ( .A1(cor_maj_109_n21), .A2(cor_maj_109_n22), .ZN(
        cor_maj_109_n17) );
  NAND2_X1 cor_maj_109_U13 ( .A1(cor_maj_109_n18), .A2(cor_maj_109_n17), .ZN(
        cor_maj_109_n19) );
  NAND2_X1 cor_maj_109_U12 ( .A1(v_1_3_0[2]), .A2(cor_maj_109_n16), .ZN(
        cor_maj_109_n14) );
  NAND2_X1 cor_maj_109_U11 ( .A1(v_1_3_0[0]), .A2(v_1_3_0[1]), .ZN(
        cor_maj_109_n15) );
  NAND2_X1 cor_maj_109_U10 ( .A1(cor_maj_109_n15), .A2(cor_maj_109_n14), .ZN(
        cor_maj_109_n20) );
  XOR2_X1 cor_maj_109_U9 ( .A(v_1_3_0[3]), .B(v_1_3_0[4]), .Z(cor_maj_109_n22)
         );
  XOR2_X1 cor_maj_109_U8 ( .A(v_1_3_0[2]), .B(cor_maj_109_n16), .Z(
        cor_maj_109_n21) );
  XOR2_X1 cor_maj_109_U7 ( .A(v_1_3_0[0]), .B(v_1_3_0[1]), .Z(cor_maj_109_n16)
         );
  OR2_X1 cor_maj_109_U6 ( .A1(cor_maj_109_n20), .A2(cor_maj_109_n19), .ZN(
        cor_maj_109_n24) );
  NAND2_X1 cor_maj_109_U5 ( .A1(cor_maj_109_n24), .A2(cor_maj_109_n23), .ZN(
        cor_maj_109_n25) );
  NAND2_X1 cor_maj_109_U4 ( .A1(cor_maj_109_n20), .A2(cor_maj_109_n19), .ZN(
        cor_maj_109_n26) );
  NAND2_X1 cor_maj_109_U3 ( .A1(cor_maj_109_n26), .A2(cor_maj_109_n25), .ZN(
        cor_maj_109_port_o) );
  XOR2_X1 cor_maj_109_U2 ( .A(cor_maj_109_n22), .B(cor_maj_109_n21), .Z(
        cor_maj_109_n23) );
  NAND2_X1 cor_maj_110_U15 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_110_n18) );
  NAND2_X1 cor_maj_110_U14 ( .A1(cor_maj_110_n21), .A2(cor_maj_110_n22), .ZN(
        cor_maj_110_n17) );
  NAND2_X1 cor_maj_110_U13 ( .A1(cor_maj_110_n18), .A2(cor_maj_110_n17), .ZN(
        cor_maj_110_n19) );
  NAND2_X1 cor_maj_110_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_110_n16), .ZN(
        cor_maj_110_n14) );
  NAND2_X1 cor_maj_110_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_110_n15) );
  NAND2_X1 cor_maj_110_U10 ( .A1(cor_maj_110_n15), .A2(cor_maj_110_n14), .ZN(
        cor_maj_110_n20) );
  XOR2_X1 cor_maj_110_U9 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_110_n22)
         );
  XOR2_X1 cor_maj_110_U8 ( .A(v_1_3_1[2]), .B(cor_maj_110_n16), .Z(
        cor_maj_110_n21) );
  XOR2_X1 cor_maj_110_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_110_n16)
         );
  OR2_X1 cor_maj_110_U6 ( .A1(cor_maj_110_n20), .A2(cor_maj_110_n19), .ZN(
        cor_maj_110_n24) );
  NAND2_X1 cor_maj_110_U5 ( .A1(cor_maj_110_n24), .A2(cor_maj_110_n23), .ZN(
        cor_maj_110_n25) );
  NAND2_X1 cor_maj_110_U4 ( .A1(cor_maj_110_n20), .A2(cor_maj_110_n19), .ZN(
        cor_maj_110_n26) );
  NAND2_X1 cor_maj_110_U3 ( .A1(cor_maj_110_n26), .A2(cor_maj_110_n25), .ZN(
        cor_maj_110_port_o) );
  XOR2_X1 cor_maj_110_U2 ( .A(cor_maj_110_n22), .B(cor_maj_110_n21), .Z(
        cor_maj_110_n23) );
  NAND2_X1 cor_maj_111_U15 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_111_n18) );
  NAND2_X1 cor_maj_111_U14 ( .A1(cor_maj_111_n21), .A2(cor_maj_111_n22), .ZN(
        cor_maj_111_n17) );
  NAND2_X1 cor_maj_111_U13 ( .A1(cor_maj_111_n18), .A2(cor_maj_111_n17), .ZN(
        cor_maj_111_n19) );
  NAND2_X1 cor_maj_111_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_111_n16), .ZN(
        cor_maj_111_n14) );
  NAND2_X1 cor_maj_111_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_111_n15) );
  NAND2_X1 cor_maj_111_U10 ( .A1(cor_maj_111_n15), .A2(cor_maj_111_n14), .ZN(
        cor_maj_111_n20) );
  XOR2_X1 cor_maj_111_U9 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_111_n22)
         );
  XOR2_X1 cor_maj_111_U8 ( .A(v_1_3_1[2]), .B(cor_maj_111_n16), .Z(
        cor_maj_111_n21) );
  XOR2_X1 cor_maj_111_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_111_n16)
         );
  OR2_X1 cor_maj_111_U6 ( .A1(cor_maj_111_n20), .A2(cor_maj_111_n19), .ZN(
        cor_maj_111_n24) );
  NAND2_X1 cor_maj_111_U5 ( .A1(cor_maj_111_n24), .A2(cor_maj_111_n23), .ZN(
        cor_maj_111_n25) );
  NAND2_X1 cor_maj_111_U4 ( .A1(cor_maj_111_n20), .A2(cor_maj_111_n19), .ZN(
        cor_maj_111_n26) );
  NAND2_X1 cor_maj_111_U3 ( .A1(cor_maj_111_n26), .A2(cor_maj_111_n25), .ZN(
        cor_maj_111_port_o) );
  XOR2_X1 cor_maj_111_U2 ( .A(cor_maj_111_n22), .B(cor_maj_111_n21), .Z(
        cor_maj_111_n23) );
  NAND2_X1 cor_maj_112_U15 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_112_n18) );
  NAND2_X1 cor_maj_112_U14 ( .A1(cor_maj_112_n21), .A2(cor_maj_112_n22), .ZN(
        cor_maj_112_n17) );
  NAND2_X1 cor_maj_112_U13 ( .A1(cor_maj_112_n18), .A2(cor_maj_112_n17), .ZN(
        cor_maj_112_n19) );
  NAND2_X1 cor_maj_112_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_112_n16), .ZN(
        cor_maj_112_n14) );
  NAND2_X1 cor_maj_112_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_112_n15) );
  NAND2_X1 cor_maj_112_U10 ( .A1(cor_maj_112_n15), .A2(cor_maj_112_n14), .ZN(
        cor_maj_112_n20) );
  XOR2_X1 cor_maj_112_U9 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_112_n22)
         );
  XOR2_X1 cor_maj_112_U8 ( .A(v_1_3_1[2]), .B(cor_maj_112_n16), .Z(
        cor_maj_112_n21) );
  XOR2_X1 cor_maj_112_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_112_n16)
         );
  OR2_X1 cor_maj_112_U6 ( .A1(cor_maj_112_n20), .A2(cor_maj_112_n19), .ZN(
        cor_maj_112_n24) );
  NAND2_X1 cor_maj_112_U5 ( .A1(cor_maj_112_n24), .A2(cor_maj_112_n23), .ZN(
        cor_maj_112_n25) );
  NAND2_X1 cor_maj_112_U4 ( .A1(cor_maj_112_n20), .A2(cor_maj_112_n19), .ZN(
        cor_maj_112_n26) );
  NAND2_X1 cor_maj_112_U3 ( .A1(cor_maj_112_n26), .A2(cor_maj_112_n25), .ZN(
        cor_maj_112_port_o) );
  XOR2_X1 cor_maj_112_U2 ( .A(cor_maj_112_n22), .B(cor_maj_112_n21), .Z(
        cor_maj_112_n23) );
  NAND2_X1 cor_maj_113_U15 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_113_n18) );
  NAND2_X1 cor_maj_113_U14 ( .A1(cor_maj_113_n21), .A2(cor_maj_113_n22), .ZN(
        cor_maj_113_n17) );
  NAND2_X1 cor_maj_113_U13 ( .A1(cor_maj_113_n18), .A2(cor_maj_113_n17), .ZN(
        cor_maj_113_n19) );
  NAND2_X1 cor_maj_113_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_113_n16), .ZN(
        cor_maj_113_n14) );
  NAND2_X1 cor_maj_113_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_113_n15) );
  NAND2_X1 cor_maj_113_U10 ( .A1(cor_maj_113_n15), .A2(cor_maj_113_n14), .ZN(
        cor_maj_113_n20) );
  XOR2_X1 cor_maj_113_U9 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_113_n22)
         );
  XOR2_X1 cor_maj_113_U8 ( .A(v_1_3_1[2]), .B(cor_maj_113_n16), .Z(
        cor_maj_113_n21) );
  XOR2_X1 cor_maj_113_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_113_n16)
         );
  OR2_X1 cor_maj_113_U6 ( .A1(cor_maj_113_n20), .A2(cor_maj_113_n19), .ZN(
        cor_maj_113_n24) );
  NAND2_X1 cor_maj_113_U5 ( .A1(cor_maj_113_n24), .A2(cor_maj_113_n23), .ZN(
        cor_maj_113_n25) );
  NAND2_X1 cor_maj_113_U4 ( .A1(cor_maj_113_n20), .A2(cor_maj_113_n19), .ZN(
        cor_maj_113_n26) );
  NAND2_X1 cor_maj_113_U3 ( .A1(cor_maj_113_n26), .A2(cor_maj_113_n25), .ZN(
        cor_maj_113_port_o) );
  XOR2_X1 cor_maj_113_U2 ( .A(cor_maj_113_n22), .B(cor_maj_113_n21), .Z(
        cor_maj_113_n23) );
  NAND2_X1 cor_maj_114_U15 ( .A1(v_1_3_1[3]), .A2(v_1_3_1[4]), .ZN(
        cor_maj_114_n18) );
  NAND2_X1 cor_maj_114_U14 ( .A1(cor_maj_114_n21), .A2(cor_maj_114_n22), .ZN(
        cor_maj_114_n17) );
  NAND2_X1 cor_maj_114_U13 ( .A1(cor_maj_114_n18), .A2(cor_maj_114_n17), .ZN(
        cor_maj_114_n19) );
  NAND2_X1 cor_maj_114_U12 ( .A1(v_1_3_1[2]), .A2(cor_maj_114_n16), .ZN(
        cor_maj_114_n14) );
  NAND2_X1 cor_maj_114_U11 ( .A1(v_1_3_1[0]), .A2(v_1_3_1[1]), .ZN(
        cor_maj_114_n15) );
  NAND2_X1 cor_maj_114_U10 ( .A1(cor_maj_114_n15), .A2(cor_maj_114_n14), .ZN(
        cor_maj_114_n20) );
  XOR2_X1 cor_maj_114_U9 ( .A(v_1_3_1[3]), .B(v_1_3_1[4]), .Z(cor_maj_114_n22)
         );
  XOR2_X1 cor_maj_114_U8 ( .A(v_1_3_1[2]), .B(cor_maj_114_n16), .Z(
        cor_maj_114_n21) );
  XOR2_X1 cor_maj_114_U7 ( .A(v_1_3_1[0]), .B(v_1_3_1[1]), .Z(cor_maj_114_n16)
         );
  OR2_X1 cor_maj_114_U6 ( .A1(cor_maj_114_n20), .A2(cor_maj_114_n19), .ZN(
        cor_maj_114_n24) );
  NAND2_X1 cor_maj_114_U5 ( .A1(cor_maj_114_n24), .A2(cor_maj_114_n23), .ZN(
        cor_maj_114_n25) );
  NAND2_X1 cor_maj_114_U4 ( .A1(cor_maj_114_n20), .A2(cor_maj_114_n19), .ZN(
        cor_maj_114_n26) );
  NAND2_X1 cor_maj_114_U3 ( .A1(cor_maj_114_n26), .A2(cor_maj_114_n25), .ZN(
        cor_maj_114_port_o) );
  XOR2_X1 cor_maj_114_U2 ( .A(cor_maj_114_n22), .B(cor_maj_114_n21), .Z(
        cor_maj_114_n23) );
  NAND2_X1 cor_maj_115_U15 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_115_n18) );
  NAND2_X1 cor_maj_115_U14 ( .A1(cor_maj_115_n21), .A2(cor_maj_115_n22), .ZN(
        cor_maj_115_n17) );
  NAND2_X1 cor_maj_115_U13 ( .A1(cor_maj_115_n18), .A2(cor_maj_115_n17), .ZN(
        cor_maj_115_n19) );
  NAND2_X1 cor_maj_115_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_115_n16), .ZN(
        cor_maj_115_n14) );
  NAND2_X1 cor_maj_115_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_115_n15) );
  NAND2_X1 cor_maj_115_U10 ( .A1(cor_maj_115_n15), .A2(cor_maj_115_n14), .ZN(
        cor_maj_115_n20) );
  XOR2_X1 cor_maj_115_U9 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_115_n22)
         );
  XOR2_X1 cor_maj_115_U8 ( .A(v_1_3_2[2]), .B(cor_maj_115_n16), .Z(
        cor_maj_115_n21) );
  XOR2_X1 cor_maj_115_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_115_n16)
         );
  OR2_X1 cor_maj_115_U6 ( .A1(cor_maj_115_n20), .A2(cor_maj_115_n19), .ZN(
        cor_maj_115_n24) );
  NAND2_X1 cor_maj_115_U5 ( .A1(cor_maj_115_n24), .A2(cor_maj_115_n23), .ZN(
        cor_maj_115_n25) );
  NAND2_X1 cor_maj_115_U4 ( .A1(cor_maj_115_n20), .A2(cor_maj_115_n19), .ZN(
        cor_maj_115_n26) );
  NAND2_X1 cor_maj_115_U3 ( .A1(cor_maj_115_n26), .A2(cor_maj_115_n25), .ZN(
        cor_maj_115_port_o) );
  XOR2_X1 cor_maj_115_U2 ( .A(cor_maj_115_n22), .B(cor_maj_115_n21), .Z(
        cor_maj_115_n23) );
  NAND2_X1 cor_maj_116_U15 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_116_n18) );
  NAND2_X1 cor_maj_116_U14 ( .A1(cor_maj_116_n21), .A2(cor_maj_116_n22), .ZN(
        cor_maj_116_n17) );
  NAND2_X1 cor_maj_116_U13 ( .A1(cor_maj_116_n18), .A2(cor_maj_116_n17), .ZN(
        cor_maj_116_n19) );
  NAND2_X1 cor_maj_116_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_116_n16), .ZN(
        cor_maj_116_n14) );
  NAND2_X1 cor_maj_116_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_116_n15) );
  NAND2_X1 cor_maj_116_U10 ( .A1(cor_maj_116_n15), .A2(cor_maj_116_n14), .ZN(
        cor_maj_116_n20) );
  XOR2_X1 cor_maj_116_U9 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_116_n22)
         );
  XOR2_X1 cor_maj_116_U8 ( .A(v_1_3_2[2]), .B(cor_maj_116_n16), .Z(
        cor_maj_116_n21) );
  XOR2_X1 cor_maj_116_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_116_n16)
         );
  OR2_X1 cor_maj_116_U6 ( .A1(cor_maj_116_n20), .A2(cor_maj_116_n19), .ZN(
        cor_maj_116_n24) );
  NAND2_X1 cor_maj_116_U5 ( .A1(cor_maj_116_n24), .A2(cor_maj_116_n23), .ZN(
        cor_maj_116_n25) );
  NAND2_X1 cor_maj_116_U4 ( .A1(cor_maj_116_n20), .A2(cor_maj_116_n19), .ZN(
        cor_maj_116_n26) );
  NAND2_X1 cor_maj_116_U3 ( .A1(cor_maj_116_n26), .A2(cor_maj_116_n25), .ZN(
        cor_maj_116_port_o) );
  XOR2_X1 cor_maj_116_U2 ( .A(cor_maj_116_n22), .B(cor_maj_116_n21), .Z(
        cor_maj_116_n23) );
  NAND2_X1 cor_maj_117_U15 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_117_n18) );
  NAND2_X1 cor_maj_117_U14 ( .A1(cor_maj_117_n21), .A2(cor_maj_117_n22), .ZN(
        cor_maj_117_n17) );
  NAND2_X1 cor_maj_117_U13 ( .A1(cor_maj_117_n18), .A2(cor_maj_117_n17), .ZN(
        cor_maj_117_n19) );
  NAND2_X1 cor_maj_117_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_117_n16), .ZN(
        cor_maj_117_n14) );
  NAND2_X1 cor_maj_117_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_117_n15) );
  NAND2_X1 cor_maj_117_U10 ( .A1(cor_maj_117_n15), .A2(cor_maj_117_n14), .ZN(
        cor_maj_117_n20) );
  XOR2_X1 cor_maj_117_U9 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_117_n22)
         );
  XOR2_X1 cor_maj_117_U8 ( .A(v_1_3_2[2]), .B(cor_maj_117_n16), .Z(
        cor_maj_117_n21) );
  XOR2_X1 cor_maj_117_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_117_n16)
         );
  OR2_X1 cor_maj_117_U6 ( .A1(cor_maj_117_n20), .A2(cor_maj_117_n19), .ZN(
        cor_maj_117_n24) );
  NAND2_X1 cor_maj_117_U5 ( .A1(cor_maj_117_n24), .A2(cor_maj_117_n23), .ZN(
        cor_maj_117_n25) );
  NAND2_X1 cor_maj_117_U4 ( .A1(cor_maj_117_n20), .A2(cor_maj_117_n19), .ZN(
        cor_maj_117_n26) );
  NAND2_X1 cor_maj_117_U3 ( .A1(cor_maj_117_n26), .A2(cor_maj_117_n25), .ZN(
        cor_maj_117_port_o) );
  XOR2_X1 cor_maj_117_U2 ( .A(cor_maj_117_n22), .B(cor_maj_117_n21), .Z(
        cor_maj_117_n23) );
  NAND2_X1 cor_maj_118_U15 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_118_n18) );
  NAND2_X1 cor_maj_118_U14 ( .A1(cor_maj_118_n21), .A2(cor_maj_118_n22), .ZN(
        cor_maj_118_n17) );
  NAND2_X1 cor_maj_118_U13 ( .A1(cor_maj_118_n18), .A2(cor_maj_118_n17), .ZN(
        cor_maj_118_n19) );
  NAND2_X1 cor_maj_118_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_118_n16), .ZN(
        cor_maj_118_n14) );
  NAND2_X1 cor_maj_118_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_118_n15) );
  NAND2_X1 cor_maj_118_U10 ( .A1(cor_maj_118_n15), .A2(cor_maj_118_n14), .ZN(
        cor_maj_118_n20) );
  XOR2_X1 cor_maj_118_U9 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_118_n22)
         );
  XOR2_X1 cor_maj_118_U8 ( .A(v_1_3_2[2]), .B(cor_maj_118_n16), .Z(
        cor_maj_118_n21) );
  XOR2_X1 cor_maj_118_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_118_n16)
         );
  OR2_X1 cor_maj_118_U6 ( .A1(cor_maj_118_n20), .A2(cor_maj_118_n19), .ZN(
        cor_maj_118_n24) );
  NAND2_X1 cor_maj_118_U5 ( .A1(cor_maj_118_n24), .A2(cor_maj_118_n23), .ZN(
        cor_maj_118_n25) );
  NAND2_X1 cor_maj_118_U4 ( .A1(cor_maj_118_n20), .A2(cor_maj_118_n19), .ZN(
        cor_maj_118_n26) );
  NAND2_X1 cor_maj_118_U3 ( .A1(cor_maj_118_n26), .A2(cor_maj_118_n25), .ZN(
        cor_maj_118_port_o) );
  XOR2_X1 cor_maj_118_U2 ( .A(cor_maj_118_n22), .B(cor_maj_118_n21), .Z(
        cor_maj_118_n23) );
  NAND2_X1 cor_maj_119_U15 ( .A1(v_1_3_2[3]), .A2(v_1_3_2[4]), .ZN(
        cor_maj_119_n18) );
  NAND2_X1 cor_maj_119_U14 ( .A1(cor_maj_119_n21), .A2(cor_maj_119_n22), .ZN(
        cor_maj_119_n17) );
  NAND2_X1 cor_maj_119_U13 ( .A1(cor_maj_119_n18), .A2(cor_maj_119_n17), .ZN(
        cor_maj_119_n19) );
  NAND2_X1 cor_maj_119_U12 ( .A1(v_1_3_2[2]), .A2(cor_maj_119_n16), .ZN(
        cor_maj_119_n14) );
  NAND2_X1 cor_maj_119_U11 ( .A1(v_1_3_2[0]), .A2(v_1_3_2[1]), .ZN(
        cor_maj_119_n15) );
  NAND2_X1 cor_maj_119_U10 ( .A1(cor_maj_119_n15), .A2(cor_maj_119_n14), .ZN(
        cor_maj_119_n20) );
  XOR2_X1 cor_maj_119_U9 ( .A(v_1_3_2[3]), .B(v_1_3_2[4]), .Z(cor_maj_119_n22)
         );
  XOR2_X1 cor_maj_119_U8 ( .A(v_1_3_2[2]), .B(cor_maj_119_n16), .Z(
        cor_maj_119_n21) );
  XOR2_X1 cor_maj_119_U7 ( .A(v_1_3_2[0]), .B(v_1_3_2[1]), .Z(cor_maj_119_n16)
         );
  OR2_X1 cor_maj_119_U6 ( .A1(cor_maj_119_n20), .A2(cor_maj_119_n19), .ZN(
        cor_maj_119_n24) );
  NAND2_X1 cor_maj_119_U5 ( .A1(cor_maj_119_n24), .A2(cor_maj_119_n23), .ZN(
        cor_maj_119_n25) );
  NAND2_X1 cor_maj_119_U4 ( .A1(cor_maj_119_n20), .A2(cor_maj_119_n19), .ZN(
        cor_maj_119_n26) );
  NAND2_X1 cor_maj_119_U3 ( .A1(cor_maj_119_n26), .A2(cor_maj_119_n25), .ZN(
        cor_maj_119_port_o) );
  XOR2_X1 cor_maj_119_U2 ( .A(cor_maj_119_n22), .B(cor_maj_119_n21), .Z(
        cor_maj_119_n23) );
  XOR2_X1 simpleXor_60_U1 ( .A(n_zz_io_c_0_4[1]), .B(u_0_1[0]), .Z(
        simpleXor_60_port_z) );
  XOR2_X1 simpleXor_61_U1 ( .A(n_zz_io_c_0_4[2]), .B(u_0_2[0]), .Z(
        simpleXor_61_port_z) );
  XOR2_X1 simpleXor_62_U1 ( .A(n_zz_io_c_0_4[3]), .B(u_0_3[0]), .Z(
        simpleXor_62_port_z) );
  XOR2_X1 simpleXor_63_U1 ( .A(n_zz_io_c_1_4[1]), .B(u_1_0[0]), .Z(
        simpleXor_63_port_z) );
  XOR2_X1 simpleXor_64_U1 ( .A(n_zz_io_c_1_4[2]), .B(u_1_2[0]), .Z(
        simpleXor_64_port_z) );
  XOR2_X1 simpleXor_65_U1 ( .A(n_zz_io_c_1_4[3]), .B(u_1_3[0]), .Z(
        simpleXor_65_port_z) );
  XOR2_X1 simpleXor_66_U1 ( .A(n_zz_io_c_2_4[1]), .B(u_2_0[0]), .Z(
        simpleXor_66_port_z) );
  XOR2_X1 simpleXor_67_U1 ( .A(n_zz_io_c_2_4[2]), .B(u_2_1[0]), .Z(
        simpleXor_67_port_z) );
  XOR2_X1 simpleXor_68_U1 ( .A(n_zz_io_c_2_4[3]), .B(u_2_3[0]), .Z(
        simpleXor_68_port_z) );
  XOR2_X1 simpleXor_69_U1 ( .A(n_zz_io_c_3_4[1]), .B(u_3_0[0]), .Z(
        simpleXor_69_port_z) );
  XOR2_X1 simpleXor_70_U1 ( .A(n_zz_io_c_3_4[2]), .B(u_3_1[0]), .Z(
        simpleXor_70_port_z) );
  XOR2_X1 simpleXor_71_U1 ( .A(n_zz_io_c_3_4[3]), .B(u_3_2[0]), .Z(
        simpleXor_71_port_z) );
  XOR2_X1 simpleXor_72_U1 ( .A(n_zz_io_c_0_9[1]), .B(u_0_1[1]), .Z(
        simpleXor_72_port_z) );
  XOR2_X1 simpleXor_73_U1 ( .A(n_zz_io_c_0_9[2]), .B(u_0_2[1]), .Z(
        simpleXor_73_port_z) );
  XOR2_X1 simpleXor_74_U1 ( .A(n_zz_io_c_0_9[3]), .B(u_0_3[1]), .Z(
        simpleXor_74_port_z) );
  XOR2_X1 simpleXor_75_U1 ( .A(n_zz_io_c_1_9[1]), .B(u_1_0[1]), .Z(
        simpleXor_75_port_z) );
  XOR2_X1 simpleXor_76_U1 ( .A(n_zz_io_c_1_9[2]), .B(u_1_2[1]), .Z(
        simpleXor_76_port_z) );
  XOR2_X1 simpleXor_77_U1 ( .A(n_zz_io_c_1_9[3]), .B(u_1_3[1]), .Z(
        simpleXor_77_port_z) );
  XOR2_X1 simpleXor_78_U1 ( .A(n_zz_io_c_2_9[1]), .B(u_2_0[1]), .Z(
        simpleXor_78_port_z) );
  XOR2_X1 simpleXor_79_U1 ( .A(n_zz_io_c_2_9[2]), .B(u_2_1[1]), .Z(
        simpleXor_79_port_z) );
  XOR2_X1 simpleXor_80_U1 ( .A(n_zz_io_c_2_9[3]), .B(u_2_3[1]), .Z(
        simpleXor_80_port_z) );
  XOR2_X1 simpleXor_81_U1 ( .A(n_zz_io_c_3_9[1]), .B(u_3_0[1]), .Z(
        simpleXor_81_port_z) );
  XOR2_X1 simpleXor_82_U1 ( .A(n_zz_io_c_3_9[2]), .B(u_3_1[1]), .Z(
        simpleXor_82_port_z) );
  XOR2_X1 simpleXor_83_U1 ( .A(n_zz_io_c_3_9[3]), .B(u_3_2[1]), .Z(
        simpleXor_83_port_z) );
  XOR2_X1 simpleXor_84_U1 ( .A(n_zz_io_c_0_14[1]), .B(u_0_1[2]), .Z(
        simpleXor_84_port_z) );
  XOR2_X1 simpleXor_85_U1 ( .A(n_zz_io_c_0_14[2]), .B(u_0_2[2]), .Z(
        simpleXor_85_port_z) );
  XOR2_X1 simpleXor_86_U1 ( .A(n_zz_io_c_0_14[3]), .B(u_0_3[2]), .Z(
        simpleXor_86_port_z) );
  XOR2_X1 simpleXor_87_U1 ( .A(n_zz_io_c_1_14[1]), .B(u_1_0[2]), .Z(
        simpleXor_87_port_z) );
  XOR2_X1 simpleXor_88_U1 ( .A(n_zz_io_c_1_14[2]), .B(u_1_2[2]), .Z(
        simpleXor_88_port_z) );
  XOR2_X1 simpleXor_89_U1 ( .A(n_zz_io_c_1_14[3]), .B(u_1_3[2]), .Z(
        simpleXor_89_port_z) );
  XOR2_X1 simpleXor_90_U1 ( .A(n_zz_io_c_2_14[1]), .B(u_2_0[2]), .Z(
        simpleXor_90_port_z) );
  XOR2_X1 simpleXor_91_U1 ( .A(n_zz_io_c_2_14[2]), .B(u_2_1[2]), .Z(
        simpleXor_91_port_z) );
  XOR2_X1 simpleXor_92_U1 ( .A(n_zz_io_c_2_14[3]), .B(u_2_3[2]), .Z(
        simpleXor_92_port_z) );
  XOR2_X1 simpleXor_93_U1 ( .A(n_zz_io_c_3_14[1]), .B(u_3_0[2]), .Z(
        simpleXor_93_port_z) );
  XOR2_X1 simpleXor_94_U1 ( .A(n_zz_io_c_3_14[2]), .B(u_3_1[2]), .Z(
        simpleXor_94_port_z) );
  XOR2_X1 simpleXor_95_U1 ( .A(n_zz_io_c_3_14[3]), .B(u_3_2[2]), .Z(
        simpleXor_95_port_z) );
  XOR2_X1 simpleXor_96_U1 ( .A(n_zz_io_c_0_19[1]), .B(u_0_1[3]), .Z(
        simpleXor_96_port_z) );
  XOR2_X1 simpleXor_97_U1 ( .A(n_zz_io_c_0_19[2]), .B(u_0_2[3]), .Z(
        simpleXor_97_port_z) );
  XOR2_X1 simpleXor_98_U1 ( .A(n_zz_io_c_0_19[3]), .B(u_0_3[3]), .Z(
        simpleXor_98_port_z) );
  XOR2_X1 simpleXor_99_U1 ( .A(n_zz_io_c_1_19[1]), .B(u_1_0[3]), .Z(
        simpleXor_99_port_z) );
  XOR2_X1 simpleXor_100_U1 ( .A(n_zz_io_c_1_19[2]), .B(u_1_2[3]), .Z(
        simpleXor_100_port_z) );
  XOR2_X1 simpleXor_101_U1 ( .A(n_zz_io_c_1_19[3]), .B(u_1_3[3]), .Z(
        simpleXor_101_port_z) );
  XOR2_X1 simpleXor_102_U1 ( .A(n_zz_io_c_2_19[1]), .B(u_2_0[3]), .Z(
        simpleXor_102_port_z) );
  XOR2_X1 simpleXor_103_U1 ( .A(n_zz_io_c_2_19[2]), .B(u_2_1[3]), .Z(
        simpleXor_103_port_z) );
  XOR2_X1 simpleXor_104_U1 ( .A(n_zz_io_c_2_19[3]), .B(u_2_3[3]), .Z(
        simpleXor_104_port_z) );
  XOR2_X1 simpleXor_105_U1 ( .A(n_zz_io_c_3_19[1]), .B(u_3_0[3]), .Z(
        simpleXor_105_port_z) );
  XOR2_X1 simpleXor_106_U1 ( .A(n_zz_io_c_3_19[2]), .B(u_3_1[3]), .Z(
        simpleXor_106_port_z) );
  XOR2_X1 simpleXor_107_U1 ( .A(n_zz_io_c_3_19[3]), .B(u_3_2[3]), .Z(
        simpleXor_107_port_z) );
  XOR2_X1 simpleXor_108_U1 ( .A(n_zz_io_c_0_24[1]), .B(u_0_1[4]), .Z(
        simpleXor_108_port_z) );
  XOR2_X1 simpleXor_109_U1 ( .A(n_zz_io_c_0_24[2]), .B(u_0_2[4]), .Z(
        simpleXor_109_port_z) );
  XOR2_X1 simpleXor_110_U1 ( .A(n_zz_io_c_0_24[3]), .B(u_0_3[4]), .Z(
        simpleXor_110_port_z) );
  XOR2_X1 simpleXor_111_U1 ( .A(n_zz_io_c_1_24[1]), .B(u_1_0[4]), .Z(
        simpleXor_111_port_z) );
  XOR2_X1 simpleXor_112_U1 ( .A(n_zz_io_c_1_24[2]), .B(u_1_2[4]), .Z(
        simpleXor_112_port_z) );
  XOR2_X1 simpleXor_113_U1 ( .A(n_zz_io_c_1_24[3]), .B(u_1_3[4]), .Z(
        simpleXor_113_port_z) );
  XOR2_X1 simpleXor_114_U1 ( .A(n_zz_io_c_2_24[1]), .B(u_2_0[4]), .Z(
        simpleXor_114_port_z) );
  XOR2_X1 simpleXor_115_U1 ( .A(n_zz_io_c_2_24[2]), .B(u_2_1[4]), .Z(
        simpleXor_115_port_z) );
  XOR2_X1 simpleXor_116_U1 ( .A(n_zz_io_c_2_24[3]), .B(u_2_3[4]), .Z(
        simpleXor_116_port_z) );
  XOR2_X1 simpleXor_117_U1 ( .A(n_zz_io_c_3_24[1]), .B(u_3_0[4]), .Z(
        simpleXor_117_port_z) );
  XOR2_X1 simpleXor_118_U1 ( .A(n_zz_io_c_3_24[2]), .B(u_3_1[4]), .Z(
        simpleXor_118_port_z) );
  XOR2_X1 simpleXor_119_U1 ( .A(n_zz_io_c_3_24[3]), .B(u_3_2[4]), .Z(
        simpleXor_119_port_z) );
endmodule

