
module And_gate ( clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, 
        clock_6, reset_0, reset_1, reset_2, reset_3, reset_4, reset_5, reset_6, 
        io_i0_s0_d0, io_i0_s0_d1, io_i0_s0_d2, io_i0_s0_d3, io_i0_s0_d4, 
        io_i0_s0_d5, io_i0_s0_d6, io_i0_s1_d0, io_i0_s1_d1, io_i0_s1_d2, 
        io_i0_s1_d3, io_i0_s1_d4, io_i0_s1_d5, io_i0_s1_d6, io_i0_s2_d0, 
        io_i0_s2_d1, io_i0_s2_d2, io_i0_s2_d3, io_i0_s2_d4, io_i0_s2_d5, 
        io_i0_s2_d6, io_i0_s3_d0, io_i0_s3_d1, io_i0_s3_d2, io_i0_s3_d3, 
        io_i0_s3_d4, io_i0_s3_d5, io_i0_s3_d6, io_i1_s0_d0, io_i1_s0_d1, 
        io_i1_s0_d2, io_i1_s0_d3, io_i1_s0_d4, io_i1_s0_d5, io_i1_s0_d6, 
        io_i1_s1_d0, io_i1_s1_d1, io_i1_s1_d2, io_i1_s1_d3, io_i1_s1_d4, 
        io_i1_s1_d5, io_i1_s1_d6, io_i1_s2_d0, io_i1_s2_d1, io_i1_s2_d2, 
        io_i1_s2_d3, io_i1_s2_d4, io_i1_s2_d5, io_i1_s2_d6, io_i1_s3_d0, 
        io_i1_s3_d1, io_i1_s3_d2, io_i1_s3_d3, io_i1_s3_d4, io_i1_s3_d5, 
        io_i1_s3_d6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, 
        p_rand_5, p_rand_6, p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11, 
        io_o0_s0_d0, io_o0_s0_d1, io_o0_s0_d2, io_o0_s0_d3, io_o0_s0_d4, 
        io_o0_s0_d5, io_o0_s0_d6, io_o0_s1_d0, io_o0_s1_d1, io_o0_s1_d2, 
        io_o0_s1_d3, io_o0_s1_d4, io_o0_s1_d5, io_o0_s1_d6, io_o0_s2_d0, 
        io_o0_s2_d1, io_o0_s2_d2, io_o0_s2_d3, io_o0_s2_d4, io_o0_s2_d5, 
        io_o0_s2_d6, io_o0_s3_d0, io_o0_s3_d1, io_o0_s3_d2, io_o0_s3_d3, 
        io_o0_s3_d4, io_o0_s3_d5, io_o0_s3_d6 );
  input clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, clock_6, reset_0,
         reset_1, reset_2, reset_3, reset_4, reset_5, reset_6, io_i0_s0_d0,
         io_i0_s0_d1, io_i0_s0_d2, io_i0_s0_d3, io_i0_s0_d4, io_i0_s0_d5,
         io_i0_s0_d6, io_i0_s1_d0, io_i0_s1_d1, io_i0_s1_d2, io_i0_s1_d3,
         io_i0_s1_d4, io_i0_s1_d5, io_i0_s1_d6, io_i0_s2_d0, io_i0_s2_d1,
         io_i0_s2_d2, io_i0_s2_d3, io_i0_s2_d4, io_i0_s2_d5, io_i0_s2_d6,
         io_i0_s3_d0, io_i0_s3_d1, io_i0_s3_d2, io_i0_s3_d3, io_i0_s3_d4,
         io_i0_s3_d5, io_i0_s3_d6, io_i1_s0_d0, io_i1_s0_d1, io_i1_s0_d2,
         io_i1_s0_d3, io_i1_s0_d4, io_i1_s0_d5, io_i1_s0_d6, io_i1_s1_d0,
         io_i1_s1_d1, io_i1_s1_d2, io_i1_s1_d3, io_i1_s1_d4, io_i1_s1_d5,
         io_i1_s1_d6, io_i1_s2_d0, io_i1_s2_d1, io_i1_s2_d2, io_i1_s2_d3,
         io_i1_s2_d4, io_i1_s2_d5, io_i1_s2_d6, io_i1_s3_d0, io_i1_s3_d1,
         io_i1_s3_d2, io_i1_s3_d3, io_i1_s3_d4, io_i1_s3_d5, io_i1_s3_d6,
         p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4, p_rand_5, p_rand_6,
         p_rand_7, p_rand_8, p_rand_9, p_rand_10, p_rand_11;
  output io_o0_s0_d0, io_o0_s0_d1, io_o0_s0_d2, io_o0_s0_d3, io_o0_s0_d4,
         io_o0_s0_d5, io_o0_s0_d6, io_o0_s1_d0, io_o0_s1_d1, io_o0_s1_d2,
         io_o0_s1_d3, io_o0_s1_d4, io_o0_s1_d5, io_o0_s1_d6, io_o0_s2_d0,
         io_o0_s2_d1, io_o0_s2_d2, io_o0_s2_d3, io_o0_s2_d4, io_o0_s2_d5,
         io_o0_s2_d6, io_o0_s3_d0, io_o0_s3_d1, io_o0_s3_d2, io_o0_s3_d3,
         io_o0_s3_d4, io_o0_s3_d5, io_o0_s3_d6;
  wire   n_xor_module_1_res, n_xor_module_2_res, n_xor_module_3_res,
         n_xor_module_4_res, n_xor_module_5_res, n_xor_module_6_res,
         n_xor_module_7_res, n_xor_module_8_res, n_xor_module_9_res,
         n_xor_module_10_res, n_xor_module_11_res, n_xor_module_12_res,
         n_xor_module_13_res, n_xor_module_14_res, n_xor_module_15_res,
         n_xor_module_16_res, n_xor_module_17_res, n_xor_module_18_res,
         n_xor_module_19_res, n_xor_module_20_res, n_xor_module_21_res,
         n_xor_module_22_res, n_xor_module_23_res, n_xor_module_24_res,
         n_xor_module_25_res, n_xor_module_26_res, n_xor_module_27_res,
         n_xor_module_28_res, n_xor_module_29_res, n_xor_module_30_res,
         n_xor_module_31_res, n_xor_module_32_res, n_xor_module_33_res,
         n_xor_module_34_res, n_xor_module_35_res, n_xor_module_36_res,
         n_xor_module_37_res, n_xor_module_38_res, n_xor_module_39_res,
         n_xor_module_40_res, n_xor_module_41_res, n_xor_module_42_res,
         n_xor_module_43_res, n_xor_module_44_res, n_xor_module_45_res,
         n_xor_module_46_res, n_xor_module_47_res, n_xor_module_48_res,
         n_xor_module_49_res, n_xor_module_50_res, n_xor_module_51_res,
         n_xor_module_52_res, n_xor_module_53_res, n_xor_module_54_res,
         n_xor_module_55_res, n_xor_module_56_res, n_xor_module_57_res,
         n_xor_module_58_res, n_xor_module_59_res, n_xor_module_60_res,
         n_xor_module_61_res, n_xor_module_62_res, n_xor_module_63_res,
         n_xor_module_64_res, n_xor_module_65_res, n_xor_module_66_res,
         n_xor_module_67_res, n_xor_module_68_res, n_xor_module_69_res,
         n_xor_module_70_res, n_xor_module_71_res, n_xor_module_72_res,
         n_xor_module_73_res, n_xor_module_74_res, n_xor_module_75_res,
         n_xor_module_76_res, n_xor_module_77_res, n_xor_module_78_res,
         n_xor_module_79_res, n_xor_module_80_res, n_xor_module_81_res,
         n_xor_module_82_res, n_xor_module_83_res, n_xor_module_84_res,
         n_majority7_module_0_res, n_reg_module_1_res,
         n_majority7_module_1_res, n_reg_module_2_res,
         n_majority7_module_2_res, n_reg_module_3_res,
         n_majority7_module_3_res, n_reg_module_4_res,
         n_majority7_module_4_res, n_reg_module_5_res,
         n_majority7_module_5_res, n_reg_module_6_res,
         n_majority7_module_6_res, n_reg_module_7_res,
         n_majority7_module_7_res, n_reg_module_8_res,
         n_majority7_module_8_res, n_reg_module_9_res,
         n_majority7_module_9_res, n_reg_module_10_res,
         n_majority7_module_10_res, n_reg_module_11_res,
         n_majority7_module_11_res, n_reg_module_12_res,
         n_majority7_module_12_res, n_reg_module_13_res,
         n_majority7_module_13_res, n_reg_module_14_res,
         n_majority7_module_14_res, n_reg_module_15_res,
         n_majority7_module_15_res, n_reg_module_16_res,
         n_majority7_module_16_res, n_reg_module_17_res,
         n_majority7_module_17_res, n_reg_module_18_res,
         n_majority7_module_18_res, n_reg_module_19_res,
         n_majority7_module_19_res, n_reg_module_20_res,
         n_majority7_module_20_res, n_reg_module_21_res,
         n_majority7_module_21_res, n_reg_module_22_res,
         n_majority7_module_22_res, n_reg_module_23_res,
         n_majority7_module_23_res, n_reg_module_24_res,
         n_majority7_module_24_res, n_reg_module_25_res,
         n_majority7_module_25_res, n_reg_module_26_res,
         n_majority7_module_26_res, n_reg_module_27_res,
         n_majority7_module_27_res, n_reg_module_28_res, n_and_module_1_res,
         n_and_module_2_res, n_xor_module_85_res, n_and_module_3_res,
         n_xor_module_86_res, n_and_module_4_res, n_xor_module_87_res,
         n_and_module_5_res, n_xor_module_88_res, n_and_module_6_res,
         n_and_module_7_res, n_xor_module_89_res, n_and_module_8_res,
         n_xor_module_90_res, n_and_module_9_res, n_xor_module_91_res,
         n_and_module_10_res, n_xor_module_92_res, n_and_module_11_res,
         n_and_module_12_res, n_xor_module_93_res, n_and_module_13_res,
         n_xor_module_94_res, n_and_module_14_res, n_xor_module_95_res,
         n_and_module_15_res, n_xor_module_96_res, n_and_module_16_res,
         n_and_module_17_res, n_and_module_18_res, n_xor_module_97_res,
         n_and_module_19_res, n_xor_module_98_res, n_and_module_20_res,
         n_xor_module_99_res, n_and_module_21_res, n_xor_module_100_res,
         n_and_module_22_res, n_and_module_23_res, n_xor_module_101_res,
         n_and_module_24_res, n_xor_module_102_res, n_and_module_25_res,
         n_xor_module_103_res, n_and_module_26_res, n_xor_module_104_res,
         n_and_module_27_res, n_and_module_28_res, n_xor_module_105_res,
         n_and_module_29_res, n_xor_module_106_res, n_and_module_30_res,
         n_xor_module_107_res, n_and_module_31_res, n_xor_module_108_res,
         n_and_module_32_res, n_and_module_33_res, n_and_module_34_res,
         n_xor_module_109_res, n_and_module_35_res, n_xor_module_110_res,
         n_and_module_36_res, n_xor_module_111_res, n_and_module_37_res,
         n_xor_module_112_res, n_and_module_38_res, n_and_module_39_res,
         n_xor_module_113_res, n_and_module_40_res, n_xor_module_114_res,
         n_and_module_41_res, n_xor_module_115_res, n_and_module_42_res,
         n_xor_module_116_res, n_and_module_43_res, n_and_module_44_res,
         n_xor_module_117_res, n_and_module_45_res, n_xor_module_118_res,
         n_and_module_46_res, n_xor_module_119_res, n_and_module_47_res,
         n_xor_module_120_res, n_and_module_48_res, n_and_module_49_res,
         n_and_module_50_res, n_xor_module_121_res, n_and_module_51_res,
         n_xor_module_122_res, n_and_module_52_res, n_xor_module_123_res,
         n_and_module_53_res, n_xor_module_124_res, n_and_module_54_res,
         n_and_module_55_res, n_xor_module_125_res, n_and_module_56_res,
         n_xor_module_126_res, n_and_module_57_res, n_xor_module_127_res,
         n_and_module_58_res, n_xor_module_128_res, n_and_module_59_res,
         n_and_module_60_res, n_xor_module_129_res, n_and_module_61_res,
         n_xor_module_130_res, n_and_module_62_res, n_xor_module_131_res,
         n_and_module_63_res, n_xor_module_132_res, n_and_module_64_res,
         n_and_module_65_res, n_and_module_66_res, n_xor_module_133_res,
         n_and_module_67_res, n_xor_module_134_res, n_and_module_68_res,
         n_xor_module_135_res, n_and_module_69_res, n_xor_module_136_res,
         n_and_module_70_res, n_and_module_71_res, n_xor_module_137_res,
         n_and_module_72_res, n_xor_module_138_res, n_and_module_73_res,
         n_xor_module_139_res, n_and_module_74_res, n_xor_module_140_res,
         n_and_module_75_res, n_and_module_76_res, n_xor_module_141_res,
         n_and_module_77_res, n_xor_module_142_res, n_and_module_78_res,
         n_xor_module_143_res, n_and_module_79_res, n_xor_module_144_res,
         n_and_module_80_res, n_and_module_81_res, n_and_module_82_res,
         n_xor_module_145_res, n_and_module_83_res, n_xor_module_146_res,
         n_and_module_84_res, n_xor_module_147_res, n_and_module_85_res,
         n_xor_module_148_res, n_and_module_86_res, n_and_module_87_res,
         n_xor_module_149_res, n_and_module_88_res, n_xor_module_150_res,
         n_and_module_89_res, n_xor_module_151_res, n_and_module_90_res,
         n_xor_module_152_res, n_and_module_91_res, n_and_module_92_res,
         n_xor_module_153_res, n_and_module_93_res, n_xor_module_154_res,
         n_and_module_94_res, n_xor_module_155_res, n_and_module_95_res,
         n_xor_module_156_res, n_and_module_96_res, n_and_module_97_res,
         n_and_module_98_res, n_xor_module_157_res, n_and_module_99_res,
         n_xor_module_158_res, n_and_module_100_res, n_xor_module_159_res,
         n_and_module_101_res, n_xor_module_160_res, n_and_module_102_res,
         n_and_module_103_res, n_xor_module_161_res, n_and_module_104_res,
         n_xor_module_162_res, n_and_module_105_res, n_xor_module_163_res,
         n_and_module_106_res, n_xor_module_164_res, n_and_module_107_res,
         n_and_module_108_res, n_xor_module_165_res, n_and_module_109_res,
         n_xor_module_166_res, n_and_module_110_res, n_xor_module_167_res,
         n_and_module_111_res, n_xor_module_168_res, n_and_module_112_res,
         n_reg_module_29_res, n_majority7_module_28_res, n_reg_module_30_res,
         n_majority7_module_29_res, n_reg_module_31_res,
         n_majority7_module_30_res, n_reg_module_32_res,
         n_majority7_module_31_res, n_reg_module_33_res, n_reg_module_34_res,
         n_majority7_module_32_res, n_reg_module_35_res,
         n_majority7_module_33_res, n_reg_module_36_res,
         n_majority7_module_34_res, n_reg_module_37_res,
         n_majority7_module_35_res, n_reg_module_38_res, n_reg_module_39_res,
         n_majority7_module_36_res, n_reg_module_40_res,
         n_majority7_module_37_res, n_reg_module_41_res,
         n_majority7_module_38_res, n_reg_module_42_res,
         n_majority7_module_39_res, n_reg_module_43_res, n_reg_module_44_res,
         n_reg_module_45_res, n_majority7_module_40_res, n_reg_module_46_res,
         n_majority7_module_41_res, n_reg_module_47_res,
         n_majority7_module_42_res, n_reg_module_48_res,
         n_majority7_module_43_res, n_reg_module_49_res, n_reg_module_50_res,
         n_majority7_module_44_res, n_reg_module_51_res,
         n_majority7_module_45_res, n_reg_module_52_res,
         n_majority7_module_46_res, n_reg_module_53_res,
         n_majority7_module_47_res, n_reg_module_54_res, n_reg_module_55_res,
         n_majority7_module_48_res, n_reg_module_56_res,
         n_majority7_module_49_res, n_reg_module_57_res,
         n_majority7_module_50_res, n_reg_module_58_res,
         n_majority7_module_51_res, n_reg_module_59_res, n_reg_module_60_res,
         n_reg_module_61_res, n_majority7_module_52_res, n_reg_module_62_res,
         n_majority7_module_53_res, n_reg_module_63_res,
         n_majority7_module_54_res, n_reg_module_64_res,
         n_majority7_module_55_res, n_reg_module_65_res, n_reg_module_66_res,
         n_majority7_module_56_res, n_reg_module_67_res,
         n_majority7_module_57_res, n_reg_module_68_res,
         n_majority7_module_58_res, n_reg_module_69_res,
         n_majority7_module_59_res, n_reg_module_70_res, n_reg_module_71_res,
         n_majority7_module_60_res, n_reg_module_72_res,
         n_majority7_module_61_res, n_reg_module_73_res,
         n_majority7_module_62_res, n_reg_module_74_res,
         n_majority7_module_63_res, n_reg_module_75_res, n_reg_module_76_res,
         n_reg_module_77_res, n_majority7_module_64_res, n_reg_module_78_res,
         n_majority7_module_65_res, n_reg_module_79_res,
         n_majority7_module_66_res, n_reg_module_80_res,
         n_majority7_module_67_res, n_reg_module_81_res, n_reg_module_82_res,
         n_majority7_module_68_res, n_reg_module_83_res,
         n_majority7_module_69_res, n_reg_module_84_res,
         n_majority7_module_70_res, n_reg_module_85_res,
         n_majority7_module_71_res, n_reg_module_86_res, n_reg_module_87_res,
         n_majority7_module_72_res, n_reg_module_88_res,
         n_majority7_module_73_res, n_reg_module_89_res,
         n_majority7_module_74_res, n_reg_module_90_res,
         n_majority7_module_75_res, n_reg_module_91_res, n_reg_module_92_res,
         n_reg_module_93_res, n_majority7_module_76_res, n_reg_module_94_res,
         n_majority7_module_77_res, n_reg_module_95_res,
         n_majority7_module_78_res, n_reg_module_96_res,
         n_majority7_module_79_res, n_reg_module_97_res, n_reg_module_98_res,
         n_majority7_module_80_res, n_reg_module_99_res,
         n_majority7_module_81_res, n_reg_module_100_res,
         n_majority7_module_82_res, n_reg_module_101_res,
         n_majority7_module_83_res, n_reg_module_102_res, n_reg_module_103_res,
         n_majority7_module_84_res, n_reg_module_104_res,
         n_majority7_module_85_res, n_reg_module_105_res,
         n_majority7_module_86_res, n_reg_module_106_res,
         n_majority7_module_87_res, n_reg_module_107_res, n_reg_module_108_res,
         n_reg_module_109_res, n_majority7_module_88_res, n_reg_module_110_res,
         n_majority7_module_89_res, n_reg_module_111_res,
         n_majority7_module_90_res, n_reg_module_112_res,
         n_majority7_module_91_res, n_reg_module_113_res, n_reg_module_114_res,
         n_majority7_module_92_res, n_reg_module_115_res,
         n_majority7_module_93_res, n_reg_module_116_res,
         n_majority7_module_94_res, n_reg_module_117_res,
         n_majority7_module_95_res, n_reg_module_118_res, n_reg_module_119_res,
         n_majority7_module_96_res, n_reg_module_120_res,
         n_majority7_module_97_res, n_reg_module_121_res,
         n_majority7_module_98_res, n_reg_module_122_res,
         n_majority7_module_99_res, n_reg_module_123_res, n_reg_module_124_res,
         n_reg_module_125_res, n_majority7_module_100_res,
         n_reg_module_126_res, n_majority7_module_101_res,
         n_reg_module_127_res, n_majority7_module_102_res,
         n_reg_module_128_res, n_majority7_module_103_res,
         n_reg_module_129_res, n_reg_module_130_res,
         n_majority7_module_104_res, n_reg_module_131_res,
         n_majority7_module_105_res, n_reg_module_132_res,
         n_majority7_module_106_res, n_reg_module_133_res,
         n_majority7_module_107_res, n_reg_module_134_res,
         n_reg_module_135_res, n_majority7_module_108_res,
         n_reg_module_136_res, n_majority7_module_109_res,
         n_reg_module_137_res, n_majority7_module_110_res,
         n_reg_module_138_res, n_majority7_module_111_res,
         n_reg_module_139_res, n_reg_module_140_res, n_xor_module_169_res,
         n_xor_module_170_res, n_xor_module_172_res, n_xor_module_173_res,
         n_xor_module_175_res, n_xor_module_176_res, n_xor_module_178_res,
         n_xor_module_179_res, n_xor_module_181_res, n_xor_module_182_res,
         n_xor_module_184_res, n_xor_module_185_res, n_xor_module_187_res,
         n_xor_module_188_res, n_xor_module_190_res, n_xor_module_191_res,
         n_xor_module_193_res, n_xor_module_194_res, n_xor_module_196_res,
         n_xor_module_197_res, n_xor_module_199_res, n_xor_module_200_res,
         n_xor_module_202_res, n_xor_module_203_res, n_xor_module_205_res,
         n_xor_module_206_res, n_xor_module_208_res, n_xor_module_209_res,
         n_xor_module_211_res, n_xor_module_212_res, n_xor_module_214_res,
         n_xor_module_215_res, n_xor_module_217_res, n_xor_module_218_res,
         n_xor_module_220_res, n_xor_module_221_res, n_xor_module_223_res,
         n_xor_module_224_res, n_xor_module_226_res, n_xor_module_227_res,
         n_xor_module_229_res, n_xor_module_230_res, n_xor_module_232_res,
         n_xor_module_233_res, n_xor_module_235_res, n_xor_module_236_res,
         n_xor_module_238_res, n_xor_module_239_res, n_xor_module_241_res,
         n_xor_module_242_res, n_xor_module_244_res, n_xor_module_245_res,
         n_xor_module_247_res, n_xor_module_248_res, n_xor_module_250_res,
         n_xor_module_251_res, n_majority7_module_0__and_module_10_res,
         n_majority7_module_0__or_module_11_res,
         n_majority7_module_0__and_module_9_res,
         n_majority7_module_0__or_module_10_res,
         n_majority7_module_0__or_module_9_res,
         n_majority7_module_0__and_module_8_res,
         n_majority7_module_0__or_module_8_res,
         n_majority7_module_0__and_module_7_res,
         n_majority7_module_0__or_module_7_res,
         n_majority7_module_0__or_module_6_res,
         n_majority7_module_0__and_module_6_res,
         n_majority7_module_0__or_module_5_res,
         n_majority7_module_0__and_module_5_res,
         n_majority7_module_0__or_module_4_res,
         n_majority7_module_0__and_module_4_res,
         n_majority7_module_0__or_module_3_res,
         n_majority7_module_0__and_module_3_res,
         n_majority7_module_0__or_module_2_res,
         n_majority7_module_0__and_module_2_res,
         n_majority7_module_0__or_module_1_res,
         n_majority7_module_0__and_module_1_res,
         n_majority7_module_1__and_module_10_res,
         n_majority7_module_1__or_module_11_res,
         n_majority7_module_1__and_module_9_res,
         n_majority7_module_1__or_module_10_res,
         n_majority7_module_1__or_module_9_res,
         n_majority7_module_1__and_module_8_res,
         n_majority7_module_1__or_module_8_res,
         n_majority7_module_1__and_module_7_res,
         n_majority7_module_1__or_module_7_res,
         n_majority7_module_1__or_module_6_res,
         n_majority7_module_1__and_module_6_res,
         n_majority7_module_1__or_module_5_res,
         n_majority7_module_1__and_module_5_res,
         n_majority7_module_1__or_module_4_res,
         n_majority7_module_1__and_module_4_res,
         n_majority7_module_1__or_module_3_res,
         n_majority7_module_1__and_module_3_res,
         n_majority7_module_1__or_module_2_res,
         n_majority7_module_1__and_module_2_res,
         n_majority7_module_1__or_module_1_res,
         n_majority7_module_1__and_module_1_res,
         n_majority7_module_2__and_module_10_res,
         n_majority7_module_2__or_module_11_res,
         n_majority7_module_2__and_module_9_res,
         n_majority7_module_2__or_module_10_res,
         n_majority7_module_2__or_module_9_res,
         n_majority7_module_2__and_module_8_res,
         n_majority7_module_2__or_module_8_res,
         n_majority7_module_2__and_module_7_res,
         n_majority7_module_2__or_module_7_res,
         n_majority7_module_2__or_module_6_res,
         n_majority7_module_2__and_module_6_res,
         n_majority7_module_2__or_module_5_res,
         n_majority7_module_2__and_module_5_res,
         n_majority7_module_2__or_module_4_res,
         n_majority7_module_2__and_module_4_res,
         n_majority7_module_2__or_module_3_res,
         n_majority7_module_2__and_module_3_res,
         n_majority7_module_2__or_module_2_res,
         n_majority7_module_2__and_module_2_res,
         n_majority7_module_2__or_module_1_res,
         n_majority7_module_2__and_module_1_res,
         n_majority7_module_3__and_module_10_res,
         n_majority7_module_3__or_module_11_res,
         n_majority7_module_3__and_module_9_res,
         n_majority7_module_3__or_module_10_res,
         n_majority7_module_3__or_module_9_res,
         n_majority7_module_3__and_module_8_res,
         n_majority7_module_3__or_module_8_res,
         n_majority7_module_3__and_module_7_res,
         n_majority7_module_3__or_module_7_res,
         n_majority7_module_3__or_module_6_res,
         n_majority7_module_3__and_module_6_res,
         n_majority7_module_3__or_module_5_res,
         n_majority7_module_3__and_module_5_res,
         n_majority7_module_3__or_module_4_res,
         n_majority7_module_3__and_module_4_res,
         n_majority7_module_3__or_module_3_res,
         n_majority7_module_3__and_module_3_res,
         n_majority7_module_3__or_module_2_res,
         n_majority7_module_3__and_module_2_res,
         n_majority7_module_3__or_module_1_res,
         n_majority7_module_3__and_module_1_res,
         n_majority7_module_4__and_module_10_res,
         n_majority7_module_4__or_module_11_res,
         n_majority7_module_4__and_module_9_res,
         n_majority7_module_4__or_module_10_res,
         n_majority7_module_4__or_module_9_res,
         n_majority7_module_4__and_module_8_res,
         n_majority7_module_4__or_module_8_res,
         n_majority7_module_4__and_module_7_res,
         n_majority7_module_4__or_module_7_res,
         n_majority7_module_4__or_module_6_res,
         n_majority7_module_4__and_module_6_res,
         n_majority7_module_4__or_module_5_res,
         n_majority7_module_4__and_module_5_res,
         n_majority7_module_4__or_module_4_res,
         n_majority7_module_4__and_module_4_res,
         n_majority7_module_4__or_module_3_res,
         n_majority7_module_4__and_module_3_res,
         n_majority7_module_4__or_module_2_res,
         n_majority7_module_4__and_module_2_res,
         n_majority7_module_4__or_module_1_res,
         n_majority7_module_4__and_module_1_res,
         n_majority7_module_5__and_module_10_res,
         n_majority7_module_5__or_module_11_res,
         n_majority7_module_5__and_module_9_res,
         n_majority7_module_5__or_module_10_res,
         n_majority7_module_5__or_module_9_res,
         n_majority7_module_5__and_module_8_res,
         n_majority7_module_5__or_module_8_res,
         n_majority7_module_5__and_module_7_res,
         n_majority7_module_5__or_module_7_res,
         n_majority7_module_5__or_module_6_res,
         n_majority7_module_5__and_module_6_res,
         n_majority7_module_5__or_module_5_res,
         n_majority7_module_5__and_module_5_res,
         n_majority7_module_5__or_module_4_res,
         n_majority7_module_5__and_module_4_res,
         n_majority7_module_5__or_module_3_res,
         n_majority7_module_5__and_module_3_res,
         n_majority7_module_5__or_module_2_res,
         n_majority7_module_5__and_module_2_res,
         n_majority7_module_5__or_module_1_res,
         n_majority7_module_5__and_module_1_res,
         n_majority7_module_6__and_module_10_res,
         n_majority7_module_6__or_module_11_res,
         n_majority7_module_6__and_module_9_res,
         n_majority7_module_6__or_module_10_res,
         n_majority7_module_6__or_module_9_res,
         n_majority7_module_6__and_module_8_res,
         n_majority7_module_6__or_module_8_res,
         n_majority7_module_6__and_module_7_res,
         n_majority7_module_6__or_module_7_res,
         n_majority7_module_6__or_module_6_res,
         n_majority7_module_6__and_module_6_res,
         n_majority7_module_6__or_module_5_res,
         n_majority7_module_6__and_module_5_res,
         n_majority7_module_6__or_module_4_res,
         n_majority7_module_6__and_module_4_res,
         n_majority7_module_6__or_module_3_res,
         n_majority7_module_6__and_module_3_res,
         n_majority7_module_6__or_module_2_res,
         n_majority7_module_6__and_module_2_res,
         n_majority7_module_6__or_module_1_res,
         n_majority7_module_6__and_module_1_res,
         n_majority7_module_7__and_module_10_res,
         n_majority7_module_7__or_module_11_res,
         n_majority7_module_7__and_module_9_res,
         n_majority7_module_7__or_module_10_res,
         n_majority7_module_7__or_module_9_res,
         n_majority7_module_7__and_module_8_res,
         n_majority7_module_7__or_module_8_res,
         n_majority7_module_7__and_module_7_res,
         n_majority7_module_7__or_module_7_res,
         n_majority7_module_7__or_module_6_res,
         n_majority7_module_7__and_module_6_res,
         n_majority7_module_7__or_module_5_res,
         n_majority7_module_7__and_module_5_res,
         n_majority7_module_7__or_module_4_res,
         n_majority7_module_7__and_module_4_res,
         n_majority7_module_7__or_module_3_res,
         n_majority7_module_7__and_module_3_res,
         n_majority7_module_7__or_module_2_res,
         n_majority7_module_7__and_module_2_res,
         n_majority7_module_7__or_module_1_res,
         n_majority7_module_7__and_module_1_res,
         n_majority7_module_8__and_module_10_res,
         n_majority7_module_8__or_module_11_res,
         n_majority7_module_8__and_module_9_res,
         n_majority7_module_8__or_module_10_res,
         n_majority7_module_8__or_module_9_res,
         n_majority7_module_8__and_module_8_res,
         n_majority7_module_8__or_module_8_res,
         n_majority7_module_8__and_module_7_res,
         n_majority7_module_8__or_module_7_res,
         n_majority7_module_8__or_module_6_res,
         n_majority7_module_8__and_module_6_res,
         n_majority7_module_8__or_module_5_res,
         n_majority7_module_8__and_module_5_res,
         n_majority7_module_8__or_module_4_res,
         n_majority7_module_8__and_module_4_res,
         n_majority7_module_8__or_module_3_res,
         n_majority7_module_8__and_module_3_res,
         n_majority7_module_8__or_module_2_res,
         n_majority7_module_8__and_module_2_res,
         n_majority7_module_8__or_module_1_res,
         n_majority7_module_8__and_module_1_res,
         n_majority7_module_9__and_module_10_res,
         n_majority7_module_9__or_module_11_res,
         n_majority7_module_9__and_module_9_res,
         n_majority7_module_9__or_module_10_res,
         n_majority7_module_9__or_module_9_res,
         n_majority7_module_9__and_module_8_res,
         n_majority7_module_9__or_module_8_res,
         n_majority7_module_9__and_module_7_res,
         n_majority7_module_9__or_module_7_res,
         n_majority7_module_9__or_module_6_res,
         n_majority7_module_9__and_module_6_res,
         n_majority7_module_9__or_module_5_res,
         n_majority7_module_9__and_module_5_res,
         n_majority7_module_9__or_module_4_res,
         n_majority7_module_9__and_module_4_res,
         n_majority7_module_9__or_module_3_res,
         n_majority7_module_9__and_module_3_res,
         n_majority7_module_9__or_module_2_res,
         n_majority7_module_9__and_module_2_res,
         n_majority7_module_9__or_module_1_res,
         n_majority7_module_9__and_module_1_res,
         n_majority7_module_10__and_module_10_res,
         n_majority7_module_10__or_module_11_res,
         n_majority7_module_10__and_module_9_res,
         n_majority7_module_10__or_module_10_res,
         n_majority7_module_10__or_module_9_res,
         n_majority7_module_10__and_module_8_res,
         n_majority7_module_10__or_module_8_res,
         n_majority7_module_10__and_module_7_res,
         n_majority7_module_10__or_module_7_res,
         n_majority7_module_10__or_module_6_res,
         n_majority7_module_10__and_module_6_res,
         n_majority7_module_10__or_module_5_res,
         n_majority7_module_10__and_module_5_res,
         n_majority7_module_10__or_module_4_res,
         n_majority7_module_10__and_module_4_res,
         n_majority7_module_10__or_module_3_res,
         n_majority7_module_10__and_module_3_res,
         n_majority7_module_10__or_module_2_res,
         n_majority7_module_10__and_module_2_res,
         n_majority7_module_10__or_module_1_res,
         n_majority7_module_10__and_module_1_res,
         n_majority7_module_11__and_module_10_res,
         n_majority7_module_11__or_module_11_res,
         n_majority7_module_11__and_module_9_res,
         n_majority7_module_11__or_module_10_res,
         n_majority7_module_11__or_module_9_res,
         n_majority7_module_11__and_module_8_res,
         n_majority7_module_11__or_module_8_res,
         n_majority7_module_11__and_module_7_res,
         n_majority7_module_11__or_module_7_res,
         n_majority7_module_11__or_module_6_res,
         n_majority7_module_11__and_module_6_res,
         n_majority7_module_11__or_module_5_res,
         n_majority7_module_11__and_module_5_res,
         n_majority7_module_11__or_module_4_res,
         n_majority7_module_11__and_module_4_res,
         n_majority7_module_11__or_module_3_res,
         n_majority7_module_11__and_module_3_res,
         n_majority7_module_11__or_module_2_res,
         n_majority7_module_11__and_module_2_res,
         n_majority7_module_11__or_module_1_res,
         n_majority7_module_11__and_module_1_res,
         n_majority7_module_12__and_module_10_res,
         n_majority7_module_12__or_module_11_res,
         n_majority7_module_12__and_module_9_res,
         n_majority7_module_12__or_module_10_res,
         n_majority7_module_12__or_module_9_res,
         n_majority7_module_12__and_module_8_res,
         n_majority7_module_12__or_module_8_res,
         n_majority7_module_12__and_module_7_res,
         n_majority7_module_12__or_module_7_res,
         n_majority7_module_12__or_module_6_res,
         n_majority7_module_12__and_module_6_res,
         n_majority7_module_12__or_module_5_res,
         n_majority7_module_12__and_module_5_res,
         n_majority7_module_12__or_module_4_res,
         n_majority7_module_12__and_module_4_res,
         n_majority7_module_12__or_module_3_res,
         n_majority7_module_12__and_module_3_res,
         n_majority7_module_12__or_module_2_res,
         n_majority7_module_12__and_module_2_res,
         n_majority7_module_12__or_module_1_res,
         n_majority7_module_12__and_module_1_res,
         n_majority7_module_13__and_module_10_res,
         n_majority7_module_13__or_module_11_res,
         n_majority7_module_13__and_module_9_res,
         n_majority7_module_13__or_module_10_res,
         n_majority7_module_13__or_module_9_res,
         n_majority7_module_13__and_module_8_res,
         n_majority7_module_13__or_module_8_res,
         n_majority7_module_13__and_module_7_res,
         n_majority7_module_13__or_module_7_res,
         n_majority7_module_13__or_module_6_res,
         n_majority7_module_13__and_module_6_res,
         n_majority7_module_13__or_module_5_res,
         n_majority7_module_13__and_module_5_res,
         n_majority7_module_13__or_module_4_res,
         n_majority7_module_13__and_module_4_res,
         n_majority7_module_13__or_module_3_res,
         n_majority7_module_13__and_module_3_res,
         n_majority7_module_13__or_module_2_res,
         n_majority7_module_13__and_module_2_res,
         n_majority7_module_13__or_module_1_res,
         n_majority7_module_13__and_module_1_res,
         n_majority7_module_14__and_module_10_res,
         n_majority7_module_14__or_module_11_res,
         n_majority7_module_14__and_module_9_res,
         n_majority7_module_14__or_module_10_res,
         n_majority7_module_14__or_module_9_res,
         n_majority7_module_14__and_module_8_res,
         n_majority7_module_14__or_module_8_res,
         n_majority7_module_14__and_module_7_res,
         n_majority7_module_14__or_module_7_res,
         n_majority7_module_14__or_module_6_res,
         n_majority7_module_14__and_module_6_res,
         n_majority7_module_14__or_module_5_res,
         n_majority7_module_14__and_module_5_res,
         n_majority7_module_14__or_module_4_res,
         n_majority7_module_14__and_module_4_res,
         n_majority7_module_14__or_module_3_res,
         n_majority7_module_14__and_module_3_res,
         n_majority7_module_14__or_module_2_res,
         n_majority7_module_14__and_module_2_res,
         n_majority7_module_14__or_module_1_res,
         n_majority7_module_14__and_module_1_res,
         n_majority7_module_15__and_module_10_res,
         n_majority7_module_15__or_module_11_res,
         n_majority7_module_15__and_module_9_res,
         n_majority7_module_15__or_module_10_res,
         n_majority7_module_15__or_module_9_res,
         n_majority7_module_15__and_module_8_res,
         n_majority7_module_15__or_module_8_res,
         n_majority7_module_15__and_module_7_res,
         n_majority7_module_15__or_module_7_res,
         n_majority7_module_15__or_module_6_res,
         n_majority7_module_15__and_module_6_res,
         n_majority7_module_15__or_module_5_res,
         n_majority7_module_15__and_module_5_res,
         n_majority7_module_15__or_module_4_res,
         n_majority7_module_15__and_module_4_res,
         n_majority7_module_15__or_module_3_res,
         n_majority7_module_15__and_module_3_res,
         n_majority7_module_15__or_module_2_res,
         n_majority7_module_15__and_module_2_res,
         n_majority7_module_15__or_module_1_res,
         n_majority7_module_15__and_module_1_res,
         n_majority7_module_16__and_module_10_res,
         n_majority7_module_16__or_module_11_res,
         n_majority7_module_16__and_module_9_res,
         n_majority7_module_16__or_module_10_res,
         n_majority7_module_16__or_module_9_res,
         n_majority7_module_16__and_module_8_res,
         n_majority7_module_16__or_module_8_res,
         n_majority7_module_16__and_module_7_res,
         n_majority7_module_16__or_module_7_res,
         n_majority7_module_16__or_module_6_res,
         n_majority7_module_16__and_module_6_res,
         n_majority7_module_16__or_module_5_res,
         n_majority7_module_16__and_module_5_res,
         n_majority7_module_16__or_module_4_res,
         n_majority7_module_16__and_module_4_res,
         n_majority7_module_16__or_module_3_res,
         n_majority7_module_16__and_module_3_res,
         n_majority7_module_16__or_module_2_res,
         n_majority7_module_16__and_module_2_res,
         n_majority7_module_16__or_module_1_res,
         n_majority7_module_16__and_module_1_res,
         n_majority7_module_17__and_module_10_res,
         n_majority7_module_17__or_module_11_res,
         n_majority7_module_17__and_module_9_res,
         n_majority7_module_17__or_module_10_res,
         n_majority7_module_17__or_module_9_res,
         n_majority7_module_17__and_module_8_res,
         n_majority7_module_17__or_module_8_res,
         n_majority7_module_17__and_module_7_res,
         n_majority7_module_17__or_module_7_res,
         n_majority7_module_17__or_module_6_res,
         n_majority7_module_17__and_module_6_res,
         n_majority7_module_17__or_module_5_res,
         n_majority7_module_17__and_module_5_res,
         n_majority7_module_17__or_module_4_res,
         n_majority7_module_17__and_module_4_res,
         n_majority7_module_17__or_module_3_res,
         n_majority7_module_17__and_module_3_res,
         n_majority7_module_17__or_module_2_res,
         n_majority7_module_17__and_module_2_res,
         n_majority7_module_17__or_module_1_res,
         n_majority7_module_17__and_module_1_res,
         n_majority7_module_18__and_module_10_res,
         n_majority7_module_18__or_module_11_res,
         n_majority7_module_18__and_module_9_res,
         n_majority7_module_18__or_module_10_res,
         n_majority7_module_18__or_module_9_res,
         n_majority7_module_18__and_module_8_res,
         n_majority7_module_18__or_module_8_res,
         n_majority7_module_18__and_module_7_res,
         n_majority7_module_18__or_module_7_res,
         n_majority7_module_18__or_module_6_res,
         n_majority7_module_18__and_module_6_res,
         n_majority7_module_18__or_module_5_res,
         n_majority7_module_18__and_module_5_res,
         n_majority7_module_18__or_module_4_res,
         n_majority7_module_18__and_module_4_res,
         n_majority7_module_18__or_module_3_res,
         n_majority7_module_18__and_module_3_res,
         n_majority7_module_18__or_module_2_res,
         n_majority7_module_18__and_module_2_res,
         n_majority7_module_18__or_module_1_res,
         n_majority7_module_18__and_module_1_res,
         n_majority7_module_19__and_module_10_res,
         n_majority7_module_19__or_module_11_res,
         n_majority7_module_19__and_module_9_res,
         n_majority7_module_19__or_module_10_res,
         n_majority7_module_19__or_module_9_res,
         n_majority7_module_19__and_module_8_res,
         n_majority7_module_19__or_module_8_res,
         n_majority7_module_19__and_module_7_res,
         n_majority7_module_19__or_module_7_res,
         n_majority7_module_19__or_module_6_res,
         n_majority7_module_19__and_module_6_res,
         n_majority7_module_19__or_module_5_res,
         n_majority7_module_19__and_module_5_res,
         n_majority7_module_19__or_module_4_res,
         n_majority7_module_19__and_module_4_res,
         n_majority7_module_19__or_module_3_res,
         n_majority7_module_19__and_module_3_res,
         n_majority7_module_19__or_module_2_res,
         n_majority7_module_19__and_module_2_res,
         n_majority7_module_19__or_module_1_res,
         n_majority7_module_19__and_module_1_res,
         n_majority7_module_20__and_module_10_res,
         n_majority7_module_20__or_module_11_res,
         n_majority7_module_20__and_module_9_res,
         n_majority7_module_20__or_module_10_res,
         n_majority7_module_20__or_module_9_res,
         n_majority7_module_20__and_module_8_res,
         n_majority7_module_20__or_module_8_res,
         n_majority7_module_20__and_module_7_res,
         n_majority7_module_20__or_module_7_res,
         n_majority7_module_20__or_module_6_res,
         n_majority7_module_20__and_module_6_res,
         n_majority7_module_20__or_module_5_res,
         n_majority7_module_20__and_module_5_res,
         n_majority7_module_20__or_module_4_res,
         n_majority7_module_20__and_module_4_res,
         n_majority7_module_20__or_module_3_res,
         n_majority7_module_20__and_module_3_res,
         n_majority7_module_20__or_module_2_res,
         n_majority7_module_20__and_module_2_res,
         n_majority7_module_20__or_module_1_res,
         n_majority7_module_20__and_module_1_res,
         n_majority7_module_21__and_module_10_res,
         n_majority7_module_21__or_module_11_res,
         n_majority7_module_21__and_module_9_res,
         n_majority7_module_21__or_module_10_res,
         n_majority7_module_21__or_module_9_res,
         n_majority7_module_21__and_module_8_res,
         n_majority7_module_21__or_module_8_res,
         n_majority7_module_21__and_module_7_res,
         n_majority7_module_21__or_module_7_res,
         n_majority7_module_21__or_module_6_res,
         n_majority7_module_21__and_module_6_res,
         n_majority7_module_21__or_module_5_res,
         n_majority7_module_21__and_module_5_res,
         n_majority7_module_21__or_module_4_res,
         n_majority7_module_21__and_module_4_res,
         n_majority7_module_21__or_module_3_res,
         n_majority7_module_21__and_module_3_res,
         n_majority7_module_21__or_module_2_res,
         n_majority7_module_21__and_module_2_res,
         n_majority7_module_21__or_module_1_res,
         n_majority7_module_21__and_module_1_res,
         n_majority7_module_22__and_module_10_res,
         n_majority7_module_22__or_module_11_res,
         n_majority7_module_22__and_module_9_res,
         n_majority7_module_22__or_module_10_res,
         n_majority7_module_22__or_module_9_res,
         n_majority7_module_22__and_module_8_res,
         n_majority7_module_22__or_module_8_res,
         n_majority7_module_22__and_module_7_res,
         n_majority7_module_22__or_module_7_res,
         n_majority7_module_22__or_module_6_res,
         n_majority7_module_22__and_module_6_res,
         n_majority7_module_22__or_module_5_res,
         n_majority7_module_22__and_module_5_res,
         n_majority7_module_22__or_module_4_res,
         n_majority7_module_22__and_module_4_res,
         n_majority7_module_22__or_module_3_res,
         n_majority7_module_22__and_module_3_res,
         n_majority7_module_22__or_module_2_res,
         n_majority7_module_22__and_module_2_res,
         n_majority7_module_22__or_module_1_res,
         n_majority7_module_22__and_module_1_res,
         n_majority7_module_23__and_module_10_res,
         n_majority7_module_23__or_module_11_res,
         n_majority7_module_23__and_module_9_res,
         n_majority7_module_23__or_module_10_res,
         n_majority7_module_23__or_module_9_res,
         n_majority7_module_23__and_module_8_res,
         n_majority7_module_23__or_module_8_res,
         n_majority7_module_23__and_module_7_res,
         n_majority7_module_23__or_module_7_res,
         n_majority7_module_23__or_module_6_res,
         n_majority7_module_23__and_module_6_res,
         n_majority7_module_23__or_module_5_res,
         n_majority7_module_23__and_module_5_res,
         n_majority7_module_23__or_module_4_res,
         n_majority7_module_23__and_module_4_res,
         n_majority7_module_23__or_module_3_res,
         n_majority7_module_23__and_module_3_res,
         n_majority7_module_23__or_module_2_res,
         n_majority7_module_23__and_module_2_res,
         n_majority7_module_23__or_module_1_res,
         n_majority7_module_23__and_module_1_res,
         n_majority7_module_24__and_module_10_res,
         n_majority7_module_24__or_module_11_res,
         n_majority7_module_24__and_module_9_res,
         n_majority7_module_24__or_module_10_res,
         n_majority7_module_24__or_module_9_res,
         n_majority7_module_24__and_module_8_res,
         n_majority7_module_24__or_module_8_res,
         n_majority7_module_24__and_module_7_res,
         n_majority7_module_24__or_module_7_res,
         n_majority7_module_24__or_module_6_res,
         n_majority7_module_24__and_module_6_res,
         n_majority7_module_24__or_module_5_res,
         n_majority7_module_24__and_module_5_res,
         n_majority7_module_24__or_module_4_res,
         n_majority7_module_24__and_module_4_res,
         n_majority7_module_24__or_module_3_res,
         n_majority7_module_24__and_module_3_res,
         n_majority7_module_24__or_module_2_res,
         n_majority7_module_24__and_module_2_res,
         n_majority7_module_24__or_module_1_res,
         n_majority7_module_24__and_module_1_res,
         n_majority7_module_25__and_module_10_res,
         n_majority7_module_25__or_module_11_res,
         n_majority7_module_25__and_module_9_res,
         n_majority7_module_25__or_module_10_res,
         n_majority7_module_25__or_module_9_res,
         n_majority7_module_25__and_module_8_res,
         n_majority7_module_25__or_module_8_res,
         n_majority7_module_25__and_module_7_res,
         n_majority7_module_25__or_module_7_res,
         n_majority7_module_25__or_module_6_res,
         n_majority7_module_25__and_module_6_res,
         n_majority7_module_25__or_module_5_res,
         n_majority7_module_25__and_module_5_res,
         n_majority7_module_25__or_module_4_res,
         n_majority7_module_25__and_module_4_res,
         n_majority7_module_25__or_module_3_res,
         n_majority7_module_25__and_module_3_res,
         n_majority7_module_25__or_module_2_res,
         n_majority7_module_25__and_module_2_res,
         n_majority7_module_25__or_module_1_res,
         n_majority7_module_25__and_module_1_res,
         n_majority7_module_26__and_module_10_res,
         n_majority7_module_26__or_module_11_res,
         n_majority7_module_26__and_module_9_res,
         n_majority7_module_26__or_module_10_res,
         n_majority7_module_26__or_module_9_res,
         n_majority7_module_26__and_module_8_res,
         n_majority7_module_26__or_module_8_res,
         n_majority7_module_26__and_module_7_res,
         n_majority7_module_26__or_module_7_res,
         n_majority7_module_26__or_module_6_res,
         n_majority7_module_26__and_module_6_res,
         n_majority7_module_26__or_module_5_res,
         n_majority7_module_26__and_module_5_res,
         n_majority7_module_26__or_module_4_res,
         n_majority7_module_26__and_module_4_res,
         n_majority7_module_26__or_module_3_res,
         n_majority7_module_26__and_module_3_res,
         n_majority7_module_26__or_module_2_res,
         n_majority7_module_26__and_module_2_res,
         n_majority7_module_26__or_module_1_res,
         n_majority7_module_26__and_module_1_res,
         n_majority7_module_27__and_module_10_res,
         n_majority7_module_27__or_module_11_res,
         n_majority7_module_27__and_module_9_res,
         n_majority7_module_27__or_module_10_res,
         n_majority7_module_27__or_module_9_res,
         n_majority7_module_27__and_module_8_res,
         n_majority7_module_27__or_module_8_res,
         n_majority7_module_27__and_module_7_res,
         n_majority7_module_27__or_module_7_res,
         n_majority7_module_27__or_module_6_res,
         n_majority7_module_27__and_module_6_res,
         n_majority7_module_27__or_module_5_res,
         n_majority7_module_27__and_module_5_res,
         n_majority7_module_27__or_module_4_res,
         n_majority7_module_27__and_module_4_res,
         n_majority7_module_27__or_module_3_res,
         n_majority7_module_27__and_module_3_res,
         n_majority7_module_27__or_module_2_res,
         n_majority7_module_27__and_module_2_res,
         n_majority7_module_27__or_module_1_res,
         n_majority7_module_27__and_module_1_res,
         n_majority7_module_28__and_module_10_res,
         n_majority7_module_28__or_module_11_res,
         n_majority7_module_28__and_module_9_res,
         n_majority7_module_28__or_module_10_res,
         n_majority7_module_28__or_module_9_res,
         n_majority7_module_28__and_module_8_res,
         n_majority7_module_28__or_module_8_res,
         n_majority7_module_28__and_module_7_res,
         n_majority7_module_28__or_module_7_res,
         n_majority7_module_28__or_module_6_res,
         n_majority7_module_28__and_module_6_res,
         n_majority7_module_28__or_module_5_res,
         n_majority7_module_28__and_module_5_res,
         n_majority7_module_28__or_module_4_res,
         n_majority7_module_28__and_module_4_res,
         n_majority7_module_28__or_module_3_res,
         n_majority7_module_28__and_module_3_res,
         n_majority7_module_28__or_module_2_res,
         n_majority7_module_28__and_module_2_res,
         n_majority7_module_28__or_module_1_res,
         n_majority7_module_28__and_module_1_res,
         n_majority7_module_29__and_module_10_res,
         n_majority7_module_29__or_module_11_res,
         n_majority7_module_29__and_module_9_res,
         n_majority7_module_29__or_module_10_res,
         n_majority7_module_29__or_module_9_res,
         n_majority7_module_29__and_module_8_res,
         n_majority7_module_29__or_module_8_res,
         n_majority7_module_29__and_module_7_res,
         n_majority7_module_29__or_module_7_res,
         n_majority7_module_29__or_module_6_res,
         n_majority7_module_29__and_module_6_res,
         n_majority7_module_29__or_module_5_res,
         n_majority7_module_29__and_module_5_res,
         n_majority7_module_29__or_module_4_res,
         n_majority7_module_29__and_module_4_res,
         n_majority7_module_29__or_module_3_res,
         n_majority7_module_29__and_module_3_res,
         n_majority7_module_29__or_module_2_res,
         n_majority7_module_29__and_module_2_res,
         n_majority7_module_29__or_module_1_res,
         n_majority7_module_29__and_module_1_res,
         n_majority7_module_30__and_module_10_res,
         n_majority7_module_30__or_module_11_res,
         n_majority7_module_30__and_module_9_res,
         n_majority7_module_30__or_module_10_res,
         n_majority7_module_30__or_module_9_res,
         n_majority7_module_30__and_module_8_res,
         n_majority7_module_30__or_module_8_res,
         n_majority7_module_30__and_module_7_res,
         n_majority7_module_30__or_module_7_res,
         n_majority7_module_30__or_module_6_res,
         n_majority7_module_30__and_module_6_res,
         n_majority7_module_30__or_module_5_res,
         n_majority7_module_30__and_module_5_res,
         n_majority7_module_30__or_module_4_res,
         n_majority7_module_30__and_module_4_res,
         n_majority7_module_30__or_module_3_res,
         n_majority7_module_30__and_module_3_res,
         n_majority7_module_30__or_module_2_res,
         n_majority7_module_30__and_module_2_res,
         n_majority7_module_30__or_module_1_res,
         n_majority7_module_30__and_module_1_res,
         n_majority7_module_31__and_module_10_res,
         n_majority7_module_31__or_module_11_res,
         n_majority7_module_31__and_module_9_res,
         n_majority7_module_31__or_module_10_res,
         n_majority7_module_31__or_module_9_res,
         n_majority7_module_31__and_module_8_res,
         n_majority7_module_31__or_module_8_res,
         n_majority7_module_31__and_module_7_res,
         n_majority7_module_31__or_module_7_res,
         n_majority7_module_31__or_module_6_res,
         n_majority7_module_31__and_module_6_res,
         n_majority7_module_31__or_module_5_res,
         n_majority7_module_31__and_module_5_res,
         n_majority7_module_31__or_module_4_res,
         n_majority7_module_31__and_module_4_res,
         n_majority7_module_31__or_module_3_res,
         n_majority7_module_31__and_module_3_res,
         n_majority7_module_31__or_module_2_res,
         n_majority7_module_31__and_module_2_res,
         n_majority7_module_31__or_module_1_res,
         n_majority7_module_31__and_module_1_res,
         n_majority7_module_32__and_module_10_res,
         n_majority7_module_32__or_module_11_res,
         n_majority7_module_32__and_module_9_res,
         n_majority7_module_32__or_module_10_res,
         n_majority7_module_32__or_module_9_res,
         n_majority7_module_32__and_module_8_res,
         n_majority7_module_32__or_module_8_res,
         n_majority7_module_32__and_module_7_res,
         n_majority7_module_32__or_module_7_res,
         n_majority7_module_32__or_module_6_res,
         n_majority7_module_32__and_module_6_res,
         n_majority7_module_32__or_module_5_res,
         n_majority7_module_32__and_module_5_res,
         n_majority7_module_32__or_module_4_res,
         n_majority7_module_32__and_module_4_res,
         n_majority7_module_32__or_module_3_res,
         n_majority7_module_32__and_module_3_res,
         n_majority7_module_32__or_module_2_res,
         n_majority7_module_32__and_module_2_res,
         n_majority7_module_32__or_module_1_res,
         n_majority7_module_32__and_module_1_res,
         n_majority7_module_33__and_module_10_res,
         n_majority7_module_33__or_module_11_res,
         n_majority7_module_33__and_module_9_res,
         n_majority7_module_33__or_module_10_res,
         n_majority7_module_33__or_module_9_res,
         n_majority7_module_33__and_module_8_res,
         n_majority7_module_33__or_module_8_res,
         n_majority7_module_33__and_module_7_res,
         n_majority7_module_33__or_module_7_res,
         n_majority7_module_33__or_module_6_res,
         n_majority7_module_33__and_module_6_res,
         n_majority7_module_33__or_module_5_res,
         n_majority7_module_33__and_module_5_res,
         n_majority7_module_33__or_module_4_res,
         n_majority7_module_33__and_module_4_res,
         n_majority7_module_33__or_module_3_res,
         n_majority7_module_33__and_module_3_res,
         n_majority7_module_33__or_module_2_res,
         n_majority7_module_33__and_module_2_res,
         n_majority7_module_33__or_module_1_res,
         n_majority7_module_33__and_module_1_res,
         n_majority7_module_34__and_module_10_res,
         n_majority7_module_34__or_module_11_res,
         n_majority7_module_34__and_module_9_res,
         n_majority7_module_34__or_module_10_res,
         n_majority7_module_34__or_module_9_res,
         n_majority7_module_34__and_module_8_res,
         n_majority7_module_34__or_module_8_res,
         n_majority7_module_34__and_module_7_res,
         n_majority7_module_34__or_module_7_res,
         n_majority7_module_34__or_module_6_res,
         n_majority7_module_34__and_module_6_res,
         n_majority7_module_34__or_module_5_res,
         n_majority7_module_34__and_module_5_res,
         n_majority7_module_34__or_module_4_res,
         n_majority7_module_34__and_module_4_res,
         n_majority7_module_34__or_module_3_res,
         n_majority7_module_34__and_module_3_res,
         n_majority7_module_34__or_module_2_res,
         n_majority7_module_34__and_module_2_res,
         n_majority7_module_34__or_module_1_res,
         n_majority7_module_34__and_module_1_res,
         n_majority7_module_35__and_module_10_res,
         n_majority7_module_35__or_module_11_res,
         n_majority7_module_35__and_module_9_res,
         n_majority7_module_35__or_module_10_res,
         n_majority7_module_35__or_module_9_res,
         n_majority7_module_35__and_module_8_res,
         n_majority7_module_35__or_module_8_res,
         n_majority7_module_35__and_module_7_res,
         n_majority7_module_35__or_module_7_res,
         n_majority7_module_35__or_module_6_res,
         n_majority7_module_35__and_module_6_res,
         n_majority7_module_35__or_module_5_res,
         n_majority7_module_35__and_module_5_res,
         n_majority7_module_35__or_module_4_res,
         n_majority7_module_35__and_module_4_res,
         n_majority7_module_35__or_module_3_res,
         n_majority7_module_35__and_module_3_res,
         n_majority7_module_35__or_module_2_res,
         n_majority7_module_35__and_module_2_res,
         n_majority7_module_35__or_module_1_res,
         n_majority7_module_35__and_module_1_res,
         n_majority7_module_36__and_module_10_res,
         n_majority7_module_36__or_module_11_res,
         n_majority7_module_36__and_module_9_res,
         n_majority7_module_36__or_module_10_res,
         n_majority7_module_36__or_module_9_res,
         n_majority7_module_36__and_module_8_res,
         n_majority7_module_36__or_module_8_res,
         n_majority7_module_36__and_module_7_res,
         n_majority7_module_36__or_module_7_res,
         n_majority7_module_36__or_module_6_res,
         n_majority7_module_36__and_module_6_res,
         n_majority7_module_36__or_module_5_res,
         n_majority7_module_36__and_module_5_res,
         n_majority7_module_36__or_module_4_res,
         n_majority7_module_36__and_module_4_res,
         n_majority7_module_36__or_module_3_res,
         n_majority7_module_36__and_module_3_res,
         n_majority7_module_36__or_module_2_res,
         n_majority7_module_36__and_module_2_res,
         n_majority7_module_36__or_module_1_res,
         n_majority7_module_36__and_module_1_res,
         n_majority7_module_37__and_module_10_res,
         n_majority7_module_37__or_module_11_res,
         n_majority7_module_37__and_module_9_res,
         n_majority7_module_37__or_module_10_res,
         n_majority7_module_37__or_module_9_res,
         n_majority7_module_37__and_module_8_res,
         n_majority7_module_37__or_module_8_res,
         n_majority7_module_37__and_module_7_res,
         n_majority7_module_37__or_module_7_res,
         n_majority7_module_37__or_module_6_res,
         n_majority7_module_37__and_module_6_res,
         n_majority7_module_37__or_module_5_res,
         n_majority7_module_37__and_module_5_res,
         n_majority7_module_37__or_module_4_res,
         n_majority7_module_37__and_module_4_res,
         n_majority7_module_37__or_module_3_res,
         n_majority7_module_37__and_module_3_res,
         n_majority7_module_37__or_module_2_res,
         n_majority7_module_37__and_module_2_res,
         n_majority7_module_37__or_module_1_res,
         n_majority7_module_37__and_module_1_res,
         n_majority7_module_38__and_module_10_res,
         n_majority7_module_38__or_module_11_res,
         n_majority7_module_38__and_module_9_res,
         n_majority7_module_38__or_module_10_res,
         n_majority7_module_38__or_module_9_res,
         n_majority7_module_38__and_module_8_res,
         n_majority7_module_38__or_module_8_res,
         n_majority7_module_38__and_module_7_res,
         n_majority7_module_38__or_module_7_res,
         n_majority7_module_38__or_module_6_res,
         n_majority7_module_38__and_module_6_res,
         n_majority7_module_38__or_module_5_res,
         n_majority7_module_38__and_module_5_res,
         n_majority7_module_38__or_module_4_res,
         n_majority7_module_38__and_module_4_res,
         n_majority7_module_38__or_module_3_res,
         n_majority7_module_38__and_module_3_res,
         n_majority7_module_38__or_module_2_res,
         n_majority7_module_38__and_module_2_res,
         n_majority7_module_38__or_module_1_res,
         n_majority7_module_38__and_module_1_res,
         n_majority7_module_39__and_module_10_res,
         n_majority7_module_39__or_module_11_res,
         n_majority7_module_39__and_module_9_res,
         n_majority7_module_39__or_module_10_res,
         n_majority7_module_39__or_module_9_res,
         n_majority7_module_39__and_module_8_res,
         n_majority7_module_39__or_module_8_res,
         n_majority7_module_39__and_module_7_res,
         n_majority7_module_39__or_module_7_res,
         n_majority7_module_39__or_module_6_res,
         n_majority7_module_39__and_module_6_res,
         n_majority7_module_39__or_module_5_res,
         n_majority7_module_39__and_module_5_res,
         n_majority7_module_39__or_module_4_res,
         n_majority7_module_39__and_module_4_res,
         n_majority7_module_39__or_module_3_res,
         n_majority7_module_39__and_module_3_res,
         n_majority7_module_39__or_module_2_res,
         n_majority7_module_39__and_module_2_res,
         n_majority7_module_39__or_module_1_res,
         n_majority7_module_39__and_module_1_res,
         n_majority7_module_40__and_module_10_res,
         n_majority7_module_40__or_module_11_res,
         n_majority7_module_40__and_module_9_res,
         n_majority7_module_40__or_module_10_res,
         n_majority7_module_40__or_module_9_res,
         n_majority7_module_40__and_module_8_res,
         n_majority7_module_40__or_module_8_res,
         n_majority7_module_40__and_module_7_res,
         n_majority7_module_40__or_module_7_res,
         n_majority7_module_40__or_module_6_res,
         n_majority7_module_40__and_module_6_res,
         n_majority7_module_40__or_module_5_res,
         n_majority7_module_40__and_module_5_res,
         n_majority7_module_40__or_module_4_res,
         n_majority7_module_40__and_module_4_res,
         n_majority7_module_40__or_module_3_res,
         n_majority7_module_40__and_module_3_res,
         n_majority7_module_40__or_module_2_res,
         n_majority7_module_40__and_module_2_res,
         n_majority7_module_40__or_module_1_res,
         n_majority7_module_40__and_module_1_res,
         n_majority7_module_41__and_module_10_res,
         n_majority7_module_41__or_module_11_res,
         n_majority7_module_41__and_module_9_res,
         n_majority7_module_41__or_module_10_res,
         n_majority7_module_41__or_module_9_res,
         n_majority7_module_41__and_module_8_res,
         n_majority7_module_41__or_module_8_res,
         n_majority7_module_41__and_module_7_res,
         n_majority7_module_41__or_module_7_res,
         n_majority7_module_41__or_module_6_res,
         n_majority7_module_41__and_module_6_res,
         n_majority7_module_41__or_module_5_res,
         n_majority7_module_41__and_module_5_res,
         n_majority7_module_41__or_module_4_res,
         n_majority7_module_41__and_module_4_res,
         n_majority7_module_41__or_module_3_res,
         n_majority7_module_41__and_module_3_res,
         n_majority7_module_41__or_module_2_res,
         n_majority7_module_41__and_module_2_res,
         n_majority7_module_41__or_module_1_res,
         n_majority7_module_41__and_module_1_res,
         n_majority7_module_42__and_module_10_res,
         n_majority7_module_42__or_module_11_res,
         n_majority7_module_42__and_module_9_res,
         n_majority7_module_42__or_module_10_res,
         n_majority7_module_42__or_module_9_res,
         n_majority7_module_42__and_module_8_res,
         n_majority7_module_42__or_module_8_res,
         n_majority7_module_42__and_module_7_res,
         n_majority7_module_42__or_module_7_res,
         n_majority7_module_42__or_module_6_res,
         n_majority7_module_42__and_module_6_res,
         n_majority7_module_42__or_module_5_res,
         n_majority7_module_42__and_module_5_res,
         n_majority7_module_42__or_module_4_res,
         n_majority7_module_42__and_module_4_res,
         n_majority7_module_42__or_module_3_res,
         n_majority7_module_42__and_module_3_res,
         n_majority7_module_42__or_module_2_res,
         n_majority7_module_42__and_module_2_res,
         n_majority7_module_42__or_module_1_res,
         n_majority7_module_42__and_module_1_res,
         n_majority7_module_43__and_module_10_res,
         n_majority7_module_43__or_module_11_res,
         n_majority7_module_43__and_module_9_res,
         n_majority7_module_43__or_module_10_res,
         n_majority7_module_43__or_module_9_res,
         n_majority7_module_43__and_module_8_res,
         n_majority7_module_43__or_module_8_res,
         n_majority7_module_43__and_module_7_res,
         n_majority7_module_43__or_module_7_res,
         n_majority7_module_43__or_module_6_res,
         n_majority7_module_43__and_module_6_res,
         n_majority7_module_43__or_module_5_res,
         n_majority7_module_43__and_module_5_res,
         n_majority7_module_43__or_module_4_res,
         n_majority7_module_43__and_module_4_res,
         n_majority7_module_43__or_module_3_res,
         n_majority7_module_43__and_module_3_res,
         n_majority7_module_43__or_module_2_res,
         n_majority7_module_43__and_module_2_res,
         n_majority7_module_43__or_module_1_res,
         n_majority7_module_43__and_module_1_res,
         n_majority7_module_44__and_module_10_res,
         n_majority7_module_44__or_module_11_res,
         n_majority7_module_44__and_module_9_res,
         n_majority7_module_44__or_module_10_res,
         n_majority7_module_44__or_module_9_res,
         n_majority7_module_44__and_module_8_res,
         n_majority7_module_44__or_module_8_res,
         n_majority7_module_44__and_module_7_res,
         n_majority7_module_44__or_module_7_res,
         n_majority7_module_44__or_module_6_res,
         n_majority7_module_44__and_module_6_res,
         n_majority7_module_44__or_module_5_res,
         n_majority7_module_44__and_module_5_res,
         n_majority7_module_44__or_module_4_res,
         n_majority7_module_44__and_module_4_res,
         n_majority7_module_44__or_module_3_res,
         n_majority7_module_44__and_module_3_res,
         n_majority7_module_44__or_module_2_res,
         n_majority7_module_44__and_module_2_res,
         n_majority7_module_44__or_module_1_res,
         n_majority7_module_44__and_module_1_res,
         n_majority7_module_45__and_module_10_res,
         n_majority7_module_45__or_module_11_res,
         n_majority7_module_45__and_module_9_res,
         n_majority7_module_45__or_module_10_res,
         n_majority7_module_45__or_module_9_res,
         n_majority7_module_45__and_module_8_res,
         n_majority7_module_45__or_module_8_res,
         n_majority7_module_45__and_module_7_res,
         n_majority7_module_45__or_module_7_res,
         n_majority7_module_45__or_module_6_res,
         n_majority7_module_45__and_module_6_res,
         n_majority7_module_45__or_module_5_res,
         n_majority7_module_45__and_module_5_res,
         n_majority7_module_45__or_module_4_res,
         n_majority7_module_45__and_module_4_res,
         n_majority7_module_45__or_module_3_res,
         n_majority7_module_45__and_module_3_res,
         n_majority7_module_45__or_module_2_res,
         n_majority7_module_45__and_module_2_res,
         n_majority7_module_45__or_module_1_res,
         n_majority7_module_45__and_module_1_res,
         n_majority7_module_46__and_module_10_res,
         n_majority7_module_46__or_module_11_res,
         n_majority7_module_46__and_module_9_res,
         n_majority7_module_46__or_module_10_res,
         n_majority7_module_46__or_module_9_res,
         n_majority7_module_46__and_module_8_res,
         n_majority7_module_46__or_module_8_res,
         n_majority7_module_46__and_module_7_res,
         n_majority7_module_46__or_module_7_res,
         n_majority7_module_46__or_module_6_res,
         n_majority7_module_46__and_module_6_res,
         n_majority7_module_46__or_module_5_res,
         n_majority7_module_46__and_module_5_res,
         n_majority7_module_46__or_module_4_res,
         n_majority7_module_46__and_module_4_res,
         n_majority7_module_46__or_module_3_res,
         n_majority7_module_46__and_module_3_res,
         n_majority7_module_46__or_module_2_res,
         n_majority7_module_46__and_module_2_res,
         n_majority7_module_46__or_module_1_res,
         n_majority7_module_46__and_module_1_res,
         n_majority7_module_47__and_module_10_res,
         n_majority7_module_47__or_module_11_res,
         n_majority7_module_47__and_module_9_res,
         n_majority7_module_47__or_module_10_res,
         n_majority7_module_47__or_module_9_res,
         n_majority7_module_47__and_module_8_res,
         n_majority7_module_47__or_module_8_res,
         n_majority7_module_47__and_module_7_res,
         n_majority7_module_47__or_module_7_res,
         n_majority7_module_47__or_module_6_res,
         n_majority7_module_47__and_module_6_res,
         n_majority7_module_47__or_module_5_res,
         n_majority7_module_47__and_module_5_res,
         n_majority7_module_47__or_module_4_res,
         n_majority7_module_47__and_module_4_res,
         n_majority7_module_47__or_module_3_res,
         n_majority7_module_47__and_module_3_res,
         n_majority7_module_47__or_module_2_res,
         n_majority7_module_47__and_module_2_res,
         n_majority7_module_47__or_module_1_res,
         n_majority7_module_47__and_module_1_res,
         n_majority7_module_48__and_module_10_res,
         n_majority7_module_48__or_module_11_res,
         n_majority7_module_48__and_module_9_res,
         n_majority7_module_48__or_module_10_res,
         n_majority7_module_48__or_module_9_res,
         n_majority7_module_48__and_module_8_res,
         n_majority7_module_48__or_module_8_res,
         n_majority7_module_48__and_module_7_res,
         n_majority7_module_48__or_module_7_res,
         n_majority7_module_48__or_module_6_res,
         n_majority7_module_48__and_module_6_res,
         n_majority7_module_48__or_module_5_res,
         n_majority7_module_48__and_module_5_res,
         n_majority7_module_48__or_module_4_res,
         n_majority7_module_48__and_module_4_res,
         n_majority7_module_48__or_module_3_res,
         n_majority7_module_48__and_module_3_res,
         n_majority7_module_48__or_module_2_res,
         n_majority7_module_48__and_module_2_res,
         n_majority7_module_48__or_module_1_res,
         n_majority7_module_48__and_module_1_res,
         n_majority7_module_49__and_module_10_res,
         n_majority7_module_49__or_module_11_res,
         n_majority7_module_49__and_module_9_res,
         n_majority7_module_49__or_module_10_res,
         n_majority7_module_49__or_module_9_res,
         n_majority7_module_49__and_module_8_res,
         n_majority7_module_49__or_module_8_res,
         n_majority7_module_49__and_module_7_res,
         n_majority7_module_49__or_module_7_res,
         n_majority7_module_49__or_module_6_res,
         n_majority7_module_49__and_module_6_res,
         n_majority7_module_49__or_module_5_res,
         n_majority7_module_49__and_module_5_res,
         n_majority7_module_49__or_module_4_res,
         n_majority7_module_49__and_module_4_res,
         n_majority7_module_49__or_module_3_res,
         n_majority7_module_49__and_module_3_res,
         n_majority7_module_49__or_module_2_res,
         n_majority7_module_49__and_module_2_res,
         n_majority7_module_49__or_module_1_res,
         n_majority7_module_49__and_module_1_res,
         n_majority7_module_50__and_module_10_res,
         n_majority7_module_50__or_module_11_res,
         n_majority7_module_50__and_module_9_res,
         n_majority7_module_50__or_module_10_res,
         n_majority7_module_50__or_module_9_res,
         n_majority7_module_50__and_module_8_res,
         n_majority7_module_50__or_module_8_res,
         n_majority7_module_50__and_module_7_res,
         n_majority7_module_50__or_module_7_res,
         n_majority7_module_50__or_module_6_res,
         n_majority7_module_50__and_module_6_res,
         n_majority7_module_50__or_module_5_res,
         n_majority7_module_50__and_module_5_res,
         n_majority7_module_50__or_module_4_res,
         n_majority7_module_50__and_module_4_res,
         n_majority7_module_50__or_module_3_res,
         n_majority7_module_50__and_module_3_res,
         n_majority7_module_50__or_module_2_res,
         n_majority7_module_50__and_module_2_res,
         n_majority7_module_50__or_module_1_res,
         n_majority7_module_50__and_module_1_res,
         n_majority7_module_51__and_module_10_res,
         n_majority7_module_51__or_module_11_res,
         n_majority7_module_51__and_module_9_res,
         n_majority7_module_51__or_module_10_res,
         n_majority7_module_51__or_module_9_res,
         n_majority7_module_51__and_module_8_res,
         n_majority7_module_51__or_module_8_res,
         n_majority7_module_51__and_module_7_res,
         n_majority7_module_51__or_module_7_res,
         n_majority7_module_51__or_module_6_res,
         n_majority7_module_51__and_module_6_res,
         n_majority7_module_51__or_module_5_res,
         n_majority7_module_51__and_module_5_res,
         n_majority7_module_51__or_module_4_res,
         n_majority7_module_51__and_module_4_res,
         n_majority7_module_51__or_module_3_res,
         n_majority7_module_51__and_module_3_res,
         n_majority7_module_51__or_module_2_res,
         n_majority7_module_51__and_module_2_res,
         n_majority7_module_51__or_module_1_res,
         n_majority7_module_51__and_module_1_res,
         n_majority7_module_52__and_module_10_res,
         n_majority7_module_52__or_module_11_res,
         n_majority7_module_52__and_module_9_res,
         n_majority7_module_52__or_module_10_res,
         n_majority7_module_52__or_module_9_res,
         n_majority7_module_52__and_module_8_res,
         n_majority7_module_52__or_module_8_res,
         n_majority7_module_52__and_module_7_res,
         n_majority7_module_52__or_module_7_res,
         n_majority7_module_52__or_module_6_res,
         n_majority7_module_52__and_module_6_res,
         n_majority7_module_52__or_module_5_res,
         n_majority7_module_52__and_module_5_res,
         n_majority7_module_52__or_module_4_res,
         n_majority7_module_52__and_module_4_res,
         n_majority7_module_52__or_module_3_res,
         n_majority7_module_52__and_module_3_res,
         n_majority7_module_52__or_module_2_res,
         n_majority7_module_52__and_module_2_res,
         n_majority7_module_52__or_module_1_res,
         n_majority7_module_52__and_module_1_res,
         n_majority7_module_53__and_module_10_res,
         n_majority7_module_53__or_module_11_res,
         n_majority7_module_53__and_module_9_res,
         n_majority7_module_53__or_module_10_res,
         n_majority7_module_53__or_module_9_res,
         n_majority7_module_53__and_module_8_res,
         n_majority7_module_53__or_module_8_res,
         n_majority7_module_53__and_module_7_res,
         n_majority7_module_53__or_module_7_res,
         n_majority7_module_53__or_module_6_res,
         n_majority7_module_53__and_module_6_res,
         n_majority7_module_53__or_module_5_res,
         n_majority7_module_53__and_module_5_res,
         n_majority7_module_53__or_module_4_res,
         n_majority7_module_53__and_module_4_res,
         n_majority7_module_53__or_module_3_res,
         n_majority7_module_53__and_module_3_res,
         n_majority7_module_53__or_module_2_res,
         n_majority7_module_53__and_module_2_res,
         n_majority7_module_53__or_module_1_res,
         n_majority7_module_53__and_module_1_res,
         n_majority7_module_54__and_module_10_res,
         n_majority7_module_54__or_module_11_res,
         n_majority7_module_54__and_module_9_res,
         n_majority7_module_54__or_module_10_res,
         n_majority7_module_54__or_module_9_res,
         n_majority7_module_54__and_module_8_res,
         n_majority7_module_54__or_module_8_res,
         n_majority7_module_54__and_module_7_res,
         n_majority7_module_54__or_module_7_res,
         n_majority7_module_54__or_module_6_res,
         n_majority7_module_54__and_module_6_res,
         n_majority7_module_54__or_module_5_res,
         n_majority7_module_54__and_module_5_res,
         n_majority7_module_54__or_module_4_res,
         n_majority7_module_54__and_module_4_res,
         n_majority7_module_54__or_module_3_res,
         n_majority7_module_54__and_module_3_res,
         n_majority7_module_54__or_module_2_res,
         n_majority7_module_54__and_module_2_res,
         n_majority7_module_54__or_module_1_res,
         n_majority7_module_54__and_module_1_res,
         n_majority7_module_55__and_module_10_res,
         n_majority7_module_55__or_module_11_res,
         n_majority7_module_55__and_module_9_res,
         n_majority7_module_55__or_module_10_res,
         n_majority7_module_55__or_module_9_res,
         n_majority7_module_55__and_module_8_res,
         n_majority7_module_55__or_module_8_res,
         n_majority7_module_55__and_module_7_res,
         n_majority7_module_55__or_module_7_res,
         n_majority7_module_55__or_module_6_res,
         n_majority7_module_55__and_module_6_res,
         n_majority7_module_55__or_module_5_res,
         n_majority7_module_55__and_module_5_res,
         n_majority7_module_55__or_module_4_res,
         n_majority7_module_55__and_module_4_res,
         n_majority7_module_55__or_module_3_res,
         n_majority7_module_55__and_module_3_res,
         n_majority7_module_55__or_module_2_res,
         n_majority7_module_55__and_module_2_res,
         n_majority7_module_55__or_module_1_res,
         n_majority7_module_55__and_module_1_res,
         n_majority7_module_56__and_module_10_res,
         n_majority7_module_56__or_module_11_res,
         n_majority7_module_56__and_module_9_res,
         n_majority7_module_56__or_module_10_res,
         n_majority7_module_56__or_module_9_res,
         n_majority7_module_56__and_module_8_res,
         n_majority7_module_56__or_module_8_res,
         n_majority7_module_56__and_module_7_res,
         n_majority7_module_56__or_module_7_res,
         n_majority7_module_56__or_module_6_res,
         n_majority7_module_56__and_module_6_res,
         n_majority7_module_56__or_module_5_res,
         n_majority7_module_56__and_module_5_res,
         n_majority7_module_56__or_module_4_res,
         n_majority7_module_56__and_module_4_res,
         n_majority7_module_56__or_module_3_res,
         n_majority7_module_56__and_module_3_res,
         n_majority7_module_56__or_module_2_res,
         n_majority7_module_56__and_module_2_res,
         n_majority7_module_56__or_module_1_res,
         n_majority7_module_56__and_module_1_res,
         n_majority7_module_57__and_module_10_res,
         n_majority7_module_57__or_module_11_res,
         n_majority7_module_57__and_module_9_res,
         n_majority7_module_57__or_module_10_res,
         n_majority7_module_57__or_module_9_res,
         n_majority7_module_57__and_module_8_res,
         n_majority7_module_57__or_module_8_res,
         n_majority7_module_57__and_module_7_res,
         n_majority7_module_57__or_module_7_res,
         n_majority7_module_57__or_module_6_res,
         n_majority7_module_57__and_module_6_res,
         n_majority7_module_57__or_module_5_res,
         n_majority7_module_57__and_module_5_res,
         n_majority7_module_57__or_module_4_res,
         n_majority7_module_57__and_module_4_res,
         n_majority7_module_57__or_module_3_res,
         n_majority7_module_57__and_module_3_res,
         n_majority7_module_57__or_module_2_res,
         n_majority7_module_57__and_module_2_res,
         n_majority7_module_57__or_module_1_res,
         n_majority7_module_57__and_module_1_res,
         n_majority7_module_58__and_module_10_res,
         n_majority7_module_58__or_module_11_res,
         n_majority7_module_58__and_module_9_res,
         n_majority7_module_58__or_module_10_res,
         n_majority7_module_58__or_module_9_res,
         n_majority7_module_58__and_module_8_res,
         n_majority7_module_58__or_module_8_res,
         n_majority7_module_58__and_module_7_res,
         n_majority7_module_58__or_module_7_res,
         n_majority7_module_58__or_module_6_res,
         n_majority7_module_58__and_module_6_res,
         n_majority7_module_58__or_module_5_res,
         n_majority7_module_58__and_module_5_res,
         n_majority7_module_58__or_module_4_res,
         n_majority7_module_58__and_module_4_res,
         n_majority7_module_58__or_module_3_res,
         n_majority7_module_58__and_module_3_res,
         n_majority7_module_58__or_module_2_res,
         n_majority7_module_58__and_module_2_res,
         n_majority7_module_58__or_module_1_res,
         n_majority7_module_58__and_module_1_res,
         n_majority7_module_59__and_module_10_res,
         n_majority7_module_59__or_module_11_res,
         n_majority7_module_59__and_module_9_res,
         n_majority7_module_59__or_module_10_res,
         n_majority7_module_59__or_module_9_res,
         n_majority7_module_59__and_module_8_res,
         n_majority7_module_59__or_module_8_res,
         n_majority7_module_59__and_module_7_res,
         n_majority7_module_59__or_module_7_res,
         n_majority7_module_59__or_module_6_res,
         n_majority7_module_59__and_module_6_res,
         n_majority7_module_59__or_module_5_res,
         n_majority7_module_59__and_module_5_res,
         n_majority7_module_59__or_module_4_res,
         n_majority7_module_59__and_module_4_res,
         n_majority7_module_59__or_module_3_res,
         n_majority7_module_59__and_module_3_res,
         n_majority7_module_59__or_module_2_res,
         n_majority7_module_59__and_module_2_res,
         n_majority7_module_59__or_module_1_res,
         n_majority7_module_59__and_module_1_res,
         n_majority7_module_60__and_module_10_res,
         n_majority7_module_60__or_module_11_res,
         n_majority7_module_60__and_module_9_res,
         n_majority7_module_60__or_module_10_res,
         n_majority7_module_60__or_module_9_res,
         n_majority7_module_60__and_module_8_res,
         n_majority7_module_60__or_module_8_res,
         n_majority7_module_60__and_module_7_res,
         n_majority7_module_60__or_module_7_res,
         n_majority7_module_60__or_module_6_res,
         n_majority7_module_60__and_module_6_res,
         n_majority7_module_60__or_module_5_res,
         n_majority7_module_60__and_module_5_res,
         n_majority7_module_60__or_module_4_res,
         n_majority7_module_60__and_module_4_res,
         n_majority7_module_60__or_module_3_res,
         n_majority7_module_60__and_module_3_res,
         n_majority7_module_60__or_module_2_res,
         n_majority7_module_60__and_module_2_res,
         n_majority7_module_60__or_module_1_res,
         n_majority7_module_60__and_module_1_res,
         n_majority7_module_61__and_module_10_res,
         n_majority7_module_61__or_module_11_res,
         n_majority7_module_61__and_module_9_res,
         n_majority7_module_61__or_module_10_res,
         n_majority7_module_61__or_module_9_res,
         n_majority7_module_61__and_module_8_res,
         n_majority7_module_61__or_module_8_res,
         n_majority7_module_61__and_module_7_res,
         n_majority7_module_61__or_module_7_res,
         n_majority7_module_61__or_module_6_res,
         n_majority7_module_61__and_module_6_res,
         n_majority7_module_61__or_module_5_res,
         n_majority7_module_61__and_module_5_res,
         n_majority7_module_61__or_module_4_res,
         n_majority7_module_61__and_module_4_res,
         n_majority7_module_61__or_module_3_res,
         n_majority7_module_61__and_module_3_res,
         n_majority7_module_61__or_module_2_res,
         n_majority7_module_61__and_module_2_res,
         n_majority7_module_61__or_module_1_res,
         n_majority7_module_61__and_module_1_res,
         n_majority7_module_62__and_module_10_res,
         n_majority7_module_62__or_module_11_res,
         n_majority7_module_62__and_module_9_res,
         n_majority7_module_62__or_module_10_res,
         n_majority7_module_62__or_module_9_res,
         n_majority7_module_62__and_module_8_res,
         n_majority7_module_62__or_module_8_res,
         n_majority7_module_62__and_module_7_res,
         n_majority7_module_62__or_module_7_res,
         n_majority7_module_62__or_module_6_res,
         n_majority7_module_62__and_module_6_res,
         n_majority7_module_62__or_module_5_res,
         n_majority7_module_62__and_module_5_res,
         n_majority7_module_62__or_module_4_res,
         n_majority7_module_62__and_module_4_res,
         n_majority7_module_62__or_module_3_res,
         n_majority7_module_62__and_module_3_res,
         n_majority7_module_62__or_module_2_res,
         n_majority7_module_62__and_module_2_res,
         n_majority7_module_62__or_module_1_res,
         n_majority7_module_62__and_module_1_res,
         n_majority7_module_63__and_module_10_res,
         n_majority7_module_63__or_module_11_res,
         n_majority7_module_63__and_module_9_res,
         n_majority7_module_63__or_module_10_res,
         n_majority7_module_63__or_module_9_res,
         n_majority7_module_63__and_module_8_res,
         n_majority7_module_63__or_module_8_res,
         n_majority7_module_63__and_module_7_res,
         n_majority7_module_63__or_module_7_res,
         n_majority7_module_63__or_module_6_res,
         n_majority7_module_63__and_module_6_res,
         n_majority7_module_63__or_module_5_res,
         n_majority7_module_63__and_module_5_res,
         n_majority7_module_63__or_module_4_res,
         n_majority7_module_63__and_module_4_res,
         n_majority7_module_63__or_module_3_res,
         n_majority7_module_63__and_module_3_res,
         n_majority7_module_63__or_module_2_res,
         n_majority7_module_63__and_module_2_res,
         n_majority7_module_63__or_module_1_res,
         n_majority7_module_63__and_module_1_res,
         n_majority7_module_64__and_module_10_res,
         n_majority7_module_64__or_module_11_res,
         n_majority7_module_64__and_module_9_res,
         n_majority7_module_64__or_module_10_res,
         n_majority7_module_64__or_module_9_res,
         n_majority7_module_64__and_module_8_res,
         n_majority7_module_64__or_module_8_res,
         n_majority7_module_64__and_module_7_res,
         n_majority7_module_64__or_module_7_res,
         n_majority7_module_64__or_module_6_res,
         n_majority7_module_64__and_module_6_res,
         n_majority7_module_64__or_module_5_res,
         n_majority7_module_64__and_module_5_res,
         n_majority7_module_64__or_module_4_res,
         n_majority7_module_64__and_module_4_res,
         n_majority7_module_64__or_module_3_res,
         n_majority7_module_64__and_module_3_res,
         n_majority7_module_64__or_module_2_res,
         n_majority7_module_64__and_module_2_res,
         n_majority7_module_64__or_module_1_res,
         n_majority7_module_64__and_module_1_res,
         n_majority7_module_65__and_module_10_res,
         n_majority7_module_65__or_module_11_res,
         n_majority7_module_65__and_module_9_res,
         n_majority7_module_65__or_module_10_res,
         n_majority7_module_65__or_module_9_res,
         n_majority7_module_65__and_module_8_res,
         n_majority7_module_65__or_module_8_res,
         n_majority7_module_65__and_module_7_res,
         n_majority7_module_65__or_module_7_res,
         n_majority7_module_65__or_module_6_res,
         n_majority7_module_65__and_module_6_res,
         n_majority7_module_65__or_module_5_res,
         n_majority7_module_65__and_module_5_res,
         n_majority7_module_65__or_module_4_res,
         n_majority7_module_65__and_module_4_res,
         n_majority7_module_65__or_module_3_res,
         n_majority7_module_65__and_module_3_res,
         n_majority7_module_65__or_module_2_res,
         n_majority7_module_65__and_module_2_res,
         n_majority7_module_65__or_module_1_res,
         n_majority7_module_65__and_module_1_res,
         n_majority7_module_66__and_module_10_res,
         n_majority7_module_66__or_module_11_res,
         n_majority7_module_66__and_module_9_res,
         n_majority7_module_66__or_module_10_res,
         n_majority7_module_66__or_module_9_res,
         n_majority7_module_66__and_module_8_res,
         n_majority7_module_66__or_module_8_res,
         n_majority7_module_66__and_module_7_res,
         n_majority7_module_66__or_module_7_res,
         n_majority7_module_66__or_module_6_res,
         n_majority7_module_66__and_module_6_res,
         n_majority7_module_66__or_module_5_res,
         n_majority7_module_66__and_module_5_res,
         n_majority7_module_66__or_module_4_res,
         n_majority7_module_66__and_module_4_res,
         n_majority7_module_66__or_module_3_res,
         n_majority7_module_66__and_module_3_res,
         n_majority7_module_66__or_module_2_res,
         n_majority7_module_66__and_module_2_res,
         n_majority7_module_66__or_module_1_res,
         n_majority7_module_66__and_module_1_res,
         n_majority7_module_67__and_module_10_res,
         n_majority7_module_67__or_module_11_res,
         n_majority7_module_67__and_module_9_res,
         n_majority7_module_67__or_module_10_res,
         n_majority7_module_67__or_module_9_res,
         n_majority7_module_67__and_module_8_res,
         n_majority7_module_67__or_module_8_res,
         n_majority7_module_67__and_module_7_res,
         n_majority7_module_67__or_module_7_res,
         n_majority7_module_67__or_module_6_res,
         n_majority7_module_67__and_module_6_res,
         n_majority7_module_67__or_module_5_res,
         n_majority7_module_67__and_module_5_res,
         n_majority7_module_67__or_module_4_res,
         n_majority7_module_67__and_module_4_res,
         n_majority7_module_67__or_module_3_res,
         n_majority7_module_67__and_module_3_res,
         n_majority7_module_67__or_module_2_res,
         n_majority7_module_67__and_module_2_res,
         n_majority7_module_67__or_module_1_res,
         n_majority7_module_67__and_module_1_res,
         n_majority7_module_68__and_module_10_res,
         n_majority7_module_68__or_module_11_res,
         n_majority7_module_68__and_module_9_res,
         n_majority7_module_68__or_module_10_res,
         n_majority7_module_68__or_module_9_res,
         n_majority7_module_68__and_module_8_res,
         n_majority7_module_68__or_module_8_res,
         n_majority7_module_68__and_module_7_res,
         n_majority7_module_68__or_module_7_res,
         n_majority7_module_68__or_module_6_res,
         n_majority7_module_68__and_module_6_res,
         n_majority7_module_68__or_module_5_res,
         n_majority7_module_68__and_module_5_res,
         n_majority7_module_68__or_module_4_res,
         n_majority7_module_68__and_module_4_res,
         n_majority7_module_68__or_module_3_res,
         n_majority7_module_68__and_module_3_res,
         n_majority7_module_68__or_module_2_res,
         n_majority7_module_68__and_module_2_res,
         n_majority7_module_68__or_module_1_res,
         n_majority7_module_68__and_module_1_res,
         n_majority7_module_69__and_module_10_res,
         n_majority7_module_69__or_module_11_res,
         n_majority7_module_69__and_module_9_res,
         n_majority7_module_69__or_module_10_res,
         n_majority7_module_69__or_module_9_res,
         n_majority7_module_69__and_module_8_res,
         n_majority7_module_69__or_module_8_res,
         n_majority7_module_69__and_module_7_res,
         n_majority7_module_69__or_module_7_res,
         n_majority7_module_69__or_module_6_res,
         n_majority7_module_69__and_module_6_res,
         n_majority7_module_69__or_module_5_res,
         n_majority7_module_69__and_module_5_res,
         n_majority7_module_69__or_module_4_res,
         n_majority7_module_69__and_module_4_res,
         n_majority7_module_69__or_module_3_res,
         n_majority7_module_69__and_module_3_res,
         n_majority7_module_69__or_module_2_res,
         n_majority7_module_69__and_module_2_res,
         n_majority7_module_69__or_module_1_res,
         n_majority7_module_69__and_module_1_res,
         n_majority7_module_70__and_module_10_res,
         n_majority7_module_70__or_module_11_res,
         n_majority7_module_70__and_module_9_res,
         n_majority7_module_70__or_module_10_res,
         n_majority7_module_70__or_module_9_res,
         n_majority7_module_70__and_module_8_res,
         n_majority7_module_70__or_module_8_res,
         n_majority7_module_70__and_module_7_res,
         n_majority7_module_70__or_module_7_res,
         n_majority7_module_70__or_module_6_res,
         n_majority7_module_70__and_module_6_res,
         n_majority7_module_70__or_module_5_res,
         n_majority7_module_70__and_module_5_res,
         n_majority7_module_70__or_module_4_res,
         n_majority7_module_70__and_module_4_res,
         n_majority7_module_70__or_module_3_res,
         n_majority7_module_70__and_module_3_res,
         n_majority7_module_70__or_module_2_res,
         n_majority7_module_70__and_module_2_res,
         n_majority7_module_70__or_module_1_res,
         n_majority7_module_70__and_module_1_res,
         n_majority7_module_71__and_module_10_res,
         n_majority7_module_71__or_module_11_res,
         n_majority7_module_71__and_module_9_res,
         n_majority7_module_71__or_module_10_res,
         n_majority7_module_71__or_module_9_res,
         n_majority7_module_71__and_module_8_res,
         n_majority7_module_71__or_module_8_res,
         n_majority7_module_71__and_module_7_res,
         n_majority7_module_71__or_module_7_res,
         n_majority7_module_71__or_module_6_res,
         n_majority7_module_71__and_module_6_res,
         n_majority7_module_71__or_module_5_res,
         n_majority7_module_71__and_module_5_res,
         n_majority7_module_71__or_module_4_res,
         n_majority7_module_71__and_module_4_res,
         n_majority7_module_71__or_module_3_res,
         n_majority7_module_71__and_module_3_res,
         n_majority7_module_71__or_module_2_res,
         n_majority7_module_71__and_module_2_res,
         n_majority7_module_71__or_module_1_res,
         n_majority7_module_71__and_module_1_res,
         n_majority7_module_72__and_module_10_res,
         n_majority7_module_72__or_module_11_res,
         n_majority7_module_72__and_module_9_res,
         n_majority7_module_72__or_module_10_res,
         n_majority7_module_72__or_module_9_res,
         n_majority7_module_72__and_module_8_res,
         n_majority7_module_72__or_module_8_res,
         n_majority7_module_72__and_module_7_res,
         n_majority7_module_72__or_module_7_res,
         n_majority7_module_72__or_module_6_res,
         n_majority7_module_72__and_module_6_res,
         n_majority7_module_72__or_module_5_res,
         n_majority7_module_72__and_module_5_res,
         n_majority7_module_72__or_module_4_res,
         n_majority7_module_72__and_module_4_res,
         n_majority7_module_72__or_module_3_res,
         n_majority7_module_72__and_module_3_res,
         n_majority7_module_72__or_module_2_res,
         n_majority7_module_72__and_module_2_res,
         n_majority7_module_72__or_module_1_res,
         n_majority7_module_72__and_module_1_res,
         n_majority7_module_73__and_module_10_res,
         n_majority7_module_73__or_module_11_res,
         n_majority7_module_73__and_module_9_res,
         n_majority7_module_73__or_module_10_res,
         n_majority7_module_73__or_module_9_res,
         n_majority7_module_73__and_module_8_res,
         n_majority7_module_73__or_module_8_res,
         n_majority7_module_73__and_module_7_res,
         n_majority7_module_73__or_module_7_res,
         n_majority7_module_73__or_module_6_res,
         n_majority7_module_73__and_module_6_res,
         n_majority7_module_73__or_module_5_res,
         n_majority7_module_73__and_module_5_res,
         n_majority7_module_73__or_module_4_res,
         n_majority7_module_73__and_module_4_res,
         n_majority7_module_73__or_module_3_res,
         n_majority7_module_73__and_module_3_res,
         n_majority7_module_73__or_module_2_res,
         n_majority7_module_73__and_module_2_res,
         n_majority7_module_73__or_module_1_res,
         n_majority7_module_73__and_module_1_res,
         n_majority7_module_74__and_module_10_res,
         n_majority7_module_74__or_module_11_res,
         n_majority7_module_74__and_module_9_res,
         n_majority7_module_74__or_module_10_res,
         n_majority7_module_74__or_module_9_res,
         n_majority7_module_74__and_module_8_res,
         n_majority7_module_74__or_module_8_res,
         n_majority7_module_74__and_module_7_res,
         n_majority7_module_74__or_module_7_res,
         n_majority7_module_74__or_module_6_res,
         n_majority7_module_74__and_module_6_res,
         n_majority7_module_74__or_module_5_res,
         n_majority7_module_74__and_module_5_res,
         n_majority7_module_74__or_module_4_res,
         n_majority7_module_74__and_module_4_res,
         n_majority7_module_74__or_module_3_res,
         n_majority7_module_74__and_module_3_res,
         n_majority7_module_74__or_module_2_res,
         n_majority7_module_74__and_module_2_res,
         n_majority7_module_74__or_module_1_res,
         n_majority7_module_74__and_module_1_res,
         n_majority7_module_75__and_module_10_res,
         n_majority7_module_75__or_module_11_res,
         n_majority7_module_75__and_module_9_res,
         n_majority7_module_75__or_module_10_res,
         n_majority7_module_75__or_module_9_res,
         n_majority7_module_75__and_module_8_res,
         n_majority7_module_75__or_module_8_res,
         n_majority7_module_75__and_module_7_res,
         n_majority7_module_75__or_module_7_res,
         n_majority7_module_75__or_module_6_res,
         n_majority7_module_75__and_module_6_res,
         n_majority7_module_75__or_module_5_res,
         n_majority7_module_75__and_module_5_res,
         n_majority7_module_75__or_module_4_res,
         n_majority7_module_75__and_module_4_res,
         n_majority7_module_75__or_module_3_res,
         n_majority7_module_75__and_module_3_res,
         n_majority7_module_75__or_module_2_res,
         n_majority7_module_75__and_module_2_res,
         n_majority7_module_75__or_module_1_res,
         n_majority7_module_75__and_module_1_res,
         n_majority7_module_76__and_module_10_res,
         n_majority7_module_76__or_module_11_res,
         n_majority7_module_76__and_module_9_res,
         n_majority7_module_76__or_module_10_res,
         n_majority7_module_76__or_module_9_res,
         n_majority7_module_76__and_module_8_res,
         n_majority7_module_76__or_module_8_res,
         n_majority7_module_76__and_module_7_res,
         n_majority7_module_76__or_module_7_res,
         n_majority7_module_76__or_module_6_res,
         n_majority7_module_76__and_module_6_res,
         n_majority7_module_76__or_module_5_res,
         n_majority7_module_76__and_module_5_res,
         n_majority7_module_76__or_module_4_res,
         n_majority7_module_76__and_module_4_res,
         n_majority7_module_76__or_module_3_res,
         n_majority7_module_76__and_module_3_res,
         n_majority7_module_76__or_module_2_res,
         n_majority7_module_76__and_module_2_res,
         n_majority7_module_76__or_module_1_res,
         n_majority7_module_76__and_module_1_res,
         n_majority7_module_77__and_module_10_res,
         n_majority7_module_77__or_module_11_res,
         n_majority7_module_77__and_module_9_res,
         n_majority7_module_77__or_module_10_res,
         n_majority7_module_77__or_module_9_res,
         n_majority7_module_77__and_module_8_res,
         n_majority7_module_77__or_module_8_res,
         n_majority7_module_77__and_module_7_res,
         n_majority7_module_77__or_module_7_res,
         n_majority7_module_77__or_module_6_res,
         n_majority7_module_77__and_module_6_res,
         n_majority7_module_77__or_module_5_res,
         n_majority7_module_77__and_module_5_res,
         n_majority7_module_77__or_module_4_res,
         n_majority7_module_77__and_module_4_res,
         n_majority7_module_77__or_module_3_res,
         n_majority7_module_77__and_module_3_res,
         n_majority7_module_77__or_module_2_res,
         n_majority7_module_77__and_module_2_res,
         n_majority7_module_77__or_module_1_res,
         n_majority7_module_77__and_module_1_res,
         n_majority7_module_78__and_module_10_res,
         n_majority7_module_78__or_module_11_res,
         n_majority7_module_78__and_module_9_res,
         n_majority7_module_78__or_module_10_res,
         n_majority7_module_78__or_module_9_res,
         n_majority7_module_78__and_module_8_res,
         n_majority7_module_78__or_module_8_res,
         n_majority7_module_78__and_module_7_res,
         n_majority7_module_78__or_module_7_res,
         n_majority7_module_78__or_module_6_res,
         n_majority7_module_78__and_module_6_res,
         n_majority7_module_78__or_module_5_res,
         n_majority7_module_78__and_module_5_res,
         n_majority7_module_78__or_module_4_res,
         n_majority7_module_78__and_module_4_res,
         n_majority7_module_78__or_module_3_res,
         n_majority7_module_78__and_module_3_res,
         n_majority7_module_78__or_module_2_res,
         n_majority7_module_78__and_module_2_res,
         n_majority7_module_78__or_module_1_res,
         n_majority7_module_78__and_module_1_res,
         n_majority7_module_79__and_module_10_res,
         n_majority7_module_79__or_module_11_res,
         n_majority7_module_79__and_module_9_res,
         n_majority7_module_79__or_module_10_res,
         n_majority7_module_79__or_module_9_res,
         n_majority7_module_79__and_module_8_res,
         n_majority7_module_79__or_module_8_res,
         n_majority7_module_79__and_module_7_res,
         n_majority7_module_79__or_module_7_res,
         n_majority7_module_79__or_module_6_res,
         n_majority7_module_79__and_module_6_res,
         n_majority7_module_79__or_module_5_res,
         n_majority7_module_79__and_module_5_res,
         n_majority7_module_79__or_module_4_res,
         n_majority7_module_79__and_module_4_res,
         n_majority7_module_79__or_module_3_res,
         n_majority7_module_79__and_module_3_res,
         n_majority7_module_79__or_module_2_res,
         n_majority7_module_79__and_module_2_res,
         n_majority7_module_79__or_module_1_res,
         n_majority7_module_79__and_module_1_res,
         n_majority7_module_80__and_module_10_res,
         n_majority7_module_80__or_module_11_res,
         n_majority7_module_80__and_module_9_res,
         n_majority7_module_80__or_module_10_res,
         n_majority7_module_80__or_module_9_res,
         n_majority7_module_80__and_module_8_res,
         n_majority7_module_80__or_module_8_res,
         n_majority7_module_80__and_module_7_res,
         n_majority7_module_80__or_module_7_res,
         n_majority7_module_80__or_module_6_res,
         n_majority7_module_80__and_module_6_res,
         n_majority7_module_80__or_module_5_res,
         n_majority7_module_80__and_module_5_res,
         n_majority7_module_80__or_module_4_res,
         n_majority7_module_80__and_module_4_res,
         n_majority7_module_80__or_module_3_res,
         n_majority7_module_80__and_module_3_res,
         n_majority7_module_80__or_module_2_res,
         n_majority7_module_80__and_module_2_res,
         n_majority7_module_80__or_module_1_res,
         n_majority7_module_80__and_module_1_res,
         n_majority7_module_81__and_module_10_res,
         n_majority7_module_81__or_module_11_res,
         n_majority7_module_81__and_module_9_res,
         n_majority7_module_81__or_module_10_res,
         n_majority7_module_81__or_module_9_res,
         n_majority7_module_81__and_module_8_res,
         n_majority7_module_81__or_module_8_res,
         n_majority7_module_81__and_module_7_res,
         n_majority7_module_81__or_module_7_res,
         n_majority7_module_81__or_module_6_res,
         n_majority7_module_81__and_module_6_res,
         n_majority7_module_81__or_module_5_res,
         n_majority7_module_81__and_module_5_res,
         n_majority7_module_81__or_module_4_res,
         n_majority7_module_81__and_module_4_res,
         n_majority7_module_81__or_module_3_res,
         n_majority7_module_81__and_module_3_res,
         n_majority7_module_81__or_module_2_res,
         n_majority7_module_81__and_module_2_res,
         n_majority7_module_81__or_module_1_res,
         n_majority7_module_81__and_module_1_res,
         n_majority7_module_82__and_module_10_res,
         n_majority7_module_82__or_module_11_res,
         n_majority7_module_82__and_module_9_res,
         n_majority7_module_82__or_module_10_res,
         n_majority7_module_82__or_module_9_res,
         n_majority7_module_82__and_module_8_res,
         n_majority7_module_82__or_module_8_res,
         n_majority7_module_82__and_module_7_res,
         n_majority7_module_82__or_module_7_res,
         n_majority7_module_82__or_module_6_res,
         n_majority7_module_82__and_module_6_res,
         n_majority7_module_82__or_module_5_res,
         n_majority7_module_82__and_module_5_res,
         n_majority7_module_82__or_module_4_res,
         n_majority7_module_82__and_module_4_res,
         n_majority7_module_82__or_module_3_res,
         n_majority7_module_82__and_module_3_res,
         n_majority7_module_82__or_module_2_res,
         n_majority7_module_82__and_module_2_res,
         n_majority7_module_82__or_module_1_res,
         n_majority7_module_82__and_module_1_res,
         n_majority7_module_83__and_module_10_res,
         n_majority7_module_83__or_module_11_res,
         n_majority7_module_83__and_module_9_res,
         n_majority7_module_83__or_module_10_res,
         n_majority7_module_83__or_module_9_res,
         n_majority7_module_83__and_module_8_res,
         n_majority7_module_83__or_module_8_res,
         n_majority7_module_83__and_module_7_res,
         n_majority7_module_83__or_module_7_res,
         n_majority7_module_83__or_module_6_res,
         n_majority7_module_83__and_module_6_res,
         n_majority7_module_83__or_module_5_res,
         n_majority7_module_83__and_module_5_res,
         n_majority7_module_83__or_module_4_res,
         n_majority7_module_83__and_module_4_res,
         n_majority7_module_83__or_module_3_res,
         n_majority7_module_83__and_module_3_res,
         n_majority7_module_83__or_module_2_res,
         n_majority7_module_83__and_module_2_res,
         n_majority7_module_83__or_module_1_res,
         n_majority7_module_83__and_module_1_res,
         n_majority7_module_84__and_module_10_res,
         n_majority7_module_84__or_module_11_res,
         n_majority7_module_84__and_module_9_res,
         n_majority7_module_84__or_module_10_res,
         n_majority7_module_84__or_module_9_res,
         n_majority7_module_84__and_module_8_res,
         n_majority7_module_84__or_module_8_res,
         n_majority7_module_84__and_module_7_res,
         n_majority7_module_84__or_module_7_res,
         n_majority7_module_84__or_module_6_res,
         n_majority7_module_84__and_module_6_res,
         n_majority7_module_84__or_module_5_res,
         n_majority7_module_84__and_module_5_res,
         n_majority7_module_84__or_module_4_res,
         n_majority7_module_84__and_module_4_res,
         n_majority7_module_84__or_module_3_res,
         n_majority7_module_84__and_module_3_res,
         n_majority7_module_84__or_module_2_res,
         n_majority7_module_84__and_module_2_res,
         n_majority7_module_84__or_module_1_res,
         n_majority7_module_84__and_module_1_res,
         n_majority7_module_85__and_module_10_res,
         n_majority7_module_85__or_module_11_res,
         n_majority7_module_85__and_module_9_res,
         n_majority7_module_85__or_module_10_res,
         n_majority7_module_85__or_module_9_res,
         n_majority7_module_85__and_module_8_res,
         n_majority7_module_85__or_module_8_res,
         n_majority7_module_85__and_module_7_res,
         n_majority7_module_85__or_module_7_res,
         n_majority7_module_85__or_module_6_res,
         n_majority7_module_85__and_module_6_res,
         n_majority7_module_85__or_module_5_res,
         n_majority7_module_85__and_module_5_res,
         n_majority7_module_85__or_module_4_res,
         n_majority7_module_85__and_module_4_res,
         n_majority7_module_85__or_module_3_res,
         n_majority7_module_85__and_module_3_res,
         n_majority7_module_85__or_module_2_res,
         n_majority7_module_85__and_module_2_res,
         n_majority7_module_85__or_module_1_res,
         n_majority7_module_85__and_module_1_res,
         n_majority7_module_86__and_module_10_res,
         n_majority7_module_86__or_module_11_res,
         n_majority7_module_86__and_module_9_res,
         n_majority7_module_86__or_module_10_res,
         n_majority7_module_86__or_module_9_res,
         n_majority7_module_86__and_module_8_res,
         n_majority7_module_86__or_module_8_res,
         n_majority7_module_86__and_module_7_res,
         n_majority7_module_86__or_module_7_res,
         n_majority7_module_86__or_module_6_res,
         n_majority7_module_86__and_module_6_res,
         n_majority7_module_86__or_module_5_res,
         n_majority7_module_86__and_module_5_res,
         n_majority7_module_86__or_module_4_res,
         n_majority7_module_86__and_module_4_res,
         n_majority7_module_86__or_module_3_res,
         n_majority7_module_86__and_module_3_res,
         n_majority7_module_86__or_module_2_res,
         n_majority7_module_86__and_module_2_res,
         n_majority7_module_86__or_module_1_res,
         n_majority7_module_86__and_module_1_res,
         n_majority7_module_87__and_module_10_res,
         n_majority7_module_87__or_module_11_res,
         n_majority7_module_87__and_module_9_res,
         n_majority7_module_87__or_module_10_res,
         n_majority7_module_87__or_module_9_res,
         n_majority7_module_87__and_module_8_res,
         n_majority7_module_87__or_module_8_res,
         n_majority7_module_87__and_module_7_res,
         n_majority7_module_87__or_module_7_res,
         n_majority7_module_87__or_module_6_res,
         n_majority7_module_87__and_module_6_res,
         n_majority7_module_87__or_module_5_res,
         n_majority7_module_87__and_module_5_res,
         n_majority7_module_87__or_module_4_res,
         n_majority7_module_87__and_module_4_res,
         n_majority7_module_87__or_module_3_res,
         n_majority7_module_87__and_module_3_res,
         n_majority7_module_87__or_module_2_res,
         n_majority7_module_87__and_module_2_res,
         n_majority7_module_87__or_module_1_res,
         n_majority7_module_87__and_module_1_res,
         n_majority7_module_88__and_module_10_res,
         n_majority7_module_88__or_module_11_res,
         n_majority7_module_88__and_module_9_res,
         n_majority7_module_88__or_module_10_res,
         n_majority7_module_88__or_module_9_res,
         n_majority7_module_88__and_module_8_res,
         n_majority7_module_88__or_module_8_res,
         n_majority7_module_88__and_module_7_res,
         n_majority7_module_88__or_module_7_res,
         n_majority7_module_88__or_module_6_res,
         n_majority7_module_88__and_module_6_res,
         n_majority7_module_88__or_module_5_res,
         n_majority7_module_88__and_module_5_res,
         n_majority7_module_88__or_module_4_res,
         n_majority7_module_88__and_module_4_res,
         n_majority7_module_88__or_module_3_res,
         n_majority7_module_88__and_module_3_res,
         n_majority7_module_88__or_module_2_res,
         n_majority7_module_88__and_module_2_res,
         n_majority7_module_88__or_module_1_res,
         n_majority7_module_88__and_module_1_res,
         n_majority7_module_89__and_module_10_res,
         n_majority7_module_89__or_module_11_res,
         n_majority7_module_89__and_module_9_res,
         n_majority7_module_89__or_module_10_res,
         n_majority7_module_89__or_module_9_res,
         n_majority7_module_89__and_module_8_res,
         n_majority7_module_89__or_module_8_res,
         n_majority7_module_89__and_module_7_res,
         n_majority7_module_89__or_module_7_res,
         n_majority7_module_89__or_module_6_res,
         n_majority7_module_89__and_module_6_res,
         n_majority7_module_89__or_module_5_res,
         n_majority7_module_89__and_module_5_res,
         n_majority7_module_89__or_module_4_res,
         n_majority7_module_89__and_module_4_res,
         n_majority7_module_89__or_module_3_res,
         n_majority7_module_89__and_module_3_res,
         n_majority7_module_89__or_module_2_res,
         n_majority7_module_89__and_module_2_res,
         n_majority7_module_89__or_module_1_res,
         n_majority7_module_89__and_module_1_res,
         n_majority7_module_90__and_module_10_res,
         n_majority7_module_90__or_module_11_res,
         n_majority7_module_90__and_module_9_res,
         n_majority7_module_90__or_module_10_res,
         n_majority7_module_90__or_module_9_res,
         n_majority7_module_90__and_module_8_res,
         n_majority7_module_90__or_module_8_res,
         n_majority7_module_90__and_module_7_res,
         n_majority7_module_90__or_module_7_res,
         n_majority7_module_90__or_module_6_res,
         n_majority7_module_90__and_module_6_res,
         n_majority7_module_90__or_module_5_res,
         n_majority7_module_90__and_module_5_res,
         n_majority7_module_90__or_module_4_res,
         n_majority7_module_90__and_module_4_res,
         n_majority7_module_90__or_module_3_res,
         n_majority7_module_90__and_module_3_res,
         n_majority7_module_90__or_module_2_res,
         n_majority7_module_90__and_module_2_res,
         n_majority7_module_90__or_module_1_res,
         n_majority7_module_90__and_module_1_res,
         n_majority7_module_91__and_module_10_res,
         n_majority7_module_91__or_module_11_res,
         n_majority7_module_91__and_module_9_res,
         n_majority7_module_91__or_module_10_res,
         n_majority7_module_91__or_module_9_res,
         n_majority7_module_91__and_module_8_res,
         n_majority7_module_91__or_module_8_res,
         n_majority7_module_91__and_module_7_res,
         n_majority7_module_91__or_module_7_res,
         n_majority7_module_91__or_module_6_res,
         n_majority7_module_91__and_module_6_res,
         n_majority7_module_91__or_module_5_res,
         n_majority7_module_91__and_module_5_res,
         n_majority7_module_91__or_module_4_res,
         n_majority7_module_91__and_module_4_res,
         n_majority7_module_91__or_module_3_res,
         n_majority7_module_91__and_module_3_res,
         n_majority7_module_91__or_module_2_res,
         n_majority7_module_91__and_module_2_res,
         n_majority7_module_91__or_module_1_res,
         n_majority7_module_91__and_module_1_res,
         n_majority7_module_92__and_module_10_res,
         n_majority7_module_92__or_module_11_res,
         n_majority7_module_92__and_module_9_res,
         n_majority7_module_92__or_module_10_res,
         n_majority7_module_92__or_module_9_res,
         n_majority7_module_92__and_module_8_res,
         n_majority7_module_92__or_module_8_res,
         n_majority7_module_92__and_module_7_res,
         n_majority7_module_92__or_module_7_res,
         n_majority7_module_92__or_module_6_res,
         n_majority7_module_92__and_module_6_res,
         n_majority7_module_92__or_module_5_res,
         n_majority7_module_92__and_module_5_res,
         n_majority7_module_92__or_module_4_res,
         n_majority7_module_92__and_module_4_res,
         n_majority7_module_92__or_module_3_res,
         n_majority7_module_92__and_module_3_res,
         n_majority7_module_92__or_module_2_res,
         n_majority7_module_92__and_module_2_res,
         n_majority7_module_92__or_module_1_res,
         n_majority7_module_92__and_module_1_res,
         n_majority7_module_93__and_module_10_res,
         n_majority7_module_93__or_module_11_res,
         n_majority7_module_93__and_module_9_res,
         n_majority7_module_93__or_module_10_res,
         n_majority7_module_93__or_module_9_res,
         n_majority7_module_93__and_module_8_res,
         n_majority7_module_93__or_module_8_res,
         n_majority7_module_93__and_module_7_res,
         n_majority7_module_93__or_module_7_res,
         n_majority7_module_93__or_module_6_res,
         n_majority7_module_93__and_module_6_res,
         n_majority7_module_93__or_module_5_res,
         n_majority7_module_93__and_module_5_res,
         n_majority7_module_93__or_module_4_res,
         n_majority7_module_93__and_module_4_res,
         n_majority7_module_93__or_module_3_res,
         n_majority7_module_93__and_module_3_res,
         n_majority7_module_93__or_module_2_res,
         n_majority7_module_93__and_module_2_res,
         n_majority7_module_93__or_module_1_res,
         n_majority7_module_93__and_module_1_res,
         n_majority7_module_94__and_module_10_res,
         n_majority7_module_94__or_module_11_res,
         n_majority7_module_94__and_module_9_res,
         n_majority7_module_94__or_module_10_res,
         n_majority7_module_94__or_module_9_res,
         n_majority7_module_94__and_module_8_res,
         n_majority7_module_94__or_module_8_res,
         n_majority7_module_94__and_module_7_res,
         n_majority7_module_94__or_module_7_res,
         n_majority7_module_94__or_module_6_res,
         n_majority7_module_94__and_module_6_res,
         n_majority7_module_94__or_module_5_res,
         n_majority7_module_94__and_module_5_res,
         n_majority7_module_94__or_module_4_res,
         n_majority7_module_94__and_module_4_res,
         n_majority7_module_94__or_module_3_res,
         n_majority7_module_94__and_module_3_res,
         n_majority7_module_94__or_module_2_res,
         n_majority7_module_94__and_module_2_res,
         n_majority7_module_94__or_module_1_res,
         n_majority7_module_94__and_module_1_res,
         n_majority7_module_95__and_module_10_res,
         n_majority7_module_95__or_module_11_res,
         n_majority7_module_95__and_module_9_res,
         n_majority7_module_95__or_module_10_res,
         n_majority7_module_95__or_module_9_res,
         n_majority7_module_95__and_module_8_res,
         n_majority7_module_95__or_module_8_res,
         n_majority7_module_95__and_module_7_res,
         n_majority7_module_95__or_module_7_res,
         n_majority7_module_95__or_module_6_res,
         n_majority7_module_95__and_module_6_res,
         n_majority7_module_95__or_module_5_res,
         n_majority7_module_95__and_module_5_res,
         n_majority7_module_95__or_module_4_res,
         n_majority7_module_95__and_module_4_res,
         n_majority7_module_95__or_module_3_res,
         n_majority7_module_95__and_module_3_res,
         n_majority7_module_95__or_module_2_res,
         n_majority7_module_95__and_module_2_res,
         n_majority7_module_95__or_module_1_res,
         n_majority7_module_95__and_module_1_res,
         n_majority7_module_96__and_module_10_res,
         n_majority7_module_96__or_module_11_res,
         n_majority7_module_96__and_module_9_res,
         n_majority7_module_96__or_module_10_res,
         n_majority7_module_96__or_module_9_res,
         n_majority7_module_96__and_module_8_res,
         n_majority7_module_96__or_module_8_res,
         n_majority7_module_96__and_module_7_res,
         n_majority7_module_96__or_module_7_res,
         n_majority7_module_96__or_module_6_res,
         n_majority7_module_96__and_module_6_res,
         n_majority7_module_96__or_module_5_res,
         n_majority7_module_96__and_module_5_res,
         n_majority7_module_96__or_module_4_res,
         n_majority7_module_96__and_module_4_res,
         n_majority7_module_96__or_module_3_res,
         n_majority7_module_96__and_module_3_res,
         n_majority7_module_96__or_module_2_res,
         n_majority7_module_96__and_module_2_res,
         n_majority7_module_96__or_module_1_res,
         n_majority7_module_96__and_module_1_res,
         n_majority7_module_97__and_module_10_res,
         n_majority7_module_97__or_module_11_res,
         n_majority7_module_97__and_module_9_res,
         n_majority7_module_97__or_module_10_res,
         n_majority7_module_97__or_module_9_res,
         n_majority7_module_97__and_module_8_res,
         n_majority7_module_97__or_module_8_res,
         n_majority7_module_97__and_module_7_res,
         n_majority7_module_97__or_module_7_res,
         n_majority7_module_97__or_module_6_res,
         n_majority7_module_97__and_module_6_res,
         n_majority7_module_97__or_module_5_res,
         n_majority7_module_97__and_module_5_res,
         n_majority7_module_97__or_module_4_res,
         n_majority7_module_97__and_module_4_res,
         n_majority7_module_97__or_module_3_res,
         n_majority7_module_97__and_module_3_res,
         n_majority7_module_97__or_module_2_res,
         n_majority7_module_97__and_module_2_res,
         n_majority7_module_97__or_module_1_res,
         n_majority7_module_97__and_module_1_res,
         n_majority7_module_98__and_module_10_res,
         n_majority7_module_98__or_module_11_res,
         n_majority7_module_98__and_module_9_res,
         n_majority7_module_98__or_module_10_res,
         n_majority7_module_98__or_module_9_res,
         n_majority7_module_98__and_module_8_res,
         n_majority7_module_98__or_module_8_res,
         n_majority7_module_98__and_module_7_res,
         n_majority7_module_98__or_module_7_res,
         n_majority7_module_98__or_module_6_res,
         n_majority7_module_98__and_module_6_res,
         n_majority7_module_98__or_module_5_res,
         n_majority7_module_98__and_module_5_res,
         n_majority7_module_98__or_module_4_res,
         n_majority7_module_98__and_module_4_res,
         n_majority7_module_98__or_module_3_res,
         n_majority7_module_98__and_module_3_res,
         n_majority7_module_98__or_module_2_res,
         n_majority7_module_98__and_module_2_res,
         n_majority7_module_98__or_module_1_res,
         n_majority7_module_98__and_module_1_res,
         n_majority7_module_99__and_module_10_res,
         n_majority7_module_99__or_module_11_res,
         n_majority7_module_99__and_module_9_res,
         n_majority7_module_99__or_module_10_res,
         n_majority7_module_99__or_module_9_res,
         n_majority7_module_99__and_module_8_res,
         n_majority7_module_99__or_module_8_res,
         n_majority7_module_99__and_module_7_res,
         n_majority7_module_99__or_module_7_res,
         n_majority7_module_99__or_module_6_res,
         n_majority7_module_99__and_module_6_res,
         n_majority7_module_99__or_module_5_res,
         n_majority7_module_99__and_module_5_res,
         n_majority7_module_99__or_module_4_res,
         n_majority7_module_99__and_module_4_res,
         n_majority7_module_99__or_module_3_res,
         n_majority7_module_99__and_module_3_res,
         n_majority7_module_99__or_module_2_res,
         n_majority7_module_99__and_module_2_res,
         n_majority7_module_99__or_module_1_res,
         n_majority7_module_99__and_module_1_res,
         n_majority7_module_100__and_module_10_res,
         n_majority7_module_100__or_module_11_res,
         n_majority7_module_100__and_module_9_res,
         n_majority7_module_100__or_module_10_res,
         n_majority7_module_100__or_module_9_res,
         n_majority7_module_100__and_module_8_res,
         n_majority7_module_100__or_module_8_res,
         n_majority7_module_100__and_module_7_res,
         n_majority7_module_100__or_module_7_res,
         n_majority7_module_100__or_module_6_res,
         n_majority7_module_100__and_module_6_res,
         n_majority7_module_100__or_module_5_res,
         n_majority7_module_100__and_module_5_res,
         n_majority7_module_100__or_module_4_res,
         n_majority7_module_100__and_module_4_res,
         n_majority7_module_100__or_module_3_res,
         n_majority7_module_100__and_module_3_res,
         n_majority7_module_100__or_module_2_res,
         n_majority7_module_100__and_module_2_res,
         n_majority7_module_100__or_module_1_res,
         n_majority7_module_100__and_module_1_res,
         n_majority7_module_101__and_module_10_res,
         n_majority7_module_101__or_module_11_res,
         n_majority7_module_101__and_module_9_res,
         n_majority7_module_101__or_module_10_res,
         n_majority7_module_101__or_module_9_res,
         n_majority7_module_101__and_module_8_res,
         n_majority7_module_101__or_module_8_res,
         n_majority7_module_101__and_module_7_res,
         n_majority7_module_101__or_module_7_res,
         n_majority7_module_101__or_module_6_res,
         n_majority7_module_101__and_module_6_res,
         n_majority7_module_101__or_module_5_res,
         n_majority7_module_101__and_module_5_res,
         n_majority7_module_101__or_module_4_res,
         n_majority7_module_101__and_module_4_res,
         n_majority7_module_101__or_module_3_res,
         n_majority7_module_101__and_module_3_res,
         n_majority7_module_101__or_module_2_res,
         n_majority7_module_101__and_module_2_res,
         n_majority7_module_101__or_module_1_res,
         n_majority7_module_101__and_module_1_res,
         n_majority7_module_102__and_module_10_res,
         n_majority7_module_102__or_module_11_res,
         n_majority7_module_102__and_module_9_res,
         n_majority7_module_102__or_module_10_res,
         n_majority7_module_102__or_module_9_res,
         n_majority7_module_102__and_module_8_res,
         n_majority7_module_102__or_module_8_res,
         n_majority7_module_102__and_module_7_res,
         n_majority7_module_102__or_module_7_res,
         n_majority7_module_102__or_module_6_res,
         n_majority7_module_102__and_module_6_res,
         n_majority7_module_102__or_module_5_res,
         n_majority7_module_102__and_module_5_res,
         n_majority7_module_102__or_module_4_res,
         n_majority7_module_102__and_module_4_res,
         n_majority7_module_102__or_module_3_res,
         n_majority7_module_102__and_module_3_res,
         n_majority7_module_102__or_module_2_res,
         n_majority7_module_102__and_module_2_res,
         n_majority7_module_102__or_module_1_res,
         n_majority7_module_102__and_module_1_res,
         n_majority7_module_103__and_module_10_res,
         n_majority7_module_103__or_module_11_res,
         n_majority7_module_103__and_module_9_res,
         n_majority7_module_103__or_module_10_res,
         n_majority7_module_103__or_module_9_res,
         n_majority7_module_103__and_module_8_res,
         n_majority7_module_103__or_module_8_res,
         n_majority7_module_103__and_module_7_res,
         n_majority7_module_103__or_module_7_res,
         n_majority7_module_103__or_module_6_res,
         n_majority7_module_103__and_module_6_res,
         n_majority7_module_103__or_module_5_res,
         n_majority7_module_103__and_module_5_res,
         n_majority7_module_103__or_module_4_res,
         n_majority7_module_103__and_module_4_res,
         n_majority7_module_103__or_module_3_res,
         n_majority7_module_103__and_module_3_res,
         n_majority7_module_103__or_module_2_res,
         n_majority7_module_103__and_module_2_res,
         n_majority7_module_103__or_module_1_res,
         n_majority7_module_103__and_module_1_res,
         n_majority7_module_104__and_module_10_res,
         n_majority7_module_104__or_module_11_res,
         n_majority7_module_104__and_module_9_res,
         n_majority7_module_104__or_module_10_res,
         n_majority7_module_104__or_module_9_res,
         n_majority7_module_104__and_module_8_res,
         n_majority7_module_104__or_module_8_res,
         n_majority7_module_104__and_module_7_res,
         n_majority7_module_104__or_module_7_res,
         n_majority7_module_104__or_module_6_res,
         n_majority7_module_104__and_module_6_res,
         n_majority7_module_104__or_module_5_res,
         n_majority7_module_104__and_module_5_res,
         n_majority7_module_104__or_module_4_res,
         n_majority7_module_104__and_module_4_res,
         n_majority7_module_104__or_module_3_res,
         n_majority7_module_104__and_module_3_res,
         n_majority7_module_104__or_module_2_res,
         n_majority7_module_104__and_module_2_res,
         n_majority7_module_104__or_module_1_res,
         n_majority7_module_104__and_module_1_res,
         n_majority7_module_105__and_module_10_res,
         n_majority7_module_105__or_module_11_res,
         n_majority7_module_105__and_module_9_res,
         n_majority7_module_105__or_module_10_res,
         n_majority7_module_105__or_module_9_res,
         n_majority7_module_105__and_module_8_res,
         n_majority7_module_105__or_module_8_res,
         n_majority7_module_105__and_module_7_res,
         n_majority7_module_105__or_module_7_res,
         n_majority7_module_105__or_module_6_res,
         n_majority7_module_105__and_module_6_res,
         n_majority7_module_105__or_module_5_res,
         n_majority7_module_105__and_module_5_res,
         n_majority7_module_105__or_module_4_res,
         n_majority7_module_105__and_module_4_res,
         n_majority7_module_105__or_module_3_res,
         n_majority7_module_105__and_module_3_res,
         n_majority7_module_105__or_module_2_res,
         n_majority7_module_105__and_module_2_res,
         n_majority7_module_105__or_module_1_res,
         n_majority7_module_105__and_module_1_res,
         n_majority7_module_106__and_module_10_res,
         n_majority7_module_106__or_module_11_res,
         n_majority7_module_106__and_module_9_res,
         n_majority7_module_106__or_module_10_res,
         n_majority7_module_106__or_module_9_res,
         n_majority7_module_106__and_module_8_res,
         n_majority7_module_106__or_module_8_res,
         n_majority7_module_106__and_module_7_res,
         n_majority7_module_106__or_module_7_res,
         n_majority7_module_106__or_module_6_res,
         n_majority7_module_106__and_module_6_res,
         n_majority7_module_106__or_module_5_res,
         n_majority7_module_106__and_module_5_res,
         n_majority7_module_106__or_module_4_res,
         n_majority7_module_106__and_module_4_res,
         n_majority7_module_106__or_module_3_res,
         n_majority7_module_106__and_module_3_res,
         n_majority7_module_106__or_module_2_res,
         n_majority7_module_106__and_module_2_res,
         n_majority7_module_106__or_module_1_res,
         n_majority7_module_106__and_module_1_res,
         n_majority7_module_107__and_module_10_res,
         n_majority7_module_107__or_module_11_res,
         n_majority7_module_107__and_module_9_res,
         n_majority7_module_107__or_module_10_res,
         n_majority7_module_107__or_module_9_res,
         n_majority7_module_107__and_module_8_res,
         n_majority7_module_107__or_module_8_res,
         n_majority7_module_107__and_module_7_res,
         n_majority7_module_107__or_module_7_res,
         n_majority7_module_107__or_module_6_res,
         n_majority7_module_107__and_module_6_res,
         n_majority7_module_107__or_module_5_res,
         n_majority7_module_107__and_module_5_res,
         n_majority7_module_107__or_module_4_res,
         n_majority7_module_107__and_module_4_res,
         n_majority7_module_107__or_module_3_res,
         n_majority7_module_107__and_module_3_res,
         n_majority7_module_107__or_module_2_res,
         n_majority7_module_107__and_module_2_res,
         n_majority7_module_107__or_module_1_res,
         n_majority7_module_107__and_module_1_res,
         n_majority7_module_108__and_module_10_res,
         n_majority7_module_108__or_module_11_res,
         n_majority7_module_108__and_module_9_res,
         n_majority7_module_108__or_module_10_res,
         n_majority7_module_108__or_module_9_res,
         n_majority7_module_108__and_module_8_res,
         n_majority7_module_108__or_module_8_res,
         n_majority7_module_108__and_module_7_res,
         n_majority7_module_108__or_module_7_res,
         n_majority7_module_108__or_module_6_res,
         n_majority7_module_108__and_module_6_res,
         n_majority7_module_108__or_module_5_res,
         n_majority7_module_108__and_module_5_res,
         n_majority7_module_108__or_module_4_res,
         n_majority7_module_108__and_module_4_res,
         n_majority7_module_108__or_module_3_res,
         n_majority7_module_108__and_module_3_res,
         n_majority7_module_108__or_module_2_res,
         n_majority7_module_108__and_module_2_res,
         n_majority7_module_108__or_module_1_res,
         n_majority7_module_108__and_module_1_res,
         n_majority7_module_109__and_module_10_res,
         n_majority7_module_109__or_module_11_res,
         n_majority7_module_109__and_module_9_res,
         n_majority7_module_109__or_module_10_res,
         n_majority7_module_109__or_module_9_res,
         n_majority7_module_109__and_module_8_res,
         n_majority7_module_109__or_module_8_res,
         n_majority7_module_109__and_module_7_res,
         n_majority7_module_109__or_module_7_res,
         n_majority7_module_109__or_module_6_res,
         n_majority7_module_109__and_module_6_res,
         n_majority7_module_109__or_module_5_res,
         n_majority7_module_109__and_module_5_res,
         n_majority7_module_109__or_module_4_res,
         n_majority7_module_109__and_module_4_res,
         n_majority7_module_109__or_module_3_res,
         n_majority7_module_109__and_module_3_res,
         n_majority7_module_109__or_module_2_res,
         n_majority7_module_109__and_module_2_res,
         n_majority7_module_109__or_module_1_res,
         n_majority7_module_109__and_module_1_res,
         n_majority7_module_110__and_module_10_res,
         n_majority7_module_110__or_module_11_res,
         n_majority7_module_110__and_module_9_res,
         n_majority7_module_110__or_module_10_res,
         n_majority7_module_110__or_module_9_res,
         n_majority7_module_110__and_module_8_res,
         n_majority7_module_110__or_module_8_res,
         n_majority7_module_110__and_module_7_res,
         n_majority7_module_110__or_module_7_res,
         n_majority7_module_110__or_module_6_res,
         n_majority7_module_110__and_module_6_res,
         n_majority7_module_110__or_module_5_res,
         n_majority7_module_110__and_module_5_res,
         n_majority7_module_110__or_module_4_res,
         n_majority7_module_110__and_module_4_res,
         n_majority7_module_110__or_module_3_res,
         n_majority7_module_110__and_module_3_res,
         n_majority7_module_110__or_module_2_res,
         n_majority7_module_110__and_module_2_res,
         n_majority7_module_110__or_module_1_res,
         n_majority7_module_110__and_module_1_res,
         n_majority7_module_111__and_module_10_res,
         n_majority7_module_111__or_module_11_res,
         n_majority7_module_111__and_module_9_res,
         n_majority7_module_111__or_module_10_res,
         n_majority7_module_111__or_module_9_res,
         n_majority7_module_111__and_module_8_res,
         n_majority7_module_111__or_module_8_res,
         n_majority7_module_111__and_module_7_res,
         n_majority7_module_111__or_module_7_res,
         n_majority7_module_111__or_module_6_res,
         n_majority7_module_111__and_module_6_res,
         n_majority7_module_111__or_module_5_res,
         n_majority7_module_111__and_module_5_res,
         n_majority7_module_111__or_module_4_res,
         n_majority7_module_111__and_module_4_res,
         n_majority7_module_111__or_module_3_res,
         n_majority7_module_111__and_module_3_res,
         n_majority7_module_111__or_module_2_res,
         n_majority7_module_111__and_module_2_res,
         n_majority7_module_111__or_module_1_res,
         n_majority7_module_111__and_module_1_res;

  XOR2_X1 u_xor_module_1_U1 ( .A(p_rand_0), .B(io_i1_s0_d0), .Z(
        n_xor_module_1_res) );
  XOR2_X1 u_xor_module_2_U1 ( .A(p_rand_1), .B(n_xor_module_1_res), .Z(
        n_xor_module_2_res) );
  XOR2_X1 u_xor_module_3_U1 ( .A(p_rand_2), .B(n_xor_module_2_res), .Z(
        n_xor_module_3_res) );
  XOR2_X1 u_xor_module_4_U1 ( .A(p_rand_0), .B(io_i1_s1_d0), .Z(
        n_xor_module_4_res) );
  XOR2_X1 u_xor_module_5_U1 ( .A(p_rand_3), .B(n_xor_module_4_res), .Z(
        n_xor_module_5_res) );
  XOR2_X1 u_xor_module_6_U1 ( .A(p_rand_4), .B(n_xor_module_5_res), .Z(
        n_xor_module_6_res) );
  XOR2_X1 u_xor_module_7_U1 ( .A(p_rand_1), .B(io_i1_s2_d0), .Z(
        n_xor_module_7_res) );
  XOR2_X1 u_xor_module_8_U1 ( .A(p_rand_3), .B(n_xor_module_7_res), .Z(
        n_xor_module_8_res) );
  XOR2_X1 u_xor_module_9_U1 ( .A(p_rand_5), .B(n_xor_module_8_res), .Z(
        n_xor_module_9_res) );
  XOR2_X1 u_xor_module_10_U1 ( .A(p_rand_2), .B(io_i1_s3_d0), .Z(
        n_xor_module_10_res) );
  XOR2_X1 u_xor_module_11_U1 ( .A(p_rand_4), .B(n_xor_module_10_res), .Z(
        n_xor_module_11_res) );
  XOR2_X1 u_xor_module_12_U1 ( .A(p_rand_5), .B(n_xor_module_11_res), .Z(
        n_xor_module_12_res) );
  XOR2_X1 u_xor_module_13_U1 ( .A(p_rand_0), .B(io_i1_s0_d1), .Z(
        n_xor_module_13_res) );
  XOR2_X1 u_xor_module_14_U1 ( .A(p_rand_1), .B(n_xor_module_13_res), .Z(
        n_xor_module_14_res) );
  XOR2_X1 u_xor_module_15_U1 ( .A(p_rand_2), .B(n_xor_module_14_res), .Z(
        n_xor_module_15_res) );
  XOR2_X1 u_xor_module_16_U1 ( .A(p_rand_0), .B(io_i1_s1_d1), .Z(
        n_xor_module_16_res) );
  XOR2_X1 u_xor_module_17_U1 ( .A(p_rand_3), .B(n_xor_module_16_res), .Z(
        n_xor_module_17_res) );
  XOR2_X1 u_xor_module_18_U1 ( .A(p_rand_4), .B(n_xor_module_17_res), .Z(
        n_xor_module_18_res) );
  XOR2_X1 u_xor_module_19_U1 ( .A(p_rand_1), .B(io_i1_s2_d1), .Z(
        n_xor_module_19_res) );
  XOR2_X1 u_xor_module_20_U1 ( .A(p_rand_3), .B(n_xor_module_19_res), .Z(
        n_xor_module_20_res) );
  XOR2_X1 u_xor_module_21_U1 ( .A(p_rand_5), .B(n_xor_module_20_res), .Z(
        n_xor_module_21_res) );
  XOR2_X1 u_xor_module_22_U1 ( .A(p_rand_2), .B(io_i1_s3_d1), .Z(
        n_xor_module_22_res) );
  XOR2_X1 u_xor_module_23_U1 ( .A(p_rand_4), .B(n_xor_module_22_res), .Z(
        n_xor_module_23_res) );
  XOR2_X1 u_xor_module_24_U1 ( .A(p_rand_5), .B(n_xor_module_23_res), .Z(
        n_xor_module_24_res) );
  XOR2_X1 u_xor_module_25_U1 ( .A(p_rand_0), .B(io_i1_s0_d2), .Z(
        n_xor_module_25_res) );
  XOR2_X1 u_xor_module_26_U1 ( .A(p_rand_1), .B(n_xor_module_25_res), .Z(
        n_xor_module_26_res) );
  XOR2_X1 u_xor_module_27_U1 ( .A(p_rand_2), .B(n_xor_module_26_res), .Z(
        n_xor_module_27_res) );
  XOR2_X1 u_xor_module_28_U1 ( .A(p_rand_0), .B(io_i1_s1_d2), .Z(
        n_xor_module_28_res) );
  XOR2_X1 u_xor_module_29_U1 ( .A(p_rand_3), .B(n_xor_module_28_res), .Z(
        n_xor_module_29_res) );
  XOR2_X1 u_xor_module_30_U1 ( .A(p_rand_4), .B(n_xor_module_29_res), .Z(
        n_xor_module_30_res) );
  XOR2_X1 u_xor_module_31_U1 ( .A(p_rand_1), .B(io_i1_s2_d2), .Z(
        n_xor_module_31_res) );
  XOR2_X1 u_xor_module_32_U1 ( .A(p_rand_3), .B(n_xor_module_31_res), .Z(
        n_xor_module_32_res) );
  XOR2_X1 u_xor_module_33_U1 ( .A(p_rand_5), .B(n_xor_module_32_res), .Z(
        n_xor_module_33_res) );
  XOR2_X1 u_xor_module_34_U1 ( .A(p_rand_2), .B(io_i1_s3_d2), .Z(
        n_xor_module_34_res) );
  XOR2_X1 u_xor_module_35_U1 ( .A(p_rand_4), .B(n_xor_module_34_res), .Z(
        n_xor_module_35_res) );
  XOR2_X1 u_xor_module_36_U1 ( .A(p_rand_5), .B(n_xor_module_35_res), .Z(
        n_xor_module_36_res) );
  XOR2_X1 u_xor_module_37_U1 ( .A(p_rand_0), .B(io_i1_s0_d3), .Z(
        n_xor_module_37_res) );
  XOR2_X1 u_xor_module_38_U1 ( .A(p_rand_1), .B(n_xor_module_37_res), .Z(
        n_xor_module_38_res) );
  XOR2_X1 u_xor_module_39_U1 ( .A(p_rand_2), .B(n_xor_module_38_res), .Z(
        n_xor_module_39_res) );
  XOR2_X1 u_xor_module_40_U1 ( .A(p_rand_0), .B(io_i1_s1_d3), .Z(
        n_xor_module_40_res) );
  XOR2_X1 u_xor_module_41_U1 ( .A(p_rand_3), .B(n_xor_module_40_res), .Z(
        n_xor_module_41_res) );
  XOR2_X1 u_xor_module_42_U1 ( .A(p_rand_4), .B(n_xor_module_41_res), .Z(
        n_xor_module_42_res) );
  XOR2_X1 u_xor_module_43_U1 ( .A(p_rand_1), .B(io_i1_s2_d3), .Z(
        n_xor_module_43_res) );
  XOR2_X1 u_xor_module_44_U1 ( .A(p_rand_3), .B(n_xor_module_43_res), .Z(
        n_xor_module_44_res) );
  XOR2_X1 u_xor_module_45_U1 ( .A(p_rand_5), .B(n_xor_module_44_res), .Z(
        n_xor_module_45_res) );
  XOR2_X1 u_xor_module_46_U1 ( .A(p_rand_2), .B(io_i1_s3_d3), .Z(
        n_xor_module_46_res) );
  XOR2_X1 u_xor_module_47_U1 ( .A(p_rand_4), .B(n_xor_module_46_res), .Z(
        n_xor_module_47_res) );
  XOR2_X1 u_xor_module_48_U1 ( .A(p_rand_5), .B(n_xor_module_47_res), .Z(
        n_xor_module_48_res) );
  XOR2_X1 u_xor_module_49_U1 ( .A(p_rand_0), .B(io_i1_s0_d4), .Z(
        n_xor_module_49_res) );
  XOR2_X1 u_xor_module_50_U1 ( .A(p_rand_1), .B(n_xor_module_49_res), .Z(
        n_xor_module_50_res) );
  XOR2_X1 u_xor_module_51_U1 ( .A(p_rand_2), .B(n_xor_module_50_res), .Z(
        n_xor_module_51_res) );
  XOR2_X1 u_xor_module_52_U1 ( .A(p_rand_0), .B(io_i1_s1_d4), .Z(
        n_xor_module_52_res) );
  XOR2_X1 u_xor_module_53_U1 ( .A(p_rand_3), .B(n_xor_module_52_res), .Z(
        n_xor_module_53_res) );
  XOR2_X1 u_xor_module_54_U1 ( .A(p_rand_4), .B(n_xor_module_53_res), .Z(
        n_xor_module_54_res) );
  XOR2_X1 u_xor_module_55_U1 ( .A(p_rand_1), .B(io_i1_s2_d4), .Z(
        n_xor_module_55_res) );
  XOR2_X1 u_xor_module_56_U1 ( .A(p_rand_3), .B(n_xor_module_55_res), .Z(
        n_xor_module_56_res) );
  XOR2_X1 u_xor_module_57_U1 ( .A(p_rand_5), .B(n_xor_module_56_res), .Z(
        n_xor_module_57_res) );
  XOR2_X1 u_xor_module_58_U1 ( .A(p_rand_2), .B(io_i1_s3_d4), .Z(
        n_xor_module_58_res) );
  XOR2_X1 u_xor_module_59_U1 ( .A(p_rand_4), .B(n_xor_module_58_res), .Z(
        n_xor_module_59_res) );
  XOR2_X1 u_xor_module_60_U1 ( .A(p_rand_5), .B(n_xor_module_59_res), .Z(
        n_xor_module_60_res) );
  XOR2_X1 u_xor_module_61_U1 ( .A(p_rand_0), .B(io_i1_s0_d5), .Z(
        n_xor_module_61_res) );
  XOR2_X1 u_xor_module_62_U1 ( .A(p_rand_1), .B(n_xor_module_61_res), .Z(
        n_xor_module_62_res) );
  XOR2_X1 u_xor_module_63_U1 ( .A(p_rand_2), .B(n_xor_module_62_res), .Z(
        n_xor_module_63_res) );
  XOR2_X1 u_xor_module_64_U1 ( .A(p_rand_0), .B(io_i1_s1_d5), .Z(
        n_xor_module_64_res) );
  XOR2_X1 u_xor_module_65_U1 ( .A(p_rand_3), .B(n_xor_module_64_res), .Z(
        n_xor_module_65_res) );
  XOR2_X1 u_xor_module_66_U1 ( .A(p_rand_4), .B(n_xor_module_65_res), .Z(
        n_xor_module_66_res) );
  XOR2_X1 u_xor_module_67_U1 ( .A(p_rand_1), .B(io_i1_s2_d5), .Z(
        n_xor_module_67_res) );
  XOR2_X1 u_xor_module_68_U1 ( .A(p_rand_3), .B(n_xor_module_67_res), .Z(
        n_xor_module_68_res) );
  XOR2_X1 u_xor_module_69_U1 ( .A(p_rand_5), .B(n_xor_module_68_res), .Z(
        n_xor_module_69_res) );
  XOR2_X1 u_xor_module_70_U1 ( .A(p_rand_2), .B(io_i1_s3_d5), .Z(
        n_xor_module_70_res) );
  XOR2_X1 u_xor_module_71_U1 ( .A(p_rand_4), .B(n_xor_module_70_res), .Z(
        n_xor_module_71_res) );
  XOR2_X1 u_xor_module_72_U1 ( .A(p_rand_5), .B(n_xor_module_71_res), .Z(
        n_xor_module_72_res) );
  XOR2_X1 u_xor_module_73_U1 ( .A(p_rand_0), .B(io_i1_s0_d6), .Z(
        n_xor_module_73_res) );
  XOR2_X1 u_xor_module_74_U1 ( .A(p_rand_1), .B(n_xor_module_73_res), .Z(
        n_xor_module_74_res) );
  XOR2_X1 u_xor_module_75_U1 ( .A(p_rand_2), .B(n_xor_module_74_res), .Z(
        n_xor_module_75_res) );
  XOR2_X1 u_xor_module_76_U1 ( .A(p_rand_0), .B(io_i1_s1_d6), .Z(
        n_xor_module_76_res) );
  XOR2_X1 u_xor_module_77_U1 ( .A(p_rand_3), .B(n_xor_module_76_res), .Z(
        n_xor_module_77_res) );
  XOR2_X1 u_xor_module_78_U1 ( .A(p_rand_4), .B(n_xor_module_77_res), .Z(
        n_xor_module_78_res) );
  XOR2_X1 u_xor_module_79_U1 ( .A(p_rand_1), .B(io_i1_s2_d6), .Z(
        n_xor_module_79_res) );
  XOR2_X1 u_xor_module_80_U1 ( .A(p_rand_3), .B(n_xor_module_79_res), .Z(
        n_xor_module_80_res) );
  XOR2_X1 u_xor_module_81_U1 ( .A(p_rand_5), .B(n_xor_module_80_res), .Z(
        n_xor_module_81_res) );
  XOR2_X1 u_xor_module_82_U1 ( .A(p_rand_2), .B(io_i1_s3_d6), .Z(
        n_xor_module_82_res) );
  XOR2_X1 u_xor_module_83_U1 ( .A(p_rand_4), .B(n_xor_module_82_res), .Z(
        n_xor_module_83_res) );
  XOR2_X1 u_xor_module_84_U1 ( .A(p_rand_5), .B(n_xor_module_83_res), .Z(
        n_xor_module_84_res) );
  AND2_X1 u_majority7_module_0__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_0__and_module_1_res)
         );
  OR2_X1 u_majority7_module_0__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_0__or_module_1_res) );
  AND2_X1 u_majority7_module_0__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_0__and_module_2_res)
         );
  OR2_X1 u_majority7_module_0__or_module_2_U1 ( .A1(n_xor_module_27_res), .A2(
        n_xor_module_39_res), .ZN(n_majority7_module_0__or_module_2_res) );
  AND2_X1 u_majority7_module_0__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_0__and_module_3_res)
         );
  OR2_X1 u_majority7_module_0__or_module_3_U1 ( .A1(n_xor_module_51_res), .A2(
        n_xor_module_63_res), .ZN(n_majority7_module_0__or_module_3_res) );
  AND2_X1 u_majority7_module_0__and_module_4_U1 ( .A1(
        n_majority7_module_0__and_module_2_res), .A2(
        n_majority7_module_0__and_module_1_res), .ZN(
        n_majority7_module_0__and_module_4_res) );
  OR2_X1 u_majority7_module_0__or_module_4_U1 ( .A1(
        n_majority7_module_0__and_module_1_res), .A2(
        n_majority7_module_0__and_module_2_res), .ZN(
        n_majority7_module_0__or_module_4_res) );
  AND2_X1 u_majority7_module_0__and_module_5_U1 ( .A1(
        n_majority7_module_0__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_0__and_module_5_res) );
  OR2_X1 u_majority7_module_0__or_module_5_U1 ( .A1(n_xor_module_15_res), .A2(
        n_majority7_module_0__and_module_3_res), .ZN(
        n_majority7_module_0__or_module_5_res) );
  AND2_X1 u_majority7_module_0__and_module_6_U1 ( .A1(
        n_majority7_module_0__or_module_1_res), .A2(
        n_majority7_module_0__or_module_2_res), .ZN(
        n_majority7_module_0__and_module_6_res) );
  OR2_X1 u_majority7_module_0__or_module_6_U1 ( .A1(
        n_majority7_module_0__or_module_2_res), .A2(
        n_majority7_module_0__or_module_1_res), .ZN(
        n_majority7_module_0__or_module_6_res) );
  OR2_X1 u_majority7_module_0__or_module_7_U1 ( .A1(
        n_majority7_module_0__and_module_4_res), .A2(
        n_majority7_module_0__and_module_5_res), .ZN(
        n_majority7_module_0__or_module_7_res) );
  AND2_X1 u_majority7_module_0__and_module_7_U1 ( .A1(
        n_majority7_module_0__or_module_3_res), .A2(
        n_majority7_module_0__or_module_4_res), .ZN(
        n_majority7_module_0__and_module_7_res) );
  OR2_X1 u_majority7_module_0__or_module_8_U1 ( .A1(
        n_majority7_module_0__or_module_4_res), .A2(
        n_majority7_module_0__or_module_3_res), .ZN(
        n_majority7_module_0__or_module_8_res) );
  AND2_X1 u_majority7_module_0__and_module_8_U1 ( .A1(
        n_majority7_module_0__or_module_5_res), .A2(
        n_majority7_module_0__and_module_6_res), .ZN(
        n_majority7_module_0__and_module_8_res) );
  OR2_X1 u_majority7_module_0__or_module_9_U1 ( .A1(
        n_majority7_module_0__and_module_6_res), .A2(
        n_majority7_module_0__or_module_5_res), .ZN(
        n_majority7_module_0__or_module_9_res) );
  OR2_X1 u_majority7_module_0__or_module_10_U1 ( .A1(
        n_majority7_module_0__or_module_7_res), .A2(
        n_majority7_module_0__and_module_7_res), .ZN(
        n_majority7_module_0__or_module_10_res) );
  AND2_X1 u_majority7_module_0__and_module_9_U1 ( .A1(
        n_majority7_module_0__or_module_6_res), .A2(
        n_majority7_module_0__or_module_9_res), .ZN(
        n_majority7_module_0__and_module_9_res) );
  OR2_X1 u_majority7_module_0__or_module_11_U1 ( .A1(
        n_majority7_module_0__or_module_10_res), .A2(
        n_majority7_module_0__and_module_8_res), .ZN(
        n_majority7_module_0__or_module_11_res) );
  AND2_X1 u_majority7_module_0__and_module_10_U1 ( .A1(
        n_majority7_module_0__or_module_8_res), .A2(
        n_majority7_module_0__and_module_9_res), .ZN(
        n_majority7_module_0__and_module_10_res) );
  AND2_X1 u_majority7_module_0__and_module_11_U1 ( .A1(
        n_majority7_module_0__and_module_10_res), .A2(
        n_majority7_module_0__or_module_11_res), .ZN(n_majority7_module_0_res)
         );
  DFF_X1 u_reg_module_1__cini_mul_v00_reg ( .D(n_majority7_module_0_res), .CK(
        clock_0), .Q(n_reg_module_1_res), .QN() );
  AND2_X1 u_majority7_module_1__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_1__and_module_1_res)
         );
  OR2_X1 u_majority7_module_1__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_1__or_module_1_res) );
  AND2_X1 u_majority7_module_1__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_1__and_module_2_res)
         );
  OR2_X1 u_majority7_module_1__or_module_2_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_1__or_module_2_res) );
  AND2_X1 u_majority7_module_1__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_1__and_module_3_res)
         );
  OR2_X1 u_majority7_module_1__or_module_3_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_66_res), .ZN(n_majority7_module_1__or_module_3_res) );
  AND2_X1 u_majority7_module_1__and_module_4_U1 ( .A1(
        n_majority7_module_1__and_module_2_res), .A2(
        n_majority7_module_1__and_module_1_res), .ZN(
        n_majority7_module_1__and_module_4_res) );
  OR2_X1 u_majority7_module_1__or_module_4_U1 ( .A1(
        n_majority7_module_1__and_module_1_res), .A2(
        n_majority7_module_1__and_module_2_res), .ZN(
        n_majority7_module_1__or_module_4_res) );
  AND2_X1 u_majority7_module_1__and_module_5_U1 ( .A1(
        n_majority7_module_1__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_1__and_module_5_res) );
  OR2_X1 u_majority7_module_1__or_module_5_U1 ( .A1(n_xor_module_18_res), .A2(
        n_majority7_module_1__and_module_3_res), .ZN(
        n_majority7_module_1__or_module_5_res) );
  AND2_X1 u_majority7_module_1__and_module_6_U1 ( .A1(
        n_majority7_module_1__or_module_1_res), .A2(
        n_majority7_module_1__or_module_2_res), .ZN(
        n_majority7_module_1__and_module_6_res) );
  OR2_X1 u_majority7_module_1__or_module_6_U1 ( .A1(
        n_majority7_module_1__or_module_2_res), .A2(
        n_majority7_module_1__or_module_1_res), .ZN(
        n_majority7_module_1__or_module_6_res) );
  OR2_X1 u_majority7_module_1__or_module_7_U1 ( .A1(
        n_majority7_module_1__and_module_4_res), .A2(
        n_majority7_module_1__and_module_5_res), .ZN(
        n_majority7_module_1__or_module_7_res) );
  AND2_X1 u_majority7_module_1__and_module_7_U1 ( .A1(
        n_majority7_module_1__or_module_3_res), .A2(
        n_majority7_module_1__or_module_4_res), .ZN(
        n_majority7_module_1__and_module_7_res) );
  OR2_X1 u_majority7_module_1__or_module_8_U1 ( .A1(
        n_majority7_module_1__or_module_4_res), .A2(
        n_majority7_module_1__or_module_3_res), .ZN(
        n_majority7_module_1__or_module_8_res) );
  AND2_X1 u_majority7_module_1__and_module_8_U1 ( .A1(
        n_majority7_module_1__or_module_5_res), .A2(
        n_majority7_module_1__and_module_6_res), .ZN(
        n_majority7_module_1__and_module_8_res) );
  OR2_X1 u_majority7_module_1__or_module_9_U1 ( .A1(
        n_majority7_module_1__and_module_6_res), .A2(
        n_majority7_module_1__or_module_5_res), .ZN(
        n_majority7_module_1__or_module_9_res) );
  OR2_X1 u_majority7_module_1__or_module_10_U1 ( .A1(
        n_majority7_module_1__or_module_7_res), .A2(
        n_majority7_module_1__and_module_7_res), .ZN(
        n_majority7_module_1__or_module_10_res) );
  AND2_X1 u_majority7_module_1__and_module_9_U1 ( .A1(
        n_majority7_module_1__or_module_6_res), .A2(
        n_majority7_module_1__or_module_9_res), .ZN(
        n_majority7_module_1__and_module_9_res) );
  OR2_X1 u_majority7_module_1__or_module_11_U1 ( .A1(
        n_majority7_module_1__or_module_10_res), .A2(
        n_majority7_module_1__and_module_8_res), .ZN(
        n_majority7_module_1__or_module_11_res) );
  AND2_X1 u_majority7_module_1__and_module_10_U1 ( .A1(
        n_majority7_module_1__or_module_8_res), .A2(
        n_majority7_module_1__and_module_9_res), .ZN(
        n_majority7_module_1__and_module_10_res) );
  AND2_X1 u_majority7_module_1__and_module_11_U1 ( .A1(
        n_majority7_module_1__and_module_10_res), .A2(
        n_majority7_module_1__or_module_11_res), .ZN(n_majority7_module_1_res)
         );
  DFF_X1 u_reg_module_2__cini_mul_v00_reg ( .D(n_majority7_module_1_res), .CK(
        clock_0), .Q(n_reg_module_2_res), .QN() );
  AND2_X1 u_majority7_module_2__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_2__and_module_1_res)
         );
  OR2_X1 u_majority7_module_2__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_2__or_module_1_res) );
  AND2_X1 u_majority7_module_2__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_2__and_module_2_res)
         );
  OR2_X1 u_majority7_module_2__or_module_2_U1 ( .A1(n_xor_module_33_res), .A2(
        n_xor_module_45_res), .ZN(n_majority7_module_2__or_module_2_res) );
  AND2_X1 u_majority7_module_2__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_2__and_module_3_res)
         );
  OR2_X1 u_majority7_module_2__or_module_3_U1 ( .A1(n_xor_module_57_res), .A2(
        n_xor_module_69_res), .ZN(n_majority7_module_2__or_module_3_res) );
  AND2_X1 u_majority7_module_2__and_module_4_U1 ( .A1(
        n_majority7_module_2__and_module_2_res), .A2(
        n_majority7_module_2__and_module_1_res), .ZN(
        n_majority7_module_2__and_module_4_res) );
  OR2_X1 u_majority7_module_2__or_module_4_U1 ( .A1(
        n_majority7_module_2__and_module_1_res), .A2(
        n_majority7_module_2__and_module_2_res), .ZN(
        n_majority7_module_2__or_module_4_res) );
  AND2_X1 u_majority7_module_2__and_module_5_U1 ( .A1(
        n_majority7_module_2__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_2__and_module_5_res) );
  OR2_X1 u_majority7_module_2__or_module_5_U1 ( .A1(n_xor_module_21_res), .A2(
        n_majority7_module_2__and_module_3_res), .ZN(
        n_majority7_module_2__or_module_5_res) );
  AND2_X1 u_majority7_module_2__and_module_6_U1 ( .A1(
        n_majority7_module_2__or_module_1_res), .A2(
        n_majority7_module_2__or_module_2_res), .ZN(
        n_majority7_module_2__and_module_6_res) );
  OR2_X1 u_majority7_module_2__or_module_6_U1 ( .A1(
        n_majority7_module_2__or_module_2_res), .A2(
        n_majority7_module_2__or_module_1_res), .ZN(
        n_majority7_module_2__or_module_6_res) );
  OR2_X1 u_majority7_module_2__or_module_7_U1 ( .A1(
        n_majority7_module_2__and_module_4_res), .A2(
        n_majority7_module_2__and_module_5_res), .ZN(
        n_majority7_module_2__or_module_7_res) );
  AND2_X1 u_majority7_module_2__and_module_7_U1 ( .A1(
        n_majority7_module_2__or_module_3_res), .A2(
        n_majority7_module_2__or_module_4_res), .ZN(
        n_majority7_module_2__and_module_7_res) );
  OR2_X1 u_majority7_module_2__or_module_8_U1 ( .A1(
        n_majority7_module_2__or_module_4_res), .A2(
        n_majority7_module_2__or_module_3_res), .ZN(
        n_majority7_module_2__or_module_8_res) );
  AND2_X1 u_majority7_module_2__and_module_8_U1 ( .A1(
        n_majority7_module_2__or_module_5_res), .A2(
        n_majority7_module_2__and_module_6_res), .ZN(
        n_majority7_module_2__and_module_8_res) );
  OR2_X1 u_majority7_module_2__or_module_9_U1 ( .A1(
        n_majority7_module_2__and_module_6_res), .A2(
        n_majority7_module_2__or_module_5_res), .ZN(
        n_majority7_module_2__or_module_9_res) );
  OR2_X1 u_majority7_module_2__or_module_10_U1 ( .A1(
        n_majority7_module_2__or_module_7_res), .A2(
        n_majority7_module_2__and_module_7_res), .ZN(
        n_majority7_module_2__or_module_10_res) );
  AND2_X1 u_majority7_module_2__and_module_9_U1 ( .A1(
        n_majority7_module_2__or_module_6_res), .A2(
        n_majority7_module_2__or_module_9_res), .ZN(
        n_majority7_module_2__and_module_9_res) );
  OR2_X1 u_majority7_module_2__or_module_11_U1 ( .A1(
        n_majority7_module_2__or_module_10_res), .A2(
        n_majority7_module_2__and_module_8_res), .ZN(
        n_majority7_module_2__or_module_11_res) );
  AND2_X1 u_majority7_module_2__and_module_10_U1 ( .A1(
        n_majority7_module_2__or_module_8_res), .A2(
        n_majority7_module_2__and_module_9_res), .ZN(
        n_majority7_module_2__and_module_10_res) );
  AND2_X1 u_majority7_module_2__and_module_11_U1 ( .A1(
        n_majority7_module_2__and_module_10_res), .A2(
        n_majority7_module_2__or_module_11_res), .ZN(n_majority7_module_2_res)
         );
  DFF_X1 u_reg_module_3__cini_mul_v00_reg ( .D(n_majority7_module_2_res), .CK(
        clock_0), .Q(n_reg_module_3_res), .QN() );
  AND2_X1 u_majority7_module_3__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_3__and_module_1_res)
         );
  OR2_X1 u_majority7_module_3__or_module_1_U1 ( .A1(n_xor_module_12_res), .A2(
        n_xor_module_84_res), .ZN(n_majority7_module_3__or_module_1_res) );
  AND2_X1 u_majority7_module_3__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_3__and_module_2_res)
         );
  OR2_X1 u_majority7_module_3__or_module_2_U1 ( .A1(n_xor_module_36_res), .A2(
        n_xor_module_48_res), .ZN(n_majority7_module_3__or_module_2_res) );
  AND2_X1 u_majority7_module_3__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_3__and_module_3_res)
         );
  OR2_X1 u_majority7_module_3__or_module_3_U1 ( .A1(n_xor_module_60_res), .A2(
        n_xor_module_72_res), .ZN(n_majority7_module_3__or_module_3_res) );
  AND2_X1 u_majority7_module_3__and_module_4_U1 ( .A1(
        n_majority7_module_3__and_module_2_res), .A2(
        n_majority7_module_3__and_module_1_res), .ZN(
        n_majority7_module_3__and_module_4_res) );
  OR2_X1 u_majority7_module_3__or_module_4_U1 ( .A1(
        n_majority7_module_3__and_module_1_res), .A2(
        n_majority7_module_3__and_module_2_res), .ZN(
        n_majority7_module_3__or_module_4_res) );
  AND2_X1 u_majority7_module_3__and_module_5_U1 ( .A1(
        n_majority7_module_3__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_3__and_module_5_res) );
  OR2_X1 u_majority7_module_3__or_module_5_U1 ( .A1(n_xor_module_24_res), .A2(
        n_majority7_module_3__and_module_3_res), .ZN(
        n_majority7_module_3__or_module_5_res) );
  AND2_X1 u_majority7_module_3__and_module_6_U1 ( .A1(
        n_majority7_module_3__or_module_1_res), .A2(
        n_majority7_module_3__or_module_2_res), .ZN(
        n_majority7_module_3__and_module_6_res) );
  OR2_X1 u_majority7_module_3__or_module_6_U1 ( .A1(
        n_majority7_module_3__or_module_2_res), .A2(
        n_majority7_module_3__or_module_1_res), .ZN(
        n_majority7_module_3__or_module_6_res) );
  OR2_X1 u_majority7_module_3__or_module_7_U1 ( .A1(
        n_majority7_module_3__and_module_4_res), .A2(
        n_majority7_module_3__and_module_5_res), .ZN(
        n_majority7_module_3__or_module_7_res) );
  AND2_X1 u_majority7_module_3__and_module_7_U1 ( .A1(
        n_majority7_module_3__or_module_3_res), .A2(
        n_majority7_module_3__or_module_4_res), .ZN(
        n_majority7_module_3__and_module_7_res) );
  OR2_X1 u_majority7_module_3__or_module_8_U1 ( .A1(
        n_majority7_module_3__or_module_4_res), .A2(
        n_majority7_module_3__or_module_3_res), .ZN(
        n_majority7_module_3__or_module_8_res) );
  AND2_X1 u_majority7_module_3__and_module_8_U1 ( .A1(
        n_majority7_module_3__or_module_5_res), .A2(
        n_majority7_module_3__and_module_6_res), .ZN(
        n_majority7_module_3__and_module_8_res) );
  OR2_X1 u_majority7_module_3__or_module_9_U1 ( .A1(
        n_majority7_module_3__and_module_6_res), .A2(
        n_majority7_module_3__or_module_5_res), .ZN(
        n_majority7_module_3__or_module_9_res) );
  OR2_X1 u_majority7_module_3__or_module_10_U1 ( .A1(
        n_majority7_module_3__or_module_7_res), .A2(
        n_majority7_module_3__and_module_7_res), .ZN(
        n_majority7_module_3__or_module_10_res) );
  AND2_X1 u_majority7_module_3__and_module_9_U1 ( .A1(
        n_majority7_module_3__or_module_6_res), .A2(
        n_majority7_module_3__or_module_9_res), .ZN(
        n_majority7_module_3__and_module_9_res) );
  OR2_X1 u_majority7_module_3__or_module_11_U1 ( .A1(
        n_majority7_module_3__or_module_10_res), .A2(
        n_majority7_module_3__and_module_8_res), .ZN(
        n_majority7_module_3__or_module_11_res) );
  AND2_X1 u_majority7_module_3__and_module_10_U1 ( .A1(
        n_majority7_module_3__or_module_8_res), .A2(
        n_majority7_module_3__and_module_9_res), .ZN(
        n_majority7_module_3__and_module_10_res) );
  AND2_X1 u_majority7_module_3__and_module_11_U1 ( .A1(
        n_majority7_module_3__and_module_10_res), .A2(
        n_majority7_module_3__or_module_11_res), .ZN(n_majority7_module_3_res)
         );
  DFF_X1 u_reg_module_4__cini_mul_v00_reg ( .D(n_majority7_module_3_res), .CK(
        clock_0), .Q(n_reg_module_4_res), .QN() );
  AND2_X1 u_majority7_module_4__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_4__and_module_1_res)
         );
  OR2_X1 u_majority7_module_4__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_4__or_module_1_res) );
  AND2_X1 u_majority7_module_4__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_4__and_module_2_res)
         );
  OR2_X1 u_majority7_module_4__or_module_2_U1 ( .A1(n_xor_module_27_res), .A2(
        n_xor_module_39_res), .ZN(n_majority7_module_4__or_module_2_res) );
  AND2_X1 u_majority7_module_4__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_4__and_module_3_res)
         );
  OR2_X1 u_majority7_module_4__or_module_3_U1 ( .A1(n_xor_module_51_res), .A2(
        n_xor_module_63_res), .ZN(n_majority7_module_4__or_module_3_res) );
  AND2_X1 u_majority7_module_4__and_module_4_U1 ( .A1(
        n_majority7_module_4__and_module_2_res), .A2(
        n_majority7_module_4__and_module_1_res), .ZN(
        n_majority7_module_4__and_module_4_res) );
  OR2_X1 u_majority7_module_4__or_module_4_U1 ( .A1(
        n_majority7_module_4__and_module_1_res), .A2(
        n_majority7_module_4__and_module_2_res), .ZN(
        n_majority7_module_4__or_module_4_res) );
  AND2_X1 u_majority7_module_4__and_module_5_U1 ( .A1(
        n_majority7_module_4__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_4__and_module_5_res) );
  OR2_X1 u_majority7_module_4__or_module_5_U1 ( .A1(n_xor_module_15_res), .A2(
        n_majority7_module_4__and_module_3_res), .ZN(
        n_majority7_module_4__or_module_5_res) );
  AND2_X1 u_majority7_module_4__and_module_6_U1 ( .A1(
        n_majority7_module_4__or_module_1_res), .A2(
        n_majority7_module_4__or_module_2_res), .ZN(
        n_majority7_module_4__and_module_6_res) );
  OR2_X1 u_majority7_module_4__or_module_6_U1 ( .A1(
        n_majority7_module_4__or_module_2_res), .A2(
        n_majority7_module_4__or_module_1_res), .ZN(
        n_majority7_module_4__or_module_6_res) );
  OR2_X1 u_majority7_module_4__or_module_7_U1 ( .A1(
        n_majority7_module_4__and_module_4_res), .A2(
        n_majority7_module_4__and_module_5_res), .ZN(
        n_majority7_module_4__or_module_7_res) );
  AND2_X1 u_majority7_module_4__and_module_7_U1 ( .A1(
        n_majority7_module_4__or_module_3_res), .A2(
        n_majority7_module_4__or_module_4_res), .ZN(
        n_majority7_module_4__and_module_7_res) );
  OR2_X1 u_majority7_module_4__or_module_8_U1 ( .A1(
        n_majority7_module_4__or_module_4_res), .A2(
        n_majority7_module_4__or_module_3_res), .ZN(
        n_majority7_module_4__or_module_8_res) );
  AND2_X1 u_majority7_module_4__and_module_8_U1 ( .A1(
        n_majority7_module_4__or_module_5_res), .A2(
        n_majority7_module_4__and_module_6_res), .ZN(
        n_majority7_module_4__and_module_8_res) );
  OR2_X1 u_majority7_module_4__or_module_9_U1 ( .A1(
        n_majority7_module_4__and_module_6_res), .A2(
        n_majority7_module_4__or_module_5_res), .ZN(
        n_majority7_module_4__or_module_9_res) );
  OR2_X1 u_majority7_module_4__or_module_10_U1 ( .A1(
        n_majority7_module_4__or_module_7_res), .A2(
        n_majority7_module_4__and_module_7_res), .ZN(
        n_majority7_module_4__or_module_10_res) );
  AND2_X1 u_majority7_module_4__and_module_9_U1 ( .A1(
        n_majority7_module_4__or_module_6_res), .A2(
        n_majority7_module_4__or_module_9_res), .ZN(
        n_majority7_module_4__and_module_9_res) );
  OR2_X1 u_majority7_module_4__or_module_11_U1 ( .A1(
        n_majority7_module_4__or_module_10_res), .A2(
        n_majority7_module_4__and_module_8_res), .ZN(
        n_majority7_module_4__or_module_11_res) );
  AND2_X1 u_majority7_module_4__and_module_10_U1 ( .A1(
        n_majority7_module_4__or_module_8_res), .A2(
        n_majority7_module_4__and_module_9_res), .ZN(
        n_majority7_module_4__and_module_10_res) );
  AND2_X1 u_majority7_module_4__and_module_11_U1 ( .A1(
        n_majority7_module_4__and_module_10_res), .A2(
        n_majority7_module_4__or_module_11_res), .ZN(n_majority7_module_4_res)
         );
  DFF_X1 u_reg_module_5__cini_mul_v00_reg ( .D(n_majority7_module_4_res), .CK(
        clock_1), .Q(n_reg_module_5_res), .QN() );
  AND2_X1 u_majority7_module_5__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_5__and_module_1_res)
         );
  OR2_X1 u_majority7_module_5__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_5__or_module_1_res) );
  AND2_X1 u_majority7_module_5__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_5__and_module_2_res)
         );
  OR2_X1 u_majority7_module_5__or_module_2_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_5__or_module_2_res) );
  AND2_X1 u_majority7_module_5__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_5__and_module_3_res)
         );
  OR2_X1 u_majority7_module_5__or_module_3_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_66_res), .ZN(n_majority7_module_5__or_module_3_res) );
  AND2_X1 u_majority7_module_5__and_module_4_U1 ( .A1(
        n_majority7_module_5__and_module_2_res), .A2(
        n_majority7_module_5__and_module_1_res), .ZN(
        n_majority7_module_5__and_module_4_res) );
  OR2_X1 u_majority7_module_5__or_module_4_U1 ( .A1(
        n_majority7_module_5__and_module_1_res), .A2(
        n_majority7_module_5__and_module_2_res), .ZN(
        n_majority7_module_5__or_module_4_res) );
  AND2_X1 u_majority7_module_5__and_module_5_U1 ( .A1(
        n_majority7_module_5__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_5__and_module_5_res) );
  OR2_X1 u_majority7_module_5__or_module_5_U1 ( .A1(n_xor_module_18_res), .A2(
        n_majority7_module_5__and_module_3_res), .ZN(
        n_majority7_module_5__or_module_5_res) );
  AND2_X1 u_majority7_module_5__and_module_6_U1 ( .A1(
        n_majority7_module_5__or_module_1_res), .A2(
        n_majority7_module_5__or_module_2_res), .ZN(
        n_majority7_module_5__and_module_6_res) );
  OR2_X1 u_majority7_module_5__or_module_6_U1 ( .A1(
        n_majority7_module_5__or_module_2_res), .A2(
        n_majority7_module_5__or_module_1_res), .ZN(
        n_majority7_module_5__or_module_6_res) );
  OR2_X1 u_majority7_module_5__or_module_7_U1 ( .A1(
        n_majority7_module_5__and_module_4_res), .A2(
        n_majority7_module_5__and_module_5_res), .ZN(
        n_majority7_module_5__or_module_7_res) );
  AND2_X1 u_majority7_module_5__and_module_7_U1 ( .A1(
        n_majority7_module_5__or_module_3_res), .A2(
        n_majority7_module_5__or_module_4_res), .ZN(
        n_majority7_module_5__and_module_7_res) );
  OR2_X1 u_majority7_module_5__or_module_8_U1 ( .A1(
        n_majority7_module_5__or_module_4_res), .A2(
        n_majority7_module_5__or_module_3_res), .ZN(
        n_majority7_module_5__or_module_8_res) );
  AND2_X1 u_majority7_module_5__and_module_8_U1 ( .A1(
        n_majority7_module_5__or_module_5_res), .A2(
        n_majority7_module_5__and_module_6_res), .ZN(
        n_majority7_module_5__and_module_8_res) );
  OR2_X1 u_majority7_module_5__or_module_9_U1 ( .A1(
        n_majority7_module_5__and_module_6_res), .A2(
        n_majority7_module_5__or_module_5_res), .ZN(
        n_majority7_module_5__or_module_9_res) );
  OR2_X1 u_majority7_module_5__or_module_10_U1 ( .A1(
        n_majority7_module_5__or_module_7_res), .A2(
        n_majority7_module_5__and_module_7_res), .ZN(
        n_majority7_module_5__or_module_10_res) );
  AND2_X1 u_majority7_module_5__and_module_9_U1 ( .A1(
        n_majority7_module_5__or_module_6_res), .A2(
        n_majority7_module_5__or_module_9_res), .ZN(
        n_majority7_module_5__and_module_9_res) );
  OR2_X1 u_majority7_module_5__or_module_11_U1 ( .A1(
        n_majority7_module_5__or_module_10_res), .A2(
        n_majority7_module_5__and_module_8_res), .ZN(
        n_majority7_module_5__or_module_11_res) );
  AND2_X1 u_majority7_module_5__and_module_10_U1 ( .A1(
        n_majority7_module_5__or_module_8_res), .A2(
        n_majority7_module_5__and_module_9_res), .ZN(
        n_majority7_module_5__and_module_10_res) );
  AND2_X1 u_majority7_module_5__and_module_11_U1 ( .A1(
        n_majority7_module_5__and_module_10_res), .A2(
        n_majority7_module_5__or_module_11_res), .ZN(n_majority7_module_5_res)
         );
  DFF_X1 u_reg_module_6__cini_mul_v00_reg ( .D(n_majority7_module_5_res), .CK(
        clock_1), .Q(n_reg_module_6_res), .QN() );
  AND2_X1 u_majority7_module_6__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_6__and_module_1_res)
         );
  OR2_X1 u_majority7_module_6__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_6__or_module_1_res) );
  AND2_X1 u_majority7_module_6__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_6__and_module_2_res)
         );
  OR2_X1 u_majority7_module_6__or_module_2_U1 ( .A1(n_xor_module_33_res), .A2(
        n_xor_module_45_res), .ZN(n_majority7_module_6__or_module_2_res) );
  AND2_X1 u_majority7_module_6__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_6__and_module_3_res)
         );
  OR2_X1 u_majority7_module_6__or_module_3_U1 ( .A1(n_xor_module_57_res), .A2(
        n_xor_module_69_res), .ZN(n_majority7_module_6__or_module_3_res) );
  AND2_X1 u_majority7_module_6__and_module_4_U1 ( .A1(
        n_majority7_module_6__and_module_2_res), .A2(
        n_majority7_module_6__and_module_1_res), .ZN(
        n_majority7_module_6__and_module_4_res) );
  OR2_X1 u_majority7_module_6__or_module_4_U1 ( .A1(
        n_majority7_module_6__and_module_1_res), .A2(
        n_majority7_module_6__and_module_2_res), .ZN(
        n_majority7_module_6__or_module_4_res) );
  AND2_X1 u_majority7_module_6__and_module_5_U1 ( .A1(
        n_majority7_module_6__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_6__and_module_5_res) );
  OR2_X1 u_majority7_module_6__or_module_5_U1 ( .A1(n_xor_module_21_res), .A2(
        n_majority7_module_6__and_module_3_res), .ZN(
        n_majority7_module_6__or_module_5_res) );
  AND2_X1 u_majority7_module_6__and_module_6_U1 ( .A1(
        n_majority7_module_6__or_module_1_res), .A2(
        n_majority7_module_6__or_module_2_res), .ZN(
        n_majority7_module_6__and_module_6_res) );
  OR2_X1 u_majority7_module_6__or_module_6_U1 ( .A1(
        n_majority7_module_6__or_module_2_res), .A2(
        n_majority7_module_6__or_module_1_res), .ZN(
        n_majority7_module_6__or_module_6_res) );
  OR2_X1 u_majority7_module_6__or_module_7_U1 ( .A1(
        n_majority7_module_6__and_module_4_res), .A2(
        n_majority7_module_6__and_module_5_res), .ZN(
        n_majority7_module_6__or_module_7_res) );
  AND2_X1 u_majority7_module_6__and_module_7_U1 ( .A1(
        n_majority7_module_6__or_module_3_res), .A2(
        n_majority7_module_6__or_module_4_res), .ZN(
        n_majority7_module_6__and_module_7_res) );
  OR2_X1 u_majority7_module_6__or_module_8_U1 ( .A1(
        n_majority7_module_6__or_module_4_res), .A2(
        n_majority7_module_6__or_module_3_res), .ZN(
        n_majority7_module_6__or_module_8_res) );
  AND2_X1 u_majority7_module_6__and_module_8_U1 ( .A1(
        n_majority7_module_6__or_module_5_res), .A2(
        n_majority7_module_6__and_module_6_res), .ZN(
        n_majority7_module_6__and_module_8_res) );
  OR2_X1 u_majority7_module_6__or_module_9_U1 ( .A1(
        n_majority7_module_6__and_module_6_res), .A2(
        n_majority7_module_6__or_module_5_res), .ZN(
        n_majority7_module_6__or_module_9_res) );
  OR2_X1 u_majority7_module_6__or_module_10_U1 ( .A1(
        n_majority7_module_6__or_module_7_res), .A2(
        n_majority7_module_6__and_module_7_res), .ZN(
        n_majority7_module_6__or_module_10_res) );
  AND2_X1 u_majority7_module_6__and_module_9_U1 ( .A1(
        n_majority7_module_6__or_module_6_res), .A2(
        n_majority7_module_6__or_module_9_res), .ZN(
        n_majority7_module_6__and_module_9_res) );
  OR2_X1 u_majority7_module_6__or_module_11_U1 ( .A1(
        n_majority7_module_6__or_module_10_res), .A2(
        n_majority7_module_6__and_module_8_res), .ZN(
        n_majority7_module_6__or_module_11_res) );
  AND2_X1 u_majority7_module_6__and_module_10_U1 ( .A1(
        n_majority7_module_6__or_module_8_res), .A2(
        n_majority7_module_6__and_module_9_res), .ZN(
        n_majority7_module_6__and_module_10_res) );
  AND2_X1 u_majority7_module_6__and_module_11_U1 ( .A1(
        n_majority7_module_6__and_module_10_res), .A2(
        n_majority7_module_6__or_module_11_res), .ZN(n_majority7_module_6_res)
         );
  DFF_X1 u_reg_module_7__cini_mul_v00_reg ( .D(n_majority7_module_6_res), .CK(
        clock_1), .Q(n_reg_module_7_res), .QN() );
  AND2_X1 u_majority7_module_7__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_7__and_module_1_res)
         );
  OR2_X1 u_majority7_module_7__or_module_1_U1 ( .A1(n_xor_module_12_res), .A2(
        n_xor_module_84_res), .ZN(n_majority7_module_7__or_module_1_res) );
  AND2_X1 u_majority7_module_7__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_7__and_module_2_res)
         );
  OR2_X1 u_majority7_module_7__or_module_2_U1 ( .A1(n_xor_module_36_res), .A2(
        n_xor_module_48_res), .ZN(n_majority7_module_7__or_module_2_res) );
  AND2_X1 u_majority7_module_7__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_7__and_module_3_res)
         );
  OR2_X1 u_majority7_module_7__or_module_3_U1 ( .A1(n_xor_module_60_res), .A2(
        n_xor_module_72_res), .ZN(n_majority7_module_7__or_module_3_res) );
  AND2_X1 u_majority7_module_7__and_module_4_U1 ( .A1(
        n_majority7_module_7__and_module_2_res), .A2(
        n_majority7_module_7__and_module_1_res), .ZN(
        n_majority7_module_7__and_module_4_res) );
  OR2_X1 u_majority7_module_7__or_module_4_U1 ( .A1(
        n_majority7_module_7__and_module_1_res), .A2(
        n_majority7_module_7__and_module_2_res), .ZN(
        n_majority7_module_7__or_module_4_res) );
  AND2_X1 u_majority7_module_7__and_module_5_U1 ( .A1(
        n_majority7_module_7__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_7__and_module_5_res) );
  OR2_X1 u_majority7_module_7__or_module_5_U1 ( .A1(n_xor_module_24_res), .A2(
        n_majority7_module_7__and_module_3_res), .ZN(
        n_majority7_module_7__or_module_5_res) );
  AND2_X1 u_majority7_module_7__and_module_6_U1 ( .A1(
        n_majority7_module_7__or_module_1_res), .A2(
        n_majority7_module_7__or_module_2_res), .ZN(
        n_majority7_module_7__and_module_6_res) );
  OR2_X1 u_majority7_module_7__or_module_6_U1 ( .A1(
        n_majority7_module_7__or_module_2_res), .A2(
        n_majority7_module_7__or_module_1_res), .ZN(
        n_majority7_module_7__or_module_6_res) );
  OR2_X1 u_majority7_module_7__or_module_7_U1 ( .A1(
        n_majority7_module_7__and_module_4_res), .A2(
        n_majority7_module_7__and_module_5_res), .ZN(
        n_majority7_module_7__or_module_7_res) );
  AND2_X1 u_majority7_module_7__and_module_7_U1 ( .A1(
        n_majority7_module_7__or_module_3_res), .A2(
        n_majority7_module_7__or_module_4_res), .ZN(
        n_majority7_module_7__and_module_7_res) );
  OR2_X1 u_majority7_module_7__or_module_8_U1 ( .A1(
        n_majority7_module_7__or_module_4_res), .A2(
        n_majority7_module_7__or_module_3_res), .ZN(
        n_majority7_module_7__or_module_8_res) );
  AND2_X1 u_majority7_module_7__and_module_8_U1 ( .A1(
        n_majority7_module_7__or_module_5_res), .A2(
        n_majority7_module_7__and_module_6_res), .ZN(
        n_majority7_module_7__and_module_8_res) );
  OR2_X1 u_majority7_module_7__or_module_9_U1 ( .A1(
        n_majority7_module_7__and_module_6_res), .A2(
        n_majority7_module_7__or_module_5_res), .ZN(
        n_majority7_module_7__or_module_9_res) );
  OR2_X1 u_majority7_module_7__or_module_10_U1 ( .A1(
        n_majority7_module_7__or_module_7_res), .A2(
        n_majority7_module_7__and_module_7_res), .ZN(
        n_majority7_module_7__or_module_10_res) );
  AND2_X1 u_majority7_module_7__and_module_9_U1 ( .A1(
        n_majority7_module_7__or_module_6_res), .A2(
        n_majority7_module_7__or_module_9_res), .ZN(
        n_majority7_module_7__and_module_9_res) );
  OR2_X1 u_majority7_module_7__or_module_11_U1 ( .A1(
        n_majority7_module_7__or_module_10_res), .A2(
        n_majority7_module_7__and_module_8_res), .ZN(
        n_majority7_module_7__or_module_11_res) );
  AND2_X1 u_majority7_module_7__and_module_10_U1 ( .A1(
        n_majority7_module_7__or_module_8_res), .A2(
        n_majority7_module_7__and_module_9_res), .ZN(
        n_majority7_module_7__and_module_10_res) );
  AND2_X1 u_majority7_module_7__and_module_11_U1 ( .A1(
        n_majority7_module_7__and_module_10_res), .A2(
        n_majority7_module_7__or_module_11_res), .ZN(n_majority7_module_7_res)
         );
  DFF_X1 u_reg_module_8__cini_mul_v00_reg ( .D(n_majority7_module_7_res), .CK(
        clock_1), .Q(n_reg_module_8_res), .QN() );
  AND2_X1 u_majority7_module_8__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_8__and_module_1_res)
         );
  OR2_X1 u_majority7_module_8__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_8__or_module_1_res) );
  AND2_X1 u_majority7_module_8__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_8__and_module_2_res)
         );
  OR2_X1 u_majority7_module_8__or_module_2_U1 ( .A1(n_xor_module_27_res), .A2(
        n_xor_module_39_res), .ZN(n_majority7_module_8__or_module_2_res) );
  AND2_X1 u_majority7_module_8__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_8__and_module_3_res)
         );
  OR2_X1 u_majority7_module_8__or_module_3_U1 ( .A1(n_xor_module_51_res), .A2(
        n_xor_module_63_res), .ZN(n_majority7_module_8__or_module_3_res) );
  AND2_X1 u_majority7_module_8__and_module_4_U1 ( .A1(
        n_majority7_module_8__and_module_2_res), .A2(
        n_majority7_module_8__and_module_1_res), .ZN(
        n_majority7_module_8__and_module_4_res) );
  OR2_X1 u_majority7_module_8__or_module_4_U1 ( .A1(
        n_majority7_module_8__and_module_1_res), .A2(
        n_majority7_module_8__and_module_2_res), .ZN(
        n_majority7_module_8__or_module_4_res) );
  AND2_X1 u_majority7_module_8__and_module_5_U1 ( .A1(
        n_majority7_module_8__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_8__and_module_5_res) );
  OR2_X1 u_majority7_module_8__or_module_5_U1 ( .A1(n_xor_module_15_res), .A2(
        n_majority7_module_8__and_module_3_res), .ZN(
        n_majority7_module_8__or_module_5_res) );
  AND2_X1 u_majority7_module_8__and_module_6_U1 ( .A1(
        n_majority7_module_8__or_module_1_res), .A2(
        n_majority7_module_8__or_module_2_res), .ZN(
        n_majority7_module_8__and_module_6_res) );
  OR2_X1 u_majority7_module_8__or_module_6_U1 ( .A1(
        n_majority7_module_8__or_module_2_res), .A2(
        n_majority7_module_8__or_module_1_res), .ZN(
        n_majority7_module_8__or_module_6_res) );
  OR2_X1 u_majority7_module_8__or_module_7_U1 ( .A1(
        n_majority7_module_8__and_module_4_res), .A2(
        n_majority7_module_8__and_module_5_res), .ZN(
        n_majority7_module_8__or_module_7_res) );
  AND2_X1 u_majority7_module_8__and_module_7_U1 ( .A1(
        n_majority7_module_8__or_module_3_res), .A2(
        n_majority7_module_8__or_module_4_res), .ZN(
        n_majority7_module_8__and_module_7_res) );
  OR2_X1 u_majority7_module_8__or_module_8_U1 ( .A1(
        n_majority7_module_8__or_module_4_res), .A2(
        n_majority7_module_8__or_module_3_res), .ZN(
        n_majority7_module_8__or_module_8_res) );
  AND2_X1 u_majority7_module_8__and_module_8_U1 ( .A1(
        n_majority7_module_8__or_module_5_res), .A2(
        n_majority7_module_8__and_module_6_res), .ZN(
        n_majority7_module_8__and_module_8_res) );
  OR2_X1 u_majority7_module_8__or_module_9_U1 ( .A1(
        n_majority7_module_8__and_module_6_res), .A2(
        n_majority7_module_8__or_module_5_res), .ZN(
        n_majority7_module_8__or_module_9_res) );
  OR2_X1 u_majority7_module_8__or_module_10_U1 ( .A1(
        n_majority7_module_8__or_module_7_res), .A2(
        n_majority7_module_8__and_module_7_res), .ZN(
        n_majority7_module_8__or_module_10_res) );
  AND2_X1 u_majority7_module_8__and_module_9_U1 ( .A1(
        n_majority7_module_8__or_module_6_res), .A2(
        n_majority7_module_8__or_module_9_res), .ZN(
        n_majority7_module_8__and_module_9_res) );
  OR2_X1 u_majority7_module_8__or_module_11_U1 ( .A1(
        n_majority7_module_8__or_module_10_res), .A2(
        n_majority7_module_8__and_module_8_res), .ZN(
        n_majority7_module_8__or_module_11_res) );
  AND2_X1 u_majority7_module_8__and_module_10_U1 ( .A1(
        n_majority7_module_8__or_module_8_res), .A2(
        n_majority7_module_8__and_module_9_res), .ZN(
        n_majority7_module_8__and_module_10_res) );
  AND2_X1 u_majority7_module_8__and_module_11_U1 ( .A1(
        n_majority7_module_8__and_module_10_res), .A2(
        n_majority7_module_8__or_module_11_res), .ZN(n_majority7_module_8_res)
         );
  DFF_X1 u_reg_module_9__cini_mul_v00_reg ( .D(n_majority7_module_8_res), .CK(
        clock_2), .Q(n_reg_module_9_res), .QN() );
  AND2_X1 u_majority7_module_9__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_9__and_module_1_res)
         );
  OR2_X1 u_majority7_module_9__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_9__or_module_1_res) );
  AND2_X1 u_majority7_module_9__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_9__and_module_2_res)
         );
  OR2_X1 u_majority7_module_9__or_module_2_U1 ( .A1(n_xor_module_30_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_9__or_module_2_res) );
  AND2_X1 u_majority7_module_9__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_9__and_module_3_res)
         );
  OR2_X1 u_majority7_module_9__or_module_3_U1 ( .A1(n_xor_module_54_res), .A2(
        n_xor_module_66_res), .ZN(n_majority7_module_9__or_module_3_res) );
  AND2_X1 u_majority7_module_9__and_module_4_U1 ( .A1(
        n_majority7_module_9__and_module_2_res), .A2(
        n_majority7_module_9__and_module_1_res), .ZN(
        n_majority7_module_9__and_module_4_res) );
  OR2_X1 u_majority7_module_9__or_module_4_U1 ( .A1(
        n_majority7_module_9__and_module_1_res), .A2(
        n_majority7_module_9__and_module_2_res), .ZN(
        n_majority7_module_9__or_module_4_res) );
  AND2_X1 u_majority7_module_9__and_module_5_U1 ( .A1(
        n_majority7_module_9__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_9__and_module_5_res) );
  OR2_X1 u_majority7_module_9__or_module_5_U1 ( .A1(n_xor_module_18_res), .A2(
        n_majority7_module_9__and_module_3_res), .ZN(
        n_majority7_module_9__or_module_5_res) );
  AND2_X1 u_majority7_module_9__and_module_6_U1 ( .A1(
        n_majority7_module_9__or_module_1_res), .A2(
        n_majority7_module_9__or_module_2_res), .ZN(
        n_majority7_module_9__and_module_6_res) );
  OR2_X1 u_majority7_module_9__or_module_6_U1 ( .A1(
        n_majority7_module_9__or_module_2_res), .A2(
        n_majority7_module_9__or_module_1_res), .ZN(
        n_majority7_module_9__or_module_6_res) );
  OR2_X1 u_majority7_module_9__or_module_7_U1 ( .A1(
        n_majority7_module_9__and_module_4_res), .A2(
        n_majority7_module_9__and_module_5_res), .ZN(
        n_majority7_module_9__or_module_7_res) );
  AND2_X1 u_majority7_module_9__and_module_7_U1 ( .A1(
        n_majority7_module_9__or_module_3_res), .A2(
        n_majority7_module_9__or_module_4_res), .ZN(
        n_majority7_module_9__and_module_7_res) );
  OR2_X1 u_majority7_module_9__or_module_8_U1 ( .A1(
        n_majority7_module_9__or_module_4_res), .A2(
        n_majority7_module_9__or_module_3_res), .ZN(
        n_majority7_module_9__or_module_8_res) );
  AND2_X1 u_majority7_module_9__and_module_8_U1 ( .A1(
        n_majority7_module_9__or_module_5_res), .A2(
        n_majority7_module_9__and_module_6_res), .ZN(
        n_majority7_module_9__and_module_8_res) );
  OR2_X1 u_majority7_module_9__or_module_9_U1 ( .A1(
        n_majority7_module_9__and_module_6_res), .A2(
        n_majority7_module_9__or_module_5_res), .ZN(
        n_majority7_module_9__or_module_9_res) );
  OR2_X1 u_majority7_module_9__or_module_10_U1 ( .A1(
        n_majority7_module_9__or_module_7_res), .A2(
        n_majority7_module_9__and_module_7_res), .ZN(
        n_majority7_module_9__or_module_10_res) );
  AND2_X1 u_majority7_module_9__and_module_9_U1 ( .A1(
        n_majority7_module_9__or_module_6_res), .A2(
        n_majority7_module_9__or_module_9_res), .ZN(
        n_majority7_module_9__and_module_9_res) );
  OR2_X1 u_majority7_module_9__or_module_11_U1 ( .A1(
        n_majority7_module_9__or_module_10_res), .A2(
        n_majority7_module_9__and_module_8_res), .ZN(
        n_majority7_module_9__or_module_11_res) );
  AND2_X1 u_majority7_module_9__and_module_10_U1 ( .A1(
        n_majority7_module_9__or_module_8_res), .A2(
        n_majority7_module_9__and_module_9_res), .ZN(
        n_majority7_module_9__and_module_10_res) );
  AND2_X1 u_majority7_module_9__and_module_11_U1 ( .A1(
        n_majority7_module_9__and_module_10_res), .A2(
        n_majority7_module_9__or_module_11_res), .ZN(n_majority7_module_9_res)
         );
  DFF_X1 u_reg_module_10__cini_mul_v00_reg ( .D(n_majority7_module_9_res), 
        .CK(clock_2), .Q(n_reg_module_10_res), .QN() );
  AND2_X1 u_majority7_module_10__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_10__and_module_1_res)
         );
  OR2_X1 u_majority7_module_10__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_10__or_module_1_res) );
  AND2_X1 u_majority7_module_10__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_10__and_module_2_res)
         );
  OR2_X1 u_majority7_module_10__or_module_2_U1 ( .A1(n_xor_module_33_res), 
        .A2(n_xor_module_45_res), .ZN(n_majority7_module_10__or_module_2_res)
         );
  AND2_X1 u_majority7_module_10__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_10__and_module_3_res)
         );
  OR2_X1 u_majority7_module_10__or_module_3_U1 ( .A1(n_xor_module_57_res), 
        .A2(n_xor_module_69_res), .ZN(n_majority7_module_10__or_module_3_res)
         );
  AND2_X1 u_majority7_module_10__and_module_4_U1 ( .A1(
        n_majority7_module_10__and_module_2_res), .A2(
        n_majority7_module_10__and_module_1_res), .ZN(
        n_majority7_module_10__and_module_4_res) );
  OR2_X1 u_majority7_module_10__or_module_4_U1 ( .A1(
        n_majority7_module_10__and_module_1_res), .A2(
        n_majority7_module_10__and_module_2_res), .ZN(
        n_majority7_module_10__or_module_4_res) );
  AND2_X1 u_majority7_module_10__and_module_5_U1 ( .A1(
        n_majority7_module_10__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_10__and_module_5_res) );
  OR2_X1 u_majority7_module_10__or_module_5_U1 ( .A1(n_xor_module_21_res), 
        .A2(n_majority7_module_10__and_module_3_res), .ZN(
        n_majority7_module_10__or_module_5_res) );
  AND2_X1 u_majority7_module_10__and_module_6_U1 ( .A1(
        n_majority7_module_10__or_module_1_res), .A2(
        n_majority7_module_10__or_module_2_res), .ZN(
        n_majority7_module_10__and_module_6_res) );
  OR2_X1 u_majority7_module_10__or_module_6_U1 ( .A1(
        n_majority7_module_10__or_module_2_res), .A2(
        n_majority7_module_10__or_module_1_res), .ZN(
        n_majority7_module_10__or_module_6_res) );
  OR2_X1 u_majority7_module_10__or_module_7_U1 ( .A1(
        n_majority7_module_10__and_module_4_res), .A2(
        n_majority7_module_10__and_module_5_res), .ZN(
        n_majority7_module_10__or_module_7_res) );
  AND2_X1 u_majority7_module_10__and_module_7_U1 ( .A1(
        n_majority7_module_10__or_module_3_res), .A2(
        n_majority7_module_10__or_module_4_res), .ZN(
        n_majority7_module_10__and_module_7_res) );
  OR2_X1 u_majority7_module_10__or_module_8_U1 ( .A1(
        n_majority7_module_10__or_module_4_res), .A2(
        n_majority7_module_10__or_module_3_res), .ZN(
        n_majority7_module_10__or_module_8_res) );
  AND2_X1 u_majority7_module_10__and_module_8_U1 ( .A1(
        n_majority7_module_10__or_module_5_res), .A2(
        n_majority7_module_10__and_module_6_res), .ZN(
        n_majority7_module_10__and_module_8_res) );
  OR2_X1 u_majority7_module_10__or_module_9_U1 ( .A1(
        n_majority7_module_10__and_module_6_res), .A2(
        n_majority7_module_10__or_module_5_res), .ZN(
        n_majority7_module_10__or_module_9_res) );
  OR2_X1 u_majority7_module_10__or_module_10_U1 ( .A1(
        n_majority7_module_10__or_module_7_res), .A2(
        n_majority7_module_10__and_module_7_res), .ZN(
        n_majority7_module_10__or_module_10_res) );
  AND2_X1 u_majority7_module_10__and_module_9_U1 ( .A1(
        n_majority7_module_10__or_module_6_res), .A2(
        n_majority7_module_10__or_module_9_res), .ZN(
        n_majority7_module_10__and_module_9_res) );
  OR2_X1 u_majority7_module_10__or_module_11_U1 ( .A1(
        n_majority7_module_10__or_module_10_res), .A2(
        n_majority7_module_10__and_module_8_res), .ZN(
        n_majority7_module_10__or_module_11_res) );
  AND2_X1 u_majority7_module_10__and_module_10_U1 ( .A1(
        n_majority7_module_10__or_module_8_res), .A2(
        n_majority7_module_10__and_module_9_res), .ZN(
        n_majority7_module_10__and_module_10_res) );
  AND2_X1 u_majority7_module_10__and_module_11_U1 ( .A1(
        n_majority7_module_10__and_module_10_res), .A2(
        n_majority7_module_10__or_module_11_res), .ZN(
        n_majority7_module_10_res) );
  DFF_X1 u_reg_module_11__cini_mul_v00_reg ( .D(n_majority7_module_10_res), 
        .CK(clock_2), .Q(n_reg_module_11_res), .QN() );
  AND2_X1 u_majority7_module_11__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_11__and_module_1_res)
         );
  OR2_X1 u_majority7_module_11__or_module_1_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_xor_module_84_res), .ZN(n_majority7_module_11__or_module_1_res)
         );
  AND2_X1 u_majority7_module_11__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_11__and_module_2_res)
         );
  OR2_X1 u_majority7_module_11__or_module_2_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_48_res), .ZN(n_majority7_module_11__or_module_2_res)
         );
  AND2_X1 u_majority7_module_11__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_11__and_module_3_res)
         );
  OR2_X1 u_majority7_module_11__or_module_3_U1 ( .A1(n_xor_module_60_res), 
        .A2(n_xor_module_72_res), .ZN(n_majority7_module_11__or_module_3_res)
         );
  AND2_X1 u_majority7_module_11__and_module_4_U1 ( .A1(
        n_majority7_module_11__and_module_2_res), .A2(
        n_majority7_module_11__and_module_1_res), .ZN(
        n_majority7_module_11__and_module_4_res) );
  OR2_X1 u_majority7_module_11__or_module_4_U1 ( .A1(
        n_majority7_module_11__and_module_1_res), .A2(
        n_majority7_module_11__and_module_2_res), .ZN(
        n_majority7_module_11__or_module_4_res) );
  AND2_X1 u_majority7_module_11__and_module_5_U1 ( .A1(
        n_majority7_module_11__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_11__and_module_5_res) );
  OR2_X1 u_majority7_module_11__or_module_5_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_majority7_module_11__and_module_3_res), .ZN(
        n_majority7_module_11__or_module_5_res) );
  AND2_X1 u_majority7_module_11__and_module_6_U1 ( .A1(
        n_majority7_module_11__or_module_1_res), .A2(
        n_majority7_module_11__or_module_2_res), .ZN(
        n_majority7_module_11__and_module_6_res) );
  OR2_X1 u_majority7_module_11__or_module_6_U1 ( .A1(
        n_majority7_module_11__or_module_2_res), .A2(
        n_majority7_module_11__or_module_1_res), .ZN(
        n_majority7_module_11__or_module_6_res) );
  OR2_X1 u_majority7_module_11__or_module_7_U1 ( .A1(
        n_majority7_module_11__and_module_4_res), .A2(
        n_majority7_module_11__and_module_5_res), .ZN(
        n_majority7_module_11__or_module_7_res) );
  AND2_X1 u_majority7_module_11__and_module_7_U1 ( .A1(
        n_majority7_module_11__or_module_3_res), .A2(
        n_majority7_module_11__or_module_4_res), .ZN(
        n_majority7_module_11__and_module_7_res) );
  OR2_X1 u_majority7_module_11__or_module_8_U1 ( .A1(
        n_majority7_module_11__or_module_4_res), .A2(
        n_majority7_module_11__or_module_3_res), .ZN(
        n_majority7_module_11__or_module_8_res) );
  AND2_X1 u_majority7_module_11__and_module_8_U1 ( .A1(
        n_majority7_module_11__or_module_5_res), .A2(
        n_majority7_module_11__and_module_6_res), .ZN(
        n_majority7_module_11__and_module_8_res) );
  OR2_X1 u_majority7_module_11__or_module_9_U1 ( .A1(
        n_majority7_module_11__and_module_6_res), .A2(
        n_majority7_module_11__or_module_5_res), .ZN(
        n_majority7_module_11__or_module_9_res) );
  OR2_X1 u_majority7_module_11__or_module_10_U1 ( .A1(
        n_majority7_module_11__or_module_7_res), .A2(
        n_majority7_module_11__and_module_7_res), .ZN(
        n_majority7_module_11__or_module_10_res) );
  AND2_X1 u_majority7_module_11__and_module_9_U1 ( .A1(
        n_majority7_module_11__or_module_6_res), .A2(
        n_majority7_module_11__or_module_9_res), .ZN(
        n_majority7_module_11__and_module_9_res) );
  OR2_X1 u_majority7_module_11__or_module_11_U1 ( .A1(
        n_majority7_module_11__or_module_10_res), .A2(
        n_majority7_module_11__and_module_8_res), .ZN(
        n_majority7_module_11__or_module_11_res) );
  AND2_X1 u_majority7_module_11__and_module_10_U1 ( .A1(
        n_majority7_module_11__or_module_8_res), .A2(
        n_majority7_module_11__and_module_9_res), .ZN(
        n_majority7_module_11__and_module_10_res) );
  AND2_X1 u_majority7_module_11__and_module_11_U1 ( .A1(
        n_majority7_module_11__and_module_10_res), .A2(
        n_majority7_module_11__or_module_11_res), .ZN(
        n_majority7_module_11_res) );
  DFF_X1 u_reg_module_12__cini_mul_v00_reg ( .D(n_majority7_module_11_res), 
        .CK(clock_2), .Q(n_reg_module_12_res), .QN() );
  AND2_X1 u_majority7_module_12__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_12__and_module_1_res)
         );
  OR2_X1 u_majority7_module_12__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_12__or_module_1_res) );
  AND2_X1 u_majority7_module_12__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_12__and_module_2_res)
         );
  OR2_X1 u_majority7_module_12__or_module_2_U1 ( .A1(n_xor_module_27_res), 
        .A2(n_xor_module_39_res), .ZN(n_majority7_module_12__or_module_2_res)
         );
  AND2_X1 u_majority7_module_12__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_12__and_module_3_res)
         );
  OR2_X1 u_majority7_module_12__or_module_3_U1 ( .A1(n_xor_module_51_res), 
        .A2(n_xor_module_63_res), .ZN(n_majority7_module_12__or_module_3_res)
         );
  AND2_X1 u_majority7_module_12__and_module_4_U1 ( .A1(
        n_majority7_module_12__and_module_2_res), .A2(
        n_majority7_module_12__and_module_1_res), .ZN(
        n_majority7_module_12__and_module_4_res) );
  OR2_X1 u_majority7_module_12__or_module_4_U1 ( .A1(
        n_majority7_module_12__and_module_1_res), .A2(
        n_majority7_module_12__and_module_2_res), .ZN(
        n_majority7_module_12__or_module_4_res) );
  AND2_X1 u_majority7_module_12__and_module_5_U1 ( .A1(
        n_majority7_module_12__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_12__and_module_5_res) );
  OR2_X1 u_majority7_module_12__or_module_5_U1 ( .A1(n_xor_module_15_res), 
        .A2(n_majority7_module_12__and_module_3_res), .ZN(
        n_majority7_module_12__or_module_5_res) );
  AND2_X1 u_majority7_module_12__and_module_6_U1 ( .A1(
        n_majority7_module_12__or_module_1_res), .A2(
        n_majority7_module_12__or_module_2_res), .ZN(
        n_majority7_module_12__and_module_6_res) );
  OR2_X1 u_majority7_module_12__or_module_6_U1 ( .A1(
        n_majority7_module_12__or_module_2_res), .A2(
        n_majority7_module_12__or_module_1_res), .ZN(
        n_majority7_module_12__or_module_6_res) );
  OR2_X1 u_majority7_module_12__or_module_7_U1 ( .A1(
        n_majority7_module_12__and_module_4_res), .A2(
        n_majority7_module_12__and_module_5_res), .ZN(
        n_majority7_module_12__or_module_7_res) );
  AND2_X1 u_majority7_module_12__and_module_7_U1 ( .A1(
        n_majority7_module_12__or_module_3_res), .A2(
        n_majority7_module_12__or_module_4_res), .ZN(
        n_majority7_module_12__and_module_7_res) );
  OR2_X1 u_majority7_module_12__or_module_8_U1 ( .A1(
        n_majority7_module_12__or_module_4_res), .A2(
        n_majority7_module_12__or_module_3_res), .ZN(
        n_majority7_module_12__or_module_8_res) );
  AND2_X1 u_majority7_module_12__and_module_8_U1 ( .A1(
        n_majority7_module_12__or_module_5_res), .A2(
        n_majority7_module_12__and_module_6_res), .ZN(
        n_majority7_module_12__and_module_8_res) );
  OR2_X1 u_majority7_module_12__or_module_9_U1 ( .A1(
        n_majority7_module_12__and_module_6_res), .A2(
        n_majority7_module_12__or_module_5_res), .ZN(
        n_majority7_module_12__or_module_9_res) );
  OR2_X1 u_majority7_module_12__or_module_10_U1 ( .A1(
        n_majority7_module_12__or_module_7_res), .A2(
        n_majority7_module_12__and_module_7_res), .ZN(
        n_majority7_module_12__or_module_10_res) );
  AND2_X1 u_majority7_module_12__and_module_9_U1 ( .A1(
        n_majority7_module_12__or_module_6_res), .A2(
        n_majority7_module_12__or_module_9_res), .ZN(
        n_majority7_module_12__and_module_9_res) );
  OR2_X1 u_majority7_module_12__or_module_11_U1 ( .A1(
        n_majority7_module_12__or_module_10_res), .A2(
        n_majority7_module_12__and_module_8_res), .ZN(
        n_majority7_module_12__or_module_11_res) );
  AND2_X1 u_majority7_module_12__and_module_10_U1 ( .A1(
        n_majority7_module_12__or_module_8_res), .A2(
        n_majority7_module_12__and_module_9_res), .ZN(
        n_majority7_module_12__and_module_10_res) );
  AND2_X1 u_majority7_module_12__and_module_11_U1 ( .A1(
        n_majority7_module_12__and_module_10_res), .A2(
        n_majority7_module_12__or_module_11_res), .ZN(
        n_majority7_module_12_res) );
  DFF_X1 u_reg_module_13__cini_mul_v00_reg ( .D(n_majority7_module_12_res), 
        .CK(clock_3), .Q(n_reg_module_13_res), .QN() );
  AND2_X1 u_majority7_module_13__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_13__and_module_1_res)
         );
  OR2_X1 u_majority7_module_13__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_13__or_module_1_res) );
  AND2_X1 u_majority7_module_13__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_13__and_module_2_res)
         );
  OR2_X1 u_majority7_module_13__or_module_2_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_42_res), .ZN(n_majority7_module_13__or_module_2_res)
         );
  AND2_X1 u_majority7_module_13__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_13__and_module_3_res)
         );
  OR2_X1 u_majority7_module_13__or_module_3_U1 ( .A1(n_xor_module_54_res), 
        .A2(n_xor_module_66_res), .ZN(n_majority7_module_13__or_module_3_res)
         );
  AND2_X1 u_majority7_module_13__and_module_4_U1 ( .A1(
        n_majority7_module_13__and_module_2_res), .A2(
        n_majority7_module_13__and_module_1_res), .ZN(
        n_majority7_module_13__and_module_4_res) );
  OR2_X1 u_majority7_module_13__or_module_4_U1 ( .A1(
        n_majority7_module_13__and_module_1_res), .A2(
        n_majority7_module_13__and_module_2_res), .ZN(
        n_majority7_module_13__or_module_4_res) );
  AND2_X1 u_majority7_module_13__and_module_5_U1 ( .A1(
        n_majority7_module_13__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_13__and_module_5_res) );
  OR2_X1 u_majority7_module_13__or_module_5_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_majority7_module_13__and_module_3_res), .ZN(
        n_majority7_module_13__or_module_5_res) );
  AND2_X1 u_majority7_module_13__and_module_6_U1 ( .A1(
        n_majority7_module_13__or_module_1_res), .A2(
        n_majority7_module_13__or_module_2_res), .ZN(
        n_majority7_module_13__and_module_6_res) );
  OR2_X1 u_majority7_module_13__or_module_6_U1 ( .A1(
        n_majority7_module_13__or_module_2_res), .A2(
        n_majority7_module_13__or_module_1_res), .ZN(
        n_majority7_module_13__or_module_6_res) );
  OR2_X1 u_majority7_module_13__or_module_7_U1 ( .A1(
        n_majority7_module_13__and_module_4_res), .A2(
        n_majority7_module_13__and_module_5_res), .ZN(
        n_majority7_module_13__or_module_7_res) );
  AND2_X1 u_majority7_module_13__and_module_7_U1 ( .A1(
        n_majority7_module_13__or_module_3_res), .A2(
        n_majority7_module_13__or_module_4_res), .ZN(
        n_majority7_module_13__and_module_7_res) );
  OR2_X1 u_majority7_module_13__or_module_8_U1 ( .A1(
        n_majority7_module_13__or_module_4_res), .A2(
        n_majority7_module_13__or_module_3_res), .ZN(
        n_majority7_module_13__or_module_8_res) );
  AND2_X1 u_majority7_module_13__and_module_8_U1 ( .A1(
        n_majority7_module_13__or_module_5_res), .A2(
        n_majority7_module_13__and_module_6_res), .ZN(
        n_majority7_module_13__and_module_8_res) );
  OR2_X1 u_majority7_module_13__or_module_9_U1 ( .A1(
        n_majority7_module_13__and_module_6_res), .A2(
        n_majority7_module_13__or_module_5_res), .ZN(
        n_majority7_module_13__or_module_9_res) );
  OR2_X1 u_majority7_module_13__or_module_10_U1 ( .A1(
        n_majority7_module_13__or_module_7_res), .A2(
        n_majority7_module_13__and_module_7_res), .ZN(
        n_majority7_module_13__or_module_10_res) );
  AND2_X1 u_majority7_module_13__and_module_9_U1 ( .A1(
        n_majority7_module_13__or_module_6_res), .A2(
        n_majority7_module_13__or_module_9_res), .ZN(
        n_majority7_module_13__and_module_9_res) );
  OR2_X1 u_majority7_module_13__or_module_11_U1 ( .A1(
        n_majority7_module_13__or_module_10_res), .A2(
        n_majority7_module_13__and_module_8_res), .ZN(
        n_majority7_module_13__or_module_11_res) );
  AND2_X1 u_majority7_module_13__and_module_10_U1 ( .A1(
        n_majority7_module_13__or_module_8_res), .A2(
        n_majority7_module_13__and_module_9_res), .ZN(
        n_majority7_module_13__and_module_10_res) );
  AND2_X1 u_majority7_module_13__and_module_11_U1 ( .A1(
        n_majority7_module_13__and_module_10_res), .A2(
        n_majority7_module_13__or_module_11_res), .ZN(
        n_majority7_module_13_res) );
  DFF_X1 u_reg_module_14__cini_mul_v00_reg ( .D(n_majority7_module_13_res), 
        .CK(clock_3), .Q(n_reg_module_14_res), .QN() );
  AND2_X1 u_majority7_module_14__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_14__and_module_1_res)
         );
  OR2_X1 u_majority7_module_14__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_14__or_module_1_res) );
  AND2_X1 u_majority7_module_14__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_14__and_module_2_res)
         );
  OR2_X1 u_majority7_module_14__or_module_2_U1 ( .A1(n_xor_module_33_res), 
        .A2(n_xor_module_45_res), .ZN(n_majority7_module_14__or_module_2_res)
         );
  AND2_X1 u_majority7_module_14__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_14__and_module_3_res)
         );
  OR2_X1 u_majority7_module_14__or_module_3_U1 ( .A1(n_xor_module_57_res), 
        .A2(n_xor_module_69_res), .ZN(n_majority7_module_14__or_module_3_res)
         );
  AND2_X1 u_majority7_module_14__and_module_4_U1 ( .A1(
        n_majority7_module_14__and_module_2_res), .A2(
        n_majority7_module_14__and_module_1_res), .ZN(
        n_majority7_module_14__and_module_4_res) );
  OR2_X1 u_majority7_module_14__or_module_4_U1 ( .A1(
        n_majority7_module_14__and_module_1_res), .A2(
        n_majority7_module_14__and_module_2_res), .ZN(
        n_majority7_module_14__or_module_4_res) );
  AND2_X1 u_majority7_module_14__and_module_5_U1 ( .A1(
        n_majority7_module_14__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_14__and_module_5_res) );
  OR2_X1 u_majority7_module_14__or_module_5_U1 ( .A1(n_xor_module_21_res), 
        .A2(n_majority7_module_14__and_module_3_res), .ZN(
        n_majority7_module_14__or_module_5_res) );
  AND2_X1 u_majority7_module_14__and_module_6_U1 ( .A1(
        n_majority7_module_14__or_module_1_res), .A2(
        n_majority7_module_14__or_module_2_res), .ZN(
        n_majority7_module_14__and_module_6_res) );
  OR2_X1 u_majority7_module_14__or_module_6_U1 ( .A1(
        n_majority7_module_14__or_module_2_res), .A2(
        n_majority7_module_14__or_module_1_res), .ZN(
        n_majority7_module_14__or_module_6_res) );
  OR2_X1 u_majority7_module_14__or_module_7_U1 ( .A1(
        n_majority7_module_14__and_module_4_res), .A2(
        n_majority7_module_14__and_module_5_res), .ZN(
        n_majority7_module_14__or_module_7_res) );
  AND2_X1 u_majority7_module_14__and_module_7_U1 ( .A1(
        n_majority7_module_14__or_module_3_res), .A2(
        n_majority7_module_14__or_module_4_res), .ZN(
        n_majority7_module_14__and_module_7_res) );
  OR2_X1 u_majority7_module_14__or_module_8_U1 ( .A1(
        n_majority7_module_14__or_module_4_res), .A2(
        n_majority7_module_14__or_module_3_res), .ZN(
        n_majority7_module_14__or_module_8_res) );
  AND2_X1 u_majority7_module_14__and_module_8_U1 ( .A1(
        n_majority7_module_14__or_module_5_res), .A2(
        n_majority7_module_14__and_module_6_res), .ZN(
        n_majority7_module_14__and_module_8_res) );
  OR2_X1 u_majority7_module_14__or_module_9_U1 ( .A1(
        n_majority7_module_14__and_module_6_res), .A2(
        n_majority7_module_14__or_module_5_res), .ZN(
        n_majority7_module_14__or_module_9_res) );
  OR2_X1 u_majority7_module_14__or_module_10_U1 ( .A1(
        n_majority7_module_14__or_module_7_res), .A2(
        n_majority7_module_14__and_module_7_res), .ZN(
        n_majority7_module_14__or_module_10_res) );
  AND2_X1 u_majority7_module_14__and_module_9_U1 ( .A1(
        n_majority7_module_14__or_module_6_res), .A2(
        n_majority7_module_14__or_module_9_res), .ZN(
        n_majority7_module_14__and_module_9_res) );
  OR2_X1 u_majority7_module_14__or_module_11_U1 ( .A1(
        n_majority7_module_14__or_module_10_res), .A2(
        n_majority7_module_14__and_module_8_res), .ZN(
        n_majority7_module_14__or_module_11_res) );
  AND2_X1 u_majority7_module_14__and_module_10_U1 ( .A1(
        n_majority7_module_14__or_module_8_res), .A2(
        n_majority7_module_14__and_module_9_res), .ZN(
        n_majority7_module_14__and_module_10_res) );
  AND2_X1 u_majority7_module_14__and_module_11_U1 ( .A1(
        n_majority7_module_14__and_module_10_res), .A2(
        n_majority7_module_14__or_module_11_res), .ZN(
        n_majority7_module_14_res) );
  DFF_X1 u_reg_module_15__cini_mul_v00_reg ( .D(n_majority7_module_14_res), 
        .CK(clock_3), .Q(n_reg_module_15_res), .QN() );
  AND2_X1 u_majority7_module_15__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_15__and_module_1_res)
         );
  OR2_X1 u_majority7_module_15__or_module_1_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_xor_module_84_res), .ZN(n_majority7_module_15__or_module_1_res)
         );
  AND2_X1 u_majority7_module_15__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_15__and_module_2_res)
         );
  OR2_X1 u_majority7_module_15__or_module_2_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_48_res), .ZN(n_majority7_module_15__or_module_2_res)
         );
  AND2_X1 u_majority7_module_15__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_15__and_module_3_res)
         );
  OR2_X1 u_majority7_module_15__or_module_3_U1 ( .A1(n_xor_module_60_res), 
        .A2(n_xor_module_72_res), .ZN(n_majority7_module_15__or_module_3_res)
         );
  AND2_X1 u_majority7_module_15__and_module_4_U1 ( .A1(
        n_majority7_module_15__and_module_2_res), .A2(
        n_majority7_module_15__and_module_1_res), .ZN(
        n_majority7_module_15__and_module_4_res) );
  OR2_X1 u_majority7_module_15__or_module_4_U1 ( .A1(
        n_majority7_module_15__and_module_1_res), .A2(
        n_majority7_module_15__and_module_2_res), .ZN(
        n_majority7_module_15__or_module_4_res) );
  AND2_X1 u_majority7_module_15__and_module_5_U1 ( .A1(
        n_majority7_module_15__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_15__and_module_5_res) );
  OR2_X1 u_majority7_module_15__or_module_5_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_majority7_module_15__and_module_3_res), .ZN(
        n_majority7_module_15__or_module_5_res) );
  AND2_X1 u_majority7_module_15__and_module_6_U1 ( .A1(
        n_majority7_module_15__or_module_1_res), .A2(
        n_majority7_module_15__or_module_2_res), .ZN(
        n_majority7_module_15__and_module_6_res) );
  OR2_X1 u_majority7_module_15__or_module_6_U1 ( .A1(
        n_majority7_module_15__or_module_2_res), .A2(
        n_majority7_module_15__or_module_1_res), .ZN(
        n_majority7_module_15__or_module_6_res) );
  OR2_X1 u_majority7_module_15__or_module_7_U1 ( .A1(
        n_majority7_module_15__and_module_4_res), .A2(
        n_majority7_module_15__and_module_5_res), .ZN(
        n_majority7_module_15__or_module_7_res) );
  AND2_X1 u_majority7_module_15__and_module_7_U1 ( .A1(
        n_majority7_module_15__or_module_3_res), .A2(
        n_majority7_module_15__or_module_4_res), .ZN(
        n_majority7_module_15__and_module_7_res) );
  OR2_X1 u_majority7_module_15__or_module_8_U1 ( .A1(
        n_majority7_module_15__or_module_4_res), .A2(
        n_majority7_module_15__or_module_3_res), .ZN(
        n_majority7_module_15__or_module_8_res) );
  AND2_X1 u_majority7_module_15__and_module_8_U1 ( .A1(
        n_majority7_module_15__or_module_5_res), .A2(
        n_majority7_module_15__and_module_6_res), .ZN(
        n_majority7_module_15__and_module_8_res) );
  OR2_X1 u_majority7_module_15__or_module_9_U1 ( .A1(
        n_majority7_module_15__and_module_6_res), .A2(
        n_majority7_module_15__or_module_5_res), .ZN(
        n_majority7_module_15__or_module_9_res) );
  OR2_X1 u_majority7_module_15__or_module_10_U1 ( .A1(
        n_majority7_module_15__or_module_7_res), .A2(
        n_majority7_module_15__and_module_7_res), .ZN(
        n_majority7_module_15__or_module_10_res) );
  AND2_X1 u_majority7_module_15__and_module_9_U1 ( .A1(
        n_majority7_module_15__or_module_6_res), .A2(
        n_majority7_module_15__or_module_9_res), .ZN(
        n_majority7_module_15__and_module_9_res) );
  OR2_X1 u_majority7_module_15__or_module_11_U1 ( .A1(
        n_majority7_module_15__or_module_10_res), .A2(
        n_majority7_module_15__and_module_8_res), .ZN(
        n_majority7_module_15__or_module_11_res) );
  AND2_X1 u_majority7_module_15__and_module_10_U1 ( .A1(
        n_majority7_module_15__or_module_8_res), .A2(
        n_majority7_module_15__and_module_9_res), .ZN(
        n_majority7_module_15__and_module_10_res) );
  AND2_X1 u_majority7_module_15__and_module_11_U1 ( .A1(
        n_majority7_module_15__and_module_10_res), .A2(
        n_majority7_module_15__or_module_11_res), .ZN(
        n_majority7_module_15_res) );
  DFF_X1 u_reg_module_16__cini_mul_v00_reg ( .D(n_majority7_module_15_res), 
        .CK(clock_3), .Q(n_reg_module_16_res), .QN() );
  AND2_X1 u_majority7_module_16__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_16__and_module_1_res)
         );
  OR2_X1 u_majority7_module_16__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_16__or_module_1_res) );
  AND2_X1 u_majority7_module_16__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_16__and_module_2_res)
         );
  OR2_X1 u_majority7_module_16__or_module_2_U1 ( .A1(n_xor_module_27_res), 
        .A2(n_xor_module_39_res), .ZN(n_majority7_module_16__or_module_2_res)
         );
  AND2_X1 u_majority7_module_16__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_16__and_module_3_res)
         );
  OR2_X1 u_majority7_module_16__or_module_3_U1 ( .A1(n_xor_module_51_res), 
        .A2(n_xor_module_63_res), .ZN(n_majority7_module_16__or_module_3_res)
         );
  AND2_X1 u_majority7_module_16__and_module_4_U1 ( .A1(
        n_majority7_module_16__and_module_2_res), .A2(
        n_majority7_module_16__and_module_1_res), .ZN(
        n_majority7_module_16__and_module_4_res) );
  OR2_X1 u_majority7_module_16__or_module_4_U1 ( .A1(
        n_majority7_module_16__and_module_1_res), .A2(
        n_majority7_module_16__and_module_2_res), .ZN(
        n_majority7_module_16__or_module_4_res) );
  AND2_X1 u_majority7_module_16__and_module_5_U1 ( .A1(
        n_majority7_module_16__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_16__and_module_5_res) );
  OR2_X1 u_majority7_module_16__or_module_5_U1 ( .A1(n_xor_module_15_res), 
        .A2(n_majority7_module_16__and_module_3_res), .ZN(
        n_majority7_module_16__or_module_5_res) );
  AND2_X1 u_majority7_module_16__and_module_6_U1 ( .A1(
        n_majority7_module_16__or_module_1_res), .A2(
        n_majority7_module_16__or_module_2_res), .ZN(
        n_majority7_module_16__and_module_6_res) );
  OR2_X1 u_majority7_module_16__or_module_6_U1 ( .A1(
        n_majority7_module_16__or_module_2_res), .A2(
        n_majority7_module_16__or_module_1_res), .ZN(
        n_majority7_module_16__or_module_6_res) );
  OR2_X1 u_majority7_module_16__or_module_7_U1 ( .A1(
        n_majority7_module_16__and_module_4_res), .A2(
        n_majority7_module_16__and_module_5_res), .ZN(
        n_majority7_module_16__or_module_7_res) );
  AND2_X1 u_majority7_module_16__and_module_7_U1 ( .A1(
        n_majority7_module_16__or_module_3_res), .A2(
        n_majority7_module_16__or_module_4_res), .ZN(
        n_majority7_module_16__and_module_7_res) );
  OR2_X1 u_majority7_module_16__or_module_8_U1 ( .A1(
        n_majority7_module_16__or_module_4_res), .A2(
        n_majority7_module_16__or_module_3_res), .ZN(
        n_majority7_module_16__or_module_8_res) );
  AND2_X1 u_majority7_module_16__and_module_8_U1 ( .A1(
        n_majority7_module_16__or_module_5_res), .A2(
        n_majority7_module_16__and_module_6_res), .ZN(
        n_majority7_module_16__and_module_8_res) );
  OR2_X1 u_majority7_module_16__or_module_9_U1 ( .A1(
        n_majority7_module_16__and_module_6_res), .A2(
        n_majority7_module_16__or_module_5_res), .ZN(
        n_majority7_module_16__or_module_9_res) );
  OR2_X1 u_majority7_module_16__or_module_10_U1 ( .A1(
        n_majority7_module_16__or_module_7_res), .A2(
        n_majority7_module_16__and_module_7_res), .ZN(
        n_majority7_module_16__or_module_10_res) );
  AND2_X1 u_majority7_module_16__and_module_9_U1 ( .A1(
        n_majority7_module_16__or_module_6_res), .A2(
        n_majority7_module_16__or_module_9_res), .ZN(
        n_majority7_module_16__and_module_9_res) );
  OR2_X1 u_majority7_module_16__or_module_11_U1 ( .A1(
        n_majority7_module_16__or_module_10_res), .A2(
        n_majority7_module_16__and_module_8_res), .ZN(
        n_majority7_module_16__or_module_11_res) );
  AND2_X1 u_majority7_module_16__and_module_10_U1 ( .A1(
        n_majority7_module_16__or_module_8_res), .A2(
        n_majority7_module_16__and_module_9_res), .ZN(
        n_majority7_module_16__and_module_10_res) );
  AND2_X1 u_majority7_module_16__and_module_11_U1 ( .A1(
        n_majority7_module_16__and_module_10_res), .A2(
        n_majority7_module_16__or_module_11_res), .ZN(
        n_majority7_module_16_res) );
  DFF_X1 u_reg_module_17__cini_mul_v00_reg ( .D(n_majority7_module_16_res), 
        .CK(clock_4), .Q(n_reg_module_17_res), .QN() );
  AND2_X1 u_majority7_module_17__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_17__and_module_1_res)
         );
  OR2_X1 u_majority7_module_17__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_17__or_module_1_res) );
  AND2_X1 u_majority7_module_17__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_17__and_module_2_res)
         );
  OR2_X1 u_majority7_module_17__or_module_2_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_42_res), .ZN(n_majority7_module_17__or_module_2_res)
         );
  AND2_X1 u_majority7_module_17__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_17__and_module_3_res)
         );
  OR2_X1 u_majority7_module_17__or_module_3_U1 ( .A1(n_xor_module_54_res), 
        .A2(n_xor_module_66_res), .ZN(n_majority7_module_17__or_module_3_res)
         );
  AND2_X1 u_majority7_module_17__and_module_4_U1 ( .A1(
        n_majority7_module_17__and_module_2_res), .A2(
        n_majority7_module_17__and_module_1_res), .ZN(
        n_majority7_module_17__and_module_4_res) );
  OR2_X1 u_majority7_module_17__or_module_4_U1 ( .A1(
        n_majority7_module_17__and_module_1_res), .A2(
        n_majority7_module_17__and_module_2_res), .ZN(
        n_majority7_module_17__or_module_4_res) );
  AND2_X1 u_majority7_module_17__and_module_5_U1 ( .A1(
        n_majority7_module_17__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_17__and_module_5_res) );
  OR2_X1 u_majority7_module_17__or_module_5_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_majority7_module_17__and_module_3_res), .ZN(
        n_majority7_module_17__or_module_5_res) );
  AND2_X1 u_majority7_module_17__and_module_6_U1 ( .A1(
        n_majority7_module_17__or_module_1_res), .A2(
        n_majority7_module_17__or_module_2_res), .ZN(
        n_majority7_module_17__and_module_6_res) );
  OR2_X1 u_majority7_module_17__or_module_6_U1 ( .A1(
        n_majority7_module_17__or_module_2_res), .A2(
        n_majority7_module_17__or_module_1_res), .ZN(
        n_majority7_module_17__or_module_6_res) );
  OR2_X1 u_majority7_module_17__or_module_7_U1 ( .A1(
        n_majority7_module_17__and_module_4_res), .A2(
        n_majority7_module_17__and_module_5_res), .ZN(
        n_majority7_module_17__or_module_7_res) );
  AND2_X1 u_majority7_module_17__and_module_7_U1 ( .A1(
        n_majority7_module_17__or_module_3_res), .A2(
        n_majority7_module_17__or_module_4_res), .ZN(
        n_majority7_module_17__and_module_7_res) );
  OR2_X1 u_majority7_module_17__or_module_8_U1 ( .A1(
        n_majority7_module_17__or_module_4_res), .A2(
        n_majority7_module_17__or_module_3_res), .ZN(
        n_majority7_module_17__or_module_8_res) );
  AND2_X1 u_majority7_module_17__and_module_8_U1 ( .A1(
        n_majority7_module_17__or_module_5_res), .A2(
        n_majority7_module_17__and_module_6_res), .ZN(
        n_majority7_module_17__and_module_8_res) );
  OR2_X1 u_majority7_module_17__or_module_9_U1 ( .A1(
        n_majority7_module_17__and_module_6_res), .A2(
        n_majority7_module_17__or_module_5_res), .ZN(
        n_majority7_module_17__or_module_9_res) );
  OR2_X1 u_majority7_module_17__or_module_10_U1 ( .A1(
        n_majority7_module_17__or_module_7_res), .A2(
        n_majority7_module_17__and_module_7_res), .ZN(
        n_majority7_module_17__or_module_10_res) );
  AND2_X1 u_majority7_module_17__and_module_9_U1 ( .A1(
        n_majority7_module_17__or_module_6_res), .A2(
        n_majority7_module_17__or_module_9_res), .ZN(
        n_majority7_module_17__and_module_9_res) );
  OR2_X1 u_majority7_module_17__or_module_11_U1 ( .A1(
        n_majority7_module_17__or_module_10_res), .A2(
        n_majority7_module_17__and_module_8_res), .ZN(
        n_majority7_module_17__or_module_11_res) );
  AND2_X1 u_majority7_module_17__and_module_10_U1 ( .A1(
        n_majority7_module_17__or_module_8_res), .A2(
        n_majority7_module_17__and_module_9_res), .ZN(
        n_majority7_module_17__and_module_10_res) );
  AND2_X1 u_majority7_module_17__and_module_11_U1 ( .A1(
        n_majority7_module_17__and_module_10_res), .A2(
        n_majority7_module_17__or_module_11_res), .ZN(
        n_majority7_module_17_res) );
  DFF_X1 u_reg_module_18__cini_mul_v00_reg ( .D(n_majority7_module_17_res), 
        .CK(clock_4), .Q(n_reg_module_18_res), .QN() );
  AND2_X1 u_majority7_module_18__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_18__and_module_1_res)
         );
  OR2_X1 u_majority7_module_18__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_18__or_module_1_res) );
  AND2_X1 u_majority7_module_18__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_18__and_module_2_res)
         );
  OR2_X1 u_majority7_module_18__or_module_2_U1 ( .A1(n_xor_module_33_res), 
        .A2(n_xor_module_45_res), .ZN(n_majority7_module_18__or_module_2_res)
         );
  AND2_X1 u_majority7_module_18__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_18__and_module_3_res)
         );
  OR2_X1 u_majority7_module_18__or_module_3_U1 ( .A1(n_xor_module_57_res), 
        .A2(n_xor_module_69_res), .ZN(n_majority7_module_18__or_module_3_res)
         );
  AND2_X1 u_majority7_module_18__and_module_4_U1 ( .A1(
        n_majority7_module_18__and_module_2_res), .A2(
        n_majority7_module_18__and_module_1_res), .ZN(
        n_majority7_module_18__and_module_4_res) );
  OR2_X1 u_majority7_module_18__or_module_4_U1 ( .A1(
        n_majority7_module_18__and_module_1_res), .A2(
        n_majority7_module_18__and_module_2_res), .ZN(
        n_majority7_module_18__or_module_4_res) );
  AND2_X1 u_majority7_module_18__and_module_5_U1 ( .A1(
        n_majority7_module_18__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_18__and_module_5_res) );
  OR2_X1 u_majority7_module_18__or_module_5_U1 ( .A1(n_xor_module_21_res), 
        .A2(n_majority7_module_18__and_module_3_res), .ZN(
        n_majority7_module_18__or_module_5_res) );
  AND2_X1 u_majority7_module_18__and_module_6_U1 ( .A1(
        n_majority7_module_18__or_module_1_res), .A2(
        n_majority7_module_18__or_module_2_res), .ZN(
        n_majority7_module_18__and_module_6_res) );
  OR2_X1 u_majority7_module_18__or_module_6_U1 ( .A1(
        n_majority7_module_18__or_module_2_res), .A2(
        n_majority7_module_18__or_module_1_res), .ZN(
        n_majority7_module_18__or_module_6_res) );
  OR2_X1 u_majority7_module_18__or_module_7_U1 ( .A1(
        n_majority7_module_18__and_module_4_res), .A2(
        n_majority7_module_18__and_module_5_res), .ZN(
        n_majority7_module_18__or_module_7_res) );
  AND2_X1 u_majority7_module_18__and_module_7_U1 ( .A1(
        n_majority7_module_18__or_module_3_res), .A2(
        n_majority7_module_18__or_module_4_res), .ZN(
        n_majority7_module_18__and_module_7_res) );
  OR2_X1 u_majority7_module_18__or_module_8_U1 ( .A1(
        n_majority7_module_18__or_module_4_res), .A2(
        n_majority7_module_18__or_module_3_res), .ZN(
        n_majority7_module_18__or_module_8_res) );
  AND2_X1 u_majority7_module_18__and_module_8_U1 ( .A1(
        n_majority7_module_18__or_module_5_res), .A2(
        n_majority7_module_18__and_module_6_res), .ZN(
        n_majority7_module_18__and_module_8_res) );
  OR2_X1 u_majority7_module_18__or_module_9_U1 ( .A1(
        n_majority7_module_18__and_module_6_res), .A2(
        n_majority7_module_18__or_module_5_res), .ZN(
        n_majority7_module_18__or_module_9_res) );
  OR2_X1 u_majority7_module_18__or_module_10_U1 ( .A1(
        n_majority7_module_18__or_module_7_res), .A2(
        n_majority7_module_18__and_module_7_res), .ZN(
        n_majority7_module_18__or_module_10_res) );
  AND2_X1 u_majority7_module_18__and_module_9_U1 ( .A1(
        n_majority7_module_18__or_module_6_res), .A2(
        n_majority7_module_18__or_module_9_res), .ZN(
        n_majority7_module_18__and_module_9_res) );
  OR2_X1 u_majority7_module_18__or_module_11_U1 ( .A1(
        n_majority7_module_18__or_module_10_res), .A2(
        n_majority7_module_18__and_module_8_res), .ZN(
        n_majority7_module_18__or_module_11_res) );
  AND2_X1 u_majority7_module_18__and_module_10_U1 ( .A1(
        n_majority7_module_18__or_module_8_res), .A2(
        n_majority7_module_18__and_module_9_res), .ZN(
        n_majority7_module_18__and_module_10_res) );
  AND2_X1 u_majority7_module_18__and_module_11_U1 ( .A1(
        n_majority7_module_18__and_module_10_res), .A2(
        n_majority7_module_18__or_module_11_res), .ZN(
        n_majority7_module_18_res) );
  DFF_X1 u_reg_module_19__cini_mul_v00_reg ( .D(n_majority7_module_18_res), 
        .CK(clock_4), .Q(n_reg_module_19_res), .QN() );
  AND2_X1 u_majority7_module_19__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_19__and_module_1_res)
         );
  OR2_X1 u_majority7_module_19__or_module_1_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_xor_module_84_res), .ZN(n_majority7_module_19__or_module_1_res)
         );
  AND2_X1 u_majority7_module_19__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_19__and_module_2_res)
         );
  OR2_X1 u_majority7_module_19__or_module_2_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_48_res), .ZN(n_majority7_module_19__or_module_2_res)
         );
  AND2_X1 u_majority7_module_19__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_19__and_module_3_res)
         );
  OR2_X1 u_majority7_module_19__or_module_3_U1 ( .A1(n_xor_module_60_res), 
        .A2(n_xor_module_72_res), .ZN(n_majority7_module_19__or_module_3_res)
         );
  AND2_X1 u_majority7_module_19__and_module_4_U1 ( .A1(
        n_majority7_module_19__and_module_2_res), .A2(
        n_majority7_module_19__and_module_1_res), .ZN(
        n_majority7_module_19__and_module_4_res) );
  OR2_X1 u_majority7_module_19__or_module_4_U1 ( .A1(
        n_majority7_module_19__and_module_1_res), .A2(
        n_majority7_module_19__and_module_2_res), .ZN(
        n_majority7_module_19__or_module_4_res) );
  AND2_X1 u_majority7_module_19__and_module_5_U1 ( .A1(
        n_majority7_module_19__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_19__and_module_5_res) );
  OR2_X1 u_majority7_module_19__or_module_5_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_majority7_module_19__and_module_3_res), .ZN(
        n_majority7_module_19__or_module_5_res) );
  AND2_X1 u_majority7_module_19__and_module_6_U1 ( .A1(
        n_majority7_module_19__or_module_1_res), .A2(
        n_majority7_module_19__or_module_2_res), .ZN(
        n_majority7_module_19__and_module_6_res) );
  OR2_X1 u_majority7_module_19__or_module_6_U1 ( .A1(
        n_majority7_module_19__or_module_2_res), .A2(
        n_majority7_module_19__or_module_1_res), .ZN(
        n_majority7_module_19__or_module_6_res) );
  OR2_X1 u_majority7_module_19__or_module_7_U1 ( .A1(
        n_majority7_module_19__and_module_4_res), .A2(
        n_majority7_module_19__and_module_5_res), .ZN(
        n_majority7_module_19__or_module_7_res) );
  AND2_X1 u_majority7_module_19__and_module_7_U1 ( .A1(
        n_majority7_module_19__or_module_3_res), .A2(
        n_majority7_module_19__or_module_4_res), .ZN(
        n_majority7_module_19__and_module_7_res) );
  OR2_X1 u_majority7_module_19__or_module_8_U1 ( .A1(
        n_majority7_module_19__or_module_4_res), .A2(
        n_majority7_module_19__or_module_3_res), .ZN(
        n_majority7_module_19__or_module_8_res) );
  AND2_X1 u_majority7_module_19__and_module_8_U1 ( .A1(
        n_majority7_module_19__or_module_5_res), .A2(
        n_majority7_module_19__and_module_6_res), .ZN(
        n_majority7_module_19__and_module_8_res) );
  OR2_X1 u_majority7_module_19__or_module_9_U1 ( .A1(
        n_majority7_module_19__and_module_6_res), .A2(
        n_majority7_module_19__or_module_5_res), .ZN(
        n_majority7_module_19__or_module_9_res) );
  OR2_X1 u_majority7_module_19__or_module_10_U1 ( .A1(
        n_majority7_module_19__or_module_7_res), .A2(
        n_majority7_module_19__and_module_7_res), .ZN(
        n_majority7_module_19__or_module_10_res) );
  AND2_X1 u_majority7_module_19__and_module_9_U1 ( .A1(
        n_majority7_module_19__or_module_6_res), .A2(
        n_majority7_module_19__or_module_9_res), .ZN(
        n_majority7_module_19__and_module_9_res) );
  OR2_X1 u_majority7_module_19__or_module_11_U1 ( .A1(
        n_majority7_module_19__or_module_10_res), .A2(
        n_majority7_module_19__and_module_8_res), .ZN(
        n_majority7_module_19__or_module_11_res) );
  AND2_X1 u_majority7_module_19__and_module_10_U1 ( .A1(
        n_majority7_module_19__or_module_8_res), .A2(
        n_majority7_module_19__and_module_9_res), .ZN(
        n_majority7_module_19__and_module_10_res) );
  AND2_X1 u_majority7_module_19__and_module_11_U1 ( .A1(
        n_majority7_module_19__and_module_10_res), .A2(
        n_majority7_module_19__or_module_11_res), .ZN(
        n_majority7_module_19_res) );
  DFF_X1 u_reg_module_20__cini_mul_v00_reg ( .D(n_majority7_module_19_res), 
        .CK(clock_4), .Q(n_reg_module_20_res), .QN() );
  AND2_X1 u_majority7_module_20__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_20__and_module_1_res)
         );
  OR2_X1 u_majority7_module_20__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_20__or_module_1_res) );
  AND2_X1 u_majority7_module_20__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_20__and_module_2_res)
         );
  OR2_X1 u_majority7_module_20__or_module_2_U1 ( .A1(n_xor_module_27_res), 
        .A2(n_xor_module_39_res), .ZN(n_majority7_module_20__or_module_2_res)
         );
  AND2_X1 u_majority7_module_20__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_20__and_module_3_res)
         );
  OR2_X1 u_majority7_module_20__or_module_3_U1 ( .A1(n_xor_module_51_res), 
        .A2(n_xor_module_63_res), .ZN(n_majority7_module_20__or_module_3_res)
         );
  AND2_X1 u_majority7_module_20__and_module_4_U1 ( .A1(
        n_majority7_module_20__and_module_2_res), .A2(
        n_majority7_module_20__and_module_1_res), .ZN(
        n_majority7_module_20__and_module_4_res) );
  OR2_X1 u_majority7_module_20__or_module_4_U1 ( .A1(
        n_majority7_module_20__and_module_1_res), .A2(
        n_majority7_module_20__and_module_2_res), .ZN(
        n_majority7_module_20__or_module_4_res) );
  AND2_X1 u_majority7_module_20__and_module_5_U1 ( .A1(
        n_majority7_module_20__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_20__and_module_5_res) );
  OR2_X1 u_majority7_module_20__or_module_5_U1 ( .A1(n_xor_module_15_res), 
        .A2(n_majority7_module_20__and_module_3_res), .ZN(
        n_majority7_module_20__or_module_5_res) );
  AND2_X1 u_majority7_module_20__and_module_6_U1 ( .A1(
        n_majority7_module_20__or_module_1_res), .A2(
        n_majority7_module_20__or_module_2_res), .ZN(
        n_majority7_module_20__and_module_6_res) );
  OR2_X1 u_majority7_module_20__or_module_6_U1 ( .A1(
        n_majority7_module_20__or_module_2_res), .A2(
        n_majority7_module_20__or_module_1_res), .ZN(
        n_majority7_module_20__or_module_6_res) );
  OR2_X1 u_majority7_module_20__or_module_7_U1 ( .A1(
        n_majority7_module_20__and_module_4_res), .A2(
        n_majority7_module_20__and_module_5_res), .ZN(
        n_majority7_module_20__or_module_7_res) );
  AND2_X1 u_majority7_module_20__and_module_7_U1 ( .A1(
        n_majority7_module_20__or_module_3_res), .A2(
        n_majority7_module_20__or_module_4_res), .ZN(
        n_majority7_module_20__and_module_7_res) );
  OR2_X1 u_majority7_module_20__or_module_8_U1 ( .A1(
        n_majority7_module_20__or_module_4_res), .A2(
        n_majority7_module_20__or_module_3_res), .ZN(
        n_majority7_module_20__or_module_8_res) );
  AND2_X1 u_majority7_module_20__and_module_8_U1 ( .A1(
        n_majority7_module_20__or_module_5_res), .A2(
        n_majority7_module_20__and_module_6_res), .ZN(
        n_majority7_module_20__and_module_8_res) );
  OR2_X1 u_majority7_module_20__or_module_9_U1 ( .A1(
        n_majority7_module_20__and_module_6_res), .A2(
        n_majority7_module_20__or_module_5_res), .ZN(
        n_majority7_module_20__or_module_9_res) );
  OR2_X1 u_majority7_module_20__or_module_10_U1 ( .A1(
        n_majority7_module_20__or_module_7_res), .A2(
        n_majority7_module_20__and_module_7_res), .ZN(
        n_majority7_module_20__or_module_10_res) );
  AND2_X1 u_majority7_module_20__and_module_9_U1 ( .A1(
        n_majority7_module_20__or_module_6_res), .A2(
        n_majority7_module_20__or_module_9_res), .ZN(
        n_majority7_module_20__and_module_9_res) );
  OR2_X1 u_majority7_module_20__or_module_11_U1 ( .A1(
        n_majority7_module_20__or_module_10_res), .A2(
        n_majority7_module_20__and_module_8_res), .ZN(
        n_majority7_module_20__or_module_11_res) );
  AND2_X1 u_majority7_module_20__and_module_10_U1 ( .A1(
        n_majority7_module_20__or_module_8_res), .A2(
        n_majority7_module_20__and_module_9_res), .ZN(
        n_majority7_module_20__and_module_10_res) );
  AND2_X1 u_majority7_module_20__and_module_11_U1 ( .A1(
        n_majority7_module_20__and_module_10_res), .A2(
        n_majority7_module_20__or_module_11_res), .ZN(
        n_majority7_module_20_res) );
  DFF_X1 u_reg_module_21__cini_mul_v00_reg ( .D(n_majority7_module_20_res), 
        .CK(clock_5), .Q(n_reg_module_21_res), .QN() );
  AND2_X1 u_majority7_module_21__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_21__and_module_1_res)
         );
  OR2_X1 u_majority7_module_21__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_21__or_module_1_res) );
  AND2_X1 u_majority7_module_21__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_21__and_module_2_res)
         );
  OR2_X1 u_majority7_module_21__or_module_2_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_42_res), .ZN(n_majority7_module_21__or_module_2_res)
         );
  AND2_X1 u_majority7_module_21__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_21__and_module_3_res)
         );
  OR2_X1 u_majority7_module_21__or_module_3_U1 ( .A1(n_xor_module_54_res), 
        .A2(n_xor_module_66_res), .ZN(n_majority7_module_21__or_module_3_res)
         );
  AND2_X1 u_majority7_module_21__and_module_4_U1 ( .A1(
        n_majority7_module_21__and_module_2_res), .A2(
        n_majority7_module_21__and_module_1_res), .ZN(
        n_majority7_module_21__and_module_4_res) );
  OR2_X1 u_majority7_module_21__or_module_4_U1 ( .A1(
        n_majority7_module_21__and_module_1_res), .A2(
        n_majority7_module_21__and_module_2_res), .ZN(
        n_majority7_module_21__or_module_4_res) );
  AND2_X1 u_majority7_module_21__and_module_5_U1 ( .A1(
        n_majority7_module_21__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_21__and_module_5_res) );
  OR2_X1 u_majority7_module_21__or_module_5_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_majority7_module_21__and_module_3_res), .ZN(
        n_majority7_module_21__or_module_5_res) );
  AND2_X1 u_majority7_module_21__and_module_6_U1 ( .A1(
        n_majority7_module_21__or_module_1_res), .A2(
        n_majority7_module_21__or_module_2_res), .ZN(
        n_majority7_module_21__and_module_6_res) );
  OR2_X1 u_majority7_module_21__or_module_6_U1 ( .A1(
        n_majority7_module_21__or_module_2_res), .A2(
        n_majority7_module_21__or_module_1_res), .ZN(
        n_majority7_module_21__or_module_6_res) );
  OR2_X1 u_majority7_module_21__or_module_7_U1 ( .A1(
        n_majority7_module_21__and_module_4_res), .A2(
        n_majority7_module_21__and_module_5_res), .ZN(
        n_majority7_module_21__or_module_7_res) );
  AND2_X1 u_majority7_module_21__and_module_7_U1 ( .A1(
        n_majority7_module_21__or_module_3_res), .A2(
        n_majority7_module_21__or_module_4_res), .ZN(
        n_majority7_module_21__and_module_7_res) );
  OR2_X1 u_majority7_module_21__or_module_8_U1 ( .A1(
        n_majority7_module_21__or_module_4_res), .A2(
        n_majority7_module_21__or_module_3_res), .ZN(
        n_majority7_module_21__or_module_8_res) );
  AND2_X1 u_majority7_module_21__and_module_8_U1 ( .A1(
        n_majority7_module_21__or_module_5_res), .A2(
        n_majority7_module_21__and_module_6_res), .ZN(
        n_majority7_module_21__and_module_8_res) );
  OR2_X1 u_majority7_module_21__or_module_9_U1 ( .A1(
        n_majority7_module_21__and_module_6_res), .A2(
        n_majority7_module_21__or_module_5_res), .ZN(
        n_majority7_module_21__or_module_9_res) );
  OR2_X1 u_majority7_module_21__or_module_10_U1 ( .A1(
        n_majority7_module_21__or_module_7_res), .A2(
        n_majority7_module_21__and_module_7_res), .ZN(
        n_majority7_module_21__or_module_10_res) );
  AND2_X1 u_majority7_module_21__and_module_9_U1 ( .A1(
        n_majority7_module_21__or_module_6_res), .A2(
        n_majority7_module_21__or_module_9_res), .ZN(
        n_majority7_module_21__and_module_9_res) );
  OR2_X1 u_majority7_module_21__or_module_11_U1 ( .A1(
        n_majority7_module_21__or_module_10_res), .A2(
        n_majority7_module_21__and_module_8_res), .ZN(
        n_majority7_module_21__or_module_11_res) );
  AND2_X1 u_majority7_module_21__and_module_10_U1 ( .A1(
        n_majority7_module_21__or_module_8_res), .A2(
        n_majority7_module_21__and_module_9_res), .ZN(
        n_majority7_module_21__and_module_10_res) );
  AND2_X1 u_majority7_module_21__and_module_11_U1 ( .A1(
        n_majority7_module_21__and_module_10_res), .A2(
        n_majority7_module_21__or_module_11_res), .ZN(
        n_majority7_module_21_res) );
  DFF_X1 u_reg_module_22__cini_mul_v00_reg ( .D(n_majority7_module_21_res), 
        .CK(clock_5), .Q(n_reg_module_22_res), .QN() );
  AND2_X1 u_majority7_module_22__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_22__and_module_1_res)
         );
  OR2_X1 u_majority7_module_22__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_22__or_module_1_res) );
  AND2_X1 u_majority7_module_22__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_22__and_module_2_res)
         );
  OR2_X1 u_majority7_module_22__or_module_2_U1 ( .A1(n_xor_module_33_res), 
        .A2(n_xor_module_45_res), .ZN(n_majority7_module_22__or_module_2_res)
         );
  AND2_X1 u_majority7_module_22__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_22__and_module_3_res)
         );
  OR2_X1 u_majority7_module_22__or_module_3_U1 ( .A1(n_xor_module_57_res), 
        .A2(n_xor_module_69_res), .ZN(n_majority7_module_22__or_module_3_res)
         );
  AND2_X1 u_majority7_module_22__and_module_4_U1 ( .A1(
        n_majority7_module_22__and_module_2_res), .A2(
        n_majority7_module_22__and_module_1_res), .ZN(
        n_majority7_module_22__and_module_4_res) );
  OR2_X1 u_majority7_module_22__or_module_4_U1 ( .A1(
        n_majority7_module_22__and_module_1_res), .A2(
        n_majority7_module_22__and_module_2_res), .ZN(
        n_majority7_module_22__or_module_4_res) );
  AND2_X1 u_majority7_module_22__and_module_5_U1 ( .A1(
        n_majority7_module_22__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_22__and_module_5_res) );
  OR2_X1 u_majority7_module_22__or_module_5_U1 ( .A1(n_xor_module_21_res), 
        .A2(n_majority7_module_22__and_module_3_res), .ZN(
        n_majority7_module_22__or_module_5_res) );
  AND2_X1 u_majority7_module_22__and_module_6_U1 ( .A1(
        n_majority7_module_22__or_module_1_res), .A2(
        n_majority7_module_22__or_module_2_res), .ZN(
        n_majority7_module_22__and_module_6_res) );
  OR2_X1 u_majority7_module_22__or_module_6_U1 ( .A1(
        n_majority7_module_22__or_module_2_res), .A2(
        n_majority7_module_22__or_module_1_res), .ZN(
        n_majority7_module_22__or_module_6_res) );
  OR2_X1 u_majority7_module_22__or_module_7_U1 ( .A1(
        n_majority7_module_22__and_module_4_res), .A2(
        n_majority7_module_22__and_module_5_res), .ZN(
        n_majority7_module_22__or_module_7_res) );
  AND2_X1 u_majority7_module_22__and_module_7_U1 ( .A1(
        n_majority7_module_22__or_module_3_res), .A2(
        n_majority7_module_22__or_module_4_res), .ZN(
        n_majority7_module_22__and_module_7_res) );
  OR2_X1 u_majority7_module_22__or_module_8_U1 ( .A1(
        n_majority7_module_22__or_module_4_res), .A2(
        n_majority7_module_22__or_module_3_res), .ZN(
        n_majority7_module_22__or_module_8_res) );
  AND2_X1 u_majority7_module_22__and_module_8_U1 ( .A1(
        n_majority7_module_22__or_module_5_res), .A2(
        n_majority7_module_22__and_module_6_res), .ZN(
        n_majority7_module_22__and_module_8_res) );
  OR2_X1 u_majority7_module_22__or_module_9_U1 ( .A1(
        n_majority7_module_22__and_module_6_res), .A2(
        n_majority7_module_22__or_module_5_res), .ZN(
        n_majority7_module_22__or_module_9_res) );
  OR2_X1 u_majority7_module_22__or_module_10_U1 ( .A1(
        n_majority7_module_22__or_module_7_res), .A2(
        n_majority7_module_22__and_module_7_res), .ZN(
        n_majority7_module_22__or_module_10_res) );
  AND2_X1 u_majority7_module_22__and_module_9_U1 ( .A1(
        n_majority7_module_22__or_module_6_res), .A2(
        n_majority7_module_22__or_module_9_res), .ZN(
        n_majority7_module_22__and_module_9_res) );
  OR2_X1 u_majority7_module_22__or_module_11_U1 ( .A1(
        n_majority7_module_22__or_module_10_res), .A2(
        n_majority7_module_22__and_module_8_res), .ZN(
        n_majority7_module_22__or_module_11_res) );
  AND2_X1 u_majority7_module_22__and_module_10_U1 ( .A1(
        n_majority7_module_22__or_module_8_res), .A2(
        n_majority7_module_22__and_module_9_res), .ZN(
        n_majority7_module_22__and_module_10_res) );
  AND2_X1 u_majority7_module_22__and_module_11_U1 ( .A1(
        n_majority7_module_22__and_module_10_res), .A2(
        n_majority7_module_22__or_module_11_res), .ZN(
        n_majority7_module_22_res) );
  DFF_X1 u_reg_module_23__cini_mul_v00_reg ( .D(n_majority7_module_22_res), 
        .CK(clock_5), .Q(n_reg_module_23_res), .QN() );
  AND2_X1 u_majority7_module_23__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_23__and_module_1_res)
         );
  OR2_X1 u_majority7_module_23__or_module_1_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_xor_module_84_res), .ZN(n_majority7_module_23__or_module_1_res)
         );
  AND2_X1 u_majority7_module_23__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_23__and_module_2_res)
         );
  OR2_X1 u_majority7_module_23__or_module_2_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_48_res), .ZN(n_majority7_module_23__or_module_2_res)
         );
  AND2_X1 u_majority7_module_23__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_23__and_module_3_res)
         );
  OR2_X1 u_majority7_module_23__or_module_3_U1 ( .A1(n_xor_module_60_res), 
        .A2(n_xor_module_72_res), .ZN(n_majority7_module_23__or_module_3_res)
         );
  AND2_X1 u_majority7_module_23__and_module_4_U1 ( .A1(
        n_majority7_module_23__and_module_2_res), .A2(
        n_majority7_module_23__and_module_1_res), .ZN(
        n_majority7_module_23__and_module_4_res) );
  OR2_X1 u_majority7_module_23__or_module_4_U1 ( .A1(
        n_majority7_module_23__and_module_1_res), .A2(
        n_majority7_module_23__and_module_2_res), .ZN(
        n_majority7_module_23__or_module_4_res) );
  AND2_X1 u_majority7_module_23__and_module_5_U1 ( .A1(
        n_majority7_module_23__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_23__and_module_5_res) );
  OR2_X1 u_majority7_module_23__or_module_5_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_majority7_module_23__and_module_3_res), .ZN(
        n_majority7_module_23__or_module_5_res) );
  AND2_X1 u_majority7_module_23__and_module_6_U1 ( .A1(
        n_majority7_module_23__or_module_1_res), .A2(
        n_majority7_module_23__or_module_2_res), .ZN(
        n_majority7_module_23__and_module_6_res) );
  OR2_X1 u_majority7_module_23__or_module_6_U1 ( .A1(
        n_majority7_module_23__or_module_2_res), .A2(
        n_majority7_module_23__or_module_1_res), .ZN(
        n_majority7_module_23__or_module_6_res) );
  OR2_X1 u_majority7_module_23__or_module_7_U1 ( .A1(
        n_majority7_module_23__and_module_4_res), .A2(
        n_majority7_module_23__and_module_5_res), .ZN(
        n_majority7_module_23__or_module_7_res) );
  AND2_X1 u_majority7_module_23__and_module_7_U1 ( .A1(
        n_majority7_module_23__or_module_3_res), .A2(
        n_majority7_module_23__or_module_4_res), .ZN(
        n_majority7_module_23__and_module_7_res) );
  OR2_X1 u_majority7_module_23__or_module_8_U1 ( .A1(
        n_majority7_module_23__or_module_4_res), .A2(
        n_majority7_module_23__or_module_3_res), .ZN(
        n_majority7_module_23__or_module_8_res) );
  AND2_X1 u_majority7_module_23__and_module_8_U1 ( .A1(
        n_majority7_module_23__or_module_5_res), .A2(
        n_majority7_module_23__and_module_6_res), .ZN(
        n_majority7_module_23__and_module_8_res) );
  OR2_X1 u_majority7_module_23__or_module_9_U1 ( .A1(
        n_majority7_module_23__and_module_6_res), .A2(
        n_majority7_module_23__or_module_5_res), .ZN(
        n_majority7_module_23__or_module_9_res) );
  OR2_X1 u_majority7_module_23__or_module_10_U1 ( .A1(
        n_majority7_module_23__or_module_7_res), .A2(
        n_majority7_module_23__and_module_7_res), .ZN(
        n_majority7_module_23__or_module_10_res) );
  AND2_X1 u_majority7_module_23__and_module_9_U1 ( .A1(
        n_majority7_module_23__or_module_6_res), .A2(
        n_majority7_module_23__or_module_9_res), .ZN(
        n_majority7_module_23__and_module_9_res) );
  OR2_X1 u_majority7_module_23__or_module_11_U1 ( .A1(
        n_majority7_module_23__or_module_10_res), .A2(
        n_majority7_module_23__and_module_8_res), .ZN(
        n_majority7_module_23__or_module_11_res) );
  AND2_X1 u_majority7_module_23__and_module_10_U1 ( .A1(
        n_majority7_module_23__or_module_8_res), .A2(
        n_majority7_module_23__and_module_9_res), .ZN(
        n_majority7_module_23__and_module_10_res) );
  AND2_X1 u_majority7_module_23__and_module_11_U1 ( .A1(
        n_majority7_module_23__and_module_10_res), .A2(
        n_majority7_module_23__or_module_11_res), .ZN(
        n_majority7_module_23_res) );
  DFF_X1 u_reg_module_24__cini_mul_v00_reg ( .D(n_majority7_module_23_res), 
        .CK(clock_5), .Q(n_reg_module_24_res), .QN() );
  AND2_X1 u_majority7_module_24__and_module_1_U1 ( .A1(n_xor_module_75_res), 
        .A2(n_xor_module_3_res), .ZN(n_majority7_module_24__and_module_1_res)
         );
  OR2_X1 u_majority7_module_24__or_module_1_U1 ( .A1(n_xor_module_3_res), .A2(
        n_xor_module_75_res), .ZN(n_majority7_module_24__or_module_1_res) );
  AND2_X1 u_majority7_module_24__and_module_2_U1 ( .A1(n_xor_module_39_res), 
        .A2(n_xor_module_27_res), .ZN(n_majority7_module_24__and_module_2_res)
         );
  OR2_X1 u_majority7_module_24__or_module_2_U1 ( .A1(n_xor_module_27_res), 
        .A2(n_xor_module_39_res), .ZN(n_majority7_module_24__or_module_2_res)
         );
  AND2_X1 u_majority7_module_24__and_module_3_U1 ( .A1(n_xor_module_63_res), 
        .A2(n_xor_module_51_res), .ZN(n_majority7_module_24__and_module_3_res)
         );
  OR2_X1 u_majority7_module_24__or_module_3_U1 ( .A1(n_xor_module_51_res), 
        .A2(n_xor_module_63_res), .ZN(n_majority7_module_24__or_module_3_res)
         );
  AND2_X1 u_majority7_module_24__and_module_4_U1 ( .A1(
        n_majority7_module_24__and_module_2_res), .A2(
        n_majority7_module_24__and_module_1_res), .ZN(
        n_majority7_module_24__and_module_4_res) );
  OR2_X1 u_majority7_module_24__or_module_4_U1 ( .A1(
        n_majority7_module_24__and_module_1_res), .A2(
        n_majority7_module_24__and_module_2_res), .ZN(
        n_majority7_module_24__or_module_4_res) );
  AND2_X1 u_majority7_module_24__and_module_5_U1 ( .A1(
        n_majority7_module_24__and_module_3_res), .A2(n_xor_module_15_res), 
        .ZN(n_majority7_module_24__and_module_5_res) );
  OR2_X1 u_majority7_module_24__or_module_5_U1 ( .A1(n_xor_module_15_res), 
        .A2(n_majority7_module_24__and_module_3_res), .ZN(
        n_majority7_module_24__or_module_5_res) );
  AND2_X1 u_majority7_module_24__and_module_6_U1 ( .A1(
        n_majority7_module_24__or_module_1_res), .A2(
        n_majority7_module_24__or_module_2_res), .ZN(
        n_majority7_module_24__and_module_6_res) );
  OR2_X1 u_majority7_module_24__or_module_6_U1 ( .A1(
        n_majority7_module_24__or_module_2_res), .A2(
        n_majority7_module_24__or_module_1_res), .ZN(
        n_majority7_module_24__or_module_6_res) );
  OR2_X1 u_majority7_module_24__or_module_7_U1 ( .A1(
        n_majority7_module_24__and_module_4_res), .A2(
        n_majority7_module_24__and_module_5_res), .ZN(
        n_majority7_module_24__or_module_7_res) );
  AND2_X1 u_majority7_module_24__and_module_7_U1 ( .A1(
        n_majority7_module_24__or_module_3_res), .A2(
        n_majority7_module_24__or_module_4_res), .ZN(
        n_majority7_module_24__and_module_7_res) );
  OR2_X1 u_majority7_module_24__or_module_8_U1 ( .A1(
        n_majority7_module_24__or_module_4_res), .A2(
        n_majority7_module_24__or_module_3_res), .ZN(
        n_majority7_module_24__or_module_8_res) );
  AND2_X1 u_majority7_module_24__and_module_8_U1 ( .A1(
        n_majority7_module_24__or_module_5_res), .A2(
        n_majority7_module_24__and_module_6_res), .ZN(
        n_majority7_module_24__and_module_8_res) );
  OR2_X1 u_majority7_module_24__or_module_9_U1 ( .A1(
        n_majority7_module_24__and_module_6_res), .A2(
        n_majority7_module_24__or_module_5_res), .ZN(
        n_majority7_module_24__or_module_9_res) );
  OR2_X1 u_majority7_module_24__or_module_10_U1 ( .A1(
        n_majority7_module_24__or_module_7_res), .A2(
        n_majority7_module_24__and_module_7_res), .ZN(
        n_majority7_module_24__or_module_10_res) );
  AND2_X1 u_majority7_module_24__and_module_9_U1 ( .A1(
        n_majority7_module_24__or_module_6_res), .A2(
        n_majority7_module_24__or_module_9_res), .ZN(
        n_majority7_module_24__and_module_9_res) );
  OR2_X1 u_majority7_module_24__or_module_11_U1 ( .A1(
        n_majority7_module_24__or_module_10_res), .A2(
        n_majority7_module_24__and_module_8_res), .ZN(
        n_majority7_module_24__or_module_11_res) );
  AND2_X1 u_majority7_module_24__and_module_10_U1 ( .A1(
        n_majority7_module_24__or_module_8_res), .A2(
        n_majority7_module_24__and_module_9_res), .ZN(
        n_majority7_module_24__and_module_10_res) );
  AND2_X1 u_majority7_module_24__and_module_11_U1 ( .A1(
        n_majority7_module_24__and_module_10_res), .A2(
        n_majority7_module_24__or_module_11_res), .ZN(
        n_majority7_module_24_res) );
  DFF_X1 u_reg_module_25__cini_mul_v00_reg ( .D(n_majority7_module_24_res), 
        .CK(clock_6), .Q(n_reg_module_25_res), .QN() );
  AND2_X1 u_majority7_module_25__and_module_1_U1 ( .A1(n_xor_module_78_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_25__and_module_1_res)
         );
  OR2_X1 u_majority7_module_25__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_78_res), .ZN(n_majority7_module_25__or_module_1_res) );
  AND2_X1 u_majority7_module_25__and_module_2_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_25__and_module_2_res)
         );
  OR2_X1 u_majority7_module_25__or_module_2_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_42_res), .ZN(n_majority7_module_25__or_module_2_res)
         );
  AND2_X1 u_majority7_module_25__and_module_3_U1 ( .A1(n_xor_module_66_res), 
        .A2(n_xor_module_54_res), .ZN(n_majority7_module_25__and_module_3_res)
         );
  OR2_X1 u_majority7_module_25__or_module_3_U1 ( .A1(n_xor_module_54_res), 
        .A2(n_xor_module_66_res), .ZN(n_majority7_module_25__or_module_3_res)
         );
  AND2_X1 u_majority7_module_25__and_module_4_U1 ( .A1(
        n_majority7_module_25__and_module_2_res), .A2(
        n_majority7_module_25__and_module_1_res), .ZN(
        n_majority7_module_25__and_module_4_res) );
  OR2_X1 u_majority7_module_25__or_module_4_U1 ( .A1(
        n_majority7_module_25__and_module_1_res), .A2(
        n_majority7_module_25__and_module_2_res), .ZN(
        n_majority7_module_25__or_module_4_res) );
  AND2_X1 u_majority7_module_25__and_module_5_U1 ( .A1(
        n_majority7_module_25__and_module_3_res), .A2(n_xor_module_18_res), 
        .ZN(n_majority7_module_25__and_module_5_res) );
  OR2_X1 u_majority7_module_25__or_module_5_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_majority7_module_25__and_module_3_res), .ZN(
        n_majority7_module_25__or_module_5_res) );
  AND2_X1 u_majority7_module_25__and_module_6_U1 ( .A1(
        n_majority7_module_25__or_module_1_res), .A2(
        n_majority7_module_25__or_module_2_res), .ZN(
        n_majority7_module_25__and_module_6_res) );
  OR2_X1 u_majority7_module_25__or_module_6_U1 ( .A1(
        n_majority7_module_25__or_module_2_res), .A2(
        n_majority7_module_25__or_module_1_res), .ZN(
        n_majority7_module_25__or_module_6_res) );
  OR2_X1 u_majority7_module_25__or_module_7_U1 ( .A1(
        n_majority7_module_25__and_module_4_res), .A2(
        n_majority7_module_25__and_module_5_res), .ZN(
        n_majority7_module_25__or_module_7_res) );
  AND2_X1 u_majority7_module_25__and_module_7_U1 ( .A1(
        n_majority7_module_25__or_module_3_res), .A2(
        n_majority7_module_25__or_module_4_res), .ZN(
        n_majority7_module_25__and_module_7_res) );
  OR2_X1 u_majority7_module_25__or_module_8_U1 ( .A1(
        n_majority7_module_25__or_module_4_res), .A2(
        n_majority7_module_25__or_module_3_res), .ZN(
        n_majority7_module_25__or_module_8_res) );
  AND2_X1 u_majority7_module_25__and_module_8_U1 ( .A1(
        n_majority7_module_25__or_module_5_res), .A2(
        n_majority7_module_25__and_module_6_res), .ZN(
        n_majority7_module_25__and_module_8_res) );
  OR2_X1 u_majority7_module_25__or_module_9_U1 ( .A1(
        n_majority7_module_25__and_module_6_res), .A2(
        n_majority7_module_25__or_module_5_res), .ZN(
        n_majority7_module_25__or_module_9_res) );
  OR2_X1 u_majority7_module_25__or_module_10_U1 ( .A1(
        n_majority7_module_25__or_module_7_res), .A2(
        n_majority7_module_25__and_module_7_res), .ZN(
        n_majority7_module_25__or_module_10_res) );
  AND2_X1 u_majority7_module_25__and_module_9_U1 ( .A1(
        n_majority7_module_25__or_module_6_res), .A2(
        n_majority7_module_25__or_module_9_res), .ZN(
        n_majority7_module_25__and_module_9_res) );
  OR2_X1 u_majority7_module_25__or_module_11_U1 ( .A1(
        n_majority7_module_25__or_module_10_res), .A2(
        n_majority7_module_25__and_module_8_res), .ZN(
        n_majority7_module_25__or_module_11_res) );
  AND2_X1 u_majority7_module_25__and_module_10_U1 ( .A1(
        n_majority7_module_25__or_module_8_res), .A2(
        n_majority7_module_25__and_module_9_res), .ZN(
        n_majority7_module_25__and_module_10_res) );
  AND2_X1 u_majority7_module_25__and_module_11_U1 ( .A1(
        n_majority7_module_25__and_module_10_res), .A2(
        n_majority7_module_25__or_module_11_res), .ZN(
        n_majority7_module_25_res) );
  DFF_X1 u_reg_module_26__cini_mul_v00_reg ( .D(n_majority7_module_25_res), 
        .CK(clock_6), .Q(n_reg_module_26_res), .QN() );
  AND2_X1 u_majority7_module_26__and_module_1_U1 ( .A1(n_xor_module_81_res), 
        .A2(n_xor_module_9_res), .ZN(n_majority7_module_26__and_module_1_res)
         );
  OR2_X1 u_majority7_module_26__or_module_1_U1 ( .A1(n_xor_module_9_res), .A2(
        n_xor_module_81_res), .ZN(n_majority7_module_26__or_module_1_res) );
  AND2_X1 u_majority7_module_26__and_module_2_U1 ( .A1(n_xor_module_45_res), 
        .A2(n_xor_module_33_res), .ZN(n_majority7_module_26__and_module_2_res)
         );
  OR2_X1 u_majority7_module_26__or_module_2_U1 ( .A1(n_xor_module_33_res), 
        .A2(n_xor_module_45_res), .ZN(n_majority7_module_26__or_module_2_res)
         );
  AND2_X1 u_majority7_module_26__and_module_3_U1 ( .A1(n_xor_module_69_res), 
        .A2(n_xor_module_57_res), .ZN(n_majority7_module_26__and_module_3_res)
         );
  OR2_X1 u_majority7_module_26__or_module_3_U1 ( .A1(n_xor_module_57_res), 
        .A2(n_xor_module_69_res), .ZN(n_majority7_module_26__or_module_3_res)
         );
  AND2_X1 u_majority7_module_26__and_module_4_U1 ( .A1(
        n_majority7_module_26__and_module_2_res), .A2(
        n_majority7_module_26__and_module_1_res), .ZN(
        n_majority7_module_26__and_module_4_res) );
  OR2_X1 u_majority7_module_26__or_module_4_U1 ( .A1(
        n_majority7_module_26__and_module_1_res), .A2(
        n_majority7_module_26__and_module_2_res), .ZN(
        n_majority7_module_26__or_module_4_res) );
  AND2_X1 u_majority7_module_26__and_module_5_U1 ( .A1(
        n_majority7_module_26__and_module_3_res), .A2(n_xor_module_21_res), 
        .ZN(n_majority7_module_26__and_module_5_res) );
  OR2_X1 u_majority7_module_26__or_module_5_U1 ( .A1(n_xor_module_21_res), 
        .A2(n_majority7_module_26__and_module_3_res), .ZN(
        n_majority7_module_26__or_module_5_res) );
  AND2_X1 u_majority7_module_26__and_module_6_U1 ( .A1(
        n_majority7_module_26__or_module_1_res), .A2(
        n_majority7_module_26__or_module_2_res), .ZN(
        n_majority7_module_26__and_module_6_res) );
  OR2_X1 u_majority7_module_26__or_module_6_U1 ( .A1(
        n_majority7_module_26__or_module_2_res), .A2(
        n_majority7_module_26__or_module_1_res), .ZN(
        n_majority7_module_26__or_module_6_res) );
  OR2_X1 u_majority7_module_26__or_module_7_U1 ( .A1(
        n_majority7_module_26__and_module_4_res), .A2(
        n_majority7_module_26__and_module_5_res), .ZN(
        n_majority7_module_26__or_module_7_res) );
  AND2_X1 u_majority7_module_26__and_module_7_U1 ( .A1(
        n_majority7_module_26__or_module_3_res), .A2(
        n_majority7_module_26__or_module_4_res), .ZN(
        n_majority7_module_26__and_module_7_res) );
  OR2_X1 u_majority7_module_26__or_module_8_U1 ( .A1(
        n_majority7_module_26__or_module_4_res), .A2(
        n_majority7_module_26__or_module_3_res), .ZN(
        n_majority7_module_26__or_module_8_res) );
  AND2_X1 u_majority7_module_26__and_module_8_U1 ( .A1(
        n_majority7_module_26__or_module_5_res), .A2(
        n_majority7_module_26__and_module_6_res), .ZN(
        n_majority7_module_26__and_module_8_res) );
  OR2_X1 u_majority7_module_26__or_module_9_U1 ( .A1(
        n_majority7_module_26__and_module_6_res), .A2(
        n_majority7_module_26__or_module_5_res), .ZN(
        n_majority7_module_26__or_module_9_res) );
  OR2_X1 u_majority7_module_26__or_module_10_U1 ( .A1(
        n_majority7_module_26__or_module_7_res), .A2(
        n_majority7_module_26__and_module_7_res), .ZN(
        n_majority7_module_26__or_module_10_res) );
  AND2_X1 u_majority7_module_26__and_module_9_U1 ( .A1(
        n_majority7_module_26__or_module_6_res), .A2(
        n_majority7_module_26__or_module_9_res), .ZN(
        n_majority7_module_26__and_module_9_res) );
  OR2_X1 u_majority7_module_26__or_module_11_U1 ( .A1(
        n_majority7_module_26__or_module_10_res), .A2(
        n_majority7_module_26__and_module_8_res), .ZN(
        n_majority7_module_26__or_module_11_res) );
  AND2_X1 u_majority7_module_26__and_module_10_U1 ( .A1(
        n_majority7_module_26__or_module_8_res), .A2(
        n_majority7_module_26__and_module_9_res), .ZN(
        n_majority7_module_26__and_module_10_res) );
  AND2_X1 u_majority7_module_26__and_module_11_U1 ( .A1(
        n_majority7_module_26__and_module_10_res), .A2(
        n_majority7_module_26__or_module_11_res), .ZN(
        n_majority7_module_26_res) );
  DFF_X1 u_reg_module_27__cini_mul_v00_reg ( .D(n_majority7_module_26_res), 
        .CK(clock_6), .Q(n_reg_module_27_res), .QN() );
  AND2_X1 u_majority7_module_27__and_module_1_U1 ( .A1(n_xor_module_84_res), 
        .A2(n_xor_module_12_res), .ZN(n_majority7_module_27__and_module_1_res)
         );
  OR2_X1 u_majority7_module_27__or_module_1_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_xor_module_84_res), .ZN(n_majority7_module_27__or_module_1_res)
         );
  AND2_X1 u_majority7_module_27__and_module_2_U1 ( .A1(n_xor_module_48_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_27__and_module_2_res)
         );
  OR2_X1 u_majority7_module_27__or_module_2_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_48_res), .ZN(n_majority7_module_27__or_module_2_res)
         );
  AND2_X1 u_majority7_module_27__and_module_3_U1 ( .A1(n_xor_module_72_res), 
        .A2(n_xor_module_60_res), .ZN(n_majority7_module_27__and_module_3_res)
         );
  OR2_X1 u_majority7_module_27__or_module_3_U1 ( .A1(n_xor_module_60_res), 
        .A2(n_xor_module_72_res), .ZN(n_majority7_module_27__or_module_3_res)
         );
  AND2_X1 u_majority7_module_27__and_module_4_U1 ( .A1(
        n_majority7_module_27__and_module_2_res), .A2(
        n_majority7_module_27__and_module_1_res), .ZN(
        n_majority7_module_27__and_module_4_res) );
  OR2_X1 u_majority7_module_27__or_module_4_U1 ( .A1(
        n_majority7_module_27__and_module_1_res), .A2(
        n_majority7_module_27__and_module_2_res), .ZN(
        n_majority7_module_27__or_module_4_res) );
  AND2_X1 u_majority7_module_27__and_module_5_U1 ( .A1(
        n_majority7_module_27__and_module_3_res), .A2(n_xor_module_24_res), 
        .ZN(n_majority7_module_27__and_module_5_res) );
  OR2_X1 u_majority7_module_27__or_module_5_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_majority7_module_27__and_module_3_res), .ZN(
        n_majority7_module_27__or_module_5_res) );
  AND2_X1 u_majority7_module_27__and_module_6_U1 ( .A1(
        n_majority7_module_27__or_module_1_res), .A2(
        n_majority7_module_27__or_module_2_res), .ZN(
        n_majority7_module_27__and_module_6_res) );
  OR2_X1 u_majority7_module_27__or_module_6_U1 ( .A1(
        n_majority7_module_27__or_module_2_res), .A2(
        n_majority7_module_27__or_module_1_res), .ZN(
        n_majority7_module_27__or_module_6_res) );
  OR2_X1 u_majority7_module_27__or_module_7_U1 ( .A1(
        n_majority7_module_27__and_module_4_res), .A2(
        n_majority7_module_27__and_module_5_res), .ZN(
        n_majority7_module_27__or_module_7_res) );
  AND2_X1 u_majority7_module_27__and_module_7_U1 ( .A1(
        n_majority7_module_27__or_module_3_res), .A2(
        n_majority7_module_27__or_module_4_res), .ZN(
        n_majority7_module_27__and_module_7_res) );
  OR2_X1 u_majority7_module_27__or_module_8_U1 ( .A1(
        n_majority7_module_27__or_module_4_res), .A2(
        n_majority7_module_27__or_module_3_res), .ZN(
        n_majority7_module_27__or_module_8_res) );
  AND2_X1 u_majority7_module_27__and_module_8_U1 ( .A1(
        n_majority7_module_27__or_module_5_res), .A2(
        n_majority7_module_27__and_module_6_res), .ZN(
        n_majority7_module_27__and_module_8_res) );
  OR2_X1 u_majority7_module_27__or_module_9_U1 ( .A1(
        n_majority7_module_27__and_module_6_res), .A2(
        n_majority7_module_27__or_module_5_res), .ZN(
        n_majority7_module_27__or_module_9_res) );
  OR2_X1 u_majority7_module_27__or_module_10_U1 ( .A1(
        n_majority7_module_27__or_module_7_res), .A2(
        n_majority7_module_27__and_module_7_res), .ZN(
        n_majority7_module_27__or_module_10_res) );
  AND2_X1 u_majority7_module_27__and_module_9_U1 ( .A1(
        n_majority7_module_27__or_module_6_res), .A2(
        n_majority7_module_27__or_module_9_res), .ZN(
        n_majority7_module_27__and_module_9_res) );
  OR2_X1 u_majority7_module_27__or_module_11_U1 ( .A1(
        n_majority7_module_27__or_module_10_res), .A2(
        n_majority7_module_27__and_module_8_res), .ZN(
        n_majority7_module_27__or_module_11_res) );
  AND2_X1 u_majority7_module_27__and_module_10_U1 ( .A1(
        n_majority7_module_27__or_module_8_res), .A2(
        n_majority7_module_27__and_module_9_res), .ZN(
        n_majority7_module_27__and_module_10_res) );
  AND2_X1 u_majority7_module_27__and_module_11_U1 ( .A1(
        n_majority7_module_27__and_module_10_res), .A2(
        n_majority7_module_27__or_module_11_res), .ZN(
        n_majority7_module_27_res) );
  DFF_X1 u_reg_module_28__cini_mul_v00_reg ( .D(n_majority7_module_27_res), 
        .CK(clock_6), .Q(n_reg_module_28_res), .QN() );
  AND2_X1 u_and_module_1_U1 ( .A1(n_reg_module_1_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_1_res) );
  AND2_X1 u_and_module_2_U1 ( .A1(n_reg_module_2_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_2_res) );
  XOR2_X1 u_xor_module_85_U1 ( .A(p_rand_6), .B(n_and_module_2_res), .Z(
        n_xor_module_85_res) );
  AND2_X1 u_and_module_3_U1 ( .A1(n_reg_module_3_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_3_res) );
  XOR2_X1 u_xor_module_86_U1 ( .A(p_rand_7), .B(n_and_module_3_res), .Z(
        n_xor_module_86_res) );
  AND2_X1 u_and_module_4_U1 ( .A1(n_reg_module_4_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_4_res) );
  XOR2_X1 u_xor_module_87_U1 ( .A(p_rand_8), .B(n_and_module_4_res), .Z(
        n_xor_module_87_res) );
  AND2_X1 u_and_module_5_U1 ( .A1(n_reg_module_1_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_5_res) );
  XOR2_X1 u_xor_module_88_U1 ( .A(p_rand_6), .B(n_and_module_5_res), .Z(
        n_xor_module_88_res) );
  AND2_X1 u_and_module_6_U1 ( .A1(n_reg_module_2_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_6_res) );
  AND2_X1 u_and_module_7_U1 ( .A1(n_reg_module_3_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_7_res) );
  XOR2_X1 u_xor_module_89_U1 ( .A(p_rand_9), .B(n_and_module_7_res), .Z(
        n_xor_module_89_res) );
  AND2_X1 u_and_module_8_U1 ( .A1(n_reg_module_4_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_8_res) );
  XOR2_X1 u_xor_module_90_U1 ( .A(p_rand_10), .B(n_and_module_8_res), .Z(
        n_xor_module_90_res) );
  AND2_X1 u_and_module_9_U1 ( .A1(n_reg_module_1_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_9_res) );
  XOR2_X1 u_xor_module_91_U1 ( .A(p_rand_7), .B(n_and_module_9_res), .Z(
        n_xor_module_91_res) );
  AND2_X1 u_and_module_10_U1 ( .A1(n_reg_module_2_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_10_res) );
  XOR2_X1 u_xor_module_92_U1 ( .A(p_rand_9), .B(n_and_module_10_res), .Z(
        n_xor_module_92_res) );
  AND2_X1 u_and_module_11_U1 ( .A1(n_reg_module_3_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_11_res) );
  AND2_X1 u_and_module_12_U1 ( .A1(n_reg_module_4_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_12_res) );
  XOR2_X1 u_xor_module_93_U1 ( .A(p_rand_11), .B(n_and_module_12_res), .Z(
        n_xor_module_93_res) );
  AND2_X1 u_and_module_13_U1 ( .A1(n_reg_module_1_res), .A2(io_i0_s3_d0), .ZN(
        n_and_module_13_res) );
  XOR2_X1 u_xor_module_94_U1 ( .A(p_rand_8), .B(n_and_module_13_res), .Z(
        n_xor_module_94_res) );
  AND2_X1 u_and_module_14_U1 ( .A1(n_reg_module_2_res), .A2(io_i0_s3_d0), .ZN(
        n_and_module_14_res) );
  XOR2_X1 u_xor_module_95_U1 ( .A(p_rand_10), .B(n_and_module_14_res), .Z(
        n_xor_module_95_res) );
  AND2_X1 u_and_module_15_U1 ( .A1(n_reg_module_3_res), .A2(io_i0_s3_d0), .ZN(
        n_and_module_15_res) );
  XOR2_X1 u_xor_module_96_U1 ( .A(p_rand_11), .B(n_and_module_15_res), .Z(
        n_xor_module_96_res) );
  AND2_X1 u_and_module_16_U1 ( .A1(n_reg_module_4_res), .A2(io_i0_s3_d0), .ZN(
        n_and_module_16_res) );
  AND2_X1 u_and_module_17_U1 ( .A1(n_reg_module_5_res), .A2(io_i0_s0_d1), .ZN(
        n_and_module_17_res) );
  AND2_X1 u_and_module_18_U1 ( .A1(n_reg_module_6_res), .A2(io_i0_s0_d1), .ZN(
        n_and_module_18_res) );
  XOR2_X1 u_xor_module_97_U1 ( .A(p_rand_6), .B(n_and_module_18_res), .Z(
        n_xor_module_97_res) );
  AND2_X1 u_and_module_19_U1 ( .A1(n_reg_module_7_res), .A2(io_i0_s0_d1), .ZN(
        n_and_module_19_res) );
  XOR2_X1 u_xor_module_98_U1 ( .A(p_rand_7), .B(n_and_module_19_res), .Z(
        n_xor_module_98_res) );
  AND2_X1 u_and_module_20_U1 ( .A1(n_reg_module_8_res), .A2(io_i0_s0_d1), .ZN(
        n_and_module_20_res) );
  XOR2_X1 u_xor_module_99_U1 ( .A(p_rand_8), .B(n_and_module_20_res), .Z(
        n_xor_module_99_res) );
  AND2_X1 u_and_module_21_U1 ( .A1(n_reg_module_5_res), .A2(io_i0_s1_d1), .ZN(
        n_and_module_21_res) );
  XOR2_X1 u_xor_module_100_U1 ( .A(p_rand_6), .B(n_and_module_21_res), .Z(
        n_xor_module_100_res) );
  AND2_X1 u_and_module_22_U1 ( .A1(n_reg_module_6_res), .A2(io_i0_s1_d1), .ZN(
        n_and_module_22_res) );
  AND2_X1 u_and_module_23_U1 ( .A1(n_reg_module_7_res), .A2(io_i0_s1_d1), .ZN(
        n_and_module_23_res) );
  XOR2_X1 u_xor_module_101_U1 ( .A(p_rand_9), .B(n_and_module_23_res), .Z(
        n_xor_module_101_res) );
  AND2_X1 u_and_module_24_U1 ( .A1(n_reg_module_8_res), .A2(io_i0_s1_d1), .ZN(
        n_and_module_24_res) );
  XOR2_X1 u_xor_module_102_U1 ( .A(p_rand_10), .B(n_and_module_24_res), .Z(
        n_xor_module_102_res) );
  AND2_X1 u_and_module_25_U1 ( .A1(n_reg_module_5_res), .A2(io_i0_s2_d1), .ZN(
        n_and_module_25_res) );
  XOR2_X1 u_xor_module_103_U1 ( .A(p_rand_7), .B(n_and_module_25_res), .Z(
        n_xor_module_103_res) );
  AND2_X1 u_and_module_26_U1 ( .A1(n_reg_module_6_res), .A2(io_i0_s2_d1), .ZN(
        n_and_module_26_res) );
  XOR2_X1 u_xor_module_104_U1 ( .A(p_rand_9), .B(n_and_module_26_res), .Z(
        n_xor_module_104_res) );
  AND2_X1 u_and_module_27_U1 ( .A1(n_reg_module_7_res), .A2(io_i0_s2_d1), .ZN(
        n_and_module_27_res) );
  AND2_X1 u_and_module_28_U1 ( .A1(n_reg_module_8_res), .A2(io_i0_s2_d1), .ZN(
        n_and_module_28_res) );
  XOR2_X1 u_xor_module_105_U1 ( .A(p_rand_11), .B(n_and_module_28_res), .Z(
        n_xor_module_105_res) );
  AND2_X1 u_and_module_29_U1 ( .A1(n_reg_module_5_res), .A2(io_i0_s3_d1), .ZN(
        n_and_module_29_res) );
  XOR2_X1 u_xor_module_106_U1 ( .A(p_rand_8), .B(n_and_module_29_res), .Z(
        n_xor_module_106_res) );
  AND2_X1 u_and_module_30_U1 ( .A1(n_reg_module_6_res), .A2(io_i0_s3_d1), .ZN(
        n_and_module_30_res) );
  XOR2_X1 u_xor_module_107_U1 ( .A(p_rand_10), .B(n_and_module_30_res), .Z(
        n_xor_module_107_res) );
  AND2_X1 u_and_module_31_U1 ( .A1(n_reg_module_7_res), .A2(io_i0_s3_d1), .ZN(
        n_and_module_31_res) );
  XOR2_X1 u_xor_module_108_U1 ( .A(p_rand_11), .B(n_and_module_31_res), .Z(
        n_xor_module_108_res) );
  AND2_X1 u_and_module_32_U1 ( .A1(n_reg_module_8_res), .A2(io_i0_s3_d1), .ZN(
        n_and_module_32_res) );
  AND2_X1 u_and_module_33_U1 ( .A1(n_reg_module_9_res), .A2(io_i0_s0_d2), .ZN(
        n_and_module_33_res) );
  AND2_X1 u_and_module_34_U1 ( .A1(n_reg_module_10_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_34_res) );
  XOR2_X1 u_xor_module_109_U1 ( .A(p_rand_6), .B(n_and_module_34_res), .Z(
        n_xor_module_109_res) );
  AND2_X1 u_and_module_35_U1 ( .A1(n_reg_module_11_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_35_res) );
  XOR2_X1 u_xor_module_110_U1 ( .A(p_rand_7), .B(n_and_module_35_res), .Z(
        n_xor_module_110_res) );
  AND2_X1 u_and_module_36_U1 ( .A1(n_reg_module_12_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_36_res) );
  XOR2_X1 u_xor_module_111_U1 ( .A(p_rand_8), .B(n_and_module_36_res), .Z(
        n_xor_module_111_res) );
  AND2_X1 u_and_module_37_U1 ( .A1(n_reg_module_9_res), .A2(io_i0_s1_d2), .ZN(
        n_and_module_37_res) );
  XOR2_X1 u_xor_module_112_U1 ( .A(p_rand_6), .B(n_and_module_37_res), .Z(
        n_xor_module_112_res) );
  AND2_X1 u_and_module_38_U1 ( .A1(n_reg_module_10_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_38_res) );
  AND2_X1 u_and_module_39_U1 ( .A1(n_reg_module_11_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_39_res) );
  XOR2_X1 u_xor_module_113_U1 ( .A(p_rand_9), .B(n_and_module_39_res), .Z(
        n_xor_module_113_res) );
  AND2_X1 u_and_module_40_U1 ( .A1(n_reg_module_12_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_40_res) );
  XOR2_X1 u_xor_module_114_U1 ( .A(p_rand_10), .B(n_and_module_40_res), .Z(
        n_xor_module_114_res) );
  AND2_X1 u_and_module_41_U1 ( .A1(n_reg_module_9_res), .A2(io_i0_s2_d2), .ZN(
        n_and_module_41_res) );
  XOR2_X1 u_xor_module_115_U1 ( .A(p_rand_7), .B(n_and_module_41_res), .Z(
        n_xor_module_115_res) );
  AND2_X1 u_and_module_42_U1 ( .A1(n_reg_module_10_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_42_res) );
  XOR2_X1 u_xor_module_116_U1 ( .A(p_rand_9), .B(n_and_module_42_res), .Z(
        n_xor_module_116_res) );
  AND2_X1 u_and_module_43_U1 ( .A1(n_reg_module_11_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_43_res) );
  AND2_X1 u_and_module_44_U1 ( .A1(n_reg_module_12_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_44_res) );
  XOR2_X1 u_xor_module_117_U1 ( .A(p_rand_11), .B(n_and_module_44_res), .Z(
        n_xor_module_117_res) );
  AND2_X1 u_and_module_45_U1 ( .A1(n_reg_module_9_res), .A2(io_i0_s3_d2), .ZN(
        n_and_module_45_res) );
  XOR2_X1 u_xor_module_118_U1 ( .A(p_rand_8), .B(n_and_module_45_res), .Z(
        n_xor_module_118_res) );
  AND2_X1 u_and_module_46_U1 ( .A1(n_reg_module_10_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_46_res) );
  XOR2_X1 u_xor_module_119_U1 ( .A(p_rand_10), .B(n_and_module_46_res), .Z(
        n_xor_module_119_res) );
  AND2_X1 u_and_module_47_U1 ( .A1(n_reg_module_11_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_47_res) );
  XOR2_X1 u_xor_module_120_U1 ( .A(p_rand_11), .B(n_and_module_47_res), .Z(
        n_xor_module_120_res) );
  AND2_X1 u_and_module_48_U1 ( .A1(n_reg_module_12_res), .A2(io_i0_s3_d2), 
        .ZN(n_and_module_48_res) );
  AND2_X1 u_and_module_49_U1 ( .A1(n_reg_module_13_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_49_res) );
  AND2_X1 u_and_module_50_U1 ( .A1(n_reg_module_14_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_50_res) );
  XOR2_X1 u_xor_module_121_U1 ( .A(p_rand_6), .B(n_and_module_50_res), .Z(
        n_xor_module_121_res) );
  AND2_X1 u_and_module_51_U1 ( .A1(n_reg_module_15_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_51_res) );
  XOR2_X1 u_xor_module_122_U1 ( .A(p_rand_7), .B(n_and_module_51_res), .Z(
        n_xor_module_122_res) );
  AND2_X1 u_and_module_52_U1 ( .A1(n_reg_module_16_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_52_res) );
  XOR2_X1 u_xor_module_123_U1 ( .A(p_rand_8), .B(n_and_module_52_res), .Z(
        n_xor_module_123_res) );
  AND2_X1 u_and_module_53_U1 ( .A1(n_reg_module_13_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_53_res) );
  XOR2_X1 u_xor_module_124_U1 ( .A(p_rand_6), .B(n_and_module_53_res), .Z(
        n_xor_module_124_res) );
  AND2_X1 u_and_module_54_U1 ( .A1(n_reg_module_14_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_54_res) );
  AND2_X1 u_and_module_55_U1 ( .A1(n_reg_module_15_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_55_res) );
  XOR2_X1 u_xor_module_125_U1 ( .A(p_rand_9), .B(n_and_module_55_res), .Z(
        n_xor_module_125_res) );
  AND2_X1 u_and_module_56_U1 ( .A1(n_reg_module_16_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_56_res) );
  XOR2_X1 u_xor_module_126_U1 ( .A(p_rand_10), .B(n_and_module_56_res), .Z(
        n_xor_module_126_res) );
  AND2_X1 u_and_module_57_U1 ( .A1(n_reg_module_13_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_57_res) );
  XOR2_X1 u_xor_module_127_U1 ( .A(p_rand_7), .B(n_and_module_57_res), .Z(
        n_xor_module_127_res) );
  AND2_X1 u_and_module_58_U1 ( .A1(n_reg_module_14_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_58_res) );
  XOR2_X1 u_xor_module_128_U1 ( .A(p_rand_9), .B(n_and_module_58_res), .Z(
        n_xor_module_128_res) );
  AND2_X1 u_and_module_59_U1 ( .A1(n_reg_module_15_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_59_res) );
  AND2_X1 u_and_module_60_U1 ( .A1(n_reg_module_16_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_60_res) );
  XOR2_X1 u_xor_module_129_U1 ( .A(p_rand_11), .B(n_and_module_60_res), .Z(
        n_xor_module_129_res) );
  AND2_X1 u_and_module_61_U1 ( .A1(n_reg_module_13_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_61_res) );
  XOR2_X1 u_xor_module_130_U1 ( .A(p_rand_8), .B(n_and_module_61_res), .Z(
        n_xor_module_130_res) );
  AND2_X1 u_and_module_62_U1 ( .A1(n_reg_module_14_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_62_res) );
  XOR2_X1 u_xor_module_131_U1 ( .A(p_rand_10), .B(n_and_module_62_res), .Z(
        n_xor_module_131_res) );
  AND2_X1 u_and_module_63_U1 ( .A1(n_reg_module_15_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_63_res) );
  XOR2_X1 u_xor_module_132_U1 ( .A(p_rand_11), .B(n_and_module_63_res), .Z(
        n_xor_module_132_res) );
  AND2_X1 u_and_module_64_U1 ( .A1(n_reg_module_16_res), .A2(io_i0_s3_d3), 
        .ZN(n_and_module_64_res) );
  AND2_X1 u_and_module_65_U1 ( .A1(n_reg_module_17_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_65_res) );
  AND2_X1 u_and_module_66_U1 ( .A1(n_reg_module_18_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_66_res) );
  XOR2_X1 u_xor_module_133_U1 ( .A(p_rand_6), .B(n_and_module_66_res), .Z(
        n_xor_module_133_res) );
  AND2_X1 u_and_module_67_U1 ( .A1(n_reg_module_19_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_67_res) );
  XOR2_X1 u_xor_module_134_U1 ( .A(p_rand_7), .B(n_and_module_67_res), .Z(
        n_xor_module_134_res) );
  AND2_X1 u_and_module_68_U1 ( .A1(n_reg_module_20_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_68_res) );
  XOR2_X1 u_xor_module_135_U1 ( .A(p_rand_8), .B(n_and_module_68_res), .Z(
        n_xor_module_135_res) );
  AND2_X1 u_and_module_69_U1 ( .A1(n_reg_module_17_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_69_res) );
  XOR2_X1 u_xor_module_136_U1 ( .A(p_rand_6), .B(n_and_module_69_res), .Z(
        n_xor_module_136_res) );
  AND2_X1 u_and_module_70_U1 ( .A1(n_reg_module_18_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_70_res) );
  AND2_X1 u_and_module_71_U1 ( .A1(n_reg_module_19_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_71_res) );
  XOR2_X1 u_xor_module_137_U1 ( .A(p_rand_9), .B(n_and_module_71_res), .Z(
        n_xor_module_137_res) );
  AND2_X1 u_and_module_72_U1 ( .A1(n_reg_module_20_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_72_res) );
  XOR2_X1 u_xor_module_138_U1 ( .A(p_rand_10), .B(n_and_module_72_res), .Z(
        n_xor_module_138_res) );
  AND2_X1 u_and_module_73_U1 ( .A1(n_reg_module_17_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_73_res) );
  XOR2_X1 u_xor_module_139_U1 ( .A(p_rand_7), .B(n_and_module_73_res), .Z(
        n_xor_module_139_res) );
  AND2_X1 u_and_module_74_U1 ( .A1(n_reg_module_18_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_74_res) );
  XOR2_X1 u_xor_module_140_U1 ( .A(p_rand_9), .B(n_and_module_74_res), .Z(
        n_xor_module_140_res) );
  AND2_X1 u_and_module_75_U1 ( .A1(n_reg_module_19_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_75_res) );
  AND2_X1 u_and_module_76_U1 ( .A1(n_reg_module_20_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_76_res) );
  XOR2_X1 u_xor_module_141_U1 ( .A(p_rand_11), .B(n_and_module_76_res), .Z(
        n_xor_module_141_res) );
  AND2_X1 u_and_module_77_U1 ( .A1(n_reg_module_17_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_77_res) );
  XOR2_X1 u_xor_module_142_U1 ( .A(p_rand_8), .B(n_and_module_77_res), .Z(
        n_xor_module_142_res) );
  AND2_X1 u_and_module_78_U1 ( .A1(n_reg_module_18_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_78_res) );
  XOR2_X1 u_xor_module_143_U1 ( .A(p_rand_10), .B(n_and_module_78_res), .Z(
        n_xor_module_143_res) );
  AND2_X1 u_and_module_79_U1 ( .A1(n_reg_module_19_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_79_res) );
  XOR2_X1 u_xor_module_144_U1 ( .A(p_rand_11), .B(n_and_module_79_res), .Z(
        n_xor_module_144_res) );
  AND2_X1 u_and_module_80_U1 ( .A1(n_reg_module_20_res), .A2(io_i0_s3_d4), 
        .ZN(n_and_module_80_res) );
  AND2_X1 u_and_module_81_U1 ( .A1(n_reg_module_21_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_81_res) );
  AND2_X1 u_and_module_82_U1 ( .A1(n_reg_module_22_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_82_res) );
  XOR2_X1 u_xor_module_145_U1 ( .A(p_rand_6), .B(n_and_module_82_res), .Z(
        n_xor_module_145_res) );
  AND2_X1 u_and_module_83_U1 ( .A1(n_reg_module_23_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_83_res) );
  XOR2_X1 u_xor_module_146_U1 ( .A(p_rand_7), .B(n_and_module_83_res), .Z(
        n_xor_module_146_res) );
  AND2_X1 u_and_module_84_U1 ( .A1(n_reg_module_24_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_84_res) );
  XOR2_X1 u_xor_module_147_U1 ( .A(p_rand_8), .B(n_and_module_84_res), .Z(
        n_xor_module_147_res) );
  AND2_X1 u_and_module_85_U1 ( .A1(n_reg_module_21_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_85_res) );
  XOR2_X1 u_xor_module_148_U1 ( .A(p_rand_6), .B(n_and_module_85_res), .Z(
        n_xor_module_148_res) );
  AND2_X1 u_and_module_86_U1 ( .A1(n_reg_module_22_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_86_res) );
  AND2_X1 u_and_module_87_U1 ( .A1(n_reg_module_23_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_87_res) );
  XOR2_X1 u_xor_module_149_U1 ( .A(p_rand_9), .B(n_and_module_87_res), .Z(
        n_xor_module_149_res) );
  AND2_X1 u_and_module_88_U1 ( .A1(n_reg_module_24_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_88_res) );
  XOR2_X1 u_xor_module_150_U1 ( .A(p_rand_10), .B(n_and_module_88_res), .Z(
        n_xor_module_150_res) );
  AND2_X1 u_and_module_89_U1 ( .A1(n_reg_module_21_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_89_res) );
  XOR2_X1 u_xor_module_151_U1 ( .A(p_rand_7), .B(n_and_module_89_res), .Z(
        n_xor_module_151_res) );
  AND2_X1 u_and_module_90_U1 ( .A1(n_reg_module_22_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_90_res) );
  XOR2_X1 u_xor_module_152_U1 ( .A(p_rand_9), .B(n_and_module_90_res), .Z(
        n_xor_module_152_res) );
  AND2_X1 u_and_module_91_U1 ( .A1(n_reg_module_23_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_91_res) );
  AND2_X1 u_and_module_92_U1 ( .A1(n_reg_module_24_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_92_res) );
  XOR2_X1 u_xor_module_153_U1 ( .A(p_rand_11), .B(n_and_module_92_res), .Z(
        n_xor_module_153_res) );
  AND2_X1 u_and_module_93_U1 ( .A1(n_reg_module_21_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_93_res) );
  XOR2_X1 u_xor_module_154_U1 ( .A(p_rand_8), .B(n_and_module_93_res), .Z(
        n_xor_module_154_res) );
  AND2_X1 u_and_module_94_U1 ( .A1(n_reg_module_22_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_94_res) );
  XOR2_X1 u_xor_module_155_U1 ( .A(p_rand_10), .B(n_and_module_94_res), .Z(
        n_xor_module_155_res) );
  AND2_X1 u_and_module_95_U1 ( .A1(n_reg_module_23_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_95_res) );
  XOR2_X1 u_xor_module_156_U1 ( .A(p_rand_11), .B(n_and_module_95_res), .Z(
        n_xor_module_156_res) );
  AND2_X1 u_and_module_96_U1 ( .A1(n_reg_module_24_res), .A2(io_i0_s3_d5), 
        .ZN(n_and_module_96_res) );
  AND2_X1 u_and_module_97_U1 ( .A1(n_reg_module_25_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_97_res) );
  AND2_X1 u_and_module_98_U1 ( .A1(n_reg_module_26_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_98_res) );
  XOR2_X1 u_xor_module_157_U1 ( .A(p_rand_6), .B(n_and_module_98_res), .Z(
        n_xor_module_157_res) );
  AND2_X1 u_and_module_99_U1 ( .A1(n_reg_module_27_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_99_res) );
  XOR2_X1 u_xor_module_158_U1 ( .A(p_rand_7), .B(n_and_module_99_res), .Z(
        n_xor_module_158_res) );
  AND2_X1 u_and_module_100_U1 ( .A1(n_reg_module_28_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_100_res) );
  XOR2_X1 u_xor_module_159_U1 ( .A(p_rand_8), .B(n_and_module_100_res), .Z(
        n_xor_module_159_res) );
  AND2_X1 u_and_module_101_U1 ( .A1(n_reg_module_25_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_101_res) );
  XOR2_X1 u_xor_module_160_U1 ( .A(p_rand_6), .B(n_and_module_101_res), .Z(
        n_xor_module_160_res) );
  AND2_X1 u_and_module_102_U1 ( .A1(n_reg_module_26_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_102_res) );
  AND2_X1 u_and_module_103_U1 ( .A1(n_reg_module_27_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_103_res) );
  XOR2_X1 u_xor_module_161_U1 ( .A(p_rand_9), .B(n_and_module_103_res), .Z(
        n_xor_module_161_res) );
  AND2_X1 u_and_module_104_U1 ( .A1(n_reg_module_28_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_104_res) );
  XOR2_X1 u_xor_module_162_U1 ( .A(p_rand_10), .B(n_and_module_104_res), .Z(
        n_xor_module_162_res) );
  AND2_X1 u_and_module_105_U1 ( .A1(n_reg_module_25_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_105_res) );
  XOR2_X1 u_xor_module_163_U1 ( .A(p_rand_7), .B(n_and_module_105_res), .Z(
        n_xor_module_163_res) );
  AND2_X1 u_and_module_106_U1 ( .A1(n_reg_module_26_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_106_res) );
  XOR2_X1 u_xor_module_164_U1 ( .A(p_rand_9), .B(n_and_module_106_res), .Z(
        n_xor_module_164_res) );
  AND2_X1 u_and_module_107_U1 ( .A1(n_reg_module_27_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_107_res) );
  AND2_X1 u_and_module_108_U1 ( .A1(n_reg_module_28_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_108_res) );
  XOR2_X1 u_xor_module_165_U1 ( .A(p_rand_11), .B(n_and_module_108_res), .Z(
        n_xor_module_165_res) );
  AND2_X1 u_and_module_109_U1 ( .A1(n_reg_module_25_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_109_res) );
  XOR2_X1 u_xor_module_166_U1 ( .A(p_rand_8), .B(n_and_module_109_res), .Z(
        n_xor_module_166_res) );
  AND2_X1 u_and_module_110_U1 ( .A1(n_reg_module_26_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_110_res) );
  XOR2_X1 u_xor_module_167_U1 ( .A(p_rand_10), .B(n_and_module_110_res), .Z(
        n_xor_module_167_res) );
  AND2_X1 u_and_module_111_U1 ( .A1(n_reg_module_27_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_111_res) );
  XOR2_X1 u_xor_module_168_U1 ( .A(p_rand_11), .B(n_and_module_111_res), .Z(
        n_xor_module_168_res) );
  AND2_X1 u_and_module_112_U1 ( .A1(n_reg_module_28_res), .A2(io_i0_s3_d6), 
        .ZN(n_and_module_112_res) );
  DFF_X1 u_reg_module_29__cini_mul_v00_reg ( .D(n_and_module_1_res), .CK(
        clock_0), .Q(n_reg_module_29_res), .QN() );
  AND2_X1 u_majority7_module_28__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_28__and_module_1_res)
         );
  OR2_X1 u_majority7_module_28__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_28__or_module_1_res)
         );
  AND2_X1 u_majority7_module_28__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(n_majority7_module_28__and_module_2_res) );
  OR2_X1 u_majority7_module_28__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_28__or_module_2_res)
         );
  AND2_X1 u_majority7_module_28__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(n_majority7_module_28__and_module_3_res) );
  OR2_X1 u_majority7_module_28__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_28__or_module_3_res)
         );
  AND2_X1 u_majority7_module_28__and_module_4_U1 ( .A1(
        n_majority7_module_28__and_module_2_res), .A2(
        n_majority7_module_28__and_module_1_res), .ZN(
        n_majority7_module_28__and_module_4_res) );
  OR2_X1 u_majority7_module_28__or_module_4_U1 ( .A1(
        n_majority7_module_28__and_module_1_res), .A2(
        n_majority7_module_28__and_module_2_res), .ZN(
        n_majority7_module_28__or_module_4_res) );
  AND2_X1 u_majority7_module_28__and_module_5_U1 ( .A1(
        n_majority7_module_28__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_28__and_module_5_res) );
  OR2_X1 u_majority7_module_28__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_28__and_module_3_res), .ZN(
        n_majority7_module_28__or_module_5_res) );
  AND2_X1 u_majority7_module_28__and_module_6_U1 ( .A1(
        n_majority7_module_28__or_module_1_res), .A2(
        n_majority7_module_28__or_module_2_res), .ZN(
        n_majority7_module_28__and_module_6_res) );
  OR2_X1 u_majority7_module_28__or_module_6_U1 ( .A1(
        n_majority7_module_28__or_module_2_res), .A2(
        n_majority7_module_28__or_module_1_res), .ZN(
        n_majority7_module_28__or_module_6_res) );
  OR2_X1 u_majority7_module_28__or_module_7_U1 ( .A1(
        n_majority7_module_28__and_module_4_res), .A2(
        n_majority7_module_28__and_module_5_res), .ZN(
        n_majority7_module_28__or_module_7_res) );
  AND2_X1 u_majority7_module_28__and_module_7_U1 ( .A1(
        n_majority7_module_28__or_module_3_res), .A2(
        n_majority7_module_28__or_module_4_res), .ZN(
        n_majority7_module_28__and_module_7_res) );
  OR2_X1 u_majority7_module_28__or_module_8_U1 ( .A1(
        n_majority7_module_28__or_module_4_res), .A2(
        n_majority7_module_28__or_module_3_res), .ZN(
        n_majority7_module_28__or_module_8_res) );
  AND2_X1 u_majority7_module_28__and_module_8_U1 ( .A1(
        n_majority7_module_28__or_module_5_res), .A2(
        n_majority7_module_28__and_module_6_res), .ZN(
        n_majority7_module_28__and_module_8_res) );
  OR2_X1 u_majority7_module_28__or_module_9_U1 ( .A1(
        n_majority7_module_28__and_module_6_res), .A2(
        n_majority7_module_28__or_module_5_res), .ZN(
        n_majority7_module_28__or_module_9_res) );
  OR2_X1 u_majority7_module_28__or_module_10_U1 ( .A1(
        n_majority7_module_28__or_module_7_res), .A2(
        n_majority7_module_28__and_module_7_res), .ZN(
        n_majority7_module_28__or_module_10_res) );
  AND2_X1 u_majority7_module_28__and_module_9_U1 ( .A1(
        n_majority7_module_28__or_module_6_res), .A2(
        n_majority7_module_28__or_module_9_res), .ZN(
        n_majority7_module_28__and_module_9_res) );
  OR2_X1 u_majority7_module_28__or_module_11_U1 ( .A1(
        n_majority7_module_28__or_module_10_res), .A2(
        n_majority7_module_28__and_module_8_res), .ZN(
        n_majority7_module_28__or_module_11_res) );
  AND2_X1 u_majority7_module_28__and_module_10_U1 ( .A1(
        n_majority7_module_28__or_module_8_res), .A2(
        n_majority7_module_28__and_module_9_res), .ZN(
        n_majority7_module_28__and_module_10_res) );
  AND2_X1 u_majority7_module_28__and_module_11_U1 ( .A1(
        n_majority7_module_28__and_module_10_res), .A2(
        n_majority7_module_28__or_module_11_res), .ZN(
        n_majority7_module_28_res) );
  DFF_X1 u_reg_module_30__cini_mul_v00_reg ( .D(n_majority7_module_28_res), 
        .CK(clock_0), .Q(n_reg_module_30_res), .QN() );
  AND2_X1 u_majority7_module_29__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_29__and_module_1_res)
         );
  OR2_X1 u_majority7_module_29__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_29__or_module_1_res)
         );
  AND2_X1 u_majority7_module_29__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(n_majority7_module_29__and_module_2_res) );
  OR2_X1 u_majority7_module_29__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_29__or_module_2_res)
         );
  AND2_X1 u_majority7_module_29__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(n_majority7_module_29__and_module_3_res) );
  OR2_X1 u_majority7_module_29__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_29__or_module_3_res)
         );
  AND2_X1 u_majority7_module_29__and_module_4_U1 ( .A1(
        n_majority7_module_29__and_module_2_res), .A2(
        n_majority7_module_29__and_module_1_res), .ZN(
        n_majority7_module_29__and_module_4_res) );
  OR2_X1 u_majority7_module_29__or_module_4_U1 ( .A1(
        n_majority7_module_29__and_module_1_res), .A2(
        n_majority7_module_29__and_module_2_res), .ZN(
        n_majority7_module_29__or_module_4_res) );
  AND2_X1 u_majority7_module_29__and_module_5_U1 ( .A1(
        n_majority7_module_29__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_29__and_module_5_res) );
  OR2_X1 u_majority7_module_29__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_29__and_module_3_res), .ZN(
        n_majority7_module_29__or_module_5_res) );
  AND2_X1 u_majority7_module_29__and_module_6_U1 ( .A1(
        n_majority7_module_29__or_module_1_res), .A2(
        n_majority7_module_29__or_module_2_res), .ZN(
        n_majority7_module_29__and_module_6_res) );
  OR2_X1 u_majority7_module_29__or_module_6_U1 ( .A1(
        n_majority7_module_29__or_module_2_res), .A2(
        n_majority7_module_29__or_module_1_res), .ZN(
        n_majority7_module_29__or_module_6_res) );
  OR2_X1 u_majority7_module_29__or_module_7_U1 ( .A1(
        n_majority7_module_29__and_module_4_res), .A2(
        n_majority7_module_29__and_module_5_res), .ZN(
        n_majority7_module_29__or_module_7_res) );
  AND2_X1 u_majority7_module_29__and_module_7_U1 ( .A1(
        n_majority7_module_29__or_module_3_res), .A2(
        n_majority7_module_29__or_module_4_res), .ZN(
        n_majority7_module_29__and_module_7_res) );
  OR2_X1 u_majority7_module_29__or_module_8_U1 ( .A1(
        n_majority7_module_29__or_module_4_res), .A2(
        n_majority7_module_29__or_module_3_res), .ZN(
        n_majority7_module_29__or_module_8_res) );
  AND2_X1 u_majority7_module_29__and_module_8_U1 ( .A1(
        n_majority7_module_29__or_module_5_res), .A2(
        n_majority7_module_29__and_module_6_res), .ZN(
        n_majority7_module_29__and_module_8_res) );
  OR2_X1 u_majority7_module_29__or_module_9_U1 ( .A1(
        n_majority7_module_29__and_module_6_res), .A2(
        n_majority7_module_29__or_module_5_res), .ZN(
        n_majority7_module_29__or_module_9_res) );
  OR2_X1 u_majority7_module_29__or_module_10_U1 ( .A1(
        n_majority7_module_29__or_module_7_res), .A2(
        n_majority7_module_29__and_module_7_res), .ZN(
        n_majority7_module_29__or_module_10_res) );
  AND2_X1 u_majority7_module_29__and_module_9_U1 ( .A1(
        n_majority7_module_29__or_module_6_res), .A2(
        n_majority7_module_29__or_module_9_res), .ZN(
        n_majority7_module_29__and_module_9_res) );
  OR2_X1 u_majority7_module_29__or_module_11_U1 ( .A1(
        n_majority7_module_29__or_module_10_res), .A2(
        n_majority7_module_29__and_module_8_res), .ZN(
        n_majority7_module_29__or_module_11_res) );
  AND2_X1 u_majority7_module_29__and_module_10_U1 ( .A1(
        n_majority7_module_29__or_module_8_res), .A2(
        n_majority7_module_29__and_module_9_res), .ZN(
        n_majority7_module_29__and_module_10_res) );
  AND2_X1 u_majority7_module_29__and_module_11_U1 ( .A1(
        n_majority7_module_29__and_module_10_res), .A2(
        n_majority7_module_29__or_module_11_res), .ZN(
        n_majority7_module_29_res) );
  DFF_X1 u_reg_module_31__cini_mul_v00_reg ( .D(n_majority7_module_29_res), 
        .CK(clock_0), .Q(n_reg_module_31_res), .QN() );
  AND2_X1 u_majority7_module_30__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_30__and_module_1_res)
         );
  OR2_X1 u_majority7_module_30__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_30__or_module_1_res)
         );
  AND2_X1 u_majority7_module_30__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(n_majority7_module_30__and_module_2_res) );
  OR2_X1 u_majority7_module_30__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_30__or_module_2_res)
         );
  AND2_X1 u_majority7_module_30__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(n_majority7_module_30__and_module_3_res) );
  OR2_X1 u_majority7_module_30__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_30__or_module_3_res)
         );
  AND2_X1 u_majority7_module_30__and_module_4_U1 ( .A1(
        n_majority7_module_30__and_module_2_res), .A2(
        n_majority7_module_30__and_module_1_res), .ZN(
        n_majority7_module_30__and_module_4_res) );
  OR2_X1 u_majority7_module_30__or_module_4_U1 ( .A1(
        n_majority7_module_30__and_module_1_res), .A2(
        n_majority7_module_30__and_module_2_res), .ZN(
        n_majority7_module_30__or_module_4_res) );
  AND2_X1 u_majority7_module_30__and_module_5_U1 ( .A1(
        n_majority7_module_30__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_30__and_module_5_res) );
  OR2_X1 u_majority7_module_30__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_30__and_module_3_res), .ZN(
        n_majority7_module_30__or_module_5_res) );
  AND2_X1 u_majority7_module_30__and_module_6_U1 ( .A1(
        n_majority7_module_30__or_module_1_res), .A2(
        n_majority7_module_30__or_module_2_res), .ZN(
        n_majority7_module_30__and_module_6_res) );
  OR2_X1 u_majority7_module_30__or_module_6_U1 ( .A1(
        n_majority7_module_30__or_module_2_res), .A2(
        n_majority7_module_30__or_module_1_res), .ZN(
        n_majority7_module_30__or_module_6_res) );
  OR2_X1 u_majority7_module_30__or_module_7_U1 ( .A1(
        n_majority7_module_30__and_module_4_res), .A2(
        n_majority7_module_30__and_module_5_res), .ZN(
        n_majority7_module_30__or_module_7_res) );
  AND2_X1 u_majority7_module_30__and_module_7_U1 ( .A1(
        n_majority7_module_30__or_module_3_res), .A2(
        n_majority7_module_30__or_module_4_res), .ZN(
        n_majority7_module_30__and_module_7_res) );
  OR2_X1 u_majority7_module_30__or_module_8_U1 ( .A1(
        n_majority7_module_30__or_module_4_res), .A2(
        n_majority7_module_30__or_module_3_res), .ZN(
        n_majority7_module_30__or_module_8_res) );
  AND2_X1 u_majority7_module_30__and_module_8_U1 ( .A1(
        n_majority7_module_30__or_module_5_res), .A2(
        n_majority7_module_30__and_module_6_res), .ZN(
        n_majority7_module_30__and_module_8_res) );
  OR2_X1 u_majority7_module_30__or_module_9_U1 ( .A1(
        n_majority7_module_30__and_module_6_res), .A2(
        n_majority7_module_30__or_module_5_res), .ZN(
        n_majority7_module_30__or_module_9_res) );
  OR2_X1 u_majority7_module_30__or_module_10_U1 ( .A1(
        n_majority7_module_30__or_module_7_res), .A2(
        n_majority7_module_30__and_module_7_res), .ZN(
        n_majority7_module_30__or_module_10_res) );
  AND2_X1 u_majority7_module_30__and_module_9_U1 ( .A1(
        n_majority7_module_30__or_module_6_res), .A2(
        n_majority7_module_30__or_module_9_res), .ZN(
        n_majority7_module_30__and_module_9_res) );
  OR2_X1 u_majority7_module_30__or_module_11_U1 ( .A1(
        n_majority7_module_30__or_module_10_res), .A2(
        n_majority7_module_30__and_module_8_res), .ZN(
        n_majority7_module_30__or_module_11_res) );
  AND2_X1 u_majority7_module_30__and_module_10_U1 ( .A1(
        n_majority7_module_30__or_module_8_res), .A2(
        n_majority7_module_30__and_module_9_res), .ZN(
        n_majority7_module_30__and_module_10_res) );
  AND2_X1 u_majority7_module_30__and_module_11_U1 ( .A1(
        n_majority7_module_30__and_module_10_res), .A2(
        n_majority7_module_30__or_module_11_res), .ZN(
        n_majority7_module_30_res) );
  DFF_X1 u_reg_module_32__cini_mul_v00_reg ( .D(n_majority7_module_30_res), 
        .CK(clock_0), .Q(n_reg_module_32_res), .QN() );
  AND2_X1 u_majority7_module_31__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_31__and_module_1_res)
         );
  OR2_X1 u_majority7_module_31__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_31__or_module_1_res)
         );
  AND2_X1 u_majority7_module_31__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(n_majority7_module_31__and_module_2_res) );
  OR2_X1 u_majority7_module_31__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_31__or_module_2_res)
         );
  AND2_X1 u_majority7_module_31__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(n_majority7_module_31__and_module_3_res) );
  OR2_X1 u_majority7_module_31__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_31__or_module_3_res)
         );
  AND2_X1 u_majority7_module_31__and_module_4_U1 ( .A1(
        n_majority7_module_31__and_module_2_res), .A2(
        n_majority7_module_31__and_module_1_res), .ZN(
        n_majority7_module_31__and_module_4_res) );
  OR2_X1 u_majority7_module_31__or_module_4_U1 ( .A1(
        n_majority7_module_31__and_module_1_res), .A2(
        n_majority7_module_31__and_module_2_res), .ZN(
        n_majority7_module_31__or_module_4_res) );
  AND2_X1 u_majority7_module_31__and_module_5_U1 ( .A1(
        n_majority7_module_31__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_31__and_module_5_res) );
  OR2_X1 u_majority7_module_31__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_31__and_module_3_res), .ZN(
        n_majority7_module_31__or_module_5_res) );
  AND2_X1 u_majority7_module_31__and_module_6_U1 ( .A1(
        n_majority7_module_31__or_module_1_res), .A2(
        n_majority7_module_31__or_module_2_res), .ZN(
        n_majority7_module_31__and_module_6_res) );
  OR2_X1 u_majority7_module_31__or_module_6_U1 ( .A1(
        n_majority7_module_31__or_module_2_res), .A2(
        n_majority7_module_31__or_module_1_res), .ZN(
        n_majority7_module_31__or_module_6_res) );
  OR2_X1 u_majority7_module_31__or_module_7_U1 ( .A1(
        n_majority7_module_31__and_module_4_res), .A2(
        n_majority7_module_31__and_module_5_res), .ZN(
        n_majority7_module_31__or_module_7_res) );
  AND2_X1 u_majority7_module_31__and_module_7_U1 ( .A1(
        n_majority7_module_31__or_module_3_res), .A2(
        n_majority7_module_31__or_module_4_res), .ZN(
        n_majority7_module_31__and_module_7_res) );
  OR2_X1 u_majority7_module_31__or_module_8_U1 ( .A1(
        n_majority7_module_31__or_module_4_res), .A2(
        n_majority7_module_31__or_module_3_res), .ZN(
        n_majority7_module_31__or_module_8_res) );
  AND2_X1 u_majority7_module_31__and_module_8_U1 ( .A1(
        n_majority7_module_31__or_module_5_res), .A2(
        n_majority7_module_31__and_module_6_res), .ZN(
        n_majority7_module_31__and_module_8_res) );
  OR2_X1 u_majority7_module_31__or_module_9_U1 ( .A1(
        n_majority7_module_31__and_module_6_res), .A2(
        n_majority7_module_31__or_module_5_res), .ZN(
        n_majority7_module_31__or_module_9_res) );
  OR2_X1 u_majority7_module_31__or_module_10_U1 ( .A1(
        n_majority7_module_31__or_module_7_res), .A2(
        n_majority7_module_31__and_module_7_res), .ZN(
        n_majority7_module_31__or_module_10_res) );
  AND2_X1 u_majority7_module_31__and_module_9_U1 ( .A1(
        n_majority7_module_31__or_module_6_res), .A2(
        n_majority7_module_31__or_module_9_res), .ZN(
        n_majority7_module_31__and_module_9_res) );
  OR2_X1 u_majority7_module_31__or_module_11_U1 ( .A1(
        n_majority7_module_31__or_module_10_res), .A2(
        n_majority7_module_31__and_module_8_res), .ZN(
        n_majority7_module_31__or_module_11_res) );
  AND2_X1 u_majority7_module_31__and_module_10_U1 ( .A1(
        n_majority7_module_31__or_module_8_res), .A2(
        n_majority7_module_31__and_module_9_res), .ZN(
        n_majority7_module_31__and_module_10_res) );
  AND2_X1 u_majority7_module_31__and_module_11_U1 ( .A1(
        n_majority7_module_31__and_module_10_res), .A2(
        n_majority7_module_31__or_module_11_res), .ZN(
        n_majority7_module_31_res) );
  DFF_X1 u_reg_module_33__cini_mul_v00_reg ( .D(n_majority7_module_31_res), 
        .CK(clock_0), .Q(n_reg_module_33_res), .QN() );
  DFF_X1 u_reg_module_34__cini_mul_v00_reg ( .D(n_and_module_6_res), .CK(
        clock_0), .Q(n_reg_module_34_res), .QN() );
  AND2_X1 u_majority7_module_32__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_32__and_module_1_res)
         );
  OR2_X1 u_majority7_module_32__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_32__or_module_1_res)
         );
  AND2_X1 u_majority7_module_32__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(n_majority7_module_32__and_module_2_res) );
  OR2_X1 u_majority7_module_32__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_32__or_module_2_res)
         );
  AND2_X1 u_majority7_module_32__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(n_majority7_module_32__and_module_3_res) );
  OR2_X1 u_majority7_module_32__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_32__or_module_3_res)
         );
  AND2_X1 u_majority7_module_32__and_module_4_U1 ( .A1(
        n_majority7_module_32__and_module_2_res), .A2(
        n_majority7_module_32__and_module_1_res), .ZN(
        n_majority7_module_32__and_module_4_res) );
  OR2_X1 u_majority7_module_32__or_module_4_U1 ( .A1(
        n_majority7_module_32__and_module_1_res), .A2(
        n_majority7_module_32__and_module_2_res), .ZN(
        n_majority7_module_32__or_module_4_res) );
  AND2_X1 u_majority7_module_32__and_module_5_U1 ( .A1(
        n_majority7_module_32__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_32__and_module_5_res) );
  OR2_X1 u_majority7_module_32__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_32__and_module_3_res), .ZN(
        n_majority7_module_32__or_module_5_res) );
  AND2_X1 u_majority7_module_32__and_module_6_U1 ( .A1(
        n_majority7_module_32__or_module_1_res), .A2(
        n_majority7_module_32__or_module_2_res), .ZN(
        n_majority7_module_32__and_module_6_res) );
  OR2_X1 u_majority7_module_32__or_module_6_U1 ( .A1(
        n_majority7_module_32__or_module_2_res), .A2(
        n_majority7_module_32__or_module_1_res), .ZN(
        n_majority7_module_32__or_module_6_res) );
  OR2_X1 u_majority7_module_32__or_module_7_U1 ( .A1(
        n_majority7_module_32__and_module_4_res), .A2(
        n_majority7_module_32__and_module_5_res), .ZN(
        n_majority7_module_32__or_module_7_res) );
  AND2_X1 u_majority7_module_32__and_module_7_U1 ( .A1(
        n_majority7_module_32__or_module_3_res), .A2(
        n_majority7_module_32__or_module_4_res), .ZN(
        n_majority7_module_32__and_module_7_res) );
  OR2_X1 u_majority7_module_32__or_module_8_U1 ( .A1(
        n_majority7_module_32__or_module_4_res), .A2(
        n_majority7_module_32__or_module_3_res), .ZN(
        n_majority7_module_32__or_module_8_res) );
  AND2_X1 u_majority7_module_32__and_module_8_U1 ( .A1(
        n_majority7_module_32__or_module_5_res), .A2(
        n_majority7_module_32__and_module_6_res), .ZN(
        n_majority7_module_32__and_module_8_res) );
  OR2_X1 u_majority7_module_32__or_module_9_U1 ( .A1(
        n_majority7_module_32__and_module_6_res), .A2(
        n_majority7_module_32__or_module_5_res), .ZN(
        n_majority7_module_32__or_module_9_res) );
  OR2_X1 u_majority7_module_32__or_module_10_U1 ( .A1(
        n_majority7_module_32__or_module_7_res), .A2(
        n_majority7_module_32__and_module_7_res), .ZN(
        n_majority7_module_32__or_module_10_res) );
  AND2_X1 u_majority7_module_32__and_module_9_U1 ( .A1(
        n_majority7_module_32__or_module_6_res), .A2(
        n_majority7_module_32__or_module_9_res), .ZN(
        n_majority7_module_32__and_module_9_res) );
  OR2_X1 u_majority7_module_32__or_module_11_U1 ( .A1(
        n_majority7_module_32__or_module_10_res), .A2(
        n_majority7_module_32__and_module_8_res), .ZN(
        n_majority7_module_32__or_module_11_res) );
  AND2_X1 u_majority7_module_32__and_module_10_U1 ( .A1(
        n_majority7_module_32__or_module_8_res), .A2(
        n_majority7_module_32__and_module_9_res), .ZN(
        n_majority7_module_32__and_module_10_res) );
  AND2_X1 u_majority7_module_32__and_module_11_U1 ( .A1(
        n_majority7_module_32__and_module_10_res), .A2(
        n_majority7_module_32__or_module_11_res), .ZN(
        n_majority7_module_32_res) );
  DFF_X1 u_reg_module_35__cini_mul_v00_reg ( .D(n_majority7_module_32_res), 
        .CK(clock_0), .Q(n_reg_module_35_res), .QN() );
  AND2_X1 u_majority7_module_33__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_33__and_module_1_res)
         );
  OR2_X1 u_majority7_module_33__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_33__or_module_1_res)
         );
  AND2_X1 u_majority7_module_33__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(n_majority7_module_33__and_module_2_res) );
  OR2_X1 u_majority7_module_33__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_33__or_module_2_res)
         );
  AND2_X1 u_majority7_module_33__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(n_majority7_module_33__and_module_3_res) );
  OR2_X1 u_majority7_module_33__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_33__or_module_3_res)
         );
  AND2_X1 u_majority7_module_33__and_module_4_U1 ( .A1(
        n_majority7_module_33__and_module_2_res), .A2(
        n_majority7_module_33__and_module_1_res), .ZN(
        n_majority7_module_33__and_module_4_res) );
  OR2_X1 u_majority7_module_33__or_module_4_U1 ( .A1(
        n_majority7_module_33__and_module_1_res), .A2(
        n_majority7_module_33__and_module_2_res), .ZN(
        n_majority7_module_33__or_module_4_res) );
  AND2_X1 u_majority7_module_33__and_module_5_U1 ( .A1(
        n_majority7_module_33__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_33__and_module_5_res) );
  OR2_X1 u_majority7_module_33__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_33__and_module_3_res), .ZN(
        n_majority7_module_33__or_module_5_res) );
  AND2_X1 u_majority7_module_33__and_module_6_U1 ( .A1(
        n_majority7_module_33__or_module_1_res), .A2(
        n_majority7_module_33__or_module_2_res), .ZN(
        n_majority7_module_33__and_module_6_res) );
  OR2_X1 u_majority7_module_33__or_module_6_U1 ( .A1(
        n_majority7_module_33__or_module_2_res), .A2(
        n_majority7_module_33__or_module_1_res), .ZN(
        n_majority7_module_33__or_module_6_res) );
  OR2_X1 u_majority7_module_33__or_module_7_U1 ( .A1(
        n_majority7_module_33__and_module_4_res), .A2(
        n_majority7_module_33__and_module_5_res), .ZN(
        n_majority7_module_33__or_module_7_res) );
  AND2_X1 u_majority7_module_33__and_module_7_U1 ( .A1(
        n_majority7_module_33__or_module_3_res), .A2(
        n_majority7_module_33__or_module_4_res), .ZN(
        n_majority7_module_33__and_module_7_res) );
  OR2_X1 u_majority7_module_33__or_module_8_U1 ( .A1(
        n_majority7_module_33__or_module_4_res), .A2(
        n_majority7_module_33__or_module_3_res), .ZN(
        n_majority7_module_33__or_module_8_res) );
  AND2_X1 u_majority7_module_33__and_module_8_U1 ( .A1(
        n_majority7_module_33__or_module_5_res), .A2(
        n_majority7_module_33__and_module_6_res), .ZN(
        n_majority7_module_33__and_module_8_res) );
  OR2_X1 u_majority7_module_33__or_module_9_U1 ( .A1(
        n_majority7_module_33__and_module_6_res), .A2(
        n_majority7_module_33__or_module_5_res), .ZN(
        n_majority7_module_33__or_module_9_res) );
  OR2_X1 u_majority7_module_33__or_module_10_U1 ( .A1(
        n_majority7_module_33__or_module_7_res), .A2(
        n_majority7_module_33__and_module_7_res), .ZN(
        n_majority7_module_33__or_module_10_res) );
  AND2_X1 u_majority7_module_33__and_module_9_U1 ( .A1(
        n_majority7_module_33__or_module_6_res), .A2(
        n_majority7_module_33__or_module_9_res), .ZN(
        n_majority7_module_33__and_module_9_res) );
  OR2_X1 u_majority7_module_33__or_module_11_U1 ( .A1(
        n_majority7_module_33__or_module_10_res), .A2(
        n_majority7_module_33__and_module_8_res), .ZN(
        n_majority7_module_33__or_module_11_res) );
  AND2_X1 u_majority7_module_33__and_module_10_U1 ( .A1(
        n_majority7_module_33__or_module_8_res), .A2(
        n_majority7_module_33__and_module_9_res), .ZN(
        n_majority7_module_33__and_module_10_res) );
  AND2_X1 u_majority7_module_33__and_module_11_U1 ( .A1(
        n_majority7_module_33__and_module_10_res), .A2(
        n_majority7_module_33__or_module_11_res), .ZN(
        n_majority7_module_33_res) );
  DFF_X1 u_reg_module_36__cini_mul_v00_reg ( .D(n_majority7_module_33_res), 
        .CK(clock_0), .Q(n_reg_module_36_res), .QN() );
  AND2_X1 u_majority7_module_34__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_34__and_module_1_res)
         );
  OR2_X1 u_majority7_module_34__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_34__or_module_1_res)
         );
  AND2_X1 u_majority7_module_34__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(n_majority7_module_34__and_module_2_res) );
  OR2_X1 u_majority7_module_34__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_34__or_module_2_res)
         );
  AND2_X1 u_majority7_module_34__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(n_majority7_module_34__and_module_3_res) );
  OR2_X1 u_majority7_module_34__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_34__or_module_3_res)
         );
  AND2_X1 u_majority7_module_34__and_module_4_U1 ( .A1(
        n_majority7_module_34__and_module_2_res), .A2(
        n_majority7_module_34__and_module_1_res), .ZN(
        n_majority7_module_34__and_module_4_res) );
  OR2_X1 u_majority7_module_34__or_module_4_U1 ( .A1(
        n_majority7_module_34__and_module_1_res), .A2(
        n_majority7_module_34__and_module_2_res), .ZN(
        n_majority7_module_34__or_module_4_res) );
  AND2_X1 u_majority7_module_34__and_module_5_U1 ( .A1(
        n_majority7_module_34__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_34__and_module_5_res) );
  OR2_X1 u_majority7_module_34__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_34__and_module_3_res), .ZN(
        n_majority7_module_34__or_module_5_res) );
  AND2_X1 u_majority7_module_34__and_module_6_U1 ( .A1(
        n_majority7_module_34__or_module_1_res), .A2(
        n_majority7_module_34__or_module_2_res), .ZN(
        n_majority7_module_34__and_module_6_res) );
  OR2_X1 u_majority7_module_34__or_module_6_U1 ( .A1(
        n_majority7_module_34__or_module_2_res), .A2(
        n_majority7_module_34__or_module_1_res), .ZN(
        n_majority7_module_34__or_module_6_res) );
  OR2_X1 u_majority7_module_34__or_module_7_U1 ( .A1(
        n_majority7_module_34__and_module_4_res), .A2(
        n_majority7_module_34__and_module_5_res), .ZN(
        n_majority7_module_34__or_module_7_res) );
  AND2_X1 u_majority7_module_34__and_module_7_U1 ( .A1(
        n_majority7_module_34__or_module_3_res), .A2(
        n_majority7_module_34__or_module_4_res), .ZN(
        n_majority7_module_34__and_module_7_res) );
  OR2_X1 u_majority7_module_34__or_module_8_U1 ( .A1(
        n_majority7_module_34__or_module_4_res), .A2(
        n_majority7_module_34__or_module_3_res), .ZN(
        n_majority7_module_34__or_module_8_res) );
  AND2_X1 u_majority7_module_34__and_module_8_U1 ( .A1(
        n_majority7_module_34__or_module_5_res), .A2(
        n_majority7_module_34__and_module_6_res), .ZN(
        n_majority7_module_34__and_module_8_res) );
  OR2_X1 u_majority7_module_34__or_module_9_U1 ( .A1(
        n_majority7_module_34__and_module_6_res), .A2(
        n_majority7_module_34__or_module_5_res), .ZN(
        n_majority7_module_34__or_module_9_res) );
  OR2_X1 u_majority7_module_34__or_module_10_U1 ( .A1(
        n_majority7_module_34__or_module_7_res), .A2(
        n_majority7_module_34__and_module_7_res), .ZN(
        n_majority7_module_34__or_module_10_res) );
  AND2_X1 u_majority7_module_34__and_module_9_U1 ( .A1(
        n_majority7_module_34__or_module_6_res), .A2(
        n_majority7_module_34__or_module_9_res), .ZN(
        n_majority7_module_34__and_module_9_res) );
  OR2_X1 u_majority7_module_34__or_module_11_U1 ( .A1(
        n_majority7_module_34__or_module_10_res), .A2(
        n_majority7_module_34__and_module_8_res), .ZN(
        n_majority7_module_34__or_module_11_res) );
  AND2_X1 u_majority7_module_34__and_module_10_U1 ( .A1(
        n_majority7_module_34__or_module_8_res), .A2(
        n_majority7_module_34__and_module_9_res), .ZN(
        n_majority7_module_34__and_module_10_res) );
  AND2_X1 u_majority7_module_34__and_module_11_U1 ( .A1(
        n_majority7_module_34__and_module_10_res), .A2(
        n_majority7_module_34__or_module_11_res), .ZN(
        n_majority7_module_34_res) );
  DFF_X1 u_reg_module_37__cini_mul_v00_reg ( .D(n_majority7_module_34_res), 
        .CK(clock_0), .Q(n_reg_module_37_res), .QN() );
  AND2_X1 u_majority7_module_35__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_35__and_module_1_res)
         );
  OR2_X1 u_majority7_module_35__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_35__or_module_1_res)
         );
  AND2_X1 u_majority7_module_35__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(n_majority7_module_35__and_module_2_res) );
  OR2_X1 u_majority7_module_35__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_35__or_module_2_res)
         );
  AND2_X1 u_majority7_module_35__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(n_majority7_module_35__and_module_3_res) );
  OR2_X1 u_majority7_module_35__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_35__or_module_3_res)
         );
  AND2_X1 u_majority7_module_35__and_module_4_U1 ( .A1(
        n_majority7_module_35__and_module_2_res), .A2(
        n_majority7_module_35__and_module_1_res), .ZN(
        n_majority7_module_35__and_module_4_res) );
  OR2_X1 u_majority7_module_35__or_module_4_U1 ( .A1(
        n_majority7_module_35__and_module_1_res), .A2(
        n_majority7_module_35__and_module_2_res), .ZN(
        n_majority7_module_35__or_module_4_res) );
  AND2_X1 u_majority7_module_35__and_module_5_U1 ( .A1(
        n_majority7_module_35__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_35__and_module_5_res) );
  OR2_X1 u_majority7_module_35__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_35__and_module_3_res), .ZN(
        n_majority7_module_35__or_module_5_res) );
  AND2_X1 u_majority7_module_35__and_module_6_U1 ( .A1(
        n_majority7_module_35__or_module_1_res), .A2(
        n_majority7_module_35__or_module_2_res), .ZN(
        n_majority7_module_35__and_module_6_res) );
  OR2_X1 u_majority7_module_35__or_module_6_U1 ( .A1(
        n_majority7_module_35__or_module_2_res), .A2(
        n_majority7_module_35__or_module_1_res), .ZN(
        n_majority7_module_35__or_module_6_res) );
  OR2_X1 u_majority7_module_35__or_module_7_U1 ( .A1(
        n_majority7_module_35__and_module_4_res), .A2(
        n_majority7_module_35__and_module_5_res), .ZN(
        n_majority7_module_35__or_module_7_res) );
  AND2_X1 u_majority7_module_35__and_module_7_U1 ( .A1(
        n_majority7_module_35__or_module_3_res), .A2(
        n_majority7_module_35__or_module_4_res), .ZN(
        n_majority7_module_35__and_module_7_res) );
  OR2_X1 u_majority7_module_35__or_module_8_U1 ( .A1(
        n_majority7_module_35__or_module_4_res), .A2(
        n_majority7_module_35__or_module_3_res), .ZN(
        n_majority7_module_35__or_module_8_res) );
  AND2_X1 u_majority7_module_35__and_module_8_U1 ( .A1(
        n_majority7_module_35__or_module_5_res), .A2(
        n_majority7_module_35__and_module_6_res), .ZN(
        n_majority7_module_35__and_module_8_res) );
  OR2_X1 u_majority7_module_35__or_module_9_U1 ( .A1(
        n_majority7_module_35__and_module_6_res), .A2(
        n_majority7_module_35__or_module_5_res), .ZN(
        n_majority7_module_35__or_module_9_res) );
  OR2_X1 u_majority7_module_35__or_module_10_U1 ( .A1(
        n_majority7_module_35__or_module_7_res), .A2(
        n_majority7_module_35__and_module_7_res), .ZN(
        n_majority7_module_35__or_module_10_res) );
  AND2_X1 u_majority7_module_35__and_module_9_U1 ( .A1(
        n_majority7_module_35__or_module_6_res), .A2(
        n_majority7_module_35__or_module_9_res), .ZN(
        n_majority7_module_35__and_module_9_res) );
  OR2_X1 u_majority7_module_35__or_module_11_U1 ( .A1(
        n_majority7_module_35__or_module_10_res), .A2(
        n_majority7_module_35__and_module_8_res), .ZN(
        n_majority7_module_35__or_module_11_res) );
  AND2_X1 u_majority7_module_35__and_module_10_U1 ( .A1(
        n_majority7_module_35__or_module_8_res), .A2(
        n_majority7_module_35__and_module_9_res), .ZN(
        n_majority7_module_35__and_module_10_res) );
  AND2_X1 u_majority7_module_35__and_module_11_U1 ( .A1(
        n_majority7_module_35__and_module_10_res), .A2(
        n_majority7_module_35__or_module_11_res), .ZN(
        n_majority7_module_35_res) );
  DFF_X1 u_reg_module_38__cini_mul_v00_reg ( .D(n_majority7_module_35_res), 
        .CK(clock_0), .Q(n_reg_module_38_res), .QN() );
  DFF_X1 u_reg_module_39__cini_mul_v00_reg ( .D(n_and_module_11_res), .CK(
        clock_0), .Q(n_reg_module_39_res), .QN() );
  AND2_X1 u_majority7_module_36__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_36__and_module_1_res)
         );
  OR2_X1 u_majority7_module_36__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_36__or_module_1_res)
         );
  AND2_X1 u_majority7_module_36__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(n_majority7_module_36__and_module_2_res) );
  OR2_X1 u_majority7_module_36__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_36__or_module_2_res)
         );
  AND2_X1 u_majority7_module_36__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(n_majority7_module_36__and_module_3_res) );
  OR2_X1 u_majority7_module_36__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_36__or_module_3_res)
         );
  AND2_X1 u_majority7_module_36__and_module_4_U1 ( .A1(
        n_majority7_module_36__and_module_2_res), .A2(
        n_majority7_module_36__and_module_1_res), .ZN(
        n_majority7_module_36__and_module_4_res) );
  OR2_X1 u_majority7_module_36__or_module_4_U1 ( .A1(
        n_majority7_module_36__and_module_1_res), .A2(
        n_majority7_module_36__and_module_2_res), .ZN(
        n_majority7_module_36__or_module_4_res) );
  AND2_X1 u_majority7_module_36__and_module_5_U1 ( .A1(
        n_majority7_module_36__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_36__and_module_5_res) );
  OR2_X1 u_majority7_module_36__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_36__and_module_3_res), .ZN(
        n_majority7_module_36__or_module_5_res) );
  AND2_X1 u_majority7_module_36__and_module_6_U1 ( .A1(
        n_majority7_module_36__or_module_1_res), .A2(
        n_majority7_module_36__or_module_2_res), .ZN(
        n_majority7_module_36__and_module_6_res) );
  OR2_X1 u_majority7_module_36__or_module_6_U1 ( .A1(
        n_majority7_module_36__or_module_2_res), .A2(
        n_majority7_module_36__or_module_1_res), .ZN(
        n_majority7_module_36__or_module_6_res) );
  OR2_X1 u_majority7_module_36__or_module_7_U1 ( .A1(
        n_majority7_module_36__and_module_4_res), .A2(
        n_majority7_module_36__and_module_5_res), .ZN(
        n_majority7_module_36__or_module_7_res) );
  AND2_X1 u_majority7_module_36__and_module_7_U1 ( .A1(
        n_majority7_module_36__or_module_3_res), .A2(
        n_majority7_module_36__or_module_4_res), .ZN(
        n_majority7_module_36__and_module_7_res) );
  OR2_X1 u_majority7_module_36__or_module_8_U1 ( .A1(
        n_majority7_module_36__or_module_4_res), .A2(
        n_majority7_module_36__or_module_3_res), .ZN(
        n_majority7_module_36__or_module_8_res) );
  AND2_X1 u_majority7_module_36__and_module_8_U1 ( .A1(
        n_majority7_module_36__or_module_5_res), .A2(
        n_majority7_module_36__and_module_6_res), .ZN(
        n_majority7_module_36__and_module_8_res) );
  OR2_X1 u_majority7_module_36__or_module_9_U1 ( .A1(
        n_majority7_module_36__and_module_6_res), .A2(
        n_majority7_module_36__or_module_5_res), .ZN(
        n_majority7_module_36__or_module_9_res) );
  OR2_X1 u_majority7_module_36__or_module_10_U1 ( .A1(
        n_majority7_module_36__or_module_7_res), .A2(
        n_majority7_module_36__and_module_7_res), .ZN(
        n_majority7_module_36__or_module_10_res) );
  AND2_X1 u_majority7_module_36__and_module_9_U1 ( .A1(
        n_majority7_module_36__or_module_6_res), .A2(
        n_majority7_module_36__or_module_9_res), .ZN(
        n_majority7_module_36__and_module_9_res) );
  OR2_X1 u_majority7_module_36__or_module_11_U1 ( .A1(
        n_majority7_module_36__or_module_10_res), .A2(
        n_majority7_module_36__and_module_8_res), .ZN(
        n_majority7_module_36__or_module_11_res) );
  AND2_X1 u_majority7_module_36__and_module_10_U1 ( .A1(
        n_majority7_module_36__or_module_8_res), .A2(
        n_majority7_module_36__and_module_9_res), .ZN(
        n_majority7_module_36__and_module_10_res) );
  AND2_X1 u_majority7_module_36__and_module_11_U1 ( .A1(
        n_majority7_module_36__and_module_10_res), .A2(
        n_majority7_module_36__or_module_11_res), .ZN(
        n_majority7_module_36_res) );
  DFF_X1 u_reg_module_40__cini_mul_v00_reg ( .D(n_majority7_module_36_res), 
        .CK(clock_0), .Q(n_reg_module_40_res), .QN() );
  AND2_X1 u_majority7_module_37__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_37__and_module_1_res)
         );
  OR2_X1 u_majority7_module_37__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_37__or_module_1_res)
         );
  AND2_X1 u_majority7_module_37__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(n_majority7_module_37__and_module_2_res) );
  OR2_X1 u_majority7_module_37__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_37__or_module_2_res)
         );
  AND2_X1 u_majority7_module_37__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(n_majority7_module_37__and_module_3_res) );
  OR2_X1 u_majority7_module_37__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_37__or_module_3_res)
         );
  AND2_X1 u_majority7_module_37__and_module_4_U1 ( .A1(
        n_majority7_module_37__and_module_2_res), .A2(
        n_majority7_module_37__and_module_1_res), .ZN(
        n_majority7_module_37__and_module_4_res) );
  OR2_X1 u_majority7_module_37__or_module_4_U1 ( .A1(
        n_majority7_module_37__and_module_1_res), .A2(
        n_majority7_module_37__and_module_2_res), .ZN(
        n_majority7_module_37__or_module_4_res) );
  AND2_X1 u_majority7_module_37__and_module_5_U1 ( .A1(
        n_majority7_module_37__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_37__and_module_5_res) );
  OR2_X1 u_majority7_module_37__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_37__and_module_3_res), .ZN(
        n_majority7_module_37__or_module_5_res) );
  AND2_X1 u_majority7_module_37__and_module_6_U1 ( .A1(
        n_majority7_module_37__or_module_1_res), .A2(
        n_majority7_module_37__or_module_2_res), .ZN(
        n_majority7_module_37__and_module_6_res) );
  OR2_X1 u_majority7_module_37__or_module_6_U1 ( .A1(
        n_majority7_module_37__or_module_2_res), .A2(
        n_majority7_module_37__or_module_1_res), .ZN(
        n_majority7_module_37__or_module_6_res) );
  OR2_X1 u_majority7_module_37__or_module_7_U1 ( .A1(
        n_majority7_module_37__and_module_4_res), .A2(
        n_majority7_module_37__and_module_5_res), .ZN(
        n_majority7_module_37__or_module_7_res) );
  AND2_X1 u_majority7_module_37__and_module_7_U1 ( .A1(
        n_majority7_module_37__or_module_3_res), .A2(
        n_majority7_module_37__or_module_4_res), .ZN(
        n_majority7_module_37__and_module_7_res) );
  OR2_X1 u_majority7_module_37__or_module_8_U1 ( .A1(
        n_majority7_module_37__or_module_4_res), .A2(
        n_majority7_module_37__or_module_3_res), .ZN(
        n_majority7_module_37__or_module_8_res) );
  AND2_X1 u_majority7_module_37__and_module_8_U1 ( .A1(
        n_majority7_module_37__or_module_5_res), .A2(
        n_majority7_module_37__and_module_6_res), .ZN(
        n_majority7_module_37__and_module_8_res) );
  OR2_X1 u_majority7_module_37__or_module_9_U1 ( .A1(
        n_majority7_module_37__and_module_6_res), .A2(
        n_majority7_module_37__or_module_5_res), .ZN(
        n_majority7_module_37__or_module_9_res) );
  OR2_X1 u_majority7_module_37__or_module_10_U1 ( .A1(
        n_majority7_module_37__or_module_7_res), .A2(
        n_majority7_module_37__and_module_7_res), .ZN(
        n_majority7_module_37__or_module_10_res) );
  AND2_X1 u_majority7_module_37__and_module_9_U1 ( .A1(
        n_majority7_module_37__or_module_6_res), .A2(
        n_majority7_module_37__or_module_9_res), .ZN(
        n_majority7_module_37__and_module_9_res) );
  OR2_X1 u_majority7_module_37__or_module_11_U1 ( .A1(
        n_majority7_module_37__or_module_10_res), .A2(
        n_majority7_module_37__and_module_8_res), .ZN(
        n_majority7_module_37__or_module_11_res) );
  AND2_X1 u_majority7_module_37__and_module_10_U1 ( .A1(
        n_majority7_module_37__or_module_8_res), .A2(
        n_majority7_module_37__and_module_9_res), .ZN(
        n_majority7_module_37__and_module_10_res) );
  AND2_X1 u_majority7_module_37__and_module_11_U1 ( .A1(
        n_majority7_module_37__and_module_10_res), .A2(
        n_majority7_module_37__or_module_11_res), .ZN(
        n_majority7_module_37_res) );
  DFF_X1 u_reg_module_41__cini_mul_v00_reg ( .D(n_majority7_module_37_res), 
        .CK(clock_0), .Q(n_reg_module_41_res), .QN() );
  AND2_X1 u_majority7_module_38__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_38__and_module_1_res)
         );
  OR2_X1 u_majority7_module_38__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_38__or_module_1_res)
         );
  AND2_X1 u_majority7_module_38__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(n_majority7_module_38__and_module_2_res) );
  OR2_X1 u_majority7_module_38__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_38__or_module_2_res)
         );
  AND2_X1 u_majority7_module_38__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(n_majority7_module_38__and_module_3_res) );
  OR2_X1 u_majority7_module_38__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_38__or_module_3_res)
         );
  AND2_X1 u_majority7_module_38__and_module_4_U1 ( .A1(
        n_majority7_module_38__and_module_2_res), .A2(
        n_majority7_module_38__and_module_1_res), .ZN(
        n_majority7_module_38__and_module_4_res) );
  OR2_X1 u_majority7_module_38__or_module_4_U1 ( .A1(
        n_majority7_module_38__and_module_1_res), .A2(
        n_majority7_module_38__and_module_2_res), .ZN(
        n_majority7_module_38__or_module_4_res) );
  AND2_X1 u_majority7_module_38__and_module_5_U1 ( .A1(
        n_majority7_module_38__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_38__and_module_5_res) );
  OR2_X1 u_majority7_module_38__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_38__and_module_3_res), .ZN(
        n_majority7_module_38__or_module_5_res) );
  AND2_X1 u_majority7_module_38__and_module_6_U1 ( .A1(
        n_majority7_module_38__or_module_1_res), .A2(
        n_majority7_module_38__or_module_2_res), .ZN(
        n_majority7_module_38__and_module_6_res) );
  OR2_X1 u_majority7_module_38__or_module_6_U1 ( .A1(
        n_majority7_module_38__or_module_2_res), .A2(
        n_majority7_module_38__or_module_1_res), .ZN(
        n_majority7_module_38__or_module_6_res) );
  OR2_X1 u_majority7_module_38__or_module_7_U1 ( .A1(
        n_majority7_module_38__and_module_4_res), .A2(
        n_majority7_module_38__and_module_5_res), .ZN(
        n_majority7_module_38__or_module_7_res) );
  AND2_X1 u_majority7_module_38__and_module_7_U1 ( .A1(
        n_majority7_module_38__or_module_3_res), .A2(
        n_majority7_module_38__or_module_4_res), .ZN(
        n_majority7_module_38__and_module_7_res) );
  OR2_X1 u_majority7_module_38__or_module_8_U1 ( .A1(
        n_majority7_module_38__or_module_4_res), .A2(
        n_majority7_module_38__or_module_3_res), .ZN(
        n_majority7_module_38__or_module_8_res) );
  AND2_X1 u_majority7_module_38__and_module_8_U1 ( .A1(
        n_majority7_module_38__or_module_5_res), .A2(
        n_majority7_module_38__and_module_6_res), .ZN(
        n_majority7_module_38__and_module_8_res) );
  OR2_X1 u_majority7_module_38__or_module_9_U1 ( .A1(
        n_majority7_module_38__and_module_6_res), .A2(
        n_majority7_module_38__or_module_5_res), .ZN(
        n_majority7_module_38__or_module_9_res) );
  OR2_X1 u_majority7_module_38__or_module_10_U1 ( .A1(
        n_majority7_module_38__or_module_7_res), .A2(
        n_majority7_module_38__and_module_7_res), .ZN(
        n_majority7_module_38__or_module_10_res) );
  AND2_X1 u_majority7_module_38__and_module_9_U1 ( .A1(
        n_majority7_module_38__or_module_6_res), .A2(
        n_majority7_module_38__or_module_9_res), .ZN(
        n_majority7_module_38__and_module_9_res) );
  OR2_X1 u_majority7_module_38__or_module_11_U1 ( .A1(
        n_majority7_module_38__or_module_10_res), .A2(
        n_majority7_module_38__and_module_8_res), .ZN(
        n_majority7_module_38__or_module_11_res) );
  AND2_X1 u_majority7_module_38__and_module_10_U1 ( .A1(
        n_majority7_module_38__or_module_8_res), .A2(
        n_majority7_module_38__and_module_9_res), .ZN(
        n_majority7_module_38__and_module_10_res) );
  AND2_X1 u_majority7_module_38__and_module_11_U1 ( .A1(
        n_majority7_module_38__and_module_10_res), .A2(
        n_majority7_module_38__or_module_11_res), .ZN(
        n_majority7_module_38_res) );
  DFF_X1 u_reg_module_42__cini_mul_v00_reg ( .D(n_majority7_module_38_res), 
        .CK(clock_0), .Q(n_reg_module_42_res), .QN() );
  AND2_X1 u_majority7_module_39__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_39__and_module_1_res)
         );
  OR2_X1 u_majority7_module_39__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_39__or_module_1_res)
         );
  AND2_X1 u_majority7_module_39__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(n_majority7_module_39__and_module_2_res) );
  OR2_X1 u_majority7_module_39__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_39__or_module_2_res)
         );
  AND2_X1 u_majority7_module_39__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(n_majority7_module_39__and_module_3_res) );
  OR2_X1 u_majority7_module_39__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_39__or_module_3_res)
         );
  AND2_X1 u_majority7_module_39__and_module_4_U1 ( .A1(
        n_majority7_module_39__and_module_2_res), .A2(
        n_majority7_module_39__and_module_1_res), .ZN(
        n_majority7_module_39__and_module_4_res) );
  OR2_X1 u_majority7_module_39__or_module_4_U1 ( .A1(
        n_majority7_module_39__and_module_1_res), .A2(
        n_majority7_module_39__and_module_2_res), .ZN(
        n_majority7_module_39__or_module_4_res) );
  AND2_X1 u_majority7_module_39__and_module_5_U1 ( .A1(
        n_majority7_module_39__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_39__and_module_5_res) );
  OR2_X1 u_majority7_module_39__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_39__and_module_3_res), .ZN(
        n_majority7_module_39__or_module_5_res) );
  AND2_X1 u_majority7_module_39__and_module_6_U1 ( .A1(
        n_majority7_module_39__or_module_1_res), .A2(
        n_majority7_module_39__or_module_2_res), .ZN(
        n_majority7_module_39__and_module_6_res) );
  OR2_X1 u_majority7_module_39__or_module_6_U1 ( .A1(
        n_majority7_module_39__or_module_2_res), .A2(
        n_majority7_module_39__or_module_1_res), .ZN(
        n_majority7_module_39__or_module_6_res) );
  OR2_X1 u_majority7_module_39__or_module_7_U1 ( .A1(
        n_majority7_module_39__and_module_4_res), .A2(
        n_majority7_module_39__and_module_5_res), .ZN(
        n_majority7_module_39__or_module_7_res) );
  AND2_X1 u_majority7_module_39__and_module_7_U1 ( .A1(
        n_majority7_module_39__or_module_3_res), .A2(
        n_majority7_module_39__or_module_4_res), .ZN(
        n_majority7_module_39__and_module_7_res) );
  OR2_X1 u_majority7_module_39__or_module_8_U1 ( .A1(
        n_majority7_module_39__or_module_4_res), .A2(
        n_majority7_module_39__or_module_3_res), .ZN(
        n_majority7_module_39__or_module_8_res) );
  AND2_X1 u_majority7_module_39__and_module_8_U1 ( .A1(
        n_majority7_module_39__or_module_5_res), .A2(
        n_majority7_module_39__and_module_6_res), .ZN(
        n_majority7_module_39__and_module_8_res) );
  OR2_X1 u_majority7_module_39__or_module_9_U1 ( .A1(
        n_majority7_module_39__and_module_6_res), .A2(
        n_majority7_module_39__or_module_5_res), .ZN(
        n_majority7_module_39__or_module_9_res) );
  OR2_X1 u_majority7_module_39__or_module_10_U1 ( .A1(
        n_majority7_module_39__or_module_7_res), .A2(
        n_majority7_module_39__and_module_7_res), .ZN(
        n_majority7_module_39__or_module_10_res) );
  AND2_X1 u_majority7_module_39__and_module_9_U1 ( .A1(
        n_majority7_module_39__or_module_6_res), .A2(
        n_majority7_module_39__or_module_9_res), .ZN(
        n_majority7_module_39__and_module_9_res) );
  OR2_X1 u_majority7_module_39__or_module_11_U1 ( .A1(
        n_majority7_module_39__or_module_10_res), .A2(
        n_majority7_module_39__and_module_8_res), .ZN(
        n_majority7_module_39__or_module_11_res) );
  AND2_X1 u_majority7_module_39__and_module_10_U1 ( .A1(
        n_majority7_module_39__or_module_8_res), .A2(
        n_majority7_module_39__and_module_9_res), .ZN(
        n_majority7_module_39__and_module_10_res) );
  AND2_X1 u_majority7_module_39__and_module_11_U1 ( .A1(
        n_majority7_module_39__and_module_10_res), .A2(
        n_majority7_module_39__or_module_11_res), .ZN(
        n_majority7_module_39_res) );
  DFF_X1 u_reg_module_43__cini_mul_v00_reg ( .D(n_majority7_module_39_res), 
        .CK(clock_0), .Q(n_reg_module_43_res), .QN() );
  DFF_X1 u_reg_module_44__cini_mul_v00_reg ( .D(n_and_module_16_res), .CK(
        clock_0), .Q(n_reg_module_44_res), .QN() );
  DFF_X1 u_reg_module_45__cini_mul_v00_reg ( .D(n_and_module_17_res), .CK(
        clock_1), .Q(n_reg_module_45_res), .QN() );
  AND2_X1 u_majority7_module_40__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_40__and_module_1_res)
         );
  OR2_X1 u_majority7_module_40__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_40__or_module_1_res)
         );
  AND2_X1 u_majority7_module_40__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(n_majority7_module_40__and_module_2_res) );
  OR2_X1 u_majority7_module_40__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_40__or_module_2_res)
         );
  AND2_X1 u_majority7_module_40__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(n_majority7_module_40__and_module_3_res) );
  OR2_X1 u_majority7_module_40__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_40__or_module_3_res)
         );
  AND2_X1 u_majority7_module_40__and_module_4_U1 ( .A1(
        n_majority7_module_40__and_module_2_res), .A2(
        n_majority7_module_40__and_module_1_res), .ZN(
        n_majority7_module_40__and_module_4_res) );
  OR2_X1 u_majority7_module_40__or_module_4_U1 ( .A1(
        n_majority7_module_40__and_module_1_res), .A2(
        n_majority7_module_40__and_module_2_res), .ZN(
        n_majority7_module_40__or_module_4_res) );
  AND2_X1 u_majority7_module_40__and_module_5_U1 ( .A1(
        n_majority7_module_40__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_40__and_module_5_res) );
  OR2_X1 u_majority7_module_40__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_40__and_module_3_res), .ZN(
        n_majority7_module_40__or_module_5_res) );
  AND2_X1 u_majority7_module_40__and_module_6_U1 ( .A1(
        n_majority7_module_40__or_module_1_res), .A2(
        n_majority7_module_40__or_module_2_res), .ZN(
        n_majority7_module_40__and_module_6_res) );
  OR2_X1 u_majority7_module_40__or_module_6_U1 ( .A1(
        n_majority7_module_40__or_module_2_res), .A2(
        n_majority7_module_40__or_module_1_res), .ZN(
        n_majority7_module_40__or_module_6_res) );
  OR2_X1 u_majority7_module_40__or_module_7_U1 ( .A1(
        n_majority7_module_40__and_module_4_res), .A2(
        n_majority7_module_40__and_module_5_res), .ZN(
        n_majority7_module_40__or_module_7_res) );
  AND2_X1 u_majority7_module_40__and_module_7_U1 ( .A1(
        n_majority7_module_40__or_module_3_res), .A2(
        n_majority7_module_40__or_module_4_res), .ZN(
        n_majority7_module_40__and_module_7_res) );
  OR2_X1 u_majority7_module_40__or_module_8_U1 ( .A1(
        n_majority7_module_40__or_module_4_res), .A2(
        n_majority7_module_40__or_module_3_res), .ZN(
        n_majority7_module_40__or_module_8_res) );
  AND2_X1 u_majority7_module_40__and_module_8_U1 ( .A1(
        n_majority7_module_40__or_module_5_res), .A2(
        n_majority7_module_40__and_module_6_res), .ZN(
        n_majority7_module_40__and_module_8_res) );
  OR2_X1 u_majority7_module_40__or_module_9_U1 ( .A1(
        n_majority7_module_40__and_module_6_res), .A2(
        n_majority7_module_40__or_module_5_res), .ZN(
        n_majority7_module_40__or_module_9_res) );
  OR2_X1 u_majority7_module_40__or_module_10_U1 ( .A1(
        n_majority7_module_40__or_module_7_res), .A2(
        n_majority7_module_40__and_module_7_res), .ZN(
        n_majority7_module_40__or_module_10_res) );
  AND2_X1 u_majority7_module_40__and_module_9_U1 ( .A1(
        n_majority7_module_40__or_module_6_res), .A2(
        n_majority7_module_40__or_module_9_res), .ZN(
        n_majority7_module_40__and_module_9_res) );
  OR2_X1 u_majority7_module_40__or_module_11_U1 ( .A1(
        n_majority7_module_40__or_module_10_res), .A2(
        n_majority7_module_40__and_module_8_res), .ZN(
        n_majority7_module_40__or_module_11_res) );
  AND2_X1 u_majority7_module_40__and_module_10_U1 ( .A1(
        n_majority7_module_40__or_module_8_res), .A2(
        n_majority7_module_40__and_module_9_res), .ZN(
        n_majority7_module_40__and_module_10_res) );
  AND2_X1 u_majority7_module_40__and_module_11_U1 ( .A1(
        n_majority7_module_40__and_module_10_res), .A2(
        n_majority7_module_40__or_module_11_res), .ZN(
        n_majority7_module_40_res) );
  DFF_X1 u_reg_module_46__cini_mul_v00_reg ( .D(n_majority7_module_40_res), 
        .CK(clock_1), .Q(n_reg_module_46_res), .QN() );
  AND2_X1 u_majority7_module_41__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_41__and_module_1_res)
         );
  OR2_X1 u_majority7_module_41__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_41__or_module_1_res)
         );
  AND2_X1 u_majority7_module_41__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(n_majority7_module_41__and_module_2_res) );
  OR2_X1 u_majority7_module_41__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_41__or_module_2_res)
         );
  AND2_X1 u_majority7_module_41__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(n_majority7_module_41__and_module_3_res) );
  OR2_X1 u_majority7_module_41__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_41__or_module_3_res)
         );
  AND2_X1 u_majority7_module_41__and_module_4_U1 ( .A1(
        n_majority7_module_41__and_module_2_res), .A2(
        n_majority7_module_41__and_module_1_res), .ZN(
        n_majority7_module_41__and_module_4_res) );
  OR2_X1 u_majority7_module_41__or_module_4_U1 ( .A1(
        n_majority7_module_41__and_module_1_res), .A2(
        n_majority7_module_41__and_module_2_res), .ZN(
        n_majority7_module_41__or_module_4_res) );
  AND2_X1 u_majority7_module_41__and_module_5_U1 ( .A1(
        n_majority7_module_41__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_41__and_module_5_res) );
  OR2_X1 u_majority7_module_41__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_41__and_module_3_res), .ZN(
        n_majority7_module_41__or_module_5_res) );
  AND2_X1 u_majority7_module_41__and_module_6_U1 ( .A1(
        n_majority7_module_41__or_module_1_res), .A2(
        n_majority7_module_41__or_module_2_res), .ZN(
        n_majority7_module_41__and_module_6_res) );
  OR2_X1 u_majority7_module_41__or_module_6_U1 ( .A1(
        n_majority7_module_41__or_module_2_res), .A2(
        n_majority7_module_41__or_module_1_res), .ZN(
        n_majority7_module_41__or_module_6_res) );
  OR2_X1 u_majority7_module_41__or_module_7_U1 ( .A1(
        n_majority7_module_41__and_module_4_res), .A2(
        n_majority7_module_41__and_module_5_res), .ZN(
        n_majority7_module_41__or_module_7_res) );
  AND2_X1 u_majority7_module_41__and_module_7_U1 ( .A1(
        n_majority7_module_41__or_module_3_res), .A2(
        n_majority7_module_41__or_module_4_res), .ZN(
        n_majority7_module_41__and_module_7_res) );
  OR2_X1 u_majority7_module_41__or_module_8_U1 ( .A1(
        n_majority7_module_41__or_module_4_res), .A2(
        n_majority7_module_41__or_module_3_res), .ZN(
        n_majority7_module_41__or_module_8_res) );
  AND2_X1 u_majority7_module_41__and_module_8_U1 ( .A1(
        n_majority7_module_41__or_module_5_res), .A2(
        n_majority7_module_41__and_module_6_res), .ZN(
        n_majority7_module_41__and_module_8_res) );
  OR2_X1 u_majority7_module_41__or_module_9_U1 ( .A1(
        n_majority7_module_41__and_module_6_res), .A2(
        n_majority7_module_41__or_module_5_res), .ZN(
        n_majority7_module_41__or_module_9_res) );
  OR2_X1 u_majority7_module_41__or_module_10_U1 ( .A1(
        n_majority7_module_41__or_module_7_res), .A2(
        n_majority7_module_41__and_module_7_res), .ZN(
        n_majority7_module_41__or_module_10_res) );
  AND2_X1 u_majority7_module_41__and_module_9_U1 ( .A1(
        n_majority7_module_41__or_module_6_res), .A2(
        n_majority7_module_41__or_module_9_res), .ZN(
        n_majority7_module_41__and_module_9_res) );
  OR2_X1 u_majority7_module_41__or_module_11_U1 ( .A1(
        n_majority7_module_41__or_module_10_res), .A2(
        n_majority7_module_41__and_module_8_res), .ZN(
        n_majority7_module_41__or_module_11_res) );
  AND2_X1 u_majority7_module_41__and_module_10_U1 ( .A1(
        n_majority7_module_41__or_module_8_res), .A2(
        n_majority7_module_41__and_module_9_res), .ZN(
        n_majority7_module_41__and_module_10_res) );
  AND2_X1 u_majority7_module_41__and_module_11_U1 ( .A1(
        n_majority7_module_41__and_module_10_res), .A2(
        n_majority7_module_41__or_module_11_res), .ZN(
        n_majority7_module_41_res) );
  DFF_X1 u_reg_module_47__cini_mul_v00_reg ( .D(n_majority7_module_41_res), 
        .CK(clock_1), .Q(n_reg_module_47_res), .QN() );
  AND2_X1 u_majority7_module_42__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_42__and_module_1_res)
         );
  OR2_X1 u_majority7_module_42__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_42__or_module_1_res)
         );
  AND2_X1 u_majority7_module_42__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(n_majority7_module_42__and_module_2_res) );
  OR2_X1 u_majority7_module_42__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_42__or_module_2_res)
         );
  AND2_X1 u_majority7_module_42__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(n_majority7_module_42__and_module_3_res) );
  OR2_X1 u_majority7_module_42__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_42__or_module_3_res)
         );
  AND2_X1 u_majority7_module_42__and_module_4_U1 ( .A1(
        n_majority7_module_42__and_module_2_res), .A2(
        n_majority7_module_42__and_module_1_res), .ZN(
        n_majority7_module_42__and_module_4_res) );
  OR2_X1 u_majority7_module_42__or_module_4_U1 ( .A1(
        n_majority7_module_42__and_module_1_res), .A2(
        n_majority7_module_42__and_module_2_res), .ZN(
        n_majority7_module_42__or_module_4_res) );
  AND2_X1 u_majority7_module_42__and_module_5_U1 ( .A1(
        n_majority7_module_42__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_42__and_module_5_res) );
  OR2_X1 u_majority7_module_42__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_42__and_module_3_res), .ZN(
        n_majority7_module_42__or_module_5_res) );
  AND2_X1 u_majority7_module_42__and_module_6_U1 ( .A1(
        n_majority7_module_42__or_module_1_res), .A2(
        n_majority7_module_42__or_module_2_res), .ZN(
        n_majority7_module_42__and_module_6_res) );
  OR2_X1 u_majority7_module_42__or_module_6_U1 ( .A1(
        n_majority7_module_42__or_module_2_res), .A2(
        n_majority7_module_42__or_module_1_res), .ZN(
        n_majority7_module_42__or_module_6_res) );
  OR2_X1 u_majority7_module_42__or_module_7_U1 ( .A1(
        n_majority7_module_42__and_module_4_res), .A2(
        n_majority7_module_42__and_module_5_res), .ZN(
        n_majority7_module_42__or_module_7_res) );
  AND2_X1 u_majority7_module_42__and_module_7_U1 ( .A1(
        n_majority7_module_42__or_module_3_res), .A2(
        n_majority7_module_42__or_module_4_res), .ZN(
        n_majority7_module_42__and_module_7_res) );
  OR2_X1 u_majority7_module_42__or_module_8_U1 ( .A1(
        n_majority7_module_42__or_module_4_res), .A2(
        n_majority7_module_42__or_module_3_res), .ZN(
        n_majority7_module_42__or_module_8_res) );
  AND2_X1 u_majority7_module_42__and_module_8_U1 ( .A1(
        n_majority7_module_42__or_module_5_res), .A2(
        n_majority7_module_42__and_module_6_res), .ZN(
        n_majority7_module_42__and_module_8_res) );
  OR2_X1 u_majority7_module_42__or_module_9_U1 ( .A1(
        n_majority7_module_42__and_module_6_res), .A2(
        n_majority7_module_42__or_module_5_res), .ZN(
        n_majority7_module_42__or_module_9_res) );
  OR2_X1 u_majority7_module_42__or_module_10_U1 ( .A1(
        n_majority7_module_42__or_module_7_res), .A2(
        n_majority7_module_42__and_module_7_res), .ZN(
        n_majority7_module_42__or_module_10_res) );
  AND2_X1 u_majority7_module_42__and_module_9_U1 ( .A1(
        n_majority7_module_42__or_module_6_res), .A2(
        n_majority7_module_42__or_module_9_res), .ZN(
        n_majority7_module_42__and_module_9_res) );
  OR2_X1 u_majority7_module_42__or_module_11_U1 ( .A1(
        n_majority7_module_42__or_module_10_res), .A2(
        n_majority7_module_42__and_module_8_res), .ZN(
        n_majority7_module_42__or_module_11_res) );
  AND2_X1 u_majority7_module_42__and_module_10_U1 ( .A1(
        n_majority7_module_42__or_module_8_res), .A2(
        n_majority7_module_42__and_module_9_res), .ZN(
        n_majority7_module_42__and_module_10_res) );
  AND2_X1 u_majority7_module_42__and_module_11_U1 ( .A1(
        n_majority7_module_42__and_module_10_res), .A2(
        n_majority7_module_42__or_module_11_res), .ZN(
        n_majority7_module_42_res) );
  DFF_X1 u_reg_module_48__cini_mul_v00_reg ( .D(n_majority7_module_42_res), 
        .CK(clock_1), .Q(n_reg_module_48_res), .QN() );
  AND2_X1 u_majority7_module_43__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_43__and_module_1_res)
         );
  OR2_X1 u_majority7_module_43__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_43__or_module_1_res)
         );
  AND2_X1 u_majority7_module_43__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(n_majority7_module_43__and_module_2_res) );
  OR2_X1 u_majority7_module_43__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_43__or_module_2_res)
         );
  AND2_X1 u_majority7_module_43__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(n_majority7_module_43__and_module_3_res) );
  OR2_X1 u_majority7_module_43__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_43__or_module_3_res)
         );
  AND2_X1 u_majority7_module_43__and_module_4_U1 ( .A1(
        n_majority7_module_43__and_module_2_res), .A2(
        n_majority7_module_43__and_module_1_res), .ZN(
        n_majority7_module_43__and_module_4_res) );
  OR2_X1 u_majority7_module_43__or_module_4_U1 ( .A1(
        n_majority7_module_43__and_module_1_res), .A2(
        n_majority7_module_43__and_module_2_res), .ZN(
        n_majority7_module_43__or_module_4_res) );
  AND2_X1 u_majority7_module_43__and_module_5_U1 ( .A1(
        n_majority7_module_43__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_43__and_module_5_res) );
  OR2_X1 u_majority7_module_43__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_43__and_module_3_res), .ZN(
        n_majority7_module_43__or_module_5_res) );
  AND2_X1 u_majority7_module_43__and_module_6_U1 ( .A1(
        n_majority7_module_43__or_module_1_res), .A2(
        n_majority7_module_43__or_module_2_res), .ZN(
        n_majority7_module_43__and_module_6_res) );
  OR2_X1 u_majority7_module_43__or_module_6_U1 ( .A1(
        n_majority7_module_43__or_module_2_res), .A2(
        n_majority7_module_43__or_module_1_res), .ZN(
        n_majority7_module_43__or_module_6_res) );
  OR2_X1 u_majority7_module_43__or_module_7_U1 ( .A1(
        n_majority7_module_43__and_module_4_res), .A2(
        n_majority7_module_43__and_module_5_res), .ZN(
        n_majority7_module_43__or_module_7_res) );
  AND2_X1 u_majority7_module_43__and_module_7_U1 ( .A1(
        n_majority7_module_43__or_module_3_res), .A2(
        n_majority7_module_43__or_module_4_res), .ZN(
        n_majority7_module_43__and_module_7_res) );
  OR2_X1 u_majority7_module_43__or_module_8_U1 ( .A1(
        n_majority7_module_43__or_module_4_res), .A2(
        n_majority7_module_43__or_module_3_res), .ZN(
        n_majority7_module_43__or_module_8_res) );
  AND2_X1 u_majority7_module_43__and_module_8_U1 ( .A1(
        n_majority7_module_43__or_module_5_res), .A2(
        n_majority7_module_43__and_module_6_res), .ZN(
        n_majority7_module_43__and_module_8_res) );
  OR2_X1 u_majority7_module_43__or_module_9_U1 ( .A1(
        n_majority7_module_43__and_module_6_res), .A2(
        n_majority7_module_43__or_module_5_res), .ZN(
        n_majority7_module_43__or_module_9_res) );
  OR2_X1 u_majority7_module_43__or_module_10_U1 ( .A1(
        n_majority7_module_43__or_module_7_res), .A2(
        n_majority7_module_43__and_module_7_res), .ZN(
        n_majority7_module_43__or_module_10_res) );
  AND2_X1 u_majority7_module_43__and_module_9_U1 ( .A1(
        n_majority7_module_43__or_module_6_res), .A2(
        n_majority7_module_43__or_module_9_res), .ZN(
        n_majority7_module_43__and_module_9_res) );
  OR2_X1 u_majority7_module_43__or_module_11_U1 ( .A1(
        n_majority7_module_43__or_module_10_res), .A2(
        n_majority7_module_43__and_module_8_res), .ZN(
        n_majority7_module_43__or_module_11_res) );
  AND2_X1 u_majority7_module_43__and_module_10_U1 ( .A1(
        n_majority7_module_43__or_module_8_res), .A2(
        n_majority7_module_43__and_module_9_res), .ZN(
        n_majority7_module_43__and_module_10_res) );
  AND2_X1 u_majority7_module_43__and_module_11_U1 ( .A1(
        n_majority7_module_43__and_module_10_res), .A2(
        n_majority7_module_43__or_module_11_res), .ZN(
        n_majority7_module_43_res) );
  DFF_X1 u_reg_module_49__cini_mul_v00_reg ( .D(n_majority7_module_43_res), 
        .CK(clock_1), .Q(n_reg_module_49_res), .QN() );
  DFF_X1 u_reg_module_50__cini_mul_v00_reg ( .D(n_and_module_22_res), .CK(
        clock_1), .Q(n_reg_module_50_res), .QN() );
  AND2_X1 u_majority7_module_44__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_44__and_module_1_res)
         );
  OR2_X1 u_majority7_module_44__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_44__or_module_1_res)
         );
  AND2_X1 u_majority7_module_44__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(n_majority7_module_44__and_module_2_res) );
  OR2_X1 u_majority7_module_44__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_44__or_module_2_res)
         );
  AND2_X1 u_majority7_module_44__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(n_majority7_module_44__and_module_3_res) );
  OR2_X1 u_majority7_module_44__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_44__or_module_3_res)
         );
  AND2_X1 u_majority7_module_44__and_module_4_U1 ( .A1(
        n_majority7_module_44__and_module_2_res), .A2(
        n_majority7_module_44__and_module_1_res), .ZN(
        n_majority7_module_44__and_module_4_res) );
  OR2_X1 u_majority7_module_44__or_module_4_U1 ( .A1(
        n_majority7_module_44__and_module_1_res), .A2(
        n_majority7_module_44__and_module_2_res), .ZN(
        n_majority7_module_44__or_module_4_res) );
  AND2_X1 u_majority7_module_44__and_module_5_U1 ( .A1(
        n_majority7_module_44__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_44__and_module_5_res) );
  OR2_X1 u_majority7_module_44__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_44__and_module_3_res), .ZN(
        n_majority7_module_44__or_module_5_res) );
  AND2_X1 u_majority7_module_44__and_module_6_U1 ( .A1(
        n_majority7_module_44__or_module_1_res), .A2(
        n_majority7_module_44__or_module_2_res), .ZN(
        n_majority7_module_44__and_module_6_res) );
  OR2_X1 u_majority7_module_44__or_module_6_U1 ( .A1(
        n_majority7_module_44__or_module_2_res), .A2(
        n_majority7_module_44__or_module_1_res), .ZN(
        n_majority7_module_44__or_module_6_res) );
  OR2_X1 u_majority7_module_44__or_module_7_U1 ( .A1(
        n_majority7_module_44__and_module_4_res), .A2(
        n_majority7_module_44__and_module_5_res), .ZN(
        n_majority7_module_44__or_module_7_res) );
  AND2_X1 u_majority7_module_44__and_module_7_U1 ( .A1(
        n_majority7_module_44__or_module_3_res), .A2(
        n_majority7_module_44__or_module_4_res), .ZN(
        n_majority7_module_44__and_module_7_res) );
  OR2_X1 u_majority7_module_44__or_module_8_U1 ( .A1(
        n_majority7_module_44__or_module_4_res), .A2(
        n_majority7_module_44__or_module_3_res), .ZN(
        n_majority7_module_44__or_module_8_res) );
  AND2_X1 u_majority7_module_44__and_module_8_U1 ( .A1(
        n_majority7_module_44__or_module_5_res), .A2(
        n_majority7_module_44__and_module_6_res), .ZN(
        n_majority7_module_44__and_module_8_res) );
  OR2_X1 u_majority7_module_44__or_module_9_U1 ( .A1(
        n_majority7_module_44__and_module_6_res), .A2(
        n_majority7_module_44__or_module_5_res), .ZN(
        n_majority7_module_44__or_module_9_res) );
  OR2_X1 u_majority7_module_44__or_module_10_U1 ( .A1(
        n_majority7_module_44__or_module_7_res), .A2(
        n_majority7_module_44__and_module_7_res), .ZN(
        n_majority7_module_44__or_module_10_res) );
  AND2_X1 u_majority7_module_44__and_module_9_U1 ( .A1(
        n_majority7_module_44__or_module_6_res), .A2(
        n_majority7_module_44__or_module_9_res), .ZN(
        n_majority7_module_44__and_module_9_res) );
  OR2_X1 u_majority7_module_44__or_module_11_U1 ( .A1(
        n_majority7_module_44__or_module_10_res), .A2(
        n_majority7_module_44__and_module_8_res), .ZN(
        n_majority7_module_44__or_module_11_res) );
  AND2_X1 u_majority7_module_44__and_module_10_U1 ( .A1(
        n_majority7_module_44__or_module_8_res), .A2(
        n_majority7_module_44__and_module_9_res), .ZN(
        n_majority7_module_44__and_module_10_res) );
  AND2_X1 u_majority7_module_44__and_module_11_U1 ( .A1(
        n_majority7_module_44__and_module_10_res), .A2(
        n_majority7_module_44__or_module_11_res), .ZN(
        n_majority7_module_44_res) );
  DFF_X1 u_reg_module_51__cini_mul_v00_reg ( .D(n_majority7_module_44_res), 
        .CK(clock_1), .Q(n_reg_module_51_res), .QN() );
  AND2_X1 u_majority7_module_45__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_45__and_module_1_res)
         );
  OR2_X1 u_majority7_module_45__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_45__or_module_1_res)
         );
  AND2_X1 u_majority7_module_45__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(n_majority7_module_45__and_module_2_res) );
  OR2_X1 u_majority7_module_45__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_45__or_module_2_res)
         );
  AND2_X1 u_majority7_module_45__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(n_majority7_module_45__and_module_3_res) );
  OR2_X1 u_majority7_module_45__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_45__or_module_3_res)
         );
  AND2_X1 u_majority7_module_45__and_module_4_U1 ( .A1(
        n_majority7_module_45__and_module_2_res), .A2(
        n_majority7_module_45__and_module_1_res), .ZN(
        n_majority7_module_45__and_module_4_res) );
  OR2_X1 u_majority7_module_45__or_module_4_U1 ( .A1(
        n_majority7_module_45__and_module_1_res), .A2(
        n_majority7_module_45__and_module_2_res), .ZN(
        n_majority7_module_45__or_module_4_res) );
  AND2_X1 u_majority7_module_45__and_module_5_U1 ( .A1(
        n_majority7_module_45__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_45__and_module_5_res) );
  OR2_X1 u_majority7_module_45__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_45__and_module_3_res), .ZN(
        n_majority7_module_45__or_module_5_res) );
  AND2_X1 u_majority7_module_45__and_module_6_U1 ( .A1(
        n_majority7_module_45__or_module_1_res), .A2(
        n_majority7_module_45__or_module_2_res), .ZN(
        n_majority7_module_45__and_module_6_res) );
  OR2_X1 u_majority7_module_45__or_module_6_U1 ( .A1(
        n_majority7_module_45__or_module_2_res), .A2(
        n_majority7_module_45__or_module_1_res), .ZN(
        n_majority7_module_45__or_module_6_res) );
  OR2_X1 u_majority7_module_45__or_module_7_U1 ( .A1(
        n_majority7_module_45__and_module_4_res), .A2(
        n_majority7_module_45__and_module_5_res), .ZN(
        n_majority7_module_45__or_module_7_res) );
  AND2_X1 u_majority7_module_45__and_module_7_U1 ( .A1(
        n_majority7_module_45__or_module_3_res), .A2(
        n_majority7_module_45__or_module_4_res), .ZN(
        n_majority7_module_45__and_module_7_res) );
  OR2_X1 u_majority7_module_45__or_module_8_U1 ( .A1(
        n_majority7_module_45__or_module_4_res), .A2(
        n_majority7_module_45__or_module_3_res), .ZN(
        n_majority7_module_45__or_module_8_res) );
  AND2_X1 u_majority7_module_45__and_module_8_U1 ( .A1(
        n_majority7_module_45__or_module_5_res), .A2(
        n_majority7_module_45__and_module_6_res), .ZN(
        n_majority7_module_45__and_module_8_res) );
  OR2_X1 u_majority7_module_45__or_module_9_U1 ( .A1(
        n_majority7_module_45__and_module_6_res), .A2(
        n_majority7_module_45__or_module_5_res), .ZN(
        n_majority7_module_45__or_module_9_res) );
  OR2_X1 u_majority7_module_45__or_module_10_U1 ( .A1(
        n_majority7_module_45__or_module_7_res), .A2(
        n_majority7_module_45__and_module_7_res), .ZN(
        n_majority7_module_45__or_module_10_res) );
  AND2_X1 u_majority7_module_45__and_module_9_U1 ( .A1(
        n_majority7_module_45__or_module_6_res), .A2(
        n_majority7_module_45__or_module_9_res), .ZN(
        n_majority7_module_45__and_module_9_res) );
  OR2_X1 u_majority7_module_45__or_module_11_U1 ( .A1(
        n_majority7_module_45__or_module_10_res), .A2(
        n_majority7_module_45__and_module_8_res), .ZN(
        n_majority7_module_45__or_module_11_res) );
  AND2_X1 u_majority7_module_45__and_module_10_U1 ( .A1(
        n_majority7_module_45__or_module_8_res), .A2(
        n_majority7_module_45__and_module_9_res), .ZN(
        n_majority7_module_45__and_module_10_res) );
  AND2_X1 u_majority7_module_45__and_module_11_U1 ( .A1(
        n_majority7_module_45__and_module_10_res), .A2(
        n_majority7_module_45__or_module_11_res), .ZN(
        n_majority7_module_45_res) );
  DFF_X1 u_reg_module_52__cini_mul_v00_reg ( .D(n_majority7_module_45_res), 
        .CK(clock_1), .Q(n_reg_module_52_res), .QN() );
  AND2_X1 u_majority7_module_46__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_46__and_module_1_res)
         );
  OR2_X1 u_majority7_module_46__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_46__or_module_1_res)
         );
  AND2_X1 u_majority7_module_46__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(n_majority7_module_46__and_module_2_res) );
  OR2_X1 u_majority7_module_46__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_46__or_module_2_res)
         );
  AND2_X1 u_majority7_module_46__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(n_majority7_module_46__and_module_3_res) );
  OR2_X1 u_majority7_module_46__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_46__or_module_3_res)
         );
  AND2_X1 u_majority7_module_46__and_module_4_U1 ( .A1(
        n_majority7_module_46__and_module_2_res), .A2(
        n_majority7_module_46__and_module_1_res), .ZN(
        n_majority7_module_46__and_module_4_res) );
  OR2_X1 u_majority7_module_46__or_module_4_U1 ( .A1(
        n_majority7_module_46__and_module_1_res), .A2(
        n_majority7_module_46__and_module_2_res), .ZN(
        n_majority7_module_46__or_module_4_res) );
  AND2_X1 u_majority7_module_46__and_module_5_U1 ( .A1(
        n_majority7_module_46__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_46__and_module_5_res) );
  OR2_X1 u_majority7_module_46__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_46__and_module_3_res), .ZN(
        n_majority7_module_46__or_module_5_res) );
  AND2_X1 u_majority7_module_46__and_module_6_U1 ( .A1(
        n_majority7_module_46__or_module_1_res), .A2(
        n_majority7_module_46__or_module_2_res), .ZN(
        n_majority7_module_46__and_module_6_res) );
  OR2_X1 u_majority7_module_46__or_module_6_U1 ( .A1(
        n_majority7_module_46__or_module_2_res), .A2(
        n_majority7_module_46__or_module_1_res), .ZN(
        n_majority7_module_46__or_module_6_res) );
  OR2_X1 u_majority7_module_46__or_module_7_U1 ( .A1(
        n_majority7_module_46__and_module_4_res), .A2(
        n_majority7_module_46__and_module_5_res), .ZN(
        n_majority7_module_46__or_module_7_res) );
  AND2_X1 u_majority7_module_46__and_module_7_U1 ( .A1(
        n_majority7_module_46__or_module_3_res), .A2(
        n_majority7_module_46__or_module_4_res), .ZN(
        n_majority7_module_46__and_module_7_res) );
  OR2_X1 u_majority7_module_46__or_module_8_U1 ( .A1(
        n_majority7_module_46__or_module_4_res), .A2(
        n_majority7_module_46__or_module_3_res), .ZN(
        n_majority7_module_46__or_module_8_res) );
  AND2_X1 u_majority7_module_46__and_module_8_U1 ( .A1(
        n_majority7_module_46__or_module_5_res), .A2(
        n_majority7_module_46__and_module_6_res), .ZN(
        n_majority7_module_46__and_module_8_res) );
  OR2_X1 u_majority7_module_46__or_module_9_U1 ( .A1(
        n_majority7_module_46__and_module_6_res), .A2(
        n_majority7_module_46__or_module_5_res), .ZN(
        n_majority7_module_46__or_module_9_res) );
  OR2_X1 u_majority7_module_46__or_module_10_U1 ( .A1(
        n_majority7_module_46__or_module_7_res), .A2(
        n_majority7_module_46__and_module_7_res), .ZN(
        n_majority7_module_46__or_module_10_res) );
  AND2_X1 u_majority7_module_46__and_module_9_U1 ( .A1(
        n_majority7_module_46__or_module_6_res), .A2(
        n_majority7_module_46__or_module_9_res), .ZN(
        n_majority7_module_46__and_module_9_res) );
  OR2_X1 u_majority7_module_46__or_module_11_U1 ( .A1(
        n_majority7_module_46__or_module_10_res), .A2(
        n_majority7_module_46__and_module_8_res), .ZN(
        n_majority7_module_46__or_module_11_res) );
  AND2_X1 u_majority7_module_46__and_module_10_U1 ( .A1(
        n_majority7_module_46__or_module_8_res), .A2(
        n_majority7_module_46__and_module_9_res), .ZN(
        n_majority7_module_46__and_module_10_res) );
  AND2_X1 u_majority7_module_46__and_module_11_U1 ( .A1(
        n_majority7_module_46__and_module_10_res), .A2(
        n_majority7_module_46__or_module_11_res), .ZN(
        n_majority7_module_46_res) );
  DFF_X1 u_reg_module_53__cini_mul_v00_reg ( .D(n_majority7_module_46_res), 
        .CK(clock_1), .Q(n_reg_module_53_res), .QN() );
  AND2_X1 u_majority7_module_47__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_47__and_module_1_res)
         );
  OR2_X1 u_majority7_module_47__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_47__or_module_1_res)
         );
  AND2_X1 u_majority7_module_47__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(n_majority7_module_47__and_module_2_res) );
  OR2_X1 u_majority7_module_47__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_47__or_module_2_res)
         );
  AND2_X1 u_majority7_module_47__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(n_majority7_module_47__and_module_3_res) );
  OR2_X1 u_majority7_module_47__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_47__or_module_3_res)
         );
  AND2_X1 u_majority7_module_47__and_module_4_U1 ( .A1(
        n_majority7_module_47__and_module_2_res), .A2(
        n_majority7_module_47__and_module_1_res), .ZN(
        n_majority7_module_47__and_module_4_res) );
  OR2_X1 u_majority7_module_47__or_module_4_U1 ( .A1(
        n_majority7_module_47__and_module_1_res), .A2(
        n_majority7_module_47__and_module_2_res), .ZN(
        n_majority7_module_47__or_module_4_res) );
  AND2_X1 u_majority7_module_47__and_module_5_U1 ( .A1(
        n_majority7_module_47__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_47__and_module_5_res) );
  OR2_X1 u_majority7_module_47__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_47__and_module_3_res), .ZN(
        n_majority7_module_47__or_module_5_res) );
  AND2_X1 u_majority7_module_47__and_module_6_U1 ( .A1(
        n_majority7_module_47__or_module_1_res), .A2(
        n_majority7_module_47__or_module_2_res), .ZN(
        n_majority7_module_47__and_module_6_res) );
  OR2_X1 u_majority7_module_47__or_module_6_U1 ( .A1(
        n_majority7_module_47__or_module_2_res), .A2(
        n_majority7_module_47__or_module_1_res), .ZN(
        n_majority7_module_47__or_module_6_res) );
  OR2_X1 u_majority7_module_47__or_module_7_U1 ( .A1(
        n_majority7_module_47__and_module_4_res), .A2(
        n_majority7_module_47__and_module_5_res), .ZN(
        n_majority7_module_47__or_module_7_res) );
  AND2_X1 u_majority7_module_47__and_module_7_U1 ( .A1(
        n_majority7_module_47__or_module_3_res), .A2(
        n_majority7_module_47__or_module_4_res), .ZN(
        n_majority7_module_47__and_module_7_res) );
  OR2_X1 u_majority7_module_47__or_module_8_U1 ( .A1(
        n_majority7_module_47__or_module_4_res), .A2(
        n_majority7_module_47__or_module_3_res), .ZN(
        n_majority7_module_47__or_module_8_res) );
  AND2_X1 u_majority7_module_47__and_module_8_U1 ( .A1(
        n_majority7_module_47__or_module_5_res), .A2(
        n_majority7_module_47__and_module_6_res), .ZN(
        n_majority7_module_47__and_module_8_res) );
  OR2_X1 u_majority7_module_47__or_module_9_U1 ( .A1(
        n_majority7_module_47__and_module_6_res), .A2(
        n_majority7_module_47__or_module_5_res), .ZN(
        n_majority7_module_47__or_module_9_res) );
  OR2_X1 u_majority7_module_47__or_module_10_U1 ( .A1(
        n_majority7_module_47__or_module_7_res), .A2(
        n_majority7_module_47__and_module_7_res), .ZN(
        n_majority7_module_47__or_module_10_res) );
  AND2_X1 u_majority7_module_47__and_module_9_U1 ( .A1(
        n_majority7_module_47__or_module_6_res), .A2(
        n_majority7_module_47__or_module_9_res), .ZN(
        n_majority7_module_47__and_module_9_res) );
  OR2_X1 u_majority7_module_47__or_module_11_U1 ( .A1(
        n_majority7_module_47__or_module_10_res), .A2(
        n_majority7_module_47__and_module_8_res), .ZN(
        n_majority7_module_47__or_module_11_res) );
  AND2_X1 u_majority7_module_47__and_module_10_U1 ( .A1(
        n_majority7_module_47__or_module_8_res), .A2(
        n_majority7_module_47__and_module_9_res), .ZN(
        n_majority7_module_47__and_module_10_res) );
  AND2_X1 u_majority7_module_47__and_module_11_U1 ( .A1(
        n_majority7_module_47__and_module_10_res), .A2(
        n_majority7_module_47__or_module_11_res), .ZN(
        n_majority7_module_47_res) );
  DFF_X1 u_reg_module_54__cini_mul_v00_reg ( .D(n_majority7_module_47_res), 
        .CK(clock_1), .Q(n_reg_module_54_res), .QN() );
  DFF_X1 u_reg_module_55__cini_mul_v00_reg ( .D(n_and_module_27_res), .CK(
        clock_1), .Q(n_reg_module_55_res), .QN() );
  AND2_X1 u_majority7_module_48__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_48__and_module_1_res)
         );
  OR2_X1 u_majority7_module_48__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_48__or_module_1_res)
         );
  AND2_X1 u_majority7_module_48__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(n_majority7_module_48__and_module_2_res) );
  OR2_X1 u_majority7_module_48__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_48__or_module_2_res)
         );
  AND2_X1 u_majority7_module_48__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(n_majority7_module_48__and_module_3_res) );
  OR2_X1 u_majority7_module_48__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_48__or_module_3_res)
         );
  AND2_X1 u_majority7_module_48__and_module_4_U1 ( .A1(
        n_majority7_module_48__and_module_2_res), .A2(
        n_majority7_module_48__and_module_1_res), .ZN(
        n_majority7_module_48__and_module_4_res) );
  OR2_X1 u_majority7_module_48__or_module_4_U1 ( .A1(
        n_majority7_module_48__and_module_1_res), .A2(
        n_majority7_module_48__and_module_2_res), .ZN(
        n_majority7_module_48__or_module_4_res) );
  AND2_X1 u_majority7_module_48__and_module_5_U1 ( .A1(
        n_majority7_module_48__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_48__and_module_5_res) );
  OR2_X1 u_majority7_module_48__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_48__and_module_3_res), .ZN(
        n_majority7_module_48__or_module_5_res) );
  AND2_X1 u_majority7_module_48__and_module_6_U1 ( .A1(
        n_majority7_module_48__or_module_1_res), .A2(
        n_majority7_module_48__or_module_2_res), .ZN(
        n_majority7_module_48__and_module_6_res) );
  OR2_X1 u_majority7_module_48__or_module_6_U1 ( .A1(
        n_majority7_module_48__or_module_2_res), .A2(
        n_majority7_module_48__or_module_1_res), .ZN(
        n_majority7_module_48__or_module_6_res) );
  OR2_X1 u_majority7_module_48__or_module_7_U1 ( .A1(
        n_majority7_module_48__and_module_4_res), .A2(
        n_majority7_module_48__and_module_5_res), .ZN(
        n_majority7_module_48__or_module_7_res) );
  AND2_X1 u_majority7_module_48__and_module_7_U1 ( .A1(
        n_majority7_module_48__or_module_3_res), .A2(
        n_majority7_module_48__or_module_4_res), .ZN(
        n_majority7_module_48__and_module_7_res) );
  OR2_X1 u_majority7_module_48__or_module_8_U1 ( .A1(
        n_majority7_module_48__or_module_4_res), .A2(
        n_majority7_module_48__or_module_3_res), .ZN(
        n_majority7_module_48__or_module_8_res) );
  AND2_X1 u_majority7_module_48__and_module_8_U1 ( .A1(
        n_majority7_module_48__or_module_5_res), .A2(
        n_majority7_module_48__and_module_6_res), .ZN(
        n_majority7_module_48__and_module_8_res) );
  OR2_X1 u_majority7_module_48__or_module_9_U1 ( .A1(
        n_majority7_module_48__and_module_6_res), .A2(
        n_majority7_module_48__or_module_5_res), .ZN(
        n_majority7_module_48__or_module_9_res) );
  OR2_X1 u_majority7_module_48__or_module_10_U1 ( .A1(
        n_majority7_module_48__or_module_7_res), .A2(
        n_majority7_module_48__and_module_7_res), .ZN(
        n_majority7_module_48__or_module_10_res) );
  AND2_X1 u_majority7_module_48__and_module_9_U1 ( .A1(
        n_majority7_module_48__or_module_6_res), .A2(
        n_majority7_module_48__or_module_9_res), .ZN(
        n_majority7_module_48__and_module_9_res) );
  OR2_X1 u_majority7_module_48__or_module_11_U1 ( .A1(
        n_majority7_module_48__or_module_10_res), .A2(
        n_majority7_module_48__and_module_8_res), .ZN(
        n_majority7_module_48__or_module_11_res) );
  AND2_X1 u_majority7_module_48__and_module_10_U1 ( .A1(
        n_majority7_module_48__or_module_8_res), .A2(
        n_majority7_module_48__and_module_9_res), .ZN(
        n_majority7_module_48__and_module_10_res) );
  AND2_X1 u_majority7_module_48__and_module_11_U1 ( .A1(
        n_majority7_module_48__and_module_10_res), .A2(
        n_majority7_module_48__or_module_11_res), .ZN(
        n_majority7_module_48_res) );
  DFF_X1 u_reg_module_56__cini_mul_v00_reg ( .D(n_majority7_module_48_res), 
        .CK(clock_1), .Q(n_reg_module_56_res), .QN() );
  AND2_X1 u_majority7_module_49__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_49__and_module_1_res)
         );
  OR2_X1 u_majority7_module_49__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_49__or_module_1_res)
         );
  AND2_X1 u_majority7_module_49__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(n_majority7_module_49__and_module_2_res) );
  OR2_X1 u_majority7_module_49__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_49__or_module_2_res)
         );
  AND2_X1 u_majority7_module_49__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(n_majority7_module_49__and_module_3_res) );
  OR2_X1 u_majority7_module_49__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_49__or_module_3_res)
         );
  AND2_X1 u_majority7_module_49__and_module_4_U1 ( .A1(
        n_majority7_module_49__and_module_2_res), .A2(
        n_majority7_module_49__and_module_1_res), .ZN(
        n_majority7_module_49__and_module_4_res) );
  OR2_X1 u_majority7_module_49__or_module_4_U1 ( .A1(
        n_majority7_module_49__and_module_1_res), .A2(
        n_majority7_module_49__and_module_2_res), .ZN(
        n_majority7_module_49__or_module_4_res) );
  AND2_X1 u_majority7_module_49__and_module_5_U1 ( .A1(
        n_majority7_module_49__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_49__and_module_5_res) );
  OR2_X1 u_majority7_module_49__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_49__and_module_3_res), .ZN(
        n_majority7_module_49__or_module_5_res) );
  AND2_X1 u_majority7_module_49__and_module_6_U1 ( .A1(
        n_majority7_module_49__or_module_1_res), .A2(
        n_majority7_module_49__or_module_2_res), .ZN(
        n_majority7_module_49__and_module_6_res) );
  OR2_X1 u_majority7_module_49__or_module_6_U1 ( .A1(
        n_majority7_module_49__or_module_2_res), .A2(
        n_majority7_module_49__or_module_1_res), .ZN(
        n_majority7_module_49__or_module_6_res) );
  OR2_X1 u_majority7_module_49__or_module_7_U1 ( .A1(
        n_majority7_module_49__and_module_4_res), .A2(
        n_majority7_module_49__and_module_5_res), .ZN(
        n_majority7_module_49__or_module_7_res) );
  AND2_X1 u_majority7_module_49__and_module_7_U1 ( .A1(
        n_majority7_module_49__or_module_3_res), .A2(
        n_majority7_module_49__or_module_4_res), .ZN(
        n_majority7_module_49__and_module_7_res) );
  OR2_X1 u_majority7_module_49__or_module_8_U1 ( .A1(
        n_majority7_module_49__or_module_4_res), .A2(
        n_majority7_module_49__or_module_3_res), .ZN(
        n_majority7_module_49__or_module_8_res) );
  AND2_X1 u_majority7_module_49__and_module_8_U1 ( .A1(
        n_majority7_module_49__or_module_5_res), .A2(
        n_majority7_module_49__and_module_6_res), .ZN(
        n_majority7_module_49__and_module_8_res) );
  OR2_X1 u_majority7_module_49__or_module_9_U1 ( .A1(
        n_majority7_module_49__and_module_6_res), .A2(
        n_majority7_module_49__or_module_5_res), .ZN(
        n_majority7_module_49__or_module_9_res) );
  OR2_X1 u_majority7_module_49__or_module_10_U1 ( .A1(
        n_majority7_module_49__or_module_7_res), .A2(
        n_majority7_module_49__and_module_7_res), .ZN(
        n_majority7_module_49__or_module_10_res) );
  AND2_X1 u_majority7_module_49__and_module_9_U1 ( .A1(
        n_majority7_module_49__or_module_6_res), .A2(
        n_majority7_module_49__or_module_9_res), .ZN(
        n_majority7_module_49__and_module_9_res) );
  OR2_X1 u_majority7_module_49__or_module_11_U1 ( .A1(
        n_majority7_module_49__or_module_10_res), .A2(
        n_majority7_module_49__and_module_8_res), .ZN(
        n_majority7_module_49__or_module_11_res) );
  AND2_X1 u_majority7_module_49__and_module_10_U1 ( .A1(
        n_majority7_module_49__or_module_8_res), .A2(
        n_majority7_module_49__and_module_9_res), .ZN(
        n_majority7_module_49__and_module_10_res) );
  AND2_X1 u_majority7_module_49__and_module_11_U1 ( .A1(
        n_majority7_module_49__and_module_10_res), .A2(
        n_majority7_module_49__or_module_11_res), .ZN(
        n_majority7_module_49_res) );
  DFF_X1 u_reg_module_57__cini_mul_v00_reg ( .D(n_majority7_module_49_res), 
        .CK(clock_1), .Q(n_reg_module_57_res), .QN() );
  AND2_X1 u_majority7_module_50__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_50__and_module_1_res)
         );
  OR2_X1 u_majority7_module_50__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_50__or_module_1_res)
         );
  AND2_X1 u_majority7_module_50__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(n_majority7_module_50__and_module_2_res) );
  OR2_X1 u_majority7_module_50__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_50__or_module_2_res)
         );
  AND2_X1 u_majority7_module_50__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(n_majority7_module_50__and_module_3_res) );
  OR2_X1 u_majority7_module_50__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_50__or_module_3_res)
         );
  AND2_X1 u_majority7_module_50__and_module_4_U1 ( .A1(
        n_majority7_module_50__and_module_2_res), .A2(
        n_majority7_module_50__and_module_1_res), .ZN(
        n_majority7_module_50__and_module_4_res) );
  OR2_X1 u_majority7_module_50__or_module_4_U1 ( .A1(
        n_majority7_module_50__and_module_1_res), .A2(
        n_majority7_module_50__and_module_2_res), .ZN(
        n_majority7_module_50__or_module_4_res) );
  AND2_X1 u_majority7_module_50__and_module_5_U1 ( .A1(
        n_majority7_module_50__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_50__and_module_5_res) );
  OR2_X1 u_majority7_module_50__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_50__and_module_3_res), .ZN(
        n_majority7_module_50__or_module_5_res) );
  AND2_X1 u_majority7_module_50__and_module_6_U1 ( .A1(
        n_majority7_module_50__or_module_1_res), .A2(
        n_majority7_module_50__or_module_2_res), .ZN(
        n_majority7_module_50__and_module_6_res) );
  OR2_X1 u_majority7_module_50__or_module_6_U1 ( .A1(
        n_majority7_module_50__or_module_2_res), .A2(
        n_majority7_module_50__or_module_1_res), .ZN(
        n_majority7_module_50__or_module_6_res) );
  OR2_X1 u_majority7_module_50__or_module_7_U1 ( .A1(
        n_majority7_module_50__and_module_4_res), .A2(
        n_majority7_module_50__and_module_5_res), .ZN(
        n_majority7_module_50__or_module_7_res) );
  AND2_X1 u_majority7_module_50__and_module_7_U1 ( .A1(
        n_majority7_module_50__or_module_3_res), .A2(
        n_majority7_module_50__or_module_4_res), .ZN(
        n_majority7_module_50__and_module_7_res) );
  OR2_X1 u_majority7_module_50__or_module_8_U1 ( .A1(
        n_majority7_module_50__or_module_4_res), .A2(
        n_majority7_module_50__or_module_3_res), .ZN(
        n_majority7_module_50__or_module_8_res) );
  AND2_X1 u_majority7_module_50__and_module_8_U1 ( .A1(
        n_majority7_module_50__or_module_5_res), .A2(
        n_majority7_module_50__and_module_6_res), .ZN(
        n_majority7_module_50__and_module_8_res) );
  OR2_X1 u_majority7_module_50__or_module_9_U1 ( .A1(
        n_majority7_module_50__and_module_6_res), .A2(
        n_majority7_module_50__or_module_5_res), .ZN(
        n_majority7_module_50__or_module_9_res) );
  OR2_X1 u_majority7_module_50__or_module_10_U1 ( .A1(
        n_majority7_module_50__or_module_7_res), .A2(
        n_majority7_module_50__and_module_7_res), .ZN(
        n_majority7_module_50__or_module_10_res) );
  AND2_X1 u_majority7_module_50__and_module_9_U1 ( .A1(
        n_majority7_module_50__or_module_6_res), .A2(
        n_majority7_module_50__or_module_9_res), .ZN(
        n_majority7_module_50__and_module_9_res) );
  OR2_X1 u_majority7_module_50__or_module_11_U1 ( .A1(
        n_majority7_module_50__or_module_10_res), .A2(
        n_majority7_module_50__and_module_8_res), .ZN(
        n_majority7_module_50__or_module_11_res) );
  AND2_X1 u_majority7_module_50__and_module_10_U1 ( .A1(
        n_majority7_module_50__or_module_8_res), .A2(
        n_majority7_module_50__and_module_9_res), .ZN(
        n_majority7_module_50__and_module_10_res) );
  AND2_X1 u_majority7_module_50__and_module_11_U1 ( .A1(
        n_majority7_module_50__and_module_10_res), .A2(
        n_majority7_module_50__or_module_11_res), .ZN(
        n_majority7_module_50_res) );
  DFF_X1 u_reg_module_58__cini_mul_v00_reg ( .D(n_majority7_module_50_res), 
        .CK(clock_1), .Q(n_reg_module_58_res), .QN() );
  AND2_X1 u_majority7_module_51__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_51__and_module_1_res)
         );
  OR2_X1 u_majority7_module_51__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_51__or_module_1_res)
         );
  AND2_X1 u_majority7_module_51__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(n_majority7_module_51__and_module_2_res) );
  OR2_X1 u_majority7_module_51__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_51__or_module_2_res)
         );
  AND2_X1 u_majority7_module_51__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(n_majority7_module_51__and_module_3_res) );
  OR2_X1 u_majority7_module_51__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_51__or_module_3_res)
         );
  AND2_X1 u_majority7_module_51__and_module_4_U1 ( .A1(
        n_majority7_module_51__and_module_2_res), .A2(
        n_majority7_module_51__and_module_1_res), .ZN(
        n_majority7_module_51__and_module_4_res) );
  OR2_X1 u_majority7_module_51__or_module_4_U1 ( .A1(
        n_majority7_module_51__and_module_1_res), .A2(
        n_majority7_module_51__and_module_2_res), .ZN(
        n_majority7_module_51__or_module_4_res) );
  AND2_X1 u_majority7_module_51__and_module_5_U1 ( .A1(
        n_majority7_module_51__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_51__and_module_5_res) );
  OR2_X1 u_majority7_module_51__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_51__and_module_3_res), .ZN(
        n_majority7_module_51__or_module_5_res) );
  AND2_X1 u_majority7_module_51__and_module_6_U1 ( .A1(
        n_majority7_module_51__or_module_1_res), .A2(
        n_majority7_module_51__or_module_2_res), .ZN(
        n_majority7_module_51__and_module_6_res) );
  OR2_X1 u_majority7_module_51__or_module_6_U1 ( .A1(
        n_majority7_module_51__or_module_2_res), .A2(
        n_majority7_module_51__or_module_1_res), .ZN(
        n_majority7_module_51__or_module_6_res) );
  OR2_X1 u_majority7_module_51__or_module_7_U1 ( .A1(
        n_majority7_module_51__and_module_4_res), .A2(
        n_majority7_module_51__and_module_5_res), .ZN(
        n_majority7_module_51__or_module_7_res) );
  AND2_X1 u_majority7_module_51__and_module_7_U1 ( .A1(
        n_majority7_module_51__or_module_3_res), .A2(
        n_majority7_module_51__or_module_4_res), .ZN(
        n_majority7_module_51__and_module_7_res) );
  OR2_X1 u_majority7_module_51__or_module_8_U1 ( .A1(
        n_majority7_module_51__or_module_4_res), .A2(
        n_majority7_module_51__or_module_3_res), .ZN(
        n_majority7_module_51__or_module_8_res) );
  AND2_X1 u_majority7_module_51__and_module_8_U1 ( .A1(
        n_majority7_module_51__or_module_5_res), .A2(
        n_majority7_module_51__and_module_6_res), .ZN(
        n_majority7_module_51__and_module_8_res) );
  OR2_X1 u_majority7_module_51__or_module_9_U1 ( .A1(
        n_majority7_module_51__and_module_6_res), .A2(
        n_majority7_module_51__or_module_5_res), .ZN(
        n_majority7_module_51__or_module_9_res) );
  OR2_X1 u_majority7_module_51__or_module_10_U1 ( .A1(
        n_majority7_module_51__or_module_7_res), .A2(
        n_majority7_module_51__and_module_7_res), .ZN(
        n_majority7_module_51__or_module_10_res) );
  AND2_X1 u_majority7_module_51__and_module_9_U1 ( .A1(
        n_majority7_module_51__or_module_6_res), .A2(
        n_majority7_module_51__or_module_9_res), .ZN(
        n_majority7_module_51__and_module_9_res) );
  OR2_X1 u_majority7_module_51__or_module_11_U1 ( .A1(
        n_majority7_module_51__or_module_10_res), .A2(
        n_majority7_module_51__and_module_8_res), .ZN(
        n_majority7_module_51__or_module_11_res) );
  AND2_X1 u_majority7_module_51__and_module_10_U1 ( .A1(
        n_majority7_module_51__or_module_8_res), .A2(
        n_majority7_module_51__and_module_9_res), .ZN(
        n_majority7_module_51__and_module_10_res) );
  AND2_X1 u_majority7_module_51__and_module_11_U1 ( .A1(
        n_majority7_module_51__and_module_10_res), .A2(
        n_majority7_module_51__or_module_11_res), .ZN(
        n_majority7_module_51_res) );
  DFF_X1 u_reg_module_59__cini_mul_v00_reg ( .D(n_majority7_module_51_res), 
        .CK(clock_1), .Q(n_reg_module_59_res), .QN() );
  DFF_X1 u_reg_module_60__cini_mul_v00_reg ( .D(n_and_module_32_res), .CK(
        clock_1), .Q(n_reg_module_60_res), .QN() );
  DFF_X1 u_reg_module_61__cini_mul_v00_reg ( .D(n_and_module_33_res), .CK(
        clock_2), .Q(n_reg_module_61_res), .QN() );
  AND2_X1 u_majority7_module_52__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_52__and_module_1_res)
         );
  OR2_X1 u_majority7_module_52__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_52__or_module_1_res)
         );
  AND2_X1 u_majority7_module_52__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(n_majority7_module_52__and_module_2_res) );
  OR2_X1 u_majority7_module_52__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_52__or_module_2_res)
         );
  AND2_X1 u_majority7_module_52__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(n_majority7_module_52__and_module_3_res) );
  OR2_X1 u_majority7_module_52__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_52__or_module_3_res)
         );
  AND2_X1 u_majority7_module_52__and_module_4_U1 ( .A1(
        n_majority7_module_52__and_module_2_res), .A2(
        n_majority7_module_52__and_module_1_res), .ZN(
        n_majority7_module_52__and_module_4_res) );
  OR2_X1 u_majority7_module_52__or_module_4_U1 ( .A1(
        n_majority7_module_52__and_module_1_res), .A2(
        n_majority7_module_52__and_module_2_res), .ZN(
        n_majority7_module_52__or_module_4_res) );
  AND2_X1 u_majority7_module_52__and_module_5_U1 ( .A1(
        n_majority7_module_52__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_52__and_module_5_res) );
  OR2_X1 u_majority7_module_52__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_52__and_module_3_res), .ZN(
        n_majority7_module_52__or_module_5_res) );
  AND2_X1 u_majority7_module_52__and_module_6_U1 ( .A1(
        n_majority7_module_52__or_module_1_res), .A2(
        n_majority7_module_52__or_module_2_res), .ZN(
        n_majority7_module_52__and_module_6_res) );
  OR2_X1 u_majority7_module_52__or_module_6_U1 ( .A1(
        n_majority7_module_52__or_module_2_res), .A2(
        n_majority7_module_52__or_module_1_res), .ZN(
        n_majority7_module_52__or_module_6_res) );
  OR2_X1 u_majority7_module_52__or_module_7_U1 ( .A1(
        n_majority7_module_52__and_module_4_res), .A2(
        n_majority7_module_52__and_module_5_res), .ZN(
        n_majority7_module_52__or_module_7_res) );
  AND2_X1 u_majority7_module_52__and_module_7_U1 ( .A1(
        n_majority7_module_52__or_module_3_res), .A2(
        n_majority7_module_52__or_module_4_res), .ZN(
        n_majority7_module_52__and_module_7_res) );
  OR2_X1 u_majority7_module_52__or_module_8_U1 ( .A1(
        n_majority7_module_52__or_module_4_res), .A2(
        n_majority7_module_52__or_module_3_res), .ZN(
        n_majority7_module_52__or_module_8_res) );
  AND2_X1 u_majority7_module_52__and_module_8_U1 ( .A1(
        n_majority7_module_52__or_module_5_res), .A2(
        n_majority7_module_52__and_module_6_res), .ZN(
        n_majority7_module_52__and_module_8_res) );
  OR2_X1 u_majority7_module_52__or_module_9_U1 ( .A1(
        n_majority7_module_52__and_module_6_res), .A2(
        n_majority7_module_52__or_module_5_res), .ZN(
        n_majority7_module_52__or_module_9_res) );
  OR2_X1 u_majority7_module_52__or_module_10_U1 ( .A1(
        n_majority7_module_52__or_module_7_res), .A2(
        n_majority7_module_52__and_module_7_res), .ZN(
        n_majority7_module_52__or_module_10_res) );
  AND2_X1 u_majority7_module_52__and_module_9_U1 ( .A1(
        n_majority7_module_52__or_module_6_res), .A2(
        n_majority7_module_52__or_module_9_res), .ZN(
        n_majority7_module_52__and_module_9_res) );
  OR2_X1 u_majority7_module_52__or_module_11_U1 ( .A1(
        n_majority7_module_52__or_module_10_res), .A2(
        n_majority7_module_52__and_module_8_res), .ZN(
        n_majority7_module_52__or_module_11_res) );
  AND2_X1 u_majority7_module_52__and_module_10_U1 ( .A1(
        n_majority7_module_52__or_module_8_res), .A2(
        n_majority7_module_52__and_module_9_res), .ZN(
        n_majority7_module_52__and_module_10_res) );
  AND2_X1 u_majority7_module_52__and_module_11_U1 ( .A1(
        n_majority7_module_52__and_module_10_res), .A2(
        n_majority7_module_52__or_module_11_res), .ZN(
        n_majority7_module_52_res) );
  DFF_X1 u_reg_module_62__cini_mul_v00_reg ( .D(n_majority7_module_52_res), 
        .CK(clock_2), .Q(n_reg_module_62_res), .QN() );
  AND2_X1 u_majority7_module_53__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_53__and_module_1_res)
         );
  OR2_X1 u_majority7_module_53__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_53__or_module_1_res)
         );
  AND2_X1 u_majority7_module_53__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(n_majority7_module_53__and_module_2_res) );
  OR2_X1 u_majority7_module_53__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_53__or_module_2_res)
         );
  AND2_X1 u_majority7_module_53__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(n_majority7_module_53__and_module_3_res) );
  OR2_X1 u_majority7_module_53__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_53__or_module_3_res)
         );
  AND2_X1 u_majority7_module_53__and_module_4_U1 ( .A1(
        n_majority7_module_53__and_module_2_res), .A2(
        n_majority7_module_53__and_module_1_res), .ZN(
        n_majority7_module_53__and_module_4_res) );
  OR2_X1 u_majority7_module_53__or_module_4_U1 ( .A1(
        n_majority7_module_53__and_module_1_res), .A2(
        n_majority7_module_53__and_module_2_res), .ZN(
        n_majority7_module_53__or_module_4_res) );
  AND2_X1 u_majority7_module_53__and_module_5_U1 ( .A1(
        n_majority7_module_53__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_53__and_module_5_res) );
  OR2_X1 u_majority7_module_53__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_53__and_module_3_res), .ZN(
        n_majority7_module_53__or_module_5_res) );
  AND2_X1 u_majority7_module_53__and_module_6_U1 ( .A1(
        n_majority7_module_53__or_module_1_res), .A2(
        n_majority7_module_53__or_module_2_res), .ZN(
        n_majority7_module_53__and_module_6_res) );
  OR2_X1 u_majority7_module_53__or_module_6_U1 ( .A1(
        n_majority7_module_53__or_module_2_res), .A2(
        n_majority7_module_53__or_module_1_res), .ZN(
        n_majority7_module_53__or_module_6_res) );
  OR2_X1 u_majority7_module_53__or_module_7_U1 ( .A1(
        n_majority7_module_53__and_module_4_res), .A2(
        n_majority7_module_53__and_module_5_res), .ZN(
        n_majority7_module_53__or_module_7_res) );
  AND2_X1 u_majority7_module_53__and_module_7_U1 ( .A1(
        n_majority7_module_53__or_module_3_res), .A2(
        n_majority7_module_53__or_module_4_res), .ZN(
        n_majority7_module_53__and_module_7_res) );
  OR2_X1 u_majority7_module_53__or_module_8_U1 ( .A1(
        n_majority7_module_53__or_module_4_res), .A2(
        n_majority7_module_53__or_module_3_res), .ZN(
        n_majority7_module_53__or_module_8_res) );
  AND2_X1 u_majority7_module_53__and_module_8_U1 ( .A1(
        n_majority7_module_53__or_module_5_res), .A2(
        n_majority7_module_53__and_module_6_res), .ZN(
        n_majority7_module_53__and_module_8_res) );
  OR2_X1 u_majority7_module_53__or_module_9_U1 ( .A1(
        n_majority7_module_53__and_module_6_res), .A2(
        n_majority7_module_53__or_module_5_res), .ZN(
        n_majority7_module_53__or_module_9_res) );
  OR2_X1 u_majority7_module_53__or_module_10_U1 ( .A1(
        n_majority7_module_53__or_module_7_res), .A2(
        n_majority7_module_53__and_module_7_res), .ZN(
        n_majority7_module_53__or_module_10_res) );
  AND2_X1 u_majority7_module_53__and_module_9_U1 ( .A1(
        n_majority7_module_53__or_module_6_res), .A2(
        n_majority7_module_53__or_module_9_res), .ZN(
        n_majority7_module_53__and_module_9_res) );
  OR2_X1 u_majority7_module_53__or_module_11_U1 ( .A1(
        n_majority7_module_53__or_module_10_res), .A2(
        n_majority7_module_53__and_module_8_res), .ZN(
        n_majority7_module_53__or_module_11_res) );
  AND2_X1 u_majority7_module_53__and_module_10_U1 ( .A1(
        n_majority7_module_53__or_module_8_res), .A2(
        n_majority7_module_53__and_module_9_res), .ZN(
        n_majority7_module_53__and_module_10_res) );
  AND2_X1 u_majority7_module_53__and_module_11_U1 ( .A1(
        n_majority7_module_53__and_module_10_res), .A2(
        n_majority7_module_53__or_module_11_res), .ZN(
        n_majority7_module_53_res) );
  DFF_X1 u_reg_module_63__cini_mul_v00_reg ( .D(n_majority7_module_53_res), 
        .CK(clock_2), .Q(n_reg_module_63_res), .QN() );
  AND2_X1 u_majority7_module_54__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_54__and_module_1_res)
         );
  OR2_X1 u_majority7_module_54__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_54__or_module_1_res)
         );
  AND2_X1 u_majority7_module_54__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(n_majority7_module_54__and_module_2_res) );
  OR2_X1 u_majority7_module_54__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_54__or_module_2_res)
         );
  AND2_X1 u_majority7_module_54__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(n_majority7_module_54__and_module_3_res) );
  OR2_X1 u_majority7_module_54__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_54__or_module_3_res)
         );
  AND2_X1 u_majority7_module_54__and_module_4_U1 ( .A1(
        n_majority7_module_54__and_module_2_res), .A2(
        n_majority7_module_54__and_module_1_res), .ZN(
        n_majority7_module_54__and_module_4_res) );
  OR2_X1 u_majority7_module_54__or_module_4_U1 ( .A1(
        n_majority7_module_54__and_module_1_res), .A2(
        n_majority7_module_54__and_module_2_res), .ZN(
        n_majority7_module_54__or_module_4_res) );
  AND2_X1 u_majority7_module_54__and_module_5_U1 ( .A1(
        n_majority7_module_54__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_54__and_module_5_res) );
  OR2_X1 u_majority7_module_54__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_54__and_module_3_res), .ZN(
        n_majority7_module_54__or_module_5_res) );
  AND2_X1 u_majority7_module_54__and_module_6_U1 ( .A1(
        n_majority7_module_54__or_module_1_res), .A2(
        n_majority7_module_54__or_module_2_res), .ZN(
        n_majority7_module_54__and_module_6_res) );
  OR2_X1 u_majority7_module_54__or_module_6_U1 ( .A1(
        n_majority7_module_54__or_module_2_res), .A2(
        n_majority7_module_54__or_module_1_res), .ZN(
        n_majority7_module_54__or_module_6_res) );
  OR2_X1 u_majority7_module_54__or_module_7_U1 ( .A1(
        n_majority7_module_54__and_module_4_res), .A2(
        n_majority7_module_54__and_module_5_res), .ZN(
        n_majority7_module_54__or_module_7_res) );
  AND2_X1 u_majority7_module_54__and_module_7_U1 ( .A1(
        n_majority7_module_54__or_module_3_res), .A2(
        n_majority7_module_54__or_module_4_res), .ZN(
        n_majority7_module_54__and_module_7_res) );
  OR2_X1 u_majority7_module_54__or_module_8_U1 ( .A1(
        n_majority7_module_54__or_module_4_res), .A2(
        n_majority7_module_54__or_module_3_res), .ZN(
        n_majority7_module_54__or_module_8_res) );
  AND2_X1 u_majority7_module_54__and_module_8_U1 ( .A1(
        n_majority7_module_54__or_module_5_res), .A2(
        n_majority7_module_54__and_module_6_res), .ZN(
        n_majority7_module_54__and_module_8_res) );
  OR2_X1 u_majority7_module_54__or_module_9_U1 ( .A1(
        n_majority7_module_54__and_module_6_res), .A2(
        n_majority7_module_54__or_module_5_res), .ZN(
        n_majority7_module_54__or_module_9_res) );
  OR2_X1 u_majority7_module_54__or_module_10_U1 ( .A1(
        n_majority7_module_54__or_module_7_res), .A2(
        n_majority7_module_54__and_module_7_res), .ZN(
        n_majority7_module_54__or_module_10_res) );
  AND2_X1 u_majority7_module_54__and_module_9_U1 ( .A1(
        n_majority7_module_54__or_module_6_res), .A2(
        n_majority7_module_54__or_module_9_res), .ZN(
        n_majority7_module_54__and_module_9_res) );
  OR2_X1 u_majority7_module_54__or_module_11_U1 ( .A1(
        n_majority7_module_54__or_module_10_res), .A2(
        n_majority7_module_54__and_module_8_res), .ZN(
        n_majority7_module_54__or_module_11_res) );
  AND2_X1 u_majority7_module_54__and_module_10_U1 ( .A1(
        n_majority7_module_54__or_module_8_res), .A2(
        n_majority7_module_54__and_module_9_res), .ZN(
        n_majority7_module_54__and_module_10_res) );
  AND2_X1 u_majority7_module_54__and_module_11_U1 ( .A1(
        n_majority7_module_54__and_module_10_res), .A2(
        n_majority7_module_54__or_module_11_res), .ZN(
        n_majority7_module_54_res) );
  DFF_X1 u_reg_module_64__cini_mul_v00_reg ( .D(n_majority7_module_54_res), 
        .CK(clock_2), .Q(n_reg_module_64_res), .QN() );
  AND2_X1 u_majority7_module_55__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_55__and_module_1_res)
         );
  OR2_X1 u_majority7_module_55__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_55__or_module_1_res)
         );
  AND2_X1 u_majority7_module_55__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(n_majority7_module_55__and_module_2_res) );
  OR2_X1 u_majority7_module_55__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_55__or_module_2_res)
         );
  AND2_X1 u_majority7_module_55__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(n_majority7_module_55__and_module_3_res) );
  OR2_X1 u_majority7_module_55__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_55__or_module_3_res)
         );
  AND2_X1 u_majority7_module_55__and_module_4_U1 ( .A1(
        n_majority7_module_55__and_module_2_res), .A2(
        n_majority7_module_55__and_module_1_res), .ZN(
        n_majority7_module_55__and_module_4_res) );
  OR2_X1 u_majority7_module_55__or_module_4_U1 ( .A1(
        n_majority7_module_55__and_module_1_res), .A2(
        n_majority7_module_55__and_module_2_res), .ZN(
        n_majority7_module_55__or_module_4_res) );
  AND2_X1 u_majority7_module_55__and_module_5_U1 ( .A1(
        n_majority7_module_55__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_55__and_module_5_res) );
  OR2_X1 u_majority7_module_55__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_55__and_module_3_res), .ZN(
        n_majority7_module_55__or_module_5_res) );
  AND2_X1 u_majority7_module_55__and_module_6_U1 ( .A1(
        n_majority7_module_55__or_module_1_res), .A2(
        n_majority7_module_55__or_module_2_res), .ZN(
        n_majority7_module_55__and_module_6_res) );
  OR2_X1 u_majority7_module_55__or_module_6_U1 ( .A1(
        n_majority7_module_55__or_module_2_res), .A2(
        n_majority7_module_55__or_module_1_res), .ZN(
        n_majority7_module_55__or_module_6_res) );
  OR2_X1 u_majority7_module_55__or_module_7_U1 ( .A1(
        n_majority7_module_55__and_module_4_res), .A2(
        n_majority7_module_55__and_module_5_res), .ZN(
        n_majority7_module_55__or_module_7_res) );
  AND2_X1 u_majority7_module_55__and_module_7_U1 ( .A1(
        n_majority7_module_55__or_module_3_res), .A2(
        n_majority7_module_55__or_module_4_res), .ZN(
        n_majority7_module_55__and_module_7_res) );
  OR2_X1 u_majority7_module_55__or_module_8_U1 ( .A1(
        n_majority7_module_55__or_module_4_res), .A2(
        n_majority7_module_55__or_module_3_res), .ZN(
        n_majority7_module_55__or_module_8_res) );
  AND2_X1 u_majority7_module_55__and_module_8_U1 ( .A1(
        n_majority7_module_55__or_module_5_res), .A2(
        n_majority7_module_55__and_module_6_res), .ZN(
        n_majority7_module_55__and_module_8_res) );
  OR2_X1 u_majority7_module_55__or_module_9_U1 ( .A1(
        n_majority7_module_55__and_module_6_res), .A2(
        n_majority7_module_55__or_module_5_res), .ZN(
        n_majority7_module_55__or_module_9_res) );
  OR2_X1 u_majority7_module_55__or_module_10_U1 ( .A1(
        n_majority7_module_55__or_module_7_res), .A2(
        n_majority7_module_55__and_module_7_res), .ZN(
        n_majority7_module_55__or_module_10_res) );
  AND2_X1 u_majority7_module_55__and_module_9_U1 ( .A1(
        n_majority7_module_55__or_module_6_res), .A2(
        n_majority7_module_55__or_module_9_res), .ZN(
        n_majority7_module_55__and_module_9_res) );
  OR2_X1 u_majority7_module_55__or_module_11_U1 ( .A1(
        n_majority7_module_55__or_module_10_res), .A2(
        n_majority7_module_55__and_module_8_res), .ZN(
        n_majority7_module_55__or_module_11_res) );
  AND2_X1 u_majority7_module_55__and_module_10_U1 ( .A1(
        n_majority7_module_55__or_module_8_res), .A2(
        n_majority7_module_55__and_module_9_res), .ZN(
        n_majority7_module_55__and_module_10_res) );
  AND2_X1 u_majority7_module_55__and_module_11_U1 ( .A1(
        n_majority7_module_55__and_module_10_res), .A2(
        n_majority7_module_55__or_module_11_res), .ZN(
        n_majority7_module_55_res) );
  DFF_X1 u_reg_module_65__cini_mul_v00_reg ( .D(n_majority7_module_55_res), 
        .CK(clock_2), .Q(n_reg_module_65_res), .QN() );
  DFF_X1 u_reg_module_66__cini_mul_v00_reg ( .D(n_and_module_38_res), .CK(
        clock_2), .Q(n_reg_module_66_res), .QN() );
  AND2_X1 u_majority7_module_56__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_56__and_module_1_res)
         );
  OR2_X1 u_majority7_module_56__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_56__or_module_1_res)
         );
  AND2_X1 u_majority7_module_56__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(n_majority7_module_56__and_module_2_res) );
  OR2_X1 u_majority7_module_56__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_56__or_module_2_res)
         );
  AND2_X1 u_majority7_module_56__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(n_majority7_module_56__and_module_3_res) );
  OR2_X1 u_majority7_module_56__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_56__or_module_3_res)
         );
  AND2_X1 u_majority7_module_56__and_module_4_U1 ( .A1(
        n_majority7_module_56__and_module_2_res), .A2(
        n_majority7_module_56__and_module_1_res), .ZN(
        n_majority7_module_56__and_module_4_res) );
  OR2_X1 u_majority7_module_56__or_module_4_U1 ( .A1(
        n_majority7_module_56__and_module_1_res), .A2(
        n_majority7_module_56__and_module_2_res), .ZN(
        n_majority7_module_56__or_module_4_res) );
  AND2_X1 u_majority7_module_56__and_module_5_U1 ( .A1(
        n_majority7_module_56__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_56__and_module_5_res) );
  OR2_X1 u_majority7_module_56__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_56__and_module_3_res), .ZN(
        n_majority7_module_56__or_module_5_res) );
  AND2_X1 u_majority7_module_56__and_module_6_U1 ( .A1(
        n_majority7_module_56__or_module_1_res), .A2(
        n_majority7_module_56__or_module_2_res), .ZN(
        n_majority7_module_56__and_module_6_res) );
  OR2_X1 u_majority7_module_56__or_module_6_U1 ( .A1(
        n_majority7_module_56__or_module_2_res), .A2(
        n_majority7_module_56__or_module_1_res), .ZN(
        n_majority7_module_56__or_module_6_res) );
  OR2_X1 u_majority7_module_56__or_module_7_U1 ( .A1(
        n_majority7_module_56__and_module_4_res), .A2(
        n_majority7_module_56__and_module_5_res), .ZN(
        n_majority7_module_56__or_module_7_res) );
  AND2_X1 u_majority7_module_56__and_module_7_U1 ( .A1(
        n_majority7_module_56__or_module_3_res), .A2(
        n_majority7_module_56__or_module_4_res), .ZN(
        n_majority7_module_56__and_module_7_res) );
  OR2_X1 u_majority7_module_56__or_module_8_U1 ( .A1(
        n_majority7_module_56__or_module_4_res), .A2(
        n_majority7_module_56__or_module_3_res), .ZN(
        n_majority7_module_56__or_module_8_res) );
  AND2_X1 u_majority7_module_56__and_module_8_U1 ( .A1(
        n_majority7_module_56__or_module_5_res), .A2(
        n_majority7_module_56__and_module_6_res), .ZN(
        n_majority7_module_56__and_module_8_res) );
  OR2_X1 u_majority7_module_56__or_module_9_U1 ( .A1(
        n_majority7_module_56__and_module_6_res), .A2(
        n_majority7_module_56__or_module_5_res), .ZN(
        n_majority7_module_56__or_module_9_res) );
  OR2_X1 u_majority7_module_56__or_module_10_U1 ( .A1(
        n_majority7_module_56__or_module_7_res), .A2(
        n_majority7_module_56__and_module_7_res), .ZN(
        n_majority7_module_56__or_module_10_res) );
  AND2_X1 u_majority7_module_56__and_module_9_U1 ( .A1(
        n_majority7_module_56__or_module_6_res), .A2(
        n_majority7_module_56__or_module_9_res), .ZN(
        n_majority7_module_56__and_module_9_res) );
  OR2_X1 u_majority7_module_56__or_module_11_U1 ( .A1(
        n_majority7_module_56__or_module_10_res), .A2(
        n_majority7_module_56__and_module_8_res), .ZN(
        n_majority7_module_56__or_module_11_res) );
  AND2_X1 u_majority7_module_56__and_module_10_U1 ( .A1(
        n_majority7_module_56__or_module_8_res), .A2(
        n_majority7_module_56__and_module_9_res), .ZN(
        n_majority7_module_56__and_module_10_res) );
  AND2_X1 u_majority7_module_56__and_module_11_U1 ( .A1(
        n_majority7_module_56__and_module_10_res), .A2(
        n_majority7_module_56__or_module_11_res), .ZN(
        n_majority7_module_56_res) );
  DFF_X1 u_reg_module_67__cini_mul_v00_reg ( .D(n_majority7_module_56_res), 
        .CK(clock_2), .Q(n_reg_module_67_res), .QN() );
  AND2_X1 u_majority7_module_57__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_57__and_module_1_res)
         );
  OR2_X1 u_majority7_module_57__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_57__or_module_1_res)
         );
  AND2_X1 u_majority7_module_57__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(n_majority7_module_57__and_module_2_res) );
  OR2_X1 u_majority7_module_57__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_57__or_module_2_res)
         );
  AND2_X1 u_majority7_module_57__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(n_majority7_module_57__and_module_3_res) );
  OR2_X1 u_majority7_module_57__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_57__or_module_3_res)
         );
  AND2_X1 u_majority7_module_57__and_module_4_U1 ( .A1(
        n_majority7_module_57__and_module_2_res), .A2(
        n_majority7_module_57__and_module_1_res), .ZN(
        n_majority7_module_57__and_module_4_res) );
  OR2_X1 u_majority7_module_57__or_module_4_U1 ( .A1(
        n_majority7_module_57__and_module_1_res), .A2(
        n_majority7_module_57__and_module_2_res), .ZN(
        n_majority7_module_57__or_module_4_res) );
  AND2_X1 u_majority7_module_57__and_module_5_U1 ( .A1(
        n_majority7_module_57__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_57__and_module_5_res) );
  OR2_X1 u_majority7_module_57__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_57__and_module_3_res), .ZN(
        n_majority7_module_57__or_module_5_res) );
  AND2_X1 u_majority7_module_57__and_module_6_U1 ( .A1(
        n_majority7_module_57__or_module_1_res), .A2(
        n_majority7_module_57__or_module_2_res), .ZN(
        n_majority7_module_57__and_module_6_res) );
  OR2_X1 u_majority7_module_57__or_module_6_U1 ( .A1(
        n_majority7_module_57__or_module_2_res), .A2(
        n_majority7_module_57__or_module_1_res), .ZN(
        n_majority7_module_57__or_module_6_res) );
  OR2_X1 u_majority7_module_57__or_module_7_U1 ( .A1(
        n_majority7_module_57__and_module_4_res), .A2(
        n_majority7_module_57__and_module_5_res), .ZN(
        n_majority7_module_57__or_module_7_res) );
  AND2_X1 u_majority7_module_57__and_module_7_U1 ( .A1(
        n_majority7_module_57__or_module_3_res), .A2(
        n_majority7_module_57__or_module_4_res), .ZN(
        n_majority7_module_57__and_module_7_res) );
  OR2_X1 u_majority7_module_57__or_module_8_U1 ( .A1(
        n_majority7_module_57__or_module_4_res), .A2(
        n_majority7_module_57__or_module_3_res), .ZN(
        n_majority7_module_57__or_module_8_res) );
  AND2_X1 u_majority7_module_57__and_module_8_U1 ( .A1(
        n_majority7_module_57__or_module_5_res), .A2(
        n_majority7_module_57__and_module_6_res), .ZN(
        n_majority7_module_57__and_module_8_res) );
  OR2_X1 u_majority7_module_57__or_module_9_U1 ( .A1(
        n_majority7_module_57__and_module_6_res), .A2(
        n_majority7_module_57__or_module_5_res), .ZN(
        n_majority7_module_57__or_module_9_res) );
  OR2_X1 u_majority7_module_57__or_module_10_U1 ( .A1(
        n_majority7_module_57__or_module_7_res), .A2(
        n_majority7_module_57__and_module_7_res), .ZN(
        n_majority7_module_57__or_module_10_res) );
  AND2_X1 u_majority7_module_57__and_module_9_U1 ( .A1(
        n_majority7_module_57__or_module_6_res), .A2(
        n_majority7_module_57__or_module_9_res), .ZN(
        n_majority7_module_57__and_module_9_res) );
  OR2_X1 u_majority7_module_57__or_module_11_U1 ( .A1(
        n_majority7_module_57__or_module_10_res), .A2(
        n_majority7_module_57__and_module_8_res), .ZN(
        n_majority7_module_57__or_module_11_res) );
  AND2_X1 u_majority7_module_57__and_module_10_U1 ( .A1(
        n_majority7_module_57__or_module_8_res), .A2(
        n_majority7_module_57__and_module_9_res), .ZN(
        n_majority7_module_57__and_module_10_res) );
  AND2_X1 u_majority7_module_57__and_module_11_U1 ( .A1(
        n_majority7_module_57__and_module_10_res), .A2(
        n_majority7_module_57__or_module_11_res), .ZN(
        n_majority7_module_57_res) );
  DFF_X1 u_reg_module_68__cini_mul_v00_reg ( .D(n_majority7_module_57_res), 
        .CK(clock_2), .Q(n_reg_module_68_res), .QN() );
  AND2_X1 u_majority7_module_58__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_58__and_module_1_res)
         );
  OR2_X1 u_majority7_module_58__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_58__or_module_1_res)
         );
  AND2_X1 u_majority7_module_58__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(n_majority7_module_58__and_module_2_res) );
  OR2_X1 u_majority7_module_58__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_58__or_module_2_res)
         );
  AND2_X1 u_majority7_module_58__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(n_majority7_module_58__and_module_3_res) );
  OR2_X1 u_majority7_module_58__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_58__or_module_3_res)
         );
  AND2_X1 u_majority7_module_58__and_module_4_U1 ( .A1(
        n_majority7_module_58__and_module_2_res), .A2(
        n_majority7_module_58__and_module_1_res), .ZN(
        n_majority7_module_58__and_module_4_res) );
  OR2_X1 u_majority7_module_58__or_module_4_U1 ( .A1(
        n_majority7_module_58__and_module_1_res), .A2(
        n_majority7_module_58__and_module_2_res), .ZN(
        n_majority7_module_58__or_module_4_res) );
  AND2_X1 u_majority7_module_58__and_module_5_U1 ( .A1(
        n_majority7_module_58__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_58__and_module_5_res) );
  OR2_X1 u_majority7_module_58__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_58__and_module_3_res), .ZN(
        n_majority7_module_58__or_module_5_res) );
  AND2_X1 u_majority7_module_58__and_module_6_U1 ( .A1(
        n_majority7_module_58__or_module_1_res), .A2(
        n_majority7_module_58__or_module_2_res), .ZN(
        n_majority7_module_58__and_module_6_res) );
  OR2_X1 u_majority7_module_58__or_module_6_U1 ( .A1(
        n_majority7_module_58__or_module_2_res), .A2(
        n_majority7_module_58__or_module_1_res), .ZN(
        n_majority7_module_58__or_module_6_res) );
  OR2_X1 u_majority7_module_58__or_module_7_U1 ( .A1(
        n_majority7_module_58__and_module_4_res), .A2(
        n_majority7_module_58__and_module_5_res), .ZN(
        n_majority7_module_58__or_module_7_res) );
  AND2_X1 u_majority7_module_58__and_module_7_U1 ( .A1(
        n_majority7_module_58__or_module_3_res), .A2(
        n_majority7_module_58__or_module_4_res), .ZN(
        n_majority7_module_58__and_module_7_res) );
  OR2_X1 u_majority7_module_58__or_module_8_U1 ( .A1(
        n_majority7_module_58__or_module_4_res), .A2(
        n_majority7_module_58__or_module_3_res), .ZN(
        n_majority7_module_58__or_module_8_res) );
  AND2_X1 u_majority7_module_58__and_module_8_U1 ( .A1(
        n_majority7_module_58__or_module_5_res), .A2(
        n_majority7_module_58__and_module_6_res), .ZN(
        n_majority7_module_58__and_module_8_res) );
  OR2_X1 u_majority7_module_58__or_module_9_U1 ( .A1(
        n_majority7_module_58__and_module_6_res), .A2(
        n_majority7_module_58__or_module_5_res), .ZN(
        n_majority7_module_58__or_module_9_res) );
  OR2_X1 u_majority7_module_58__or_module_10_U1 ( .A1(
        n_majority7_module_58__or_module_7_res), .A2(
        n_majority7_module_58__and_module_7_res), .ZN(
        n_majority7_module_58__or_module_10_res) );
  AND2_X1 u_majority7_module_58__and_module_9_U1 ( .A1(
        n_majority7_module_58__or_module_6_res), .A2(
        n_majority7_module_58__or_module_9_res), .ZN(
        n_majority7_module_58__and_module_9_res) );
  OR2_X1 u_majority7_module_58__or_module_11_U1 ( .A1(
        n_majority7_module_58__or_module_10_res), .A2(
        n_majority7_module_58__and_module_8_res), .ZN(
        n_majority7_module_58__or_module_11_res) );
  AND2_X1 u_majority7_module_58__and_module_10_U1 ( .A1(
        n_majority7_module_58__or_module_8_res), .A2(
        n_majority7_module_58__and_module_9_res), .ZN(
        n_majority7_module_58__and_module_10_res) );
  AND2_X1 u_majority7_module_58__and_module_11_U1 ( .A1(
        n_majority7_module_58__and_module_10_res), .A2(
        n_majority7_module_58__or_module_11_res), .ZN(
        n_majority7_module_58_res) );
  DFF_X1 u_reg_module_69__cini_mul_v00_reg ( .D(n_majority7_module_58_res), 
        .CK(clock_2), .Q(n_reg_module_69_res), .QN() );
  AND2_X1 u_majority7_module_59__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_59__and_module_1_res)
         );
  OR2_X1 u_majority7_module_59__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_59__or_module_1_res)
         );
  AND2_X1 u_majority7_module_59__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(n_majority7_module_59__and_module_2_res) );
  OR2_X1 u_majority7_module_59__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_59__or_module_2_res)
         );
  AND2_X1 u_majority7_module_59__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(n_majority7_module_59__and_module_3_res) );
  OR2_X1 u_majority7_module_59__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_59__or_module_3_res)
         );
  AND2_X1 u_majority7_module_59__and_module_4_U1 ( .A1(
        n_majority7_module_59__and_module_2_res), .A2(
        n_majority7_module_59__and_module_1_res), .ZN(
        n_majority7_module_59__and_module_4_res) );
  OR2_X1 u_majority7_module_59__or_module_4_U1 ( .A1(
        n_majority7_module_59__and_module_1_res), .A2(
        n_majority7_module_59__and_module_2_res), .ZN(
        n_majority7_module_59__or_module_4_res) );
  AND2_X1 u_majority7_module_59__and_module_5_U1 ( .A1(
        n_majority7_module_59__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_59__and_module_5_res) );
  OR2_X1 u_majority7_module_59__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_59__and_module_3_res), .ZN(
        n_majority7_module_59__or_module_5_res) );
  AND2_X1 u_majority7_module_59__and_module_6_U1 ( .A1(
        n_majority7_module_59__or_module_1_res), .A2(
        n_majority7_module_59__or_module_2_res), .ZN(
        n_majority7_module_59__and_module_6_res) );
  OR2_X1 u_majority7_module_59__or_module_6_U1 ( .A1(
        n_majority7_module_59__or_module_2_res), .A2(
        n_majority7_module_59__or_module_1_res), .ZN(
        n_majority7_module_59__or_module_6_res) );
  OR2_X1 u_majority7_module_59__or_module_7_U1 ( .A1(
        n_majority7_module_59__and_module_4_res), .A2(
        n_majority7_module_59__and_module_5_res), .ZN(
        n_majority7_module_59__or_module_7_res) );
  AND2_X1 u_majority7_module_59__and_module_7_U1 ( .A1(
        n_majority7_module_59__or_module_3_res), .A2(
        n_majority7_module_59__or_module_4_res), .ZN(
        n_majority7_module_59__and_module_7_res) );
  OR2_X1 u_majority7_module_59__or_module_8_U1 ( .A1(
        n_majority7_module_59__or_module_4_res), .A2(
        n_majority7_module_59__or_module_3_res), .ZN(
        n_majority7_module_59__or_module_8_res) );
  AND2_X1 u_majority7_module_59__and_module_8_U1 ( .A1(
        n_majority7_module_59__or_module_5_res), .A2(
        n_majority7_module_59__and_module_6_res), .ZN(
        n_majority7_module_59__and_module_8_res) );
  OR2_X1 u_majority7_module_59__or_module_9_U1 ( .A1(
        n_majority7_module_59__and_module_6_res), .A2(
        n_majority7_module_59__or_module_5_res), .ZN(
        n_majority7_module_59__or_module_9_res) );
  OR2_X1 u_majority7_module_59__or_module_10_U1 ( .A1(
        n_majority7_module_59__or_module_7_res), .A2(
        n_majority7_module_59__and_module_7_res), .ZN(
        n_majority7_module_59__or_module_10_res) );
  AND2_X1 u_majority7_module_59__and_module_9_U1 ( .A1(
        n_majority7_module_59__or_module_6_res), .A2(
        n_majority7_module_59__or_module_9_res), .ZN(
        n_majority7_module_59__and_module_9_res) );
  OR2_X1 u_majority7_module_59__or_module_11_U1 ( .A1(
        n_majority7_module_59__or_module_10_res), .A2(
        n_majority7_module_59__and_module_8_res), .ZN(
        n_majority7_module_59__or_module_11_res) );
  AND2_X1 u_majority7_module_59__and_module_10_U1 ( .A1(
        n_majority7_module_59__or_module_8_res), .A2(
        n_majority7_module_59__and_module_9_res), .ZN(
        n_majority7_module_59__and_module_10_res) );
  AND2_X1 u_majority7_module_59__and_module_11_U1 ( .A1(
        n_majority7_module_59__and_module_10_res), .A2(
        n_majority7_module_59__or_module_11_res), .ZN(
        n_majority7_module_59_res) );
  DFF_X1 u_reg_module_70__cini_mul_v00_reg ( .D(n_majority7_module_59_res), 
        .CK(clock_2), .Q(n_reg_module_70_res), .QN() );
  DFF_X1 u_reg_module_71__cini_mul_v00_reg ( .D(n_and_module_43_res), .CK(
        clock_2), .Q(n_reg_module_71_res), .QN() );
  AND2_X1 u_majority7_module_60__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_60__and_module_1_res)
         );
  OR2_X1 u_majority7_module_60__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_60__or_module_1_res)
         );
  AND2_X1 u_majority7_module_60__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(n_majority7_module_60__and_module_2_res) );
  OR2_X1 u_majority7_module_60__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_60__or_module_2_res)
         );
  AND2_X1 u_majority7_module_60__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(n_majority7_module_60__and_module_3_res) );
  OR2_X1 u_majority7_module_60__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_60__or_module_3_res)
         );
  AND2_X1 u_majority7_module_60__and_module_4_U1 ( .A1(
        n_majority7_module_60__and_module_2_res), .A2(
        n_majority7_module_60__and_module_1_res), .ZN(
        n_majority7_module_60__and_module_4_res) );
  OR2_X1 u_majority7_module_60__or_module_4_U1 ( .A1(
        n_majority7_module_60__and_module_1_res), .A2(
        n_majority7_module_60__and_module_2_res), .ZN(
        n_majority7_module_60__or_module_4_res) );
  AND2_X1 u_majority7_module_60__and_module_5_U1 ( .A1(
        n_majority7_module_60__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_60__and_module_5_res) );
  OR2_X1 u_majority7_module_60__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_60__and_module_3_res), .ZN(
        n_majority7_module_60__or_module_5_res) );
  AND2_X1 u_majority7_module_60__and_module_6_U1 ( .A1(
        n_majority7_module_60__or_module_1_res), .A2(
        n_majority7_module_60__or_module_2_res), .ZN(
        n_majority7_module_60__and_module_6_res) );
  OR2_X1 u_majority7_module_60__or_module_6_U1 ( .A1(
        n_majority7_module_60__or_module_2_res), .A2(
        n_majority7_module_60__or_module_1_res), .ZN(
        n_majority7_module_60__or_module_6_res) );
  OR2_X1 u_majority7_module_60__or_module_7_U1 ( .A1(
        n_majority7_module_60__and_module_4_res), .A2(
        n_majority7_module_60__and_module_5_res), .ZN(
        n_majority7_module_60__or_module_7_res) );
  AND2_X1 u_majority7_module_60__and_module_7_U1 ( .A1(
        n_majority7_module_60__or_module_3_res), .A2(
        n_majority7_module_60__or_module_4_res), .ZN(
        n_majority7_module_60__and_module_7_res) );
  OR2_X1 u_majority7_module_60__or_module_8_U1 ( .A1(
        n_majority7_module_60__or_module_4_res), .A2(
        n_majority7_module_60__or_module_3_res), .ZN(
        n_majority7_module_60__or_module_8_res) );
  AND2_X1 u_majority7_module_60__and_module_8_U1 ( .A1(
        n_majority7_module_60__or_module_5_res), .A2(
        n_majority7_module_60__and_module_6_res), .ZN(
        n_majority7_module_60__and_module_8_res) );
  OR2_X1 u_majority7_module_60__or_module_9_U1 ( .A1(
        n_majority7_module_60__and_module_6_res), .A2(
        n_majority7_module_60__or_module_5_res), .ZN(
        n_majority7_module_60__or_module_9_res) );
  OR2_X1 u_majority7_module_60__or_module_10_U1 ( .A1(
        n_majority7_module_60__or_module_7_res), .A2(
        n_majority7_module_60__and_module_7_res), .ZN(
        n_majority7_module_60__or_module_10_res) );
  AND2_X1 u_majority7_module_60__and_module_9_U1 ( .A1(
        n_majority7_module_60__or_module_6_res), .A2(
        n_majority7_module_60__or_module_9_res), .ZN(
        n_majority7_module_60__and_module_9_res) );
  OR2_X1 u_majority7_module_60__or_module_11_U1 ( .A1(
        n_majority7_module_60__or_module_10_res), .A2(
        n_majority7_module_60__and_module_8_res), .ZN(
        n_majority7_module_60__or_module_11_res) );
  AND2_X1 u_majority7_module_60__and_module_10_U1 ( .A1(
        n_majority7_module_60__or_module_8_res), .A2(
        n_majority7_module_60__and_module_9_res), .ZN(
        n_majority7_module_60__and_module_10_res) );
  AND2_X1 u_majority7_module_60__and_module_11_U1 ( .A1(
        n_majority7_module_60__and_module_10_res), .A2(
        n_majority7_module_60__or_module_11_res), .ZN(
        n_majority7_module_60_res) );
  DFF_X1 u_reg_module_72__cini_mul_v00_reg ( .D(n_majority7_module_60_res), 
        .CK(clock_2), .Q(n_reg_module_72_res), .QN() );
  AND2_X1 u_majority7_module_61__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_61__and_module_1_res)
         );
  OR2_X1 u_majority7_module_61__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_61__or_module_1_res)
         );
  AND2_X1 u_majority7_module_61__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(n_majority7_module_61__and_module_2_res) );
  OR2_X1 u_majority7_module_61__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_61__or_module_2_res)
         );
  AND2_X1 u_majority7_module_61__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(n_majority7_module_61__and_module_3_res) );
  OR2_X1 u_majority7_module_61__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_61__or_module_3_res)
         );
  AND2_X1 u_majority7_module_61__and_module_4_U1 ( .A1(
        n_majority7_module_61__and_module_2_res), .A2(
        n_majority7_module_61__and_module_1_res), .ZN(
        n_majority7_module_61__and_module_4_res) );
  OR2_X1 u_majority7_module_61__or_module_4_U1 ( .A1(
        n_majority7_module_61__and_module_1_res), .A2(
        n_majority7_module_61__and_module_2_res), .ZN(
        n_majority7_module_61__or_module_4_res) );
  AND2_X1 u_majority7_module_61__and_module_5_U1 ( .A1(
        n_majority7_module_61__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_61__and_module_5_res) );
  OR2_X1 u_majority7_module_61__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_61__and_module_3_res), .ZN(
        n_majority7_module_61__or_module_5_res) );
  AND2_X1 u_majority7_module_61__and_module_6_U1 ( .A1(
        n_majority7_module_61__or_module_1_res), .A2(
        n_majority7_module_61__or_module_2_res), .ZN(
        n_majority7_module_61__and_module_6_res) );
  OR2_X1 u_majority7_module_61__or_module_6_U1 ( .A1(
        n_majority7_module_61__or_module_2_res), .A2(
        n_majority7_module_61__or_module_1_res), .ZN(
        n_majority7_module_61__or_module_6_res) );
  OR2_X1 u_majority7_module_61__or_module_7_U1 ( .A1(
        n_majority7_module_61__and_module_4_res), .A2(
        n_majority7_module_61__and_module_5_res), .ZN(
        n_majority7_module_61__or_module_7_res) );
  AND2_X1 u_majority7_module_61__and_module_7_U1 ( .A1(
        n_majority7_module_61__or_module_3_res), .A2(
        n_majority7_module_61__or_module_4_res), .ZN(
        n_majority7_module_61__and_module_7_res) );
  OR2_X1 u_majority7_module_61__or_module_8_U1 ( .A1(
        n_majority7_module_61__or_module_4_res), .A2(
        n_majority7_module_61__or_module_3_res), .ZN(
        n_majority7_module_61__or_module_8_res) );
  AND2_X1 u_majority7_module_61__and_module_8_U1 ( .A1(
        n_majority7_module_61__or_module_5_res), .A2(
        n_majority7_module_61__and_module_6_res), .ZN(
        n_majority7_module_61__and_module_8_res) );
  OR2_X1 u_majority7_module_61__or_module_9_U1 ( .A1(
        n_majority7_module_61__and_module_6_res), .A2(
        n_majority7_module_61__or_module_5_res), .ZN(
        n_majority7_module_61__or_module_9_res) );
  OR2_X1 u_majority7_module_61__or_module_10_U1 ( .A1(
        n_majority7_module_61__or_module_7_res), .A2(
        n_majority7_module_61__and_module_7_res), .ZN(
        n_majority7_module_61__or_module_10_res) );
  AND2_X1 u_majority7_module_61__and_module_9_U1 ( .A1(
        n_majority7_module_61__or_module_6_res), .A2(
        n_majority7_module_61__or_module_9_res), .ZN(
        n_majority7_module_61__and_module_9_res) );
  OR2_X1 u_majority7_module_61__or_module_11_U1 ( .A1(
        n_majority7_module_61__or_module_10_res), .A2(
        n_majority7_module_61__and_module_8_res), .ZN(
        n_majority7_module_61__or_module_11_res) );
  AND2_X1 u_majority7_module_61__and_module_10_U1 ( .A1(
        n_majority7_module_61__or_module_8_res), .A2(
        n_majority7_module_61__and_module_9_res), .ZN(
        n_majority7_module_61__and_module_10_res) );
  AND2_X1 u_majority7_module_61__and_module_11_U1 ( .A1(
        n_majority7_module_61__and_module_10_res), .A2(
        n_majority7_module_61__or_module_11_res), .ZN(
        n_majority7_module_61_res) );
  DFF_X1 u_reg_module_73__cini_mul_v00_reg ( .D(n_majority7_module_61_res), 
        .CK(clock_2), .Q(n_reg_module_73_res), .QN() );
  AND2_X1 u_majority7_module_62__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_62__and_module_1_res)
         );
  OR2_X1 u_majority7_module_62__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_62__or_module_1_res)
         );
  AND2_X1 u_majority7_module_62__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(n_majority7_module_62__and_module_2_res) );
  OR2_X1 u_majority7_module_62__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_62__or_module_2_res)
         );
  AND2_X1 u_majority7_module_62__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(n_majority7_module_62__and_module_3_res) );
  OR2_X1 u_majority7_module_62__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_62__or_module_3_res)
         );
  AND2_X1 u_majority7_module_62__and_module_4_U1 ( .A1(
        n_majority7_module_62__and_module_2_res), .A2(
        n_majority7_module_62__and_module_1_res), .ZN(
        n_majority7_module_62__and_module_4_res) );
  OR2_X1 u_majority7_module_62__or_module_4_U1 ( .A1(
        n_majority7_module_62__and_module_1_res), .A2(
        n_majority7_module_62__and_module_2_res), .ZN(
        n_majority7_module_62__or_module_4_res) );
  AND2_X1 u_majority7_module_62__and_module_5_U1 ( .A1(
        n_majority7_module_62__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_62__and_module_5_res) );
  OR2_X1 u_majority7_module_62__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_62__and_module_3_res), .ZN(
        n_majority7_module_62__or_module_5_res) );
  AND2_X1 u_majority7_module_62__and_module_6_U1 ( .A1(
        n_majority7_module_62__or_module_1_res), .A2(
        n_majority7_module_62__or_module_2_res), .ZN(
        n_majority7_module_62__and_module_6_res) );
  OR2_X1 u_majority7_module_62__or_module_6_U1 ( .A1(
        n_majority7_module_62__or_module_2_res), .A2(
        n_majority7_module_62__or_module_1_res), .ZN(
        n_majority7_module_62__or_module_6_res) );
  OR2_X1 u_majority7_module_62__or_module_7_U1 ( .A1(
        n_majority7_module_62__and_module_4_res), .A2(
        n_majority7_module_62__and_module_5_res), .ZN(
        n_majority7_module_62__or_module_7_res) );
  AND2_X1 u_majority7_module_62__and_module_7_U1 ( .A1(
        n_majority7_module_62__or_module_3_res), .A2(
        n_majority7_module_62__or_module_4_res), .ZN(
        n_majority7_module_62__and_module_7_res) );
  OR2_X1 u_majority7_module_62__or_module_8_U1 ( .A1(
        n_majority7_module_62__or_module_4_res), .A2(
        n_majority7_module_62__or_module_3_res), .ZN(
        n_majority7_module_62__or_module_8_res) );
  AND2_X1 u_majority7_module_62__and_module_8_U1 ( .A1(
        n_majority7_module_62__or_module_5_res), .A2(
        n_majority7_module_62__and_module_6_res), .ZN(
        n_majority7_module_62__and_module_8_res) );
  OR2_X1 u_majority7_module_62__or_module_9_U1 ( .A1(
        n_majority7_module_62__and_module_6_res), .A2(
        n_majority7_module_62__or_module_5_res), .ZN(
        n_majority7_module_62__or_module_9_res) );
  OR2_X1 u_majority7_module_62__or_module_10_U1 ( .A1(
        n_majority7_module_62__or_module_7_res), .A2(
        n_majority7_module_62__and_module_7_res), .ZN(
        n_majority7_module_62__or_module_10_res) );
  AND2_X1 u_majority7_module_62__and_module_9_U1 ( .A1(
        n_majority7_module_62__or_module_6_res), .A2(
        n_majority7_module_62__or_module_9_res), .ZN(
        n_majority7_module_62__and_module_9_res) );
  OR2_X1 u_majority7_module_62__or_module_11_U1 ( .A1(
        n_majority7_module_62__or_module_10_res), .A2(
        n_majority7_module_62__and_module_8_res), .ZN(
        n_majority7_module_62__or_module_11_res) );
  AND2_X1 u_majority7_module_62__and_module_10_U1 ( .A1(
        n_majority7_module_62__or_module_8_res), .A2(
        n_majority7_module_62__and_module_9_res), .ZN(
        n_majority7_module_62__and_module_10_res) );
  AND2_X1 u_majority7_module_62__and_module_11_U1 ( .A1(
        n_majority7_module_62__and_module_10_res), .A2(
        n_majority7_module_62__or_module_11_res), .ZN(
        n_majority7_module_62_res) );
  DFF_X1 u_reg_module_74__cini_mul_v00_reg ( .D(n_majority7_module_62_res), 
        .CK(clock_2), .Q(n_reg_module_74_res), .QN() );
  AND2_X1 u_majority7_module_63__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_63__and_module_1_res)
         );
  OR2_X1 u_majority7_module_63__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_63__or_module_1_res)
         );
  AND2_X1 u_majority7_module_63__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(n_majority7_module_63__and_module_2_res) );
  OR2_X1 u_majority7_module_63__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_63__or_module_2_res)
         );
  AND2_X1 u_majority7_module_63__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(n_majority7_module_63__and_module_3_res) );
  OR2_X1 u_majority7_module_63__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_63__or_module_3_res)
         );
  AND2_X1 u_majority7_module_63__and_module_4_U1 ( .A1(
        n_majority7_module_63__and_module_2_res), .A2(
        n_majority7_module_63__and_module_1_res), .ZN(
        n_majority7_module_63__and_module_4_res) );
  OR2_X1 u_majority7_module_63__or_module_4_U1 ( .A1(
        n_majority7_module_63__and_module_1_res), .A2(
        n_majority7_module_63__and_module_2_res), .ZN(
        n_majority7_module_63__or_module_4_res) );
  AND2_X1 u_majority7_module_63__and_module_5_U1 ( .A1(
        n_majority7_module_63__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_63__and_module_5_res) );
  OR2_X1 u_majority7_module_63__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_63__and_module_3_res), .ZN(
        n_majority7_module_63__or_module_5_res) );
  AND2_X1 u_majority7_module_63__and_module_6_U1 ( .A1(
        n_majority7_module_63__or_module_1_res), .A2(
        n_majority7_module_63__or_module_2_res), .ZN(
        n_majority7_module_63__and_module_6_res) );
  OR2_X1 u_majority7_module_63__or_module_6_U1 ( .A1(
        n_majority7_module_63__or_module_2_res), .A2(
        n_majority7_module_63__or_module_1_res), .ZN(
        n_majority7_module_63__or_module_6_res) );
  OR2_X1 u_majority7_module_63__or_module_7_U1 ( .A1(
        n_majority7_module_63__and_module_4_res), .A2(
        n_majority7_module_63__and_module_5_res), .ZN(
        n_majority7_module_63__or_module_7_res) );
  AND2_X1 u_majority7_module_63__and_module_7_U1 ( .A1(
        n_majority7_module_63__or_module_3_res), .A2(
        n_majority7_module_63__or_module_4_res), .ZN(
        n_majority7_module_63__and_module_7_res) );
  OR2_X1 u_majority7_module_63__or_module_8_U1 ( .A1(
        n_majority7_module_63__or_module_4_res), .A2(
        n_majority7_module_63__or_module_3_res), .ZN(
        n_majority7_module_63__or_module_8_res) );
  AND2_X1 u_majority7_module_63__and_module_8_U1 ( .A1(
        n_majority7_module_63__or_module_5_res), .A2(
        n_majority7_module_63__and_module_6_res), .ZN(
        n_majority7_module_63__and_module_8_res) );
  OR2_X1 u_majority7_module_63__or_module_9_U1 ( .A1(
        n_majority7_module_63__and_module_6_res), .A2(
        n_majority7_module_63__or_module_5_res), .ZN(
        n_majority7_module_63__or_module_9_res) );
  OR2_X1 u_majority7_module_63__or_module_10_U1 ( .A1(
        n_majority7_module_63__or_module_7_res), .A2(
        n_majority7_module_63__and_module_7_res), .ZN(
        n_majority7_module_63__or_module_10_res) );
  AND2_X1 u_majority7_module_63__and_module_9_U1 ( .A1(
        n_majority7_module_63__or_module_6_res), .A2(
        n_majority7_module_63__or_module_9_res), .ZN(
        n_majority7_module_63__and_module_9_res) );
  OR2_X1 u_majority7_module_63__or_module_11_U1 ( .A1(
        n_majority7_module_63__or_module_10_res), .A2(
        n_majority7_module_63__and_module_8_res), .ZN(
        n_majority7_module_63__or_module_11_res) );
  AND2_X1 u_majority7_module_63__and_module_10_U1 ( .A1(
        n_majority7_module_63__or_module_8_res), .A2(
        n_majority7_module_63__and_module_9_res), .ZN(
        n_majority7_module_63__and_module_10_res) );
  AND2_X1 u_majority7_module_63__and_module_11_U1 ( .A1(
        n_majority7_module_63__and_module_10_res), .A2(
        n_majority7_module_63__or_module_11_res), .ZN(
        n_majority7_module_63_res) );
  DFF_X1 u_reg_module_75__cini_mul_v00_reg ( .D(n_majority7_module_63_res), 
        .CK(clock_2), .Q(n_reg_module_75_res), .QN() );
  DFF_X1 u_reg_module_76__cini_mul_v00_reg ( .D(n_and_module_48_res), .CK(
        clock_2), .Q(n_reg_module_76_res), .QN() );
  DFF_X1 u_reg_module_77__cini_mul_v00_reg ( .D(n_and_module_49_res), .CK(
        clock_3), .Q(n_reg_module_77_res), .QN() );
  AND2_X1 u_majority7_module_64__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_64__and_module_1_res)
         );
  OR2_X1 u_majority7_module_64__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_64__or_module_1_res)
         );
  AND2_X1 u_majority7_module_64__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(n_majority7_module_64__and_module_2_res) );
  OR2_X1 u_majority7_module_64__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_64__or_module_2_res)
         );
  AND2_X1 u_majority7_module_64__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(n_majority7_module_64__and_module_3_res) );
  OR2_X1 u_majority7_module_64__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_64__or_module_3_res)
         );
  AND2_X1 u_majority7_module_64__and_module_4_U1 ( .A1(
        n_majority7_module_64__and_module_2_res), .A2(
        n_majority7_module_64__and_module_1_res), .ZN(
        n_majority7_module_64__and_module_4_res) );
  OR2_X1 u_majority7_module_64__or_module_4_U1 ( .A1(
        n_majority7_module_64__and_module_1_res), .A2(
        n_majority7_module_64__and_module_2_res), .ZN(
        n_majority7_module_64__or_module_4_res) );
  AND2_X1 u_majority7_module_64__and_module_5_U1 ( .A1(
        n_majority7_module_64__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_64__and_module_5_res) );
  OR2_X1 u_majority7_module_64__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_64__and_module_3_res), .ZN(
        n_majority7_module_64__or_module_5_res) );
  AND2_X1 u_majority7_module_64__and_module_6_U1 ( .A1(
        n_majority7_module_64__or_module_1_res), .A2(
        n_majority7_module_64__or_module_2_res), .ZN(
        n_majority7_module_64__and_module_6_res) );
  OR2_X1 u_majority7_module_64__or_module_6_U1 ( .A1(
        n_majority7_module_64__or_module_2_res), .A2(
        n_majority7_module_64__or_module_1_res), .ZN(
        n_majority7_module_64__or_module_6_res) );
  OR2_X1 u_majority7_module_64__or_module_7_U1 ( .A1(
        n_majority7_module_64__and_module_4_res), .A2(
        n_majority7_module_64__and_module_5_res), .ZN(
        n_majority7_module_64__or_module_7_res) );
  AND2_X1 u_majority7_module_64__and_module_7_U1 ( .A1(
        n_majority7_module_64__or_module_3_res), .A2(
        n_majority7_module_64__or_module_4_res), .ZN(
        n_majority7_module_64__and_module_7_res) );
  OR2_X1 u_majority7_module_64__or_module_8_U1 ( .A1(
        n_majority7_module_64__or_module_4_res), .A2(
        n_majority7_module_64__or_module_3_res), .ZN(
        n_majority7_module_64__or_module_8_res) );
  AND2_X1 u_majority7_module_64__and_module_8_U1 ( .A1(
        n_majority7_module_64__or_module_5_res), .A2(
        n_majority7_module_64__and_module_6_res), .ZN(
        n_majority7_module_64__and_module_8_res) );
  OR2_X1 u_majority7_module_64__or_module_9_U1 ( .A1(
        n_majority7_module_64__and_module_6_res), .A2(
        n_majority7_module_64__or_module_5_res), .ZN(
        n_majority7_module_64__or_module_9_res) );
  OR2_X1 u_majority7_module_64__or_module_10_U1 ( .A1(
        n_majority7_module_64__or_module_7_res), .A2(
        n_majority7_module_64__and_module_7_res), .ZN(
        n_majority7_module_64__or_module_10_res) );
  AND2_X1 u_majority7_module_64__and_module_9_U1 ( .A1(
        n_majority7_module_64__or_module_6_res), .A2(
        n_majority7_module_64__or_module_9_res), .ZN(
        n_majority7_module_64__and_module_9_res) );
  OR2_X1 u_majority7_module_64__or_module_11_U1 ( .A1(
        n_majority7_module_64__or_module_10_res), .A2(
        n_majority7_module_64__and_module_8_res), .ZN(
        n_majority7_module_64__or_module_11_res) );
  AND2_X1 u_majority7_module_64__and_module_10_U1 ( .A1(
        n_majority7_module_64__or_module_8_res), .A2(
        n_majority7_module_64__and_module_9_res), .ZN(
        n_majority7_module_64__and_module_10_res) );
  AND2_X1 u_majority7_module_64__and_module_11_U1 ( .A1(
        n_majority7_module_64__and_module_10_res), .A2(
        n_majority7_module_64__or_module_11_res), .ZN(
        n_majority7_module_64_res) );
  DFF_X1 u_reg_module_78__cini_mul_v00_reg ( .D(n_majority7_module_64_res), 
        .CK(clock_3), .Q(n_reg_module_78_res), .QN() );
  AND2_X1 u_majority7_module_65__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_65__and_module_1_res)
         );
  OR2_X1 u_majority7_module_65__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_65__or_module_1_res)
         );
  AND2_X1 u_majority7_module_65__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(n_majority7_module_65__and_module_2_res) );
  OR2_X1 u_majority7_module_65__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_65__or_module_2_res)
         );
  AND2_X1 u_majority7_module_65__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(n_majority7_module_65__and_module_3_res) );
  OR2_X1 u_majority7_module_65__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_65__or_module_3_res)
         );
  AND2_X1 u_majority7_module_65__and_module_4_U1 ( .A1(
        n_majority7_module_65__and_module_2_res), .A2(
        n_majority7_module_65__and_module_1_res), .ZN(
        n_majority7_module_65__and_module_4_res) );
  OR2_X1 u_majority7_module_65__or_module_4_U1 ( .A1(
        n_majority7_module_65__and_module_1_res), .A2(
        n_majority7_module_65__and_module_2_res), .ZN(
        n_majority7_module_65__or_module_4_res) );
  AND2_X1 u_majority7_module_65__and_module_5_U1 ( .A1(
        n_majority7_module_65__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_65__and_module_5_res) );
  OR2_X1 u_majority7_module_65__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_65__and_module_3_res), .ZN(
        n_majority7_module_65__or_module_5_res) );
  AND2_X1 u_majority7_module_65__and_module_6_U1 ( .A1(
        n_majority7_module_65__or_module_1_res), .A2(
        n_majority7_module_65__or_module_2_res), .ZN(
        n_majority7_module_65__and_module_6_res) );
  OR2_X1 u_majority7_module_65__or_module_6_U1 ( .A1(
        n_majority7_module_65__or_module_2_res), .A2(
        n_majority7_module_65__or_module_1_res), .ZN(
        n_majority7_module_65__or_module_6_res) );
  OR2_X1 u_majority7_module_65__or_module_7_U1 ( .A1(
        n_majority7_module_65__and_module_4_res), .A2(
        n_majority7_module_65__and_module_5_res), .ZN(
        n_majority7_module_65__or_module_7_res) );
  AND2_X1 u_majority7_module_65__and_module_7_U1 ( .A1(
        n_majority7_module_65__or_module_3_res), .A2(
        n_majority7_module_65__or_module_4_res), .ZN(
        n_majority7_module_65__and_module_7_res) );
  OR2_X1 u_majority7_module_65__or_module_8_U1 ( .A1(
        n_majority7_module_65__or_module_4_res), .A2(
        n_majority7_module_65__or_module_3_res), .ZN(
        n_majority7_module_65__or_module_8_res) );
  AND2_X1 u_majority7_module_65__and_module_8_U1 ( .A1(
        n_majority7_module_65__or_module_5_res), .A2(
        n_majority7_module_65__and_module_6_res), .ZN(
        n_majority7_module_65__and_module_8_res) );
  OR2_X1 u_majority7_module_65__or_module_9_U1 ( .A1(
        n_majority7_module_65__and_module_6_res), .A2(
        n_majority7_module_65__or_module_5_res), .ZN(
        n_majority7_module_65__or_module_9_res) );
  OR2_X1 u_majority7_module_65__or_module_10_U1 ( .A1(
        n_majority7_module_65__or_module_7_res), .A2(
        n_majority7_module_65__and_module_7_res), .ZN(
        n_majority7_module_65__or_module_10_res) );
  AND2_X1 u_majority7_module_65__and_module_9_U1 ( .A1(
        n_majority7_module_65__or_module_6_res), .A2(
        n_majority7_module_65__or_module_9_res), .ZN(
        n_majority7_module_65__and_module_9_res) );
  OR2_X1 u_majority7_module_65__or_module_11_U1 ( .A1(
        n_majority7_module_65__or_module_10_res), .A2(
        n_majority7_module_65__and_module_8_res), .ZN(
        n_majority7_module_65__or_module_11_res) );
  AND2_X1 u_majority7_module_65__and_module_10_U1 ( .A1(
        n_majority7_module_65__or_module_8_res), .A2(
        n_majority7_module_65__and_module_9_res), .ZN(
        n_majority7_module_65__and_module_10_res) );
  AND2_X1 u_majority7_module_65__and_module_11_U1 ( .A1(
        n_majority7_module_65__and_module_10_res), .A2(
        n_majority7_module_65__or_module_11_res), .ZN(
        n_majority7_module_65_res) );
  DFF_X1 u_reg_module_79__cini_mul_v00_reg ( .D(n_majority7_module_65_res), 
        .CK(clock_3), .Q(n_reg_module_79_res), .QN() );
  AND2_X1 u_majority7_module_66__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_66__and_module_1_res)
         );
  OR2_X1 u_majority7_module_66__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_66__or_module_1_res)
         );
  AND2_X1 u_majority7_module_66__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(n_majority7_module_66__and_module_2_res) );
  OR2_X1 u_majority7_module_66__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_66__or_module_2_res)
         );
  AND2_X1 u_majority7_module_66__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(n_majority7_module_66__and_module_3_res) );
  OR2_X1 u_majority7_module_66__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_66__or_module_3_res)
         );
  AND2_X1 u_majority7_module_66__and_module_4_U1 ( .A1(
        n_majority7_module_66__and_module_2_res), .A2(
        n_majority7_module_66__and_module_1_res), .ZN(
        n_majority7_module_66__and_module_4_res) );
  OR2_X1 u_majority7_module_66__or_module_4_U1 ( .A1(
        n_majority7_module_66__and_module_1_res), .A2(
        n_majority7_module_66__and_module_2_res), .ZN(
        n_majority7_module_66__or_module_4_res) );
  AND2_X1 u_majority7_module_66__and_module_5_U1 ( .A1(
        n_majority7_module_66__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_66__and_module_5_res) );
  OR2_X1 u_majority7_module_66__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_66__and_module_3_res), .ZN(
        n_majority7_module_66__or_module_5_res) );
  AND2_X1 u_majority7_module_66__and_module_6_U1 ( .A1(
        n_majority7_module_66__or_module_1_res), .A2(
        n_majority7_module_66__or_module_2_res), .ZN(
        n_majority7_module_66__and_module_6_res) );
  OR2_X1 u_majority7_module_66__or_module_6_U1 ( .A1(
        n_majority7_module_66__or_module_2_res), .A2(
        n_majority7_module_66__or_module_1_res), .ZN(
        n_majority7_module_66__or_module_6_res) );
  OR2_X1 u_majority7_module_66__or_module_7_U1 ( .A1(
        n_majority7_module_66__and_module_4_res), .A2(
        n_majority7_module_66__and_module_5_res), .ZN(
        n_majority7_module_66__or_module_7_res) );
  AND2_X1 u_majority7_module_66__and_module_7_U1 ( .A1(
        n_majority7_module_66__or_module_3_res), .A2(
        n_majority7_module_66__or_module_4_res), .ZN(
        n_majority7_module_66__and_module_7_res) );
  OR2_X1 u_majority7_module_66__or_module_8_U1 ( .A1(
        n_majority7_module_66__or_module_4_res), .A2(
        n_majority7_module_66__or_module_3_res), .ZN(
        n_majority7_module_66__or_module_8_res) );
  AND2_X1 u_majority7_module_66__and_module_8_U1 ( .A1(
        n_majority7_module_66__or_module_5_res), .A2(
        n_majority7_module_66__and_module_6_res), .ZN(
        n_majority7_module_66__and_module_8_res) );
  OR2_X1 u_majority7_module_66__or_module_9_U1 ( .A1(
        n_majority7_module_66__and_module_6_res), .A2(
        n_majority7_module_66__or_module_5_res), .ZN(
        n_majority7_module_66__or_module_9_res) );
  OR2_X1 u_majority7_module_66__or_module_10_U1 ( .A1(
        n_majority7_module_66__or_module_7_res), .A2(
        n_majority7_module_66__and_module_7_res), .ZN(
        n_majority7_module_66__or_module_10_res) );
  AND2_X1 u_majority7_module_66__and_module_9_U1 ( .A1(
        n_majority7_module_66__or_module_6_res), .A2(
        n_majority7_module_66__or_module_9_res), .ZN(
        n_majority7_module_66__and_module_9_res) );
  OR2_X1 u_majority7_module_66__or_module_11_U1 ( .A1(
        n_majority7_module_66__or_module_10_res), .A2(
        n_majority7_module_66__and_module_8_res), .ZN(
        n_majority7_module_66__or_module_11_res) );
  AND2_X1 u_majority7_module_66__and_module_10_U1 ( .A1(
        n_majority7_module_66__or_module_8_res), .A2(
        n_majority7_module_66__and_module_9_res), .ZN(
        n_majority7_module_66__and_module_10_res) );
  AND2_X1 u_majority7_module_66__and_module_11_U1 ( .A1(
        n_majority7_module_66__and_module_10_res), .A2(
        n_majority7_module_66__or_module_11_res), .ZN(
        n_majority7_module_66_res) );
  DFF_X1 u_reg_module_80__cini_mul_v00_reg ( .D(n_majority7_module_66_res), 
        .CK(clock_3), .Q(n_reg_module_80_res), .QN() );
  AND2_X1 u_majority7_module_67__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_67__and_module_1_res)
         );
  OR2_X1 u_majority7_module_67__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_67__or_module_1_res)
         );
  AND2_X1 u_majority7_module_67__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(n_majority7_module_67__and_module_2_res) );
  OR2_X1 u_majority7_module_67__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_67__or_module_2_res)
         );
  AND2_X1 u_majority7_module_67__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(n_majority7_module_67__and_module_3_res) );
  OR2_X1 u_majority7_module_67__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_67__or_module_3_res)
         );
  AND2_X1 u_majority7_module_67__and_module_4_U1 ( .A1(
        n_majority7_module_67__and_module_2_res), .A2(
        n_majority7_module_67__and_module_1_res), .ZN(
        n_majority7_module_67__and_module_4_res) );
  OR2_X1 u_majority7_module_67__or_module_4_U1 ( .A1(
        n_majority7_module_67__and_module_1_res), .A2(
        n_majority7_module_67__and_module_2_res), .ZN(
        n_majority7_module_67__or_module_4_res) );
  AND2_X1 u_majority7_module_67__and_module_5_U1 ( .A1(
        n_majority7_module_67__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_67__and_module_5_res) );
  OR2_X1 u_majority7_module_67__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_67__and_module_3_res), .ZN(
        n_majority7_module_67__or_module_5_res) );
  AND2_X1 u_majority7_module_67__and_module_6_U1 ( .A1(
        n_majority7_module_67__or_module_1_res), .A2(
        n_majority7_module_67__or_module_2_res), .ZN(
        n_majority7_module_67__and_module_6_res) );
  OR2_X1 u_majority7_module_67__or_module_6_U1 ( .A1(
        n_majority7_module_67__or_module_2_res), .A2(
        n_majority7_module_67__or_module_1_res), .ZN(
        n_majority7_module_67__or_module_6_res) );
  OR2_X1 u_majority7_module_67__or_module_7_U1 ( .A1(
        n_majority7_module_67__and_module_4_res), .A2(
        n_majority7_module_67__and_module_5_res), .ZN(
        n_majority7_module_67__or_module_7_res) );
  AND2_X1 u_majority7_module_67__and_module_7_U1 ( .A1(
        n_majority7_module_67__or_module_3_res), .A2(
        n_majority7_module_67__or_module_4_res), .ZN(
        n_majority7_module_67__and_module_7_res) );
  OR2_X1 u_majority7_module_67__or_module_8_U1 ( .A1(
        n_majority7_module_67__or_module_4_res), .A2(
        n_majority7_module_67__or_module_3_res), .ZN(
        n_majority7_module_67__or_module_8_res) );
  AND2_X1 u_majority7_module_67__and_module_8_U1 ( .A1(
        n_majority7_module_67__or_module_5_res), .A2(
        n_majority7_module_67__and_module_6_res), .ZN(
        n_majority7_module_67__and_module_8_res) );
  OR2_X1 u_majority7_module_67__or_module_9_U1 ( .A1(
        n_majority7_module_67__and_module_6_res), .A2(
        n_majority7_module_67__or_module_5_res), .ZN(
        n_majority7_module_67__or_module_9_res) );
  OR2_X1 u_majority7_module_67__or_module_10_U1 ( .A1(
        n_majority7_module_67__or_module_7_res), .A2(
        n_majority7_module_67__and_module_7_res), .ZN(
        n_majority7_module_67__or_module_10_res) );
  AND2_X1 u_majority7_module_67__and_module_9_U1 ( .A1(
        n_majority7_module_67__or_module_6_res), .A2(
        n_majority7_module_67__or_module_9_res), .ZN(
        n_majority7_module_67__and_module_9_res) );
  OR2_X1 u_majority7_module_67__or_module_11_U1 ( .A1(
        n_majority7_module_67__or_module_10_res), .A2(
        n_majority7_module_67__and_module_8_res), .ZN(
        n_majority7_module_67__or_module_11_res) );
  AND2_X1 u_majority7_module_67__and_module_10_U1 ( .A1(
        n_majority7_module_67__or_module_8_res), .A2(
        n_majority7_module_67__and_module_9_res), .ZN(
        n_majority7_module_67__and_module_10_res) );
  AND2_X1 u_majority7_module_67__and_module_11_U1 ( .A1(
        n_majority7_module_67__and_module_10_res), .A2(
        n_majority7_module_67__or_module_11_res), .ZN(
        n_majority7_module_67_res) );
  DFF_X1 u_reg_module_81__cini_mul_v00_reg ( .D(n_majority7_module_67_res), 
        .CK(clock_3), .Q(n_reg_module_81_res), .QN() );
  DFF_X1 u_reg_module_82__cini_mul_v00_reg ( .D(n_and_module_54_res), .CK(
        clock_3), .Q(n_reg_module_82_res), .QN() );
  AND2_X1 u_majority7_module_68__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_68__and_module_1_res)
         );
  OR2_X1 u_majority7_module_68__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_68__or_module_1_res)
         );
  AND2_X1 u_majority7_module_68__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(n_majority7_module_68__and_module_2_res) );
  OR2_X1 u_majority7_module_68__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_68__or_module_2_res)
         );
  AND2_X1 u_majority7_module_68__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(n_majority7_module_68__and_module_3_res) );
  OR2_X1 u_majority7_module_68__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_68__or_module_3_res)
         );
  AND2_X1 u_majority7_module_68__and_module_4_U1 ( .A1(
        n_majority7_module_68__and_module_2_res), .A2(
        n_majority7_module_68__and_module_1_res), .ZN(
        n_majority7_module_68__and_module_4_res) );
  OR2_X1 u_majority7_module_68__or_module_4_U1 ( .A1(
        n_majority7_module_68__and_module_1_res), .A2(
        n_majority7_module_68__and_module_2_res), .ZN(
        n_majority7_module_68__or_module_4_res) );
  AND2_X1 u_majority7_module_68__and_module_5_U1 ( .A1(
        n_majority7_module_68__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_68__and_module_5_res) );
  OR2_X1 u_majority7_module_68__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_68__and_module_3_res), .ZN(
        n_majority7_module_68__or_module_5_res) );
  AND2_X1 u_majority7_module_68__and_module_6_U1 ( .A1(
        n_majority7_module_68__or_module_1_res), .A2(
        n_majority7_module_68__or_module_2_res), .ZN(
        n_majority7_module_68__and_module_6_res) );
  OR2_X1 u_majority7_module_68__or_module_6_U1 ( .A1(
        n_majority7_module_68__or_module_2_res), .A2(
        n_majority7_module_68__or_module_1_res), .ZN(
        n_majority7_module_68__or_module_6_res) );
  OR2_X1 u_majority7_module_68__or_module_7_U1 ( .A1(
        n_majority7_module_68__and_module_4_res), .A2(
        n_majority7_module_68__and_module_5_res), .ZN(
        n_majority7_module_68__or_module_7_res) );
  AND2_X1 u_majority7_module_68__and_module_7_U1 ( .A1(
        n_majority7_module_68__or_module_3_res), .A2(
        n_majority7_module_68__or_module_4_res), .ZN(
        n_majority7_module_68__and_module_7_res) );
  OR2_X1 u_majority7_module_68__or_module_8_U1 ( .A1(
        n_majority7_module_68__or_module_4_res), .A2(
        n_majority7_module_68__or_module_3_res), .ZN(
        n_majority7_module_68__or_module_8_res) );
  AND2_X1 u_majority7_module_68__and_module_8_U1 ( .A1(
        n_majority7_module_68__or_module_5_res), .A2(
        n_majority7_module_68__and_module_6_res), .ZN(
        n_majority7_module_68__and_module_8_res) );
  OR2_X1 u_majority7_module_68__or_module_9_U1 ( .A1(
        n_majority7_module_68__and_module_6_res), .A2(
        n_majority7_module_68__or_module_5_res), .ZN(
        n_majority7_module_68__or_module_9_res) );
  OR2_X1 u_majority7_module_68__or_module_10_U1 ( .A1(
        n_majority7_module_68__or_module_7_res), .A2(
        n_majority7_module_68__and_module_7_res), .ZN(
        n_majority7_module_68__or_module_10_res) );
  AND2_X1 u_majority7_module_68__and_module_9_U1 ( .A1(
        n_majority7_module_68__or_module_6_res), .A2(
        n_majority7_module_68__or_module_9_res), .ZN(
        n_majority7_module_68__and_module_9_res) );
  OR2_X1 u_majority7_module_68__or_module_11_U1 ( .A1(
        n_majority7_module_68__or_module_10_res), .A2(
        n_majority7_module_68__and_module_8_res), .ZN(
        n_majority7_module_68__or_module_11_res) );
  AND2_X1 u_majority7_module_68__and_module_10_U1 ( .A1(
        n_majority7_module_68__or_module_8_res), .A2(
        n_majority7_module_68__and_module_9_res), .ZN(
        n_majority7_module_68__and_module_10_res) );
  AND2_X1 u_majority7_module_68__and_module_11_U1 ( .A1(
        n_majority7_module_68__and_module_10_res), .A2(
        n_majority7_module_68__or_module_11_res), .ZN(
        n_majority7_module_68_res) );
  DFF_X1 u_reg_module_83__cini_mul_v00_reg ( .D(n_majority7_module_68_res), 
        .CK(clock_3), .Q(n_reg_module_83_res), .QN() );
  AND2_X1 u_majority7_module_69__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_69__and_module_1_res)
         );
  OR2_X1 u_majority7_module_69__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_69__or_module_1_res)
         );
  AND2_X1 u_majority7_module_69__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(n_majority7_module_69__and_module_2_res) );
  OR2_X1 u_majority7_module_69__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_69__or_module_2_res)
         );
  AND2_X1 u_majority7_module_69__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(n_majority7_module_69__and_module_3_res) );
  OR2_X1 u_majority7_module_69__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_69__or_module_3_res)
         );
  AND2_X1 u_majority7_module_69__and_module_4_U1 ( .A1(
        n_majority7_module_69__and_module_2_res), .A2(
        n_majority7_module_69__and_module_1_res), .ZN(
        n_majority7_module_69__and_module_4_res) );
  OR2_X1 u_majority7_module_69__or_module_4_U1 ( .A1(
        n_majority7_module_69__and_module_1_res), .A2(
        n_majority7_module_69__and_module_2_res), .ZN(
        n_majority7_module_69__or_module_4_res) );
  AND2_X1 u_majority7_module_69__and_module_5_U1 ( .A1(
        n_majority7_module_69__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_69__and_module_5_res) );
  OR2_X1 u_majority7_module_69__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_69__and_module_3_res), .ZN(
        n_majority7_module_69__or_module_5_res) );
  AND2_X1 u_majority7_module_69__and_module_6_U1 ( .A1(
        n_majority7_module_69__or_module_1_res), .A2(
        n_majority7_module_69__or_module_2_res), .ZN(
        n_majority7_module_69__and_module_6_res) );
  OR2_X1 u_majority7_module_69__or_module_6_U1 ( .A1(
        n_majority7_module_69__or_module_2_res), .A2(
        n_majority7_module_69__or_module_1_res), .ZN(
        n_majority7_module_69__or_module_6_res) );
  OR2_X1 u_majority7_module_69__or_module_7_U1 ( .A1(
        n_majority7_module_69__and_module_4_res), .A2(
        n_majority7_module_69__and_module_5_res), .ZN(
        n_majority7_module_69__or_module_7_res) );
  AND2_X1 u_majority7_module_69__and_module_7_U1 ( .A1(
        n_majority7_module_69__or_module_3_res), .A2(
        n_majority7_module_69__or_module_4_res), .ZN(
        n_majority7_module_69__and_module_7_res) );
  OR2_X1 u_majority7_module_69__or_module_8_U1 ( .A1(
        n_majority7_module_69__or_module_4_res), .A2(
        n_majority7_module_69__or_module_3_res), .ZN(
        n_majority7_module_69__or_module_8_res) );
  AND2_X1 u_majority7_module_69__and_module_8_U1 ( .A1(
        n_majority7_module_69__or_module_5_res), .A2(
        n_majority7_module_69__and_module_6_res), .ZN(
        n_majority7_module_69__and_module_8_res) );
  OR2_X1 u_majority7_module_69__or_module_9_U1 ( .A1(
        n_majority7_module_69__and_module_6_res), .A2(
        n_majority7_module_69__or_module_5_res), .ZN(
        n_majority7_module_69__or_module_9_res) );
  OR2_X1 u_majority7_module_69__or_module_10_U1 ( .A1(
        n_majority7_module_69__or_module_7_res), .A2(
        n_majority7_module_69__and_module_7_res), .ZN(
        n_majority7_module_69__or_module_10_res) );
  AND2_X1 u_majority7_module_69__and_module_9_U1 ( .A1(
        n_majority7_module_69__or_module_6_res), .A2(
        n_majority7_module_69__or_module_9_res), .ZN(
        n_majority7_module_69__and_module_9_res) );
  OR2_X1 u_majority7_module_69__or_module_11_U1 ( .A1(
        n_majority7_module_69__or_module_10_res), .A2(
        n_majority7_module_69__and_module_8_res), .ZN(
        n_majority7_module_69__or_module_11_res) );
  AND2_X1 u_majority7_module_69__and_module_10_U1 ( .A1(
        n_majority7_module_69__or_module_8_res), .A2(
        n_majority7_module_69__and_module_9_res), .ZN(
        n_majority7_module_69__and_module_10_res) );
  AND2_X1 u_majority7_module_69__and_module_11_U1 ( .A1(
        n_majority7_module_69__and_module_10_res), .A2(
        n_majority7_module_69__or_module_11_res), .ZN(
        n_majority7_module_69_res) );
  DFF_X1 u_reg_module_84__cini_mul_v00_reg ( .D(n_majority7_module_69_res), 
        .CK(clock_3), .Q(n_reg_module_84_res), .QN() );
  AND2_X1 u_majority7_module_70__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_70__and_module_1_res)
         );
  OR2_X1 u_majority7_module_70__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_70__or_module_1_res)
         );
  AND2_X1 u_majority7_module_70__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(n_majority7_module_70__and_module_2_res) );
  OR2_X1 u_majority7_module_70__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_70__or_module_2_res)
         );
  AND2_X1 u_majority7_module_70__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(n_majority7_module_70__and_module_3_res) );
  OR2_X1 u_majority7_module_70__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_70__or_module_3_res)
         );
  AND2_X1 u_majority7_module_70__and_module_4_U1 ( .A1(
        n_majority7_module_70__and_module_2_res), .A2(
        n_majority7_module_70__and_module_1_res), .ZN(
        n_majority7_module_70__and_module_4_res) );
  OR2_X1 u_majority7_module_70__or_module_4_U1 ( .A1(
        n_majority7_module_70__and_module_1_res), .A2(
        n_majority7_module_70__and_module_2_res), .ZN(
        n_majority7_module_70__or_module_4_res) );
  AND2_X1 u_majority7_module_70__and_module_5_U1 ( .A1(
        n_majority7_module_70__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_70__and_module_5_res) );
  OR2_X1 u_majority7_module_70__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_70__and_module_3_res), .ZN(
        n_majority7_module_70__or_module_5_res) );
  AND2_X1 u_majority7_module_70__and_module_6_U1 ( .A1(
        n_majority7_module_70__or_module_1_res), .A2(
        n_majority7_module_70__or_module_2_res), .ZN(
        n_majority7_module_70__and_module_6_res) );
  OR2_X1 u_majority7_module_70__or_module_6_U1 ( .A1(
        n_majority7_module_70__or_module_2_res), .A2(
        n_majority7_module_70__or_module_1_res), .ZN(
        n_majority7_module_70__or_module_6_res) );
  OR2_X1 u_majority7_module_70__or_module_7_U1 ( .A1(
        n_majority7_module_70__and_module_4_res), .A2(
        n_majority7_module_70__and_module_5_res), .ZN(
        n_majority7_module_70__or_module_7_res) );
  AND2_X1 u_majority7_module_70__and_module_7_U1 ( .A1(
        n_majority7_module_70__or_module_3_res), .A2(
        n_majority7_module_70__or_module_4_res), .ZN(
        n_majority7_module_70__and_module_7_res) );
  OR2_X1 u_majority7_module_70__or_module_8_U1 ( .A1(
        n_majority7_module_70__or_module_4_res), .A2(
        n_majority7_module_70__or_module_3_res), .ZN(
        n_majority7_module_70__or_module_8_res) );
  AND2_X1 u_majority7_module_70__and_module_8_U1 ( .A1(
        n_majority7_module_70__or_module_5_res), .A2(
        n_majority7_module_70__and_module_6_res), .ZN(
        n_majority7_module_70__and_module_8_res) );
  OR2_X1 u_majority7_module_70__or_module_9_U1 ( .A1(
        n_majority7_module_70__and_module_6_res), .A2(
        n_majority7_module_70__or_module_5_res), .ZN(
        n_majority7_module_70__or_module_9_res) );
  OR2_X1 u_majority7_module_70__or_module_10_U1 ( .A1(
        n_majority7_module_70__or_module_7_res), .A2(
        n_majority7_module_70__and_module_7_res), .ZN(
        n_majority7_module_70__or_module_10_res) );
  AND2_X1 u_majority7_module_70__and_module_9_U1 ( .A1(
        n_majority7_module_70__or_module_6_res), .A2(
        n_majority7_module_70__or_module_9_res), .ZN(
        n_majority7_module_70__and_module_9_res) );
  OR2_X1 u_majority7_module_70__or_module_11_U1 ( .A1(
        n_majority7_module_70__or_module_10_res), .A2(
        n_majority7_module_70__and_module_8_res), .ZN(
        n_majority7_module_70__or_module_11_res) );
  AND2_X1 u_majority7_module_70__and_module_10_U1 ( .A1(
        n_majority7_module_70__or_module_8_res), .A2(
        n_majority7_module_70__and_module_9_res), .ZN(
        n_majority7_module_70__and_module_10_res) );
  AND2_X1 u_majority7_module_70__and_module_11_U1 ( .A1(
        n_majority7_module_70__and_module_10_res), .A2(
        n_majority7_module_70__or_module_11_res), .ZN(
        n_majority7_module_70_res) );
  DFF_X1 u_reg_module_85__cini_mul_v00_reg ( .D(n_majority7_module_70_res), 
        .CK(clock_3), .Q(n_reg_module_85_res), .QN() );
  AND2_X1 u_majority7_module_71__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_71__and_module_1_res)
         );
  OR2_X1 u_majority7_module_71__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_71__or_module_1_res)
         );
  AND2_X1 u_majority7_module_71__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(n_majority7_module_71__and_module_2_res) );
  OR2_X1 u_majority7_module_71__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_71__or_module_2_res)
         );
  AND2_X1 u_majority7_module_71__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(n_majority7_module_71__and_module_3_res) );
  OR2_X1 u_majority7_module_71__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_71__or_module_3_res)
         );
  AND2_X1 u_majority7_module_71__and_module_4_U1 ( .A1(
        n_majority7_module_71__and_module_2_res), .A2(
        n_majority7_module_71__and_module_1_res), .ZN(
        n_majority7_module_71__and_module_4_res) );
  OR2_X1 u_majority7_module_71__or_module_4_U1 ( .A1(
        n_majority7_module_71__and_module_1_res), .A2(
        n_majority7_module_71__and_module_2_res), .ZN(
        n_majority7_module_71__or_module_4_res) );
  AND2_X1 u_majority7_module_71__and_module_5_U1 ( .A1(
        n_majority7_module_71__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_71__and_module_5_res) );
  OR2_X1 u_majority7_module_71__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_71__and_module_3_res), .ZN(
        n_majority7_module_71__or_module_5_res) );
  AND2_X1 u_majority7_module_71__and_module_6_U1 ( .A1(
        n_majority7_module_71__or_module_1_res), .A2(
        n_majority7_module_71__or_module_2_res), .ZN(
        n_majority7_module_71__and_module_6_res) );
  OR2_X1 u_majority7_module_71__or_module_6_U1 ( .A1(
        n_majority7_module_71__or_module_2_res), .A2(
        n_majority7_module_71__or_module_1_res), .ZN(
        n_majority7_module_71__or_module_6_res) );
  OR2_X1 u_majority7_module_71__or_module_7_U1 ( .A1(
        n_majority7_module_71__and_module_4_res), .A2(
        n_majority7_module_71__and_module_5_res), .ZN(
        n_majority7_module_71__or_module_7_res) );
  AND2_X1 u_majority7_module_71__and_module_7_U1 ( .A1(
        n_majority7_module_71__or_module_3_res), .A2(
        n_majority7_module_71__or_module_4_res), .ZN(
        n_majority7_module_71__and_module_7_res) );
  OR2_X1 u_majority7_module_71__or_module_8_U1 ( .A1(
        n_majority7_module_71__or_module_4_res), .A2(
        n_majority7_module_71__or_module_3_res), .ZN(
        n_majority7_module_71__or_module_8_res) );
  AND2_X1 u_majority7_module_71__and_module_8_U1 ( .A1(
        n_majority7_module_71__or_module_5_res), .A2(
        n_majority7_module_71__and_module_6_res), .ZN(
        n_majority7_module_71__and_module_8_res) );
  OR2_X1 u_majority7_module_71__or_module_9_U1 ( .A1(
        n_majority7_module_71__and_module_6_res), .A2(
        n_majority7_module_71__or_module_5_res), .ZN(
        n_majority7_module_71__or_module_9_res) );
  OR2_X1 u_majority7_module_71__or_module_10_U1 ( .A1(
        n_majority7_module_71__or_module_7_res), .A2(
        n_majority7_module_71__and_module_7_res), .ZN(
        n_majority7_module_71__or_module_10_res) );
  AND2_X1 u_majority7_module_71__and_module_9_U1 ( .A1(
        n_majority7_module_71__or_module_6_res), .A2(
        n_majority7_module_71__or_module_9_res), .ZN(
        n_majority7_module_71__and_module_9_res) );
  OR2_X1 u_majority7_module_71__or_module_11_U1 ( .A1(
        n_majority7_module_71__or_module_10_res), .A2(
        n_majority7_module_71__and_module_8_res), .ZN(
        n_majority7_module_71__or_module_11_res) );
  AND2_X1 u_majority7_module_71__and_module_10_U1 ( .A1(
        n_majority7_module_71__or_module_8_res), .A2(
        n_majority7_module_71__and_module_9_res), .ZN(
        n_majority7_module_71__and_module_10_res) );
  AND2_X1 u_majority7_module_71__and_module_11_U1 ( .A1(
        n_majority7_module_71__and_module_10_res), .A2(
        n_majority7_module_71__or_module_11_res), .ZN(
        n_majority7_module_71_res) );
  DFF_X1 u_reg_module_86__cini_mul_v00_reg ( .D(n_majority7_module_71_res), 
        .CK(clock_3), .Q(n_reg_module_86_res), .QN() );
  DFF_X1 u_reg_module_87__cini_mul_v00_reg ( .D(n_and_module_59_res), .CK(
        clock_3), .Q(n_reg_module_87_res), .QN() );
  AND2_X1 u_majority7_module_72__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_72__and_module_1_res)
         );
  OR2_X1 u_majority7_module_72__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_72__or_module_1_res)
         );
  AND2_X1 u_majority7_module_72__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(n_majority7_module_72__and_module_2_res) );
  OR2_X1 u_majority7_module_72__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_72__or_module_2_res)
         );
  AND2_X1 u_majority7_module_72__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(n_majority7_module_72__and_module_3_res) );
  OR2_X1 u_majority7_module_72__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_72__or_module_3_res)
         );
  AND2_X1 u_majority7_module_72__and_module_4_U1 ( .A1(
        n_majority7_module_72__and_module_2_res), .A2(
        n_majority7_module_72__and_module_1_res), .ZN(
        n_majority7_module_72__and_module_4_res) );
  OR2_X1 u_majority7_module_72__or_module_4_U1 ( .A1(
        n_majority7_module_72__and_module_1_res), .A2(
        n_majority7_module_72__and_module_2_res), .ZN(
        n_majority7_module_72__or_module_4_res) );
  AND2_X1 u_majority7_module_72__and_module_5_U1 ( .A1(
        n_majority7_module_72__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_72__and_module_5_res) );
  OR2_X1 u_majority7_module_72__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_72__and_module_3_res), .ZN(
        n_majority7_module_72__or_module_5_res) );
  AND2_X1 u_majority7_module_72__and_module_6_U1 ( .A1(
        n_majority7_module_72__or_module_1_res), .A2(
        n_majority7_module_72__or_module_2_res), .ZN(
        n_majority7_module_72__and_module_6_res) );
  OR2_X1 u_majority7_module_72__or_module_6_U1 ( .A1(
        n_majority7_module_72__or_module_2_res), .A2(
        n_majority7_module_72__or_module_1_res), .ZN(
        n_majority7_module_72__or_module_6_res) );
  OR2_X1 u_majority7_module_72__or_module_7_U1 ( .A1(
        n_majority7_module_72__and_module_4_res), .A2(
        n_majority7_module_72__and_module_5_res), .ZN(
        n_majority7_module_72__or_module_7_res) );
  AND2_X1 u_majority7_module_72__and_module_7_U1 ( .A1(
        n_majority7_module_72__or_module_3_res), .A2(
        n_majority7_module_72__or_module_4_res), .ZN(
        n_majority7_module_72__and_module_7_res) );
  OR2_X1 u_majority7_module_72__or_module_8_U1 ( .A1(
        n_majority7_module_72__or_module_4_res), .A2(
        n_majority7_module_72__or_module_3_res), .ZN(
        n_majority7_module_72__or_module_8_res) );
  AND2_X1 u_majority7_module_72__and_module_8_U1 ( .A1(
        n_majority7_module_72__or_module_5_res), .A2(
        n_majority7_module_72__and_module_6_res), .ZN(
        n_majority7_module_72__and_module_8_res) );
  OR2_X1 u_majority7_module_72__or_module_9_U1 ( .A1(
        n_majority7_module_72__and_module_6_res), .A2(
        n_majority7_module_72__or_module_5_res), .ZN(
        n_majority7_module_72__or_module_9_res) );
  OR2_X1 u_majority7_module_72__or_module_10_U1 ( .A1(
        n_majority7_module_72__or_module_7_res), .A2(
        n_majority7_module_72__and_module_7_res), .ZN(
        n_majority7_module_72__or_module_10_res) );
  AND2_X1 u_majority7_module_72__and_module_9_U1 ( .A1(
        n_majority7_module_72__or_module_6_res), .A2(
        n_majority7_module_72__or_module_9_res), .ZN(
        n_majority7_module_72__and_module_9_res) );
  OR2_X1 u_majority7_module_72__or_module_11_U1 ( .A1(
        n_majority7_module_72__or_module_10_res), .A2(
        n_majority7_module_72__and_module_8_res), .ZN(
        n_majority7_module_72__or_module_11_res) );
  AND2_X1 u_majority7_module_72__and_module_10_U1 ( .A1(
        n_majority7_module_72__or_module_8_res), .A2(
        n_majority7_module_72__and_module_9_res), .ZN(
        n_majority7_module_72__and_module_10_res) );
  AND2_X1 u_majority7_module_72__and_module_11_U1 ( .A1(
        n_majority7_module_72__and_module_10_res), .A2(
        n_majority7_module_72__or_module_11_res), .ZN(
        n_majority7_module_72_res) );
  DFF_X1 u_reg_module_88__cini_mul_v00_reg ( .D(n_majority7_module_72_res), 
        .CK(clock_3), .Q(n_reg_module_88_res), .QN() );
  AND2_X1 u_majority7_module_73__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_73__and_module_1_res)
         );
  OR2_X1 u_majority7_module_73__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_73__or_module_1_res)
         );
  AND2_X1 u_majority7_module_73__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(n_majority7_module_73__and_module_2_res) );
  OR2_X1 u_majority7_module_73__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_73__or_module_2_res)
         );
  AND2_X1 u_majority7_module_73__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(n_majority7_module_73__and_module_3_res) );
  OR2_X1 u_majority7_module_73__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_73__or_module_3_res)
         );
  AND2_X1 u_majority7_module_73__and_module_4_U1 ( .A1(
        n_majority7_module_73__and_module_2_res), .A2(
        n_majority7_module_73__and_module_1_res), .ZN(
        n_majority7_module_73__and_module_4_res) );
  OR2_X1 u_majority7_module_73__or_module_4_U1 ( .A1(
        n_majority7_module_73__and_module_1_res), .A2(
        n_majority7_module_73__and_module_2_res), .ZN(
        n_majority7_module_73__or_module_4_res) );
  AND2_X1 u_majority7_module_73__and_module_5_U1 ( .A1(
        n_majority7_module_73__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_73__and_module_5_res) );
  OR2_X1 u_majority7_module_73__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_73__and_module_3_res), .ZN(
        n_majority7_module_73__or_module_5_res) );
  AND2_X1 u_majority7_module_73__and_module_6_U1 ( .A1(
        n_majority7_module_73__or_module_1_res), .A2(
        n_majority7_module_73__or_module_2_res), .ZN(
        n_majority7_module_73__and_module_6_res) );
  OR2_X1 u_majority7_module_73__or_module_6_U1 ( .A1(
        n_majority7_module_73__or_module_2_res), .A2(
        n_majority7_module_73__or_module_1_res), .ZN(
        n_majority7_module_73__or_module_6_res) );
  OR2_X1 u_majority7_module_73__or_module_7_U1 ( .A1(
        n_majority7_module_73__and_module_4_res), .A2(
        n_majority7_module_73__and_module_5_res), .ZN(
        n_majority7_module_73__or_module_7_res) );
  AND2_X1 u_majority7_module_73__and_module_7_U1 ( .A1(
        n_majority7_module_73__or_module_3_res), .A2(
        n_majority7_module_73__or_module_4_res), .ZN(
        n_majority7_module_73__and_module_7_res) );
  OR2_X1 u_majority7_module_73__or_module_8_U1 ( .A1(
        n_majority7_module_73__or_module_4_res), .A2(
        n_majority7_module_73__or_module_3_res), .ZN(
        n_majority7_module_73__or_module_8_res) );
  AND2_X1 u_majority7_module_73__and_module_8_U1 ( .A1(
        n_majority7_module_73__or_module_5_res), .A2(
        n_majority7_module_73__and_module_6_res), .ZN(
        n_majority7_module_73__and_module_8_res) );
  OR2_X1 u_majority7_module_73__or_module_9_U1 ( .A1(
        n_majority7_module_73__and_module_6_res), .A2(
        n_majority7_module_73__or_module_5_res), .ZN(
        n_majority7_module_73__or_module_9_res) );
  OR2_X1 u_majority7_module_73__or_module_10_U1 ( .A1(
        n_majority7_module_73__or_module_7_res), .A2(
        n_majority7_module_73__and_module_7_res), .ZN(
        n_majority7_module_73__or_module_10_res) );
  AND2_X1 u_majority7_module_73__and_module_9_U1 ( .A1(
        n_majority7_module_73__or_module_6_res), .A2(
        n_majority7_module_73__or_module_9_res), .ZN(
        n_majority7_module_73__and_module_9_res) );
  OR2_X1 u_majority7_module_73__or_module_11_U1 ( .A1(
        n_majority7_module_73__or_module_10_res), .A2(
        n_majority7_module_73__and_module_8_res), .ZN(
        n_majority7_module_73__or_module_11_res) );
  AND2_X1 u_majority7_module_73__and_module_10_U1 ( .A1(
        n_majority7_module_73__or_module_8_res), .A2(
        n_majority7_module_73__and_module_9_res), .ZN(
        n_majority7_module_73__and_module_10_res) );
  AND2_X1 u_majority7_module_73__and_module_11_U1 ( .A1(
        n_majority7_module_73__and_module_10_res), .A2(
        n_majority7_module_73__or_module_11_res), .ZN(
        n_majority7_module_73_res) );
  DFF_X1 u_reg_module_89__cini_mul_v00_reg ( .D(n_majority7_module_73_res), 
        .CK(clock_3), .Q(n_reg_module_89_res), .QN() );
  AND2_X1 u_majority7_module_74__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_74__and_module_1_res)
         );
  OR2_X1 u_majority7_module_74__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_74__or_module_1_res)
         );
  AND2_X1 u_majority7_module_74__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(n_majority7_module_74__and_module_2_res) );
  OR2_X1 u_majority7_module_74__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_74__or_module_2_res)
         );
  AND2_X1 u_majority7_module_74__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(n_majority7_module_74__and_module_3_res) );
  OR2_X1 u_majority7_module_74__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_74__or_module_3_res)
         );
  AND2_X1 u_majority7_module_74__and_module_4_U1 ( .A1(
        n_majority7_module_74__and_module_2_res), .A2(
        n_majority7_module_74__and_module_1_res), .ZN(
        n_majority7_module_74__and_module_4_res) );
  OR2_X1 u_majority7_module_74__or_module_4_U1 ( .A1(
        n_majority7_module_74__and_module_1_res), .A2(
        n_majority7_module_74__and_module_2_res), .ZN(
        n_majority7_module_74__or_module_4_res) );
  AND2_X1 u_majority7_module_74__and_module_5_U1 ( .A1(
        n_majority7_module_74__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_74__and_module_5_res) );
  OR2_X1 u_majority7_module_74__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_74__and_module_3_res), .ZN(
        n_majority7_module_74__or_module_5_res) );
  AND2_X1 u_majority7_module_74__and_module_6_U1 ( .A1(
        n_majority7_module_74__or_module_1_res), .A2(
        n_majority7_module_74__or_module_2_res), .ZN(
        n_majority7_module_74__and_module_6_res) );
  OR2_X1 u_majority7_module_74__or_module_6_U1 ( .A1(
        n_majority7_module_74__or_module_2_res), .A2(
        n_majority7_module_74__or_module_1_res), .ZN(
        n_majority7_module_74__or_module_6_res) );
  OR2_X1 u_majority7_module_74__or_module_7_U1 ( .A1(
        n_majority7_module_74__and_module_4_res), .A2(
        n_majority7_module_74__and_module_5_res), .ZN(
        n_majority7_module_74__or_module_7_res) );
  AND2_X1 u_majority7_module_74__and_module_7_U1 ( .A1(
        n_majority7_module_74__or_module_3_res), .A2(
        n_majority7_module_74__or_module_4_res), .ZN(
        n_majority7_module_74__and_module_7_res) );
  OR2_X1 u_majority7_module_74__or_module_8_U1 ( .A1(
        n_majority7_module_74__or_module_4_res), .A2(
        n_majority7_module_74__or_module_3_res), .ZN(
        n_majority7_module_74__or_module_8_res) );
  AND2_X1 u_majority7_module_74__and_module_8_U1 ( .A1(
        n_majority7_module_74__or_module_5_res), .A2(
        n_majority7_module_74__and_module_6_res), .ZN(
        n_majority7_module_74__and_module_8_res) );
  OR2_X1 u_majority7_module_74__or_module_9_U1 ( .A1(
        n_majority7_module_74__and_module_6_res), .A2(
        n_majority7_module_74__or_module_5_res), .ZN(
        n_majority7_module_74__or_module_9_res) );
  OR2_X1 u_majority7_module_74__or_module_10_U1 ( .A1(
        n_majority7_module_74__or_module_7_res), .A2(
        n_majority7_module_74__and_module_7_res), .ZN(
        n_majority7_module_74__or_module_10_res) );
  AND2_X1 u_majority7_module_74__and_module_9_U1 ( .A1(
        n_majority7_module_74__or_module_6_res), .A2(
        n_majority7_module_74__or_module_9_res), .ZN(
        n_majority7_module_74__and_module_9_res) );
  OR2_X1 u_majority7_module_74__or_module_11_U1 ( .A1(
        n_majority7_module_74__or_module_10_res), .A2(
        n_majority7_module_74__and_module_8_res), .ZN(
        n_majority7_module_74__or_module_11_res) );
  AND2_X1 u_majority7_module_74__and_module_10_U1 ( .A1(
        n_majority7_module_74__or_module_8_res), .A2(
        n_majority7_module_74__and_module_9_res), .ZN(
        n_majority7_module_74__and_module_10_res) );
  AND2_X1 u_majority7_module_74__and_module_11_U1 ( .A1(
        n_majority7_module_74__and_module_10_res), .A2(
        n_majority7_module_74__or_module_11_res), .ZN(
        n_majority7_module_74_res) );
  DFF_X1 u_reg_module_90__cini_mul_v00_reg ( .D(n_majority7_module_74_res), 
        .CK(clock_3), .Q(n_reg_module_90_res), .QN() );
  AND2_X1 u_majority7_module_75__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_75__and_module_1_res)
         );
  OR2_X1 u_majority7_module_75__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_75__or_module_1_res)
         );
  AND2_X1 u_majority7_module_75__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(n_majority7_module_75__and_module_2_res) );
  OR2_X1 u_majority7_module_75__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_75__or_module_2_res)
         );
  AND2_X1 u_majority7_module_75__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(n_majority7_module_75__and_module_3_res) );
  OR2_X1 u_majority7_module_75__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_75__or_module_3_res)
         );
  AND2_X1 u_majority7_module_75__and_module_4_U1 ( .A1(
        n_majority7_module_75__and_module_2_res), .A2(
        n_majority7_module_75__and_module_1_res), .ZN(
        n_majority7_module_75__and_module_4_res) );
  OR2_X1 u_majority7_module_75__or_module_4_U1 ( .A1(
        n_majority7_module_75__and_module_1_res), .A2(
        n_majority7_module_75__and_module_2_res), .ZN(
        n_majority7_module_75__or_module_4_res) );
  AND2_X1 u_majority7_module_75__and_module_5_U1 ( .A1(
        n_majority7_module_75__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_75__and_module_5_res) );
  OR2_X1 u_majority7_module_75__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_75__and_module_3_res), .ZN(
        n_majority7_module_75__or_module_5_res) );
  AND2_X1 u_majority7_module_75__and_module_6_U1 ( .A1(
        n_majority7_module_75__or_module_1_res), .A2(
        n_majority7_module_75__or_module_2_res), .ZN(
        n_majority7_module_75__and_module_6_res) );
  OR2_X1 u_majority7_module_75__or_module_6_U1 ( .A1(
        n_majority7_module_75__or_module_2_res), .A2(
        n_majority7_module_75__or_module_1_res), .ZN(
        n_majority7_module_75__or_module_6_res) );
  OR2_X1 u_majority7_module_75__or_module_7_U1 ( .A1(
        n_majority7_module_75__and_module_4_res), .A2(
        n_majority7_module_75__and_module_5_res), .ZN(
        n_majority7_module_75__or_module_7_res) );
  AND2_X1 u_majority7_module_75__and_module_7_U1 ( .A1(
        n_majority7_module_75__or_module_3_res), .A2(
        n_majority7_module_75__or_module_4_res), .ZN(
        n_majority7_module_75__and_module_7_res) );
  OR2_X1 u_majority7_module_75__or_module_8_U1 ( .A1(
        n_majority7_module_75__or_module_4_res), .A2(
        n_majority7_module_75__or_module_3_res), .ZN(
        n_majority7_module_75__or_module_8_res) );
  AND2_X1 u_majority7_module_75__and_module_8_U1 ( .A1(
        n_majority7_module_75__or_module_5_res), .A2(
        n_majority7_module_75__and_module_6_res), .ZN(
        n_majority7_module_75__and_module_8_res) );
  OR2_X1 u_majority7_module_75__or_module_9_U1 ( .A1(
        n_majority7_module_75__and_module_6_res), .A2(
        n_majority7_module_75__or_module_5_res), .ZN(
        n_majority7_module_75__or_module_9_res) );
  OR2_X1 u_majority7_module_75__or_module_10_U1 ( .A1(
        n_majority7_module_75__or_module_7_res), .A2(
        n_majority7_module_75__and_module_7_res), .ZN(
        n_majority7_module_75__or_module_10_res) );
  AND2_X1 u_majority7_module_75__and_module_9_U1 ( .A1(
        n_majority7_module_75__or_module_6_res), .A2(
        n_majority7_module_75__or_module_9_res), .ZN(
        n_majority7_module_75__and_module_9_res) );
  OR2_X1 u_majority7_module_75__or_module_11_U1 ( .A1(
        n_majority7_module_75__or_module_10_res), .A2(
        n_majority7_module_75__and_module_8_res), .ZN(
        n_majority7_module_75__or_module_11_res) );
  AND2_X1 u_majority7_module_75__and_module_10_U1 ( .A1(
        n_majority7_module_75__or_module_8_res), .A2(
        n_majority7_module_75__and_module_9_res), .ZN(
        n_majority7_module_75__and_module_10_res) );
  AND2_X1 u_majority7_module_75__and_module_11_U1 ( .A1(
        n_majority7_module_75__and_module_10_res), .A2(
        n_majority7_module_75__or_module_11_res), .ZN(
        n_majority7_module_75_res) );
  DFF_X1 u_reg_module_91__cini_mul_v00_reg ( .D(n_majority7_module_75_res), 
        .CK(clock_3), .Q(n_reg_module_91_res), .QN() );
  DFF_X1 u_reg_module_92__cini_mul_v00_reg ( .D(n_and_module_64_res), .CK(
        clock_3), .Q(n_reg_module_92_res), .QN() );
  DFF_X1 u_reg_module_93__cini_mul_v00_reg ( .D(n_and_module_65_res), .CK(
        clock_4), .Q(n_reg_module_93_res), .QN() );
  AND2_X1 u_majority7_module_76__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_76__and_module_1_res)
         );
  OR2_X1 u_majority7_module_76__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_76__or_module_1_res)
         );
  AND2_X1 u_majority7_module_76__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(n_majority7_module_76__and_module_2_res) );
  OR2_X1 u_majority7_module_76__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_76__or_module_2_res)
         );
  AND2_X1 u_majority7_module_76__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(n_majority7_module_76__and_module_3_res) );
  OR2_X1 u_majority7_module_76__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_76__or_module_3_res)
         );
  AND2_X1 u_majority7_module_76__and_module_4_U1 ( .A1(
        n_majority7_module_76__and_module_2_res), .A2(
        n_majority7_module_76__and_module_1_res), .ZN(
        n_majority7_module_76__and_module_4_res) );
  OR2_X1 u_majority7_module_76__or_module_4_U1 ( .A1(
        n_majority7_module_76__and_module_1_res), .A2(
        n_majority7_module_76__and_module_2_res), .ZN(
        n_majority7_module_76__or_module_4_res) );
  AND2_X1 u_majority7_module_76__and_module_5_U1 ( .A1(
        n_majority7_module_76__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_76__and_module_5_res) );
  OR2_X1 u_majority7_module_76__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_76__and_module_3_res), .ZN(
        n_majority7_module_76__or_module_5_res) );
  AND2_X1 u_majority7_module_76__and_module_6_U1 ( .A1(
        n_majority7_module_76__or_module_1_res), .A2(
        n_majority7_module_76__or_module_2_res), .ZN(
        n_majority7_module_76__and_module_6_res) );
  OR2_X1 u_majority7_module_76__or_module_6_U1 ( .A1(
        n_majority7_module_76__or_module_2_res), .A2(
        n_majority7_module_76__or_module_1_res), .ZN(
        n_majority7_module_76__or_module_6_res) );
  OR2_X1 u_majority7_module_76__or_module_7_U1 ( .A1(
        n_majority7_module_76__and_module_4_res), .A2(
        n_majority7_module_76__and_module_5_res), .ZN(
        n_majority7_module_76__or_module_7_res) );
  AND2_X1 u_majority7_module_76__and_module_7_U1 ( .A1(
        n_majority7_module_76__or_module_3_res), .A2(
        n_majority7_module_76__or_module_4_res), .ZN(
        n_majority7_module_76__and_module_7_res) );
  OR2_X1 u_majority7_module_76__or_module_8_U1 ( .A1(
        n_majority7_module_76__or_module_4_res), .A2(
        n_majority7_module_76__or_module_3_res), .ZN(
        n_majority7_module_76__or_module_8_res) );
  AND2_X1 u_majority7_module_76__and_module_8_U1 ( .A1(
        n_majority7_module_76__or_module_5_res), .A2(
        n_majority7_module_76__and_module_6_res), .ZN(
        n_majority7_module_76__and_module_8_res) );
  OR2_X1 u_majority7_module_76__or_module_9_U1 ( .A1(
        n_majority7_module_76__and_module_6_res), .A2(
        n_majority7_module_76__or_module_5_res), .ZN(
        n_majority7_module_76__or_module_9_res) );
  OR2_X1 u_majority7_module_76__or_module_10_U1 ( .A1(
        n_majority7_module_76__or_module_7_res), .A2(
        n_majority7_module_76__and_module_7_res), .ZN(
        n_majority7_module_76__or_module_10_res) );
  AND2_X1 u_majority7_module_76__and_module_9_U1 ( .A1(
        n_majority7_module_76__or_module_6_res), .A2(
        n_majority7_module_76__or_module_9_res), .ZN(
        n_majority7_module_76__and_module_9_res) );
  OR2_X1 u_majority7_module_76__or_module_11_U1 ( .A1(
        n_majority7_module_76__or_module_10_res), .A2(
        n_majority7_module_76__and_module_8_res), .ZN(
        n_majority7_module_76__or_module_11_res) );
  AND2_X1 u_majority7_module_76__and_module_10_U1 ( .A1(
        n_majority7_module_76__or_module_8_res), .A2(
        n_majority7_module_76__and_module_9_res), .ZN(
        n_majority7_module_76__and_module_10_res) );
  AND2_X1 u_majority7_module_76__and_module_11_U1 ( .A1(
        n_majority7_module_76__and_module_10_res), .A2(
        n_majority7_module_76__or_module_11_res), .ZN(
        n_majority7_module_76_res) );
  DFF_X1 u_reg_module_94__cini_mul_v00_reg ( .D(n_majority7_module_76_res), 
        .CK(clock_4), .Q(n_reg_module_94_res), .QN() );
  AND2_X1 u_majority7_module_77__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_77__and_module_1_res)
         );
  OR2_X1 u_majority7_module_77__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_77__or_module_1_res)
         );
  AND2_X1 u_majority7_module_77__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(n_majority7_module_77__and_module_2_res) );
  OR2_X1 u_majority7_module_77__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_77__or_module_2_res)
         );
  AND2_X1 u_majority7_module_77__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(n_majority7_module_77__and_module_3_res) );
  OR2_X1 u_majority7_module_77__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_77__or_module_3_res)
         );
  AND2_X1 u_majority7_module_77__and_module_4_U1 ( .A1(
        n_majority7_module_77__and_module_2_res), .A2(
        n_majority7_module_77__and_module_1_res), .ZN(
        n_majority7_module_77__and_module_4_res) );
  OR2_X1 u_majority7_module_77__or_module_4_U1 ( .A1(
        n_majority7_module_77__and_module_1_res), .A2(
        n_majority7_module_77__and_module_2_res), .ZN(
        n_majority7_module_77__or_module_4_res) );
  AND2_X1 u_majority7_module_77__and_module_5_U1 ( .A1(
        n_majority7_module_77__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_77__and_module_5_res) );
  OR2_X1 u_majority7_module_77__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_77__and_module_3_res), .ZN(
        n_majority7_module_77__or_module_5_res) );
  AND2_X1 u_majority7_module_77__and_module_6_U1 ( .A1(
        n_majority7_module_77__or_module_1_res), .A2(
        n_majority7_module_77__or_module_2_res), .ZN(
        n_majority7_module_77__and_module_6_res) );
  OR2_X1 u_majority7_module_77__or_module_6_U1 ( .A1(
        n_majority7_module_77__or_module_2_res), .A2(
        n_majority7_module_77__or_module_1_res), .ZN(
        n_majority7_module_77__or_module_6_res) );
  OR2_X1 u_majority7_module_77__or_module_7_U1 ( .A1(
        n_majority7_module_77__and_module_4_res), .A2(
        n_majority7_module_77__and_module_5_res), .ZN(
        n_majority7_module_77__or_module_7_res) );
  AND2_X1 u_majority7_module_77__and_module_7_U1 ( .A1(
        n_majority7_module_77__or_module_3_res), .A2(
        n_majority7_module_77__or_module_4_res), .ZN(
        n_majority7_module_77__and_module_7_res) );
  OR2_X1 u_majority7_module_77__or_module_8_U1 ( .A1(
        n_majority7_module_77__or_module_4_res), .A2(
        n_majority7_module_77__or_module_3_res), .ZN(
        n_majority7_module_77__or_module_8_res) );
  AND2_X1 u_majority7_module_77__and_module_8_U1 ( .A1(
        n_majority7_module_77__or_module_5_res), .A2(
        n_majority7_module_77__and_module_6_res), .ZN(
        n_majority7_module_77__and_module_8_res) );
  OR2_X1 u_majority7_module_77__or_module_9_U1 ( .A1(
        n_majority7_module_77__and_module_6_res), .A2(
        n_majority7_module_77__or_module_5_res), .ZN(
        n_majority7_module_77__or_module_9_res) );
  OR2_X1 u_majority7_module_77__or_module_10_U1 ( .A1(
        n_majority7_module_77__or_module_7_res), .A2(
        n_majority7_module_77__and_module_7_res), .ZN(
        n_majority7_module_77__or_module_10_res) );
  AND2_X1 u_majority7_module_77__and_module_9_U1 ( .A1(
        n_majority7_module_77__or_module_6_res), .A2(
        n_majority7_module_77__or_module_9_res), .ZN(
        n_majority7_module_77__and_module_9_res) );
  OR2_X1 u_majority7_module_77__or_module_11_U1 ( .A1(
        n_majority7_module_77__or_module_10_res), .A2(
        n_majority7_module_77__and_module_8_res), .ZN(
        n_majority7_module_77__or_module_11_res) );
  AND2_X1 u_majority7_module_77__and_module_10_U1 ( .A1(
        n_majority7_module_77__or_module_8_res), .A2(
        n_majority7_module_77__and_module_9_res), .ZN(
        n_majority7_module_77__and_module_10_res) );
  AND2_X1 u_majority7_module_77__and_module_11_U1 ( .A1(
        n_majority7_module_77__and_module_10_res), .A2(
        n_majority7_module_77__or_module_11_res), .ZN(
        n_majority7_module_77_res) );
  DFF_X1 u_reg_module_95__cini_mul_v00_reg ( .D(n_majority7_module_77_res), 
        .CK(clock_4), .Q(n_reg_module_95_res), .QN() );
  AND2_X1 u_majority7_module_78__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_78__and_module_1_res)
         );
  OR2_X1 u_majority7_module_78__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_78__or_module_1_res)
         );
  AND2_X1 u_majority7_module_78__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(n_majority7_module_78__and_module_2_res) );
  OR2_X1 u_majority7_module_78__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_78__or_module_2_res)
         );
  AND2_X1 u_majority7_module_78__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(n_majority7_module_78__and_module_3_res) );
  OR2_X1 u_majority7_module_78__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_78__or_module_3_res)
         );
  AND2_X1 u_majority7_module_78__and_module_4_U1 ( .A1(
        n_majority7_module_78__and_module_2_res), .A2(
        n_majority7_module_78__and_module_1_res), .ZN(
        n_majority7_module_78__and_module_4_res) );
  OR2_X1 u_majority7_module_78__or_module_4_U1 ( .A1(
        n_majority7_module_78__and_module_1_res), .A2(
        n_majority7_module_78__and_module_2_res), .ZN(
        n_majority7_module_78__or_module_4_res) );
  AND2_X1 u_majority7_module_78__and_module_5_U1 ( .A1(
        n_majority7_module_78__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_78__and_module_5_res) );
  OR2_X1 u_majority7_module_78__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_78__and_module_3_res), .ZN(
        n_majority7_module_78__or_module_5_res) );
  AND2_X1 u_majority7_module_78__and_module_6_U1 ( .A1(
        n_majority7_module_78__or_module_1_res), .A2(
        n_majority7_module_78__or_module_2_res), .ZN(
        n_majority7_module_78__and_module_6_res) );
  OR2_X1 u_majority7_module_78__or_module_6_U1 ( .A1(
        n_majority7_module_78__or_module_2_res), .A2(
        n_majority7_module_78__or_module_1_res), .ZN(
        n_majority7_module_78__or_module_6_res) );
  OR2_X1 u_majority7_module_78__or_module_7_U1 ( .A1(
        n_majority7_module_78__and_module_4_res), .A2(
        n_majority7_module_78__and_module_5_res), .ZN(
        n_majority7_module_78__or_module_7_res) );
  AND2_X1 u_majority7_module_78__and_module_7_U1 ( .A1(
        n_majority7_module_78__or_module_3_res), .A2(
        n_majority7_module_78__or_module_4_res), .ZN(
        n_majority7_module_78__and_module_7_res) );
  OR2_X1 u_majority7_module_78__or_module_8_U1 ( .A1(
        n_majority7_module_78__or_module_4_res), .A2(
        n_majority7_module_78__or_module_3_res), .ZN(
        n_majority7_module_78__or_module_8_res) );
  AND2_X1 u_majority7_module_78__and_module_8_U1 ( .A1(
        n_majority7_module_78__or_module_5_res), .A2(
        n_majority7_module_78__and_module_6_res), .ZN(
        n_majority7_module_78__and_module_8_res) );
  OR2_X1 u_majority7_module_78__or_module_9_U1 ( .A1(
        n_majority7_module_78__and_module_6_res), .A2(
        n_majority7_module_78__or_module_5_res), .ZN(
        n_majority7_module_78__or_module_9_res) );
  OR2_X1 u_majority7_module_78__or_module_10_U1 ( .A1(
        n_majority7_module_78__or_module_7_res), .A2(
        n_majority7_module_78__and_module_7_res), .ZN(
        n_majority7_module_78__or_module_10_res) );
  AND2_X1 u_majority7_module_78__and_module_9_U1 ( .A1(
        n_majority7_module_78__or_module_6_res), .A2(
        n_majority7_module_78__or_module_9_res), .ZN(
        n_majority7_module_78__and_module_9_res) );
  OR2_X1 u_majority7_module_78__or_module_11_U1 ( .A1(
        n_majority7_module_78__or_module_10_res), .A2(
        n_majority7_module_78__and_module_8_res), .ZN(
        n_majority7_module_78__or_module_11_res) );
  AND2_X1 u_majority7_module_78__and_module_10_U1 ( .A1(
        n_majority7_module_78__or_module_8_res), .A2(
        n_majority7_module_78__and_module_9_res), .ZN(
        n_majority7_module_78__and_module_10_res) );
  AND2_X1 u_majority7_module_78__and_module_11_U1 ( .A1(
        n_majority7_module_78__and_module_10_res), .A2(
        n_majority7_module_78__or_module_11_res), .ZN(
        n_majority7_module_78_res) );
  DFF_X1 u_reg_module_96__cini_mul_v00_reg ( .D(n_majority7_module_78_res), 
        .CK(clock_4), .Q(n_reg_module_96_res), .QN() );
  AND2_X1 u_majority7_module_79__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_79__and_module_1_res)
         );
  OR2_X1 u_majority7_module_79__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_79__or_module_1_res)
         );
  AND2_X1 u_majority7_module_79__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(n_majority7_module_79__and_module_2_res) );
  OR2_X1 u_majority7_module_79__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_79__or_module_2_res)
         );
  AND2_X1 u_majority7_module_79__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(n_majority7_module_79__and_module_3_res) );
  OR2_X1 u_majority7_module_79__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_79__or_module_3_res)
         );
  AND2_X1 u_majority7_module_79__and_module_4_U1 ( .A1(
        n_majority7_module_79__and_module_2_res), .A2(
        n_majority7_module_79__and_module_1_res), .ZN(
        n_majority7_module_79__and_module_4_res) );
  OR2_X1 u_majority7_module_79__or_module_4_U1 ( .A1(
        n_majority7_module_79__and_module_1_res), .A2(
        n_majority7_module_79__and_module_2_res), .ZN(
        n_majority7_module_79__or_module_4_res) );
  AND2_X1 u_majority7_module_79__and_module_5_U1 ( .A1(
        n_majority7_module_79__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_79__and_module_5_res) );
  OR2_X1 u_majority7_module_79__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_79__and_module_3_res), .ZN(
        n_majority7_module_79__or_module_5_res) );
  AND2_X1 u_majority7_module_79__and_module_6_U1 ( .A1(
        n_majority7_module_79__or_module_1_res), .A2(
        n_majority7_module_79__or_module_2_res), .ZN(
        n_majority7_module_79__and_module_6_res) );
  OR2_X1 u_majority7_module_79__or_module_6_U1 ( .A1(
        n_majority7_module_79__or_module_2_res), .A2(
        n_majority7_module_79__or_module_1_res), .ZN(
        n_majority7_module_79__or_module_6_res) );
  OR2_X1 u_majority7_module_79__or_module_7_U1 ( .A1(
        n_majority7_module_79__and_module_4_res), .A2(
        n_majority7_module_79__and_module_5_res), .ZN(
        n_majority7_module_79__or_module_7_res) );
  AND2_X1 u_majority7_module_79__and_module_7_U1 ( .A1(
        n_majority7_module_79__or_module_3_res), .A2(
        n_majority7_module_79__or_module_4_res), .ZN(
        n_majority7_module_79__and_module_7_res) );
  OR2_X1 u_majority7_module_79__or_module_8_U1 ( .A1(
        n_majority7_module_79__or_module_4_res), .A2(
        n_majority7_module_79__or_module_3_res), .ZN(
        n_majority7_module_79__or_module_8_res) );
  AND2_X1 u_majority7_module_79__and_module_8_U1 ( .A1(
        n_majority7_module_79__or_module_5_res), .A2(
        n_majority7_module_79__and_module_6_res), .ZN(
        n_majority7_module_79__and_module_8_res) );
  OR2_X1 u_majority7_module_79__or_module_9_U1 ( .A1(
        n_majority7_module_79__and_module_6_res), .A2(
        n_majority7_module_79__or_module_5_res), .ZN(
        n_majority7_module_79__or_module_9_res) );
  OR2_X1 u_majority7_module_79__or_module_10_U1 ( .A1(
        n_majority7_module_79__or_module_7_res), .A2(
        n_majority7_module_79__and_module_7_res), .ZN(
        n_majority7_module_79__or_module_10_res) );
  AND2_X1 u_majority7_module_79__and_module_9_U1 ( .A1(
        n_majority7_module_79__or_module_6_res), .A2(
        n_majority7_module_79__or_module_9_res), .ZN(
        n_majority7_module_79__and_module_9_res) );
  OR2_X1 u_majority7_module_79__or_module_11_U1 ( .A1(
        n_majority7_module_79__or_module_10_res), .A2(
        n_majority7_module_79__and_module_8_res), .ZN(
        n_majority7_module_79__or_module_11_res) );
  AND2_X1 u_majority7_module_79__and_module_10_U1 ( .A1(
        n_majority7_module_79__or_module_8_res), .A2(
        n_majority7_module_79__and_module_9_res), .ZN(
        n_majority7_module_79__and_module_10_res) );
  AND2_X1 u_majority7_module_79__and_module_11_U1 ( .A1(
        n_majority7_module_79__and_module_10_res), .A2(
        n_majority7_module_79__or_module_11_res), .ZN(
        n_majority7_module_79_res) );
  DFF_X1 u_reg_module_97__cini_mul_v00_reg ( .D(n_majority7_module_79_res), 
        .CK(clock_4), .Q(n_reg_module_97_res), .QN() );
  DFF_X1 u_reg_module_98__cini_mul_v00_reg ( .D(n_and_module_70_res), .CK(
        clock_4), .Q(n_reg_module_98_res), .QN() );
  AND2_X1 u_majority7_module_80__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_80__and_module_1_res)
         );
  OR2_X1 u_majority7_module_80__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_80__or_module_1_res)
         );
  AND2_X1 u_majority7_module_80__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(n_majority7_module_80__and_module_2_res) );
  OR2_X1 u_majority7_module_80__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_80__or_module_2_res)
         );
  AND2_X1 u_majority7_module_80__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(n_majority7_module_80__and_module_3_res) );
  OR2_X1 u_majority7_module_80__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_80__or_module_3_res)
         );
  AND2_X1 u_majority7_module_80__and_module_4_U1 ( .A1(
        n_majority7_module_80__and_module_2_res), .A2(
        n_majority7_module_80__and_module_1_res), .ZN(
        n_majority7_module_80__and_module_4_res) );
  OR2_X1 u_majority7_module_80__or_module_4_U1 ( .A1(
        n_majority7_module_80__and_module_1_res), .A2(
        n_majority7_module_80__and_module_2_res), .ZN(
        n_majority7_module_80__or_module_4_res) );
  AND2_X1 u_majority7_module_80__and_module_5_U1 ( .A1(
        n_majority7_module_80__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_80__and_module_5_res) );
  OR2_X1 u_majority7_module_80__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_80__and_module_3_res), .ZN(
        n_majority7_module_80__or_module_5_res) );
  AND2_X1 u_majority7_module_80__and_module_6_U1 ( .A1(
        n_majority7_module_80__or_module_1_res), .A2(
        n_majority7_module_80__or_module_2_res), .ZN(
        n_majority7_module_80__and_module_6_res) );
  OR2_X1 u_majority7_module_80__or_module_6_U1 ( .A1(
        n_majority7_module_80__or_module_2_res), .A2(
        n_majority7_module_80__or_module_1_res), .ZN(
        n_majority7_module_80__or_module_6_res) );
  OR2_X1 u_majority7_module_80__or_module_7_U1 ( .A1(
        n_majority7_module_80__and_module_4_res), .A2(
        n_majority7_module_80__and_module_5_res), .ZN(
        n_majority7_module_80__or_module_7_res) );
  AND2_X1 u_majority7_module_80__and_module_7_U1 ( .A1(
        n_majority7_module_80__or_module_3_res), .A2(
        n_majority7_module_80__or_module_4_res), .ZN(
        n_majority7_module_80__and_module_7_res) );
  OR2_X1 u_majority7_module_80__or_module_8_U1 ( .A1(
        n_majority7_module_80__or_module_4_res), .A2(
        n_majority7_module_80__or_module_3_res), .ZN(
        n_majority7_module_80__or_module_8_res) );
  AND2_X1 u_majority7_module_80__and_module_8_U1 ( .A1(
        n_majority7_module_80__or_module_5_res), .A2(
        n_majority7_module_80__and_module_6_res), .ZN(
        n_majority7_module_80__and_module_8_res) );
  OR2_X1 u_majority7_module_80__or_module_9_U1 ( .A1(
        n_majority7_module_80__and_module_6_res), .A2(
        n_majority7_module_80__or_module_5_res), .ZN(
        n_majority7_module_80__or_module_9_res) );
  OR2_X1 u_majority7_module_80__or_module_10_U1 ( .A1(
        n_majority7_module_80__or_module_7_res), .A2(
        n_majority7_module_80__and_module_7_res), .ZN(
        n_majority7_module_80__or_module_10_res) );
  AND2_X1 u_majority7_module_80__and_module_9_U1 ( .A1(
        n_majority7_module_80__or_module_6_res), .A2(
        n_majority7_module_80__or_module_9_res), .ZN(
        n_majority7_module_80__and_module_9_res) );
  OR2_X1 u_majority7_module_80__or_module_11_U1 ( .A1(
        n_majority7_module_80__or_module_10_res), .A2(
        n_majority7_module_80__and_module_8_res), .ZN(
        n_majority7_module_80__or_module_11_res) );
  AND2_X1 u_majority7_module_80__and_module_10_U1 ( .A1(
        n_majority7_module_80__or_module_8_res), .A2(
        n_majority7_module_80__and_module_9_res), .ZN(
        n_majority7_module_80__and_module_10_res) );
  AND2_X1 u_majority7_module_80__and_module_11_U1 ( .A1(
        n_majority7_module_80__and_module_10_res), .A2(
        n_majority7_module_80__or_module_11_res), .ZN(
        n_majority7_module_80_res) );
  DFF_X1 u_reg_module_99__cini_mul_v00_reg ( .D(n_majority7_module_80_res), 
        .CK(clock_4), .Q(n_reg_module_99_res), .QN() );
  AND2_X1 u_majority7_module_81__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_81__and_module_1_res)
         );
  OR2_X1 u_majority7_module_81__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_81__or_module_1_res)
         );
  AND2_X1 u_majority7_module_81__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(n_majority7_module_81__and_module_2_res) );
  OR2_X1 u_majority7_module_81__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_81__or_module_2_res)
         );
  AND2_X1 u_majority7_module_81__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(n_majority7_module_81__and_module_3_res) );
  OR2_X1 u_majority7_module_81__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_81__or_module_3_res)
         );
  AND2_X1 u_majority7_module_81__and_module_4_U1 ( .A1(
        n_majority7_module_81__and_module_2_res), .A2(
        n_majority7_module_81__and_module_1_res), .ZN(
        n_majority7_module_81__and_module_4_res) );
  OR2_X1 u_majority7_module_81__or_module_4_U1 ( .A1(
        n_majority7_module_81__and_module_1_res), .A2(
        n_majority7_module_81__and_module_2_res), .ZN(
        n_majority7_module_81__or_module_4_res) );
  AND2_X1 u_majority7_module_81__and_module_5_U1 ( .A1(
        n_majority7_module_81__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_81__and_module_5_res) );
  OR2_X1 u_majority7_module_81__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_81__and_module_3_res), .ZN(
        n_majority7_module_81__or_module_5_res) );
  AND2_X1 u_majority7_module_81__and_module_6_U1 ( .A1(
        n_majority7_module_81__or_module_1_res), .A2(
        n_majority7_module_81__or_module_2_res), .ZN(
        n_majority7_module_81__and_module_6_res) );
  OR2_X1 u_majority7_module_81__or_module_6_U1 ( .A1(
        n_majority7_module_81__or_module_2_res), .A2(
        n_majority7_module_81__or_module_1_res), .ZN(
        n_majority7_module_81__or_module_6_res) );
  OR2_X1 u_majority7_module_81__or_module_7_U1 ( .A1(
        n_majority7_module_81__and_module_4_res), .A2(
        n_majority7_module_81__and_module_5_res), .ZN(
        n_majority7_module_81__or_module_7_res) );
  AND2_X1 u_majority7_module_81__and_module_7_U1 ( .A1(
        n_majority7_module_81__or_module_3_res), .A2(
        n_majority7_module_81__or_module_4_res), .ZN(
        n_majority7_module_81__and_module_7_res) );
  OR2_X1 u_majority7_module_81__or_module_8_U1 ( .A1(
        n_majority7_module_81__or_module_4_res), .A2(
        n_majority7_module_81__or_module_3_res), .ZN(
        n_majority7_module_81__or_module_8_res) );
  AND2_X1 u_majority7_module_81__and_module_8_U1 ( .A1(
        n_majority7_module_81__or_module_5_res), .A2(
        n_majority7_module_81__and_module_6_res), .ZN(
        n_majority7_module_81__and_module_8_res) );
  OR2_X1 u_majority7_module_81__or_module_9_U1 ( .A1(
        n_majority7_module_81__and_module_6_res), .A2(
        n_majority7_module_81__or_module_5_res), .ZN(
        n_majority7_module_81__or_module_9_res) );
  OR2_X1 u_majority7_module_81__or_module_10_U1 ( .A1(
        n_majority7_module_81__or_module_7_res), .A2(
        n_majority7_module_81__and_module_7_res), .ZN(
        n_majority7_module_81__or_module_10_res) );
  AND2_X1 u_majority7_module_81__and_module_9_U1 ( .A1(
        n_majority7_module_81__or_module_6_res), .A2(
        n_majority7_module_81__or_module_9_res), .ZN(
        n_majority7_module_81__and_module_9_res) );
  OR2_X1 u_majority7_module_81__or_module_11_U1 ( .A1(
        n_majority7_module_81__or_module_10_res), .A2(
        n_majority7_module_81__and_module_8_res), .ZN(
        n_majority7_module_81__or_module_11_res) );
  AND2_X1 u_majority7_module_81__and_module_10_U1 ( .A1(
        n_majority7_module_81__or_module_8_res), .A2(
        n_majority7_module_81__and_module_9_res), .ZN(
        n_majority7_module_81__and_module_10_res) );
  AND2_X1 u_majority7_module_81__and_module_11_U1 ( .A1(
        n_majority7_module_81__and_module_10_res), .A2(
        n_majority7_module_81__or_module_11_res), .ZN(
        n_majority7_module_81_res) );
  DFF_X1 u_reg_module_100__cini_mul_v00_reg ( .D(n_majority7_module_81_res), 
        .CK(clock_4), .Q(n_reg_module_100_res), .QN() );
  AND2_X1 u_majority7_module_82__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_82__and_module_1_res)
         );
  OR2_X1 u_majority7_module_82__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_82__or_module_1_res)
         );
  AND2_X1 u_majority7_module_82__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(n_majority7_module_82__and_module_2_res) );
  OR2_X1 u_majority7_module_82__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_82__or_module_2_res)
         );
  AND2_X1 u_majority7_module_82__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(n_majority7_module_82__and_module_3_res) );
  OR2_X1 u_majority7_module_82__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_82__or_module_3_res)
         );
  AND2_X1 u_majority7_module_82__and_module_4_U1 ( .A1(
        n_majority7_module_82__and_module_2_res), .A2(
        n_majority7_module_82__and_module_1_res), .ZN(
        n_majority7_module_82__and_module_4_res) );
  OR2_X1 u_majority7_module_82__or_module_4_U1 ( .A1(
        n_majority7_module_82__and_module_1_res), .A2(
        n_majority7_module_82__and_module_2_res), .ZN(
        n_majority7_module_82__or_module_4_res) );
  AND2_X1 u_majority7_module_82__and_module_5_U1 ( .A1(
        n_majority7_module_82__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_82__and_module_5_res) );
  OR2_X1 u_majority7_module_82__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_82__and_module_3_res), .ZN(
        n_majority7_module_82__or_module_5_res) );
  AND2_X1 u_majority7_module_82__and_module_6_U1 ( .A1(
        n_majority7_module_82__or_module_1_res), .A2(
        n_majority7_module_82__or_module_2_res), .ZN(
        n_majority7_module_82__and_module_6_res) );
  OR2_X1 u_majority7_module_82__or_module_6_U1 ( .A1(
        n_majority7_module_82__or_module_2_res), .A2(
        n_majority7_module_82__or_module_1_res), .ZN(
        n_majority7_module_82__or_module_6_res) );
  OR2_X1 u_majority7_module_82__or_module_7_U1 ( .A1(
        n_majority7_module_82__and_module_4_res), .A2(
        n_majority7_module_82__and_module_5_res), .ZN(
        n_majority7_module_82__or_module_7_res) );
  AND2_X1 u_majority7_module_82__and_module_7_U1 ( .A1(
        n_majority7_module_82__or_module_3_res), .A2(
        n_majority7_module_82__or_module_4_res), .ZN(
        n_majority7_module_82__and_module_7_res) );
  OR2_X1 u_majority7_module_82__or_module_8_U1 ( .A1(
        n_majority7_module_82__or_module_4_res), .A2(
        n_majority7_module_82__or_module_3_res), .ZN(
        n_majority7_module_82__or_module_8_res) );
  AND2_X1 u_majority7_module_82__and_module_8_U1 ( .A1(
        n_majority7_module_82__or_module_5_res), .A2(
        n_majority7_module_82__and_module_6_res), .ZN(
        n_majority7_module_82__and_module_8_res) );
  OR2_X1 u_majority7_module_82__or_module_9_U1 ( .A1(
        n_majority7_module_82__and_module_6_res), .A2(
        n_majority7_module_82__or_module_5_res), .ZN(
        n_majority7_module_82__or_module_9_res) );
  OR2_X1 u_majority7_module_82__or_module_10_U1 ( .A1(
        n_majority7_module_82__or_module_7_res), .A2(
        n_majority7_module_82__and_module_7_res), .ZN(
        n_majority7_module_82__or_module_10_res) );
  AND2_X1 u_majority7_module_82__and_module_9_U1 ( .A1(
        n_majority7_module_82__or_module_6_res), .A2(
        n_majority7_module_82__or_module_9_res), .ZN(
        n_majority7_module_82__and_module_9_res) );
  OR2_X1 u_majority7_module_82__or_module_11_U1 ( .A1(
        n_majority7_module_82__or_module_10_res), .A2(
        n_majority7_module_82__and_module_8_res), .ZN(
        n_majority7_module_82__or_module_11_res) );
  AND2_X1 u_majority7_module_82__and_module_10_U1 ( .A1(
        n_majority7_module_82__or_module_8_res), .A2(
        n_majority7_module_82__and_module_9_res), .ZN(
        n_majority7_module_82__and_module_10_res) );
  AND2_X1 u_majority7_module_82__and_module_11_U1 ( .A1(
        n_majority7_module_82__and_module_10_res), .A2(
        n_majority7_module_82__or_module_11_res), .ZN(
        n_majority7_module_82_res) );
  DFF_X1 u_reg_module_101__cini_mul_v00_reg ( .D(n_majority7_module_82_res), 
        .CK(clock_4), .Q(n_reg_module_101_res), .QN() );
  AND2_X1 u_majority7_module_83__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_83__and_module_1_res)
         );
  OR2_X1 u_majority7_module_83__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_83__or_module_1_res)
         );
  AND2_X1 u_majority7_module_83__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(n_majority7_module_83__and_module_2_res) );
  OR2_X1 u_majority7_module_83__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_83__or_module_2_res)
         );
  AND2_X1 u_majority7_module_83__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(n_majority7_module_83__and_module_3_res) );
  OR2_X1 u_majority7_module_83__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_83__or_module_3_res)
         );
  AND2_X1 u_majority7_module_83__and_module_4_U1 ( .A1(
        n_majority7_module_83__and_module_2_res), .A2(
        n_majority7_module_83__and_module_1_res), .ZN(
        n_majority7_module_83__and_module_4_res) );
  OR2_X1 u_majority7_module_83__or_module_4_U1 ( .A1(
        n_majority7_module_83__and_module_1_res), .A2(
        n_majority7_module_83__and_module_2_res), .ZN(
        n_majority7_module_83__or_module_4_res) );
  AND2_X1 u_majority7_module_83__and_module_5_U1 ( .A1(
        n_majority7_module_83__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_83__and_module_5_res) );
  OR2_X1 u_majority7_module_83__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_83__and_module_3_res), .ZN(
        n_majority7_module_83__or_module_5_res) );
  AND2_X1 u_majority7_module_83__and_module_6_U1 ( .A1(
        n_majority7_module_83__or_module_1_res), .A2(
        n_majority7_module_83__or_module_2_res), .ZN(
        n_majority7_module_83__and_module_6_res) );
  OR2_X1 u_majority7_module_83__or_module_6_U1 ( .A1(
        n_majority7_module_83__or_module_2_res), .A2(
        n_majority7_module_83__or_module_1_res), .ZN(
        n_majority7_module_83__or_module_6_res) );
  OR2_X1 u_majority7_module_83__or_module_7_U1 ( .A1(
        n_majority7_module_83__and_module_4_res), .A2(
        n_majority7_module_83__and_module_5_res), .ZN(
        n_majority7_module_83__or_module_7_res) );
  AND2_X1 u_majority7_module_83__and_module_7_U1 ( .A1(
        n_majority7_module_83__or_module_3_res), .A2(
        n_majority7_module_83__or_module_4_res), .ZN(
        n_majority7_module_83__and_module_7_res) );
  OR2_X1 u_majority7_module_83__or_module_8_U1 ( .A1(
        n_majority7_module_83__or_module_4_res), .A2(
        n_majority7_module_83__or_module_3_res), .ZN(
        n_majority7_module_83__or_module_8_res) );
  AND2_X1 u_majority7_module_83__and_module_8_U1 ( .A1(
        n_majority7_module_83__or_module_5_res), .A2(
        n_majority7_module_83__and_module_6_res), .ZN(
        n_majority7_module_83__and_module_8_res) );
  OR2_X1 u_majority7_module_83__or_module_9_U1 ( .A1(
        n_majority7_module_83__and_module_6_res), .A2(
        n_majority7_module_83__or_module_5_res), .ZN(
        n_majority7_module_83__or_module_9_res) );
  OR2_X1 u_majority7_module_83__or_module_10_U1 ( .A1(
        n_majority7_module_83__or_module_7_res), .A2(
        n_majority7_module_83__and_module_7_res), .ZN(
        n_majority7_module_83__or_module_10_res) );
  AND2_X1 u_majority7_module_83__and_module_9_U1 ( .A1(
        n_majority7_module_83__or_module_6_res), .A2(
        n_majority7_module_83__or_module_9_res), .ZN(
        n_majority7_module_83__and_module_9_res) );
  OR2_X1 u_majority7_module_83__or_module_11_U1 ( .A1(
        n_majority7_module_83__or_module_10_res), .A2(
        n_majority7_module_83__and_module_8_res), .ZN(
        n_majority7_module_83__or_module_11_res) );
  AND2_X1 u_majority7_module_83__and_module_10_U1 ( .A1(
        n_majority7_module_83__or_module_8_res), .A2(
        n_majority7_module_83__and_module_9_res), .ZN(
        n_majority7_module_83__and_module_10_res) );
  AND2_X1 u_majority7_module_83__and_module_11_U1 ( .A1(
        n_majority7_module_83__and_module_10_res), .A2(
        n_majority7_module_83__or_module_11_res), .ZN(
        n_majority7_module_83_res) );
  DFF_X1 u_reg_module_102__cini_mul_v00_reg ( .D(n_majority7_module_83_res), 
        .CK(clock_4), .Q(n_reg_module_102_res), .QN() );
  DFF_X1 u_reg_module_103__cini_mul_v00_reg ( .D(n_and_module_75_res), .CK(
        clock_4), .Q(n_reg_module_103_res), .QN() );
  AND2_X1 u_majority7_module_84__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_84__and_module_1_res)
         );
  OR2_X1 u_majority7_module_84__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_84__or_module_1_res)
         );
  AND2_X1 u_majority7_module_84__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(n_majority7_module_84__and_module_2_res) );
  OR2_X1 u_majority7_module_84__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_84__or_module_2_res)
         );
  AND2_X1 u_majority7_module_84__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(n_majority7_module_84__and_module_3_res) );
  OR2_X1 u_majority7_module_84__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_84__or_module_3_res)
         );
  AND2_X1 u_majority7_module_84__and_module_4_U1 ( .A1(
        n_majority7_module_84__and_module_2_res), .A2(
        n_majority7_module_84__and_module_1_res), .ZN(
        n_majority7_module_84__and_module_4_res) );
  OR2_X1 u_majority7_module_84__or_module_4_U1 ( .A1(
        n_majority7_module_84__and_module_1_res), .A2(
        n_majority7_module_84__and_module_2_res), .ZN(
        n_majority7_module_84__or_module_4_res) );
  AND2_X1 u_majority7_module_84__and_module_5_U1 ( .A1(
        n_majority7_module_84__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_84__and_module_5_res) );
  OR2_X1 u_majority7_module_84__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_84__and_module_3_res), .ZN(
        n_majority7_module_84__or_module_5_res) );
  AND2_X1 u_majority7_module_84__and_module_6_U1 ( .A1(
        n_majority7_module_84__or_module_1_res), .A2(
        n_majority7_module_84__or_module_2_res), .ZN(
        n_majority7_module_84__and_module_6_res) );
  OR2_X1 u_majority7_module_84__or_module_6_U1 ( .A1(
        n_majority7_module_84__or_module_2_res), .A2(
        n_majority7_module_84__or_module_1_res), .ZN(
        n_majority7_module_84__or_module_6_res) );
  OR2_X1 u_majority7_module_84__or_module_7_U1 ( .A1(
        n_majority7_module_84__and_module_4_res), .A2(
        n_majority7_module_84__and_module_5_res), .ZN(
        n_majority7_module_84__or_module_7_res) );
  AND2_X1 u_majority7_module_84__and_module_7_U1 ( .A1(
        n_majority7_module_84__or_module_3_res), .A2(
        n_majority7_module_84__or_module_4_res), .ZN(
        n_majority7_module_84__and_module_7_res) );
  OR2_X1 u_majority7_module_84__or_module_8_U1 ( .A1(
        n_majority7_module_84__or_module_4_res), .A2(
        n_majority7_module_84__or_module_3_res), .ZN(
        n_majority7_module_84__or_module_8_res) );
  AND2_X1 u_majority7_module_84__and_module_8_U1 ( .A1(
        n_majority7_module_84__or_module_5_res), .A2(
        n_majority7_module_84__and_module_6_res), .ZN(
        n_majority7_module_84__and_module_8_res) );
  OR2_X1 u_majority7_module_84__or_module_9_U1 ( .A1(
        n_majority7_module_84__and_module_6_res), .A2(
        n_majority7_module_84__or_module_5_res), .ZN(
        n_majority7_module_84__or_module_9_res) );
  OR2_X1 u_majority7_module_84__or_module_10_U1 ( .A1(
        n_majority7_module_84__or_module_7_res), .A2(
        n_majority7_module_84__and_module_7_res), .ZN(
        n_majority7_module_84__or_module_10_res) );
  AND2_X1 u_majority7_module_84__and_module_9_U1 ( .A1(
        n_majority7_module_84__or_module_6_res), .A2(
        n_majority7_module_84__or_module_9_res), .ZN(
        n_majority7_module_84__and_module_9_res) );
  OR2_X1 u_majority7_module_84__or_module_11_U1 ( .A1(
        n_majority7_module_84__or_module_10_res), .A2(
        n_majority7_module_84__and_module_8_res), .ZN(
        n_majority7_module_84__or_module_11_res) );
  AND2_X1 u_majority7_module_84__and_module_10_U1 ( .A1(
        n_majority7_module_84__or_module_8_res), .A2(
        n_majority7_module_84__and_module_9_res), .ZN(
        n_majority7_module_84__and_module_10_res) );
  AND2_X1 u_majority7_module_84__and_module_11_U1 ( .A1(
        n_majority7_module_84__and_module_10_res), .A2(
        n_majority7_module_84__or_module_11_res), .ZN(
        n_majority7_module_84_res) );
  DFF_X1 u_reg_module_104__cini_mul_v00_reg ( .D(n_majority7_module_84_res), 
        .CK(clock_4), .Q(n_reg_module_104_res), .QN() );
  AND2_X1 u_majority7_module_85__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_85__and_module_1_res)
         );
  OR2_X1 u_majority7_module_85__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_85__or_module_1_res)
         );
  AND2_X1 u_majority7_module_85__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(n_majority7_module_85__and_module_2_res) );
  OR2_X1 u_majority7_module_85__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_85__or_module_2_res)
         );
  AND2_X1 u_majority7_module_85__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(n_majority7_module_85__and_module_3_res) );
  OR2_X1 u_majority7_module_85__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_85__or_module_3_res)
         );
  AND2_X1 u_majority7_module_85__and_module_4_U1 ( .A1(
        n_majority7_module_85__and_module_2_res), .A2(
        n_majority7_module_85__and_module_1_res), .ZN(
        n_majority7_module_85__and_module_4_res) );
  OR2_X1 u_majority7_module_85__or_module_4_U1 ( .A1(
        n_majority7_module_85__and_module_1_res), .A2(
        n_majority7_module_85__and_module_2_res), .ZN(
        n_majority7_module_85__or_module_4_res) );
  AND2_X1 u_majority7_module_85__and_module_5_U1 ( .A1(
        n_majority7_module_85__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_85__and_module_5_res) );
  OR2_X1 u_majority7_module_85__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_85__and_module_3_res), .ZN(
        n_majority7_module_85__or_module_5_res) );
  AND2_X1 u_majority7_module_85__and_module_6_U1 ( .A1(
        n_majority7_module_85__or_module_1_res), .A2(
        n_majority7_module_85__or_module_2_res), .ZN(
        n_majority7_module_85__and_module_6_res) );
  OR2_X1 u_majority7_module_85__or_module_6_U1 ( .A1(
        n_majority7_module_85__or_module_2_res), .A2(
        n_majority7_module_85__or_module_1_res), .ZN(
        n_majority7_module_85__or_module_6_res) );
  OR2_X1 u_majority7_module_85__or_module_7_U1 ( .A1(
        n_majority7_module_85__and_module_4_res), .A2(
        n_majority7_module_85__and_module_5_res), .ZN(
        n_majority7_module_85__or_module_7_res) );
  AND2_X1 u_majority7_module_85__and_module_7_U1 ( .A1(
        n_majority7_module_85__or_module_3_res), .A2(
        n_majority7_module_85__or_module_4_res), .ZN(
        n_majority7_module_85__and_module_7_res) );
  OR2_X1 u_majority7_module_85__or_module_8_U1 ( .A1(
        n_majority7_module_85__or_module_4_res), .A2(
        n_majority7_module_85__or_module_3_res), .ZN(
        n_majority7_module_85__or_module_8_res) );
  AND2_X1 u_majority7_module_85__and_module_8_U1 ( .A1(
        n_majority7_module_85__or_module_5_res), .A2(
        n_majority7_module_85__and_module_6_res), .ZN(
        n_majority7_module_85__and_module_8_res) );
  OR2_X1 u_majority7_module_85__or_module_9_U1 ( .A1(
        n_majority7_module_85__and_module_6_res), .A2(
        n_majority7_module_85__or_module_5_res), .ZN(
        n_majority7_module_85__or_module_9_res) );
  OR2_X1 u_majority7_module_85__or_module_10_U1 ( .A1(
        n_majority7_module_85__or_module_7_res), .A2(
        n_majority7_module_85__and_module_7_res), .ZN(
        n_majority7_module_85__or_module_10_res) );
  AND2_X1 u_majority7_module_85__and_module_9_U1 ( .A1(
        n_majority7_module_85__or_module_6_res), .A2(
        n_majority7_module_85__or_module_9_res), .ZN(
        n_majority7_module_85__and_module_9_res) );
  OR2_X1 u_majority7_module_85__or_module_11_U1 ( .A1(
        n_majority7_module_85__or_module_10_res), .A2(
        n_majority7_module_85__and_module_8_res), .ZN(
        n_majority7_module_85__or_module_11_res) );
  AND2_X1 u_majority7_module_85__and_module_10_U1 ( .A1(
        n_majority7_module_85__or_module_8_res), .A2(
        n_majority7_module_85__and_module_9_res), .ZN(
        n_majority7_module_85__and_module_10_res) );
  AND2_X1 u_majority7_module_85__and_module_11_U1 ( .A1(
        n_majority7_module_85__and_module_10_res), .A2(
        n_majority7_module_85__or_module_11_res), .ZN(
        n_majority7_module_85_res) );
  DFF_X1 u_reg_module_105__cini_mul_v00_reg ( .D(n_majority7_module_85_res), 
        .CK(clock_4), .Q(n_reg_module_105_res), .QN() );
  AND2_X1 u_majority7_module_86__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_86__and_module_1_res)
         );
  OR2_X1 u_majority7_module_86__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_86__or_module_1_res)
         );
  AND2_X1 u_majority7_module_86__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(n_majority7_module_86__and_module_2_res) );
  OR2_X1 u_majority7_module_86__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_86__or_module_2_res)
         );
  AND2_X1 u_majority7_module_86__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(n_majority7_module_86__and_module_3_res) );
  OR2_X1 u_majority7_module_86__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_86__or_module_3_res)
         );
  AND2_X1 u_majority7_module_86__and_module_4_U1 ( .A1(
        n_majority7_module_86__and_module_2_res), .A2(
        n_majority7_module_86__and_module_1_res), .ZN(
        n_majority7_module_86__and_module_4_res) );
  OR2_X1 u_majority7_module_86__or_module_4_U1 ( .A1(
        n_majority7_module_86__and_module_1_res), .A2(
        n_majority7_module_86__and_module_2_res), .ZN(
        n_majority7_module_86__or_module_4_res) );
  AND2_X1 u_majority7_module_86__and_module_5_U1 ( .A1(
        n_majority7_module_86__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_86__and_module_5_res) );
  OR2_X1 u_majority7_module_86__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_86__and_module_3_res), .ZN(
        n_majority7_module_86__or_module_5_res) );
  AND2_X1 u_majority7_module_86__and_module_6_U1 ( .A1(
        n_majority7_module_86__or_module_1_res), .A2(
        n_majority7_module_86__or_module_2_res), .ZN(
        n_majority7_module_86__and_module_6_res) );
  OR2_X1 u_majority7_module_86__or_module_6_U1 ( .A1(
        n_majority7_module_86__or_module_2_res), .A2(
        n_majority7_module_86__or_module_1_res), .ZN(
        n_majority7_module_86__or_module_6_res) );
  OR2_X1 u_majority7_module_86__or_module_7_U1 ( .A1(
        n_majority7_module_86__and_module_4_res), .A2(
        n_majority7_module_86__and_module_5_res), .ZN(
        n_majority7_module_86__or_module_7_res) );
  AND2_X1 u_majority7_module_86__and_module_7_U1 ( .A1(
        n_majority7_module_86__or_module_3_res), .A2(
        n_majority7_module_86__or_module_4_res), .ZN(
        n_majority7_module_86__and_module_7_res) );
  OR2_X1 u_majority7_module_86__or_module_8_U1 ( .A1(
        n_majority7_module_86__or_module_4_res), .A2(
        n_majority7_module_86__or_module_3_res), .ZN(
        n_majority7_module_86__or_module_8_res) );
  AND2_X1 u_majority7_module_86__and_module_8_U1 ( .A1(
        n_majority7_module_86__or_module_5_res), .A2(
        n_majority7_module_86__and_module_6_res), .ZN(
        n_majority7_module_86__and_module_8_res) );
  OR2_X1 u_majority7_module_86__or_module_9_U1 ( .A1(
        n_majority7_module_86__and_module_6_res), .A2(
        n_majority7_module_86__or_module_5_res), .ZN(
        n_majority7_module_86__or_module_9_res) );
  OR2_X1 u_majority7_module_86__or_module_10_U1 ( .A1(
        n_majority7_module_86__or_module_7_res), .A2(
        n_majority7_module_86__and_module_7_res), .ZN(
        n_majority7_module_86__or_module_10_res) );
  AND2_X1 u_majority7_module_86__and_module_9_U1 ( .A1(
        n_majority7_module_86__or_module_6_res), .A2(
        n_majority7_module_86__or_module_9_res), .ZN(
        n_majority7_module_86__and_module_9_res) );
  OR2_X1 u_majority7_module_86__or_module_11_U1 ( .A1(
        n_majority7_module_86__or_module_10_res), .A2(
        n_majority7_module_86__and_module_8_res), .ZN(
        n_majority7_module_86__or_module_11_res) );
  AND2_X1 u_majority7_module_86__and_module_10_U1 ( .A1(
        n_majority7_module_86__or_module_8_res), .A2(
        n_majority7_module_86__and_module_9_res), .ZN(
        n_majority7_module_86__and_module_10_res) );
  AND2_X1 u_majority7_module_86__and_module_11_U1 ( .A1(
        n_majority7_module_86__and_module_10_res), .A2(
        n_majority7_module_86__or_module_11_res), .ZN(
        n_majority7_module_86_res) );
  DFF_X1 u_reg_module_106__cini_mul_v00_reg ( .D(n_majority7_module_86_res), 
        .CK(clock_4), .Q(n_reg_module_106_res), .QN() );
  AND2_X1 u_majority7_module_87__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_87__and_module_1_res)
         );
  OR2_X1 u_majority7_module_87__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_87__or_module_1_res)
         );
  AND2_X1 u_majority7_module_87__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(n_majority7_module_87__and_module_2_res) );
  OR2_X1 u_majority7_module_87__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_87__or_module_2_res)
         );
  AND2_X1 u_majority7_module_87__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(n_majority7_module_87__and_module_3_res) );
  OR2_X1 u_majority7_module_87__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_87__or_module_3_res)
         );
  AND2_X1 u_majority7_module_87__and_module_4_U1 ( .A1(
        n_majority7_module_87__and_module_2_res), .A2(
        n_majority7_module_87__and_module_1_res), .ZN(
        n_majority7_module_87__and_module_4_res) );
  OR2_X1 u_majority7_module_87__or_module_4_U1 ( .A1(
        n_majority7_module_87__and_module_1_res), .A2(
        n_majority7_module_87__and_module_2_res), .ZN(
        n_majority7_module_87__or_module_4_res) );
  AND2_X1 u_majority7_module_87__and_module_5_U1 ( .A1(
        n_majority7_module_87__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_87__and_module_5_res) );
  OR2_X1 u_majority7_module_87__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_87__and_module_3_res), .ZN(
        n_majority7_module_87__or_module_5_res) );
  AND2_X1 u_majority7_module_87__and_module_6_U1 ( .A1(
        n_majority7_module_87__or_module_1_res), .A2(
        n_majority7_module_87__or_module_2_res), .ZN(
        n_majority7_module_87__and_module_6_res) );
  OR2_X1 u_majority7_module_87__or_module_6_U1 ( .A1(
        n_majority7_module_87__or_module_2_res), .A2(
        n_majority7_module_87__or_module_1_res), .ZN(
        n_majority7_module_87__or_module_6_res) );
  OR2_X1 u_majority7_module_87__or_module_7_U1 ( .A1(
        n_majority7_module_87__and_module_4_res), .A2(
        n_majority7_module_87__and_module_5_res), .ZN(
        n_majority7_module_87__or_module_7_res) );
  AND2_X1 u_majority7_module_87__and_module_7_U1 ( .A1(
        n_majority7_module_87__or_module_3_res), .A2(
        n_majority7_module_87__or_module_4_res), .ZN(
        n_majority7_module_87__and_module_7_res) );
  OR2_X1 u_majority7_module_87__or_module_8_U1 ( .A1(
        n_majority7_module_87__or_module_4_res), .A2(
        n_majority7_module_87__or_module_3_res), .ZN(
        n_majority7_module_87__or_module_8_res) );
  AND2_X1 u_majority7_module_87__and_module_8_U1 ( .A1(
        n_majority7_module_87__or_module_5_res), .A2(
        n_majority7_module_87__and_module_6_res), .ZN(
        n_majority7_module_87__and_module_8_res) );
  OR2_X1 u_majority7_module_87__or_module_9_U1 ( .A1(
        n_majority7_module_87__and_module_6_res), .A2(
        n_majority7_module_87__or_module_5_res), .ZN(
        n_majority7_module_87__or_module_9_res) );
  OR2_X1 u_majority7_module_87__or_module_10_U1 ( .A1(
        n_majority7_module_87__or_module_7_res), .A2(
        n_majority7_module_87__and_module_7_res), .ZN(
        n_majority7_module_87__or_module_10_res) );
  AND2_X1 u_majority7_module_87__and_module_9_U1 ( .A1(
        n_majority7_module_87__or_module_6_res), .A2(
        n_majority7_module_87__or_module_9_res), .ZN(
        n_majority7_module_87__and_module_9_res) );
  OR2_X1 u_majority7_module_87__or_module_11_U1 ( .A1(
        n_majority7_module_87__or_module_10_res), .A2(
        n_majority7_module_87__and_module_8_res), .ZN(
        n_majority7_module_87__or_module_11_res) );
  AND2_X1 u_majority7_module_87__and_module_10_U1 ( .A1(
        n_majority7_module_87__or_module_8_res), .A2(
        n_majority7_module_87__and_module_9_res), .ZN(
        n_majority7_module_87__and_module_10_res) );
  AND2_X1 u_majority7_module_87__and_module_11_U1 ( .A1(
        n_majority7_module_87__and_module_10_res), .A2(
        n_majority7_module_87__or_module_11_res), .ZN(
        n_majority7_module_87_res) );
  DFF_X1 u_reg_module_107__cini_mul_v00_reg ( .D(n_majority7_module_87_res), 
        .CK(clock_4), .Q(n_reg_module_107_res), .QN() );
  DFF_X1 u_reg_module_108__cini_mul_v00_reg ( .D(n_and_module_80_res), .CK(
        clock_4), .Q(n_reg_module_108_res), .QN() );
  DFF_X1 u_reg_module_109__cini_mul_v00_reg ( .D(n_and_module_81_res), .CK(
        clock_5), .Q(n_reg_module_109_res), .QN() );
  AND2_X1 u_majority7_module_88__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_88__and_module_1_res)
         );
  OR2_X1 u_majority7_module_88__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_88__or_module_1_res)
         );
  AND2_X1 u_majority7_module_88__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(n_majority7_module_88__and_module_2_res) );
  OR2_X1 u_majority7_module_88__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_88__or_module_2_res)
         );
  AND2_X1 u_majority7_module_88__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(n_majority7_module_88__and_module_3_res) );
  OR2_X1 u_majority7_module_88__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_88__or_module_3_res)
         );
  AND2_X1 u_majority7_module_88__and_module_4_U1 ( .A1(
        n_majority7_module_88__and_module_2_res), .A2(
        n_majority7_module_88__and_module_1_res), .ZN(
        n_majority7_module_88__and_module_4_res) );
  OR2_X1 u_majority7_module_88__or_module_4_U1 ( .A1(
        n_majority7_module_88__and_module_1_res), .A2(
        n_majority7_module_88__and_module_2_res), .ZN(
        n_majority7_module_88__or_module_4_res) );
  AND2_X1 u_majority7_module_88__and_module_5_U1 ( .A1(
        n_majority7_module_88__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_88__and_module_5_res) );
  OR2_X1 u_majority7_module_88__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_88__and_module_3_res), .ZN(
        n_majority7_module_88__or_module_5_res) );
  AND2_X1 u_majority7_module_88__and_module_6_U1 ( .A1(
        n_majority7_module_88__or_module_1_res), .A2(
        n_majority7_module_88__or_module_2_res), .ZN(
        n_majority7_module_88__and_module_6_res) );
  OR2_X1 u_majority7_module_88__or_module_6_U1 ( .A1(
        n_majority7_module_88__or_module_2_res), .A2(
        n_majority7_module_88__or_module_1_res), .ZN(
        n_majority7_module_88__or_module_6_res) );
  OR2_X1 u_majority7_module_88__or_module_7_U1 ( .A1(
        n_majority7_module_88__and_module_4_res), .A2(
        n_majority7_module_88__and_module_5_res), .ZN(
        n_majority7_module_88__or_module_7_res) );
  AND2_X1 u_majority7_module_88__and_module_7_U1 ( .A1(
        n_majority7_module_88__or_module_3_res), .A2(
        n_majority7_module_88__or_module_4_res), .ZN(
        n_majority7_module_88__and_module_7_res) );
  OR2_X1 u_majority7_module_88__or_module_8_U1 ( .A1(
        n_majority7_module_88__or_module_4_res), .A2(
        n_majority7_module_88__or_module_3_res), .ZN(
        n_majority7_module_88__or_module_8_res) );
  AND2_X1 u_majority7_module_88__and_module_8_U1 ( .A1(
        n_majority7_module_88__or_module_5_res), .A2(
        n_majority7_module_88__and_module_6_res), .ZN(
        n_majority7_module_88__and_module_8_res) );
  OR2_X1 u_majority7_module_88__or_module_9_U1 ( .A1(
        n_majority7_module_88__and_module_6_res), .A2(
        n_majority7_module_88__or_module_5_res), .ZN(
        n_majority7_module_88__or_module_9_res) );
  OR2_X1 u_majority7_module_88__or_module_10_U1 ( .A1(
        n_majority7_module_88__or_module_7_res), .A2(
        n_majority7_module_88__and_module_7_res), .ZN(
        n_majority7_module_88__or_module_10_res) );
  AND2_X1 u_majority7_module_88__and_module_9_U1 ( .A1(
        n_majority7_module_88__or_module_6_res), .A2(
        n_majority7_module_88__or_module_9_res), .ZN(
        n_majority7_module_88__and_module_9_res) );
  OR2_X1 u_majority7_module_88__or_module_11_U1 ( .A1(
        n_majority7_module_88__or_module_10_res), .A2(
        n_majority7_module_88__and_module_8_res), .ZN(
        n_majority7_module_88__or_module_11_res) );
  AND2_X1 u_majority7_module_88__and_module_10_U1 ( .A1(
        n_majority7_module_88__or_module_8_res), .A2(
        n_majority7_module_88__and_module_9_res), .ZN(
        n_majority7_module_88__and_module_10_res) );
  AND2_X1 u_majority7_module_88__and_module_11_U1 ( .A1(
        n_majority7_module_88__and_module_10_res), .A2(
        n_majority7_module_88__or_module_11_res), .ZN(
        n_majority7_module_88_res) );
  DFF_X1 u_reg_module_110__cini_mul_v00_reg ( .D(n_majority7_module_88_res), 
        .CK(clock_5), .Q(n_reg_module_110_res), .QN() );
  AND2_X1 u_majority7_module_89__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_89__and_module_1_res)
         );
  OR2_X1 u_majority7_module_89__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_89__or_module_1_res)
         );
  AND2_X1 u_majority7_module_89__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(n_majority7_module_89__and_module_2_res) );
  OR2_X1 u_majority7_module_89__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_89__or_module_2_res)
         );
  AND2_X1 u_majority7_module_89__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(n_majority7_module_89__and_module_3_res) );
  OR2_X1 u_majority7_module_89__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_89__or_module_3_res)
         );
  AND2_X1 u_majority7_module_89__and_module_4_U1 ( .A1(
        n_majority7_module_89__and_module_2_res), .A2(
        n_majority7_module_89__and_module_1_res), .ZN(
        n_majority7_module_89__and_module_4_res) );
  OR2_X1 u_majority7_module_89__or_module_4_U1 ( .A1(
        n_majority7_module_89__and_module_1_res), .A2(
        n_majority7_module_89__and_module_2_res), .ZN(
        n_majority7_module_89__or_module_4_res) );
  AND2_X1 u_majority7_module_89__and_module_5_U1 ( .A1(
        n_majority7_module_89__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_89__and_module_5_res) );
  OR2_X1 u_majority7_module_89__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_89__and_module_3_res), .ZN(
        n_majority7_module_89__or_module_5_res) );
  AND2_X1 u_majority7_module_89__and_module_6_U1 ( .A1(
        n_majority7_module_89__or_module_1_res), .A2(
        n_majority7_module_89__or_module_2_res), .ZN(
        n_majority7_module_89__and_module_6_res) );
  OR2_X1 u_majority7_module_89__or_module_6_U1 ( .A1(
        n_majority7_module_89__or_module_2_res), .A2(
        n_majority7_module_89__or_module_1_res), .ZN(
        n_majority7_module_89__or_module_6_res) );
  OR2_X1 u_majority7_module_89__or_module_7_U1 ( .A1(
        n_majority7_module_89__and_module_4_res), .A2(
        n_majority7_module_89__and_module_5_res), .ZN(
        n_majority7_module_89__or_module_7_res) );
  AND2_X1 u_majority7_module_89__and_module_7_U1 ( .A1(
        n_majority7_module_89__or_module_3_res), .A2(
        n_majority7_module_89__or_module_4_res), .ZN(
        n_majority7_module_89__and_module_7_res) );
  OR2_X1 u_majority7_module_89__or_module_8_U1 ( .A1(
        n_majority7_module_89__or_module_4_res), .A2(
        n_majority7_module_89__or_module_3_res), .ZN(
        n_majority7_module_89__or_module_8_res) );
  AND2_X1 u_majority7_module_89__and_module_8_U1 ( .A1(
        n_majority7_module_89__or_module_5_res), .A2(
        n_majority7_module_89__and_module_6_res), .ZN(
        n_majority7_module_89__and_module_8_res) );
  OR2_X1 u_majority7_module_89__or_module_9_U1 ( .A1(
        n_majority7_module_89__and_module_6_res), .A2(
        n_majority7_module_89__or_module_5_res), .ZN(
        n_majority7_module_89__or_module_9_res) );
  OR2_X1 u_majority7_module_89__or_module_10_U1 ( .A1(
        n_majority7_module_89__or_module_7_res), .A2(
        n_majority7_module_89__and_module_7_res), .ZN(
        n_majority7_module_89__or_module_10_res) );
  AND2_X1 u_majority7_module_89__and_module_9_U1 ( .A1(
        n_majority7_module_89__or_module_6_res), .A2(
        n_majority7_module_89__or_module_9_res), .ZN(
        n_majority7_module_89__and_module_9_res) );
  OR2_X1 u_majority7_module_89__or_module_11_U1 ( .A1(
        n_majority7_module_89__or_module_10_res), .A2(
        n_majority7_module_89__and_module_8_res), .ZN(
        n_majority7_module_89__or_module_11_res) );
  AND2_X1 u_majority7_module_89__and_module_10_U1 ( .A1(
        n_majority7_module_89__or_module_8_res), .A2(
        n_majority7_module_89__and_module_9_res), .ZN(
        n_majority7_module_89__and_module_10_res) );
  AND2_X1 u_majority7_module_89__and_module_11_U1 ( .A1(
        n_majority7_module_89__and_module_10_res), .A2(
        n_majority7_module_89__or_module_11_res), .ZN(
        n_majority7_module_89_res) );
  DFF_X1 u_reg_module_111__cini_mul_v00_reg ( .D(n_majority7_module_89_res), 
        .CK(clock_5), .Q(n_reg_module_111_res), .QN() );
  AND2_X1 u_majority7_module_90__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_90__and_module_1_res)
         );
  OR2_X1 u_majority7_module_90__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_90__or_module_1_res)
         );
  AND2_X1 u_majority7_module_90__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(n_majority7_module_90__and_module_2_res) );
  OR2_X1 u_majority7_module_90__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_90__or_module_2_res)
         );
  AND2_X1 u_majority7_module_90__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(n_majority7_module_90__and_module_3_res) );
  OR2_X1 u_majority7_module_90__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_90__or_module_3_res)
         );
  AND2_X1 u_majority7_module_90__and_module_4_U1 ( .A1(
        n_majority7_module_90__and_module_2_res), .A2(
        n_majority7_module_90__and_module_1_res), .ZN(
        n_majority7_module_90__and_module_4_res) );
  OR2_X1 u_majority7_module_90__or_module_4_U1 ( .A1(
        n_majority7_module_90__and_module_1_res), .A2(
        n_majority7_module_90__and_module_2_res), .ZN(
        n_majority7_module_90__or_module_4_res) );
  AND2_X1 u_majority7_module_90__and_module_5_U1 ( .A1(
        n_majority7_module_90__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_90__and_module_5_res) );
  OR2_X1 u_majority7_module_90__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_90__and_module_3_res), .ZN(
        n_majority7_module_90__or_module_5_res) );
  AND2_X1 u_majority7_module_90__and_module_6_U1 ( .A1(
        n_majority7_module_90__or_module_1_res), .A2(
        n_majority7_module_90__or_module_2_res), .ZN(
        n_majority7_module_90__and_module_6_res) );
  OR2_X1 u_majority7_module_90__or_module_6_U1 ( .A1(
        n_majority7_module_90__or_module_2_res), .A2(
        n_majority7_module_90__or_module_1_res), .ZN(
        n_majority7_module_90__or_module_6_res) );
  OR2_X1 u_majority7_module_90__or_module_7_U1 ( .A1(
        n_majority7_module_90__and_module_4_res), .A2(
        n_majority7_module_90__and_module_5_res), .ZN(
        n_majority7_module_90__or_module_7_res) );
  AND2_X1 u_majority7_module_90__and_module_7_U1 ( .A1(
        n_majority7_module_90__or_module_3_res), .A2(
        n_majority7_module_90__or_module_4_res), .ZN(
        n_majority7_module_90__and_module_7_res) );
  OR2_X1 u_majority7_module_90__or_module_8_U1 ( .A1(
        n_majority7_module_90__or_module_4_res), .A2(
        n_majority7_module_90__or_module_3_res), .ZN(
        n_majority7_module_90__or_module_8_res) );
  AND2_X1 u_majority7_module_90__and_module_8_U1 ( .A1(
        n_majority7_module_90__or_module_5_res), .A2(
        n_majority7_module_90__and_module_6_res), .ZN(
        n_majority7_module_90__and_module_8_res) );
  OR2_X1 u_majority7_module_90__or_module_9_U1 ( .A1(
        n_majority7_module_90__and_module_6_res), .A2(
        n_majority7_module_90__or_module_5_res), .ZN(
        n_majority7_module_90__or_module_9_res) );
  OR2_X1 u_majority7_module_90__or_module_10_U1 ( .A1(
        n_majority7_module_90__or_module_7_res), .A2(
        n_majority7_module_90__and_module_7_res), .ZN(
        n_majority7_module_90__or_module_10_res) );
  AND2_X1 u_majority7_module_90__and_module_9_U1 ( .A1(
        n_majority7_module_90__or_module_6_res), .A2(
        n_majority7_module_90__or_module_9_res), .ZN(
        n_majority7_module_90__and_module_9_res) );
  OR2_X1 u_majority7_module_90__or_module_11_U1 ( .A1(
        n_majority7_module_90__or_module_10_res), .A2(
        n_majority7_module_90__and_module_8_res), .ZN(
        n_majority7_module_90__or_module_11_res) );
  AND2_X1 u_majority7_module_90__and_module_10_U1 ( .A1(
        n_majority7_module_90__or_module_8_res), .A2(
        n_majority7_module_90__and_module_9_res), .ZN(
        n_majority7_module_90__and_module_10_res) );
  AND2_X1 u_majority7_module_90__and_module_11_U1 ( .A1(
        n_majority7_module_90__and_module_10_res), .A2(
        n_majority7_module_90__or_module_11_res), .ZN(
        n_majority7_module_90_res) );
  DFF_X1 u_reg_module_112__cini_mul_v00_reg ( .D(n_majority7_module_90_res), 
        .CK(clock_5), .Q(n_reg_module_112_res), .QN() );
  AND2_X1 u_majority7_module_91__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_91__and_module_1_res)
         );
  OR2_X1 u_majority7_module_91__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_91__or_module_1_res)
         );
  AND2_X1 u_majority7_module_91__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(n_majority7_module_91__and_module_2_res) );
  OR2_X1 u_majority7_module_91__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_91__or_module_2_res)
         );
  AND2_X1 u_majority7_module_91__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(n_majority7_module_91__and_module_3_res) );
  OR2_X1 u_majority7_module_91__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_91__or_module_3_res)
         );
  AND2_X1 u_majority7_module_91__and_module_4_U1 ( .A1(
        n_majority7_module_91__and_module_2_res), .A2(
        n_majority7_module_91__and_module_1_res), .ZN(
        n_majority7_module_91__and_module_4_res) );
  OR2_X1 u_majority7_module_91__or_module_4_U1 ( .A1(
        n_majority7_module_91__and_module_1_res), .A2(
        n_majority7_module_91__and_module_2_res), .ZN(
        n_majority7_module_91__or_module_4_res) );
  AND2_X1 u_majority7_module_91__and_module_5_U1 ( .A1(
        n_majority7_module_91__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_91__and_module_5_res) );
  OR2_X1 u_majority7_module_91__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_91__and_module_3_res), .ZN(
        n_majority7_module_91__or_module_5_res) );
  AND2_X1 u_majority7_module_91__and_module_6_U1 ( .A1(
        n_majority7_module_91__or_module_1_res), .A2(
        n_majority7_module_91__or_module_2_res), .ZN(
        n_majority7_module_91__and_module_6_res) );
  OR2_X1 u_majority7_module_91__or_module_6_U1 ( .A1(
        n_majority7_module_91__or_module_2_res), .A2(
        n_majority7_module_91__or_module_1_res), .ZN(
        n_majority7_module_91__or_module_6_res) );
  OR2_X1 u_majority7_module_91__or_module_7_U1 ( .A1(
        n_majority7_module_91__and_module_4_res), .A2(
        n_majority7_module_91__and_module_5_res), .ZN(
        n_majority7_module_91__or_module_7_res) );
  AND2_X1 u_majority7_module_91__and_module_7_U1 ( .A1(
        n_majority7_module_91__or_module_3_res), .A2(
        n_majority7_module_91__or_module_4_res), .ZN(
        n_majority7_module_91__and_module_7_res) );
  OR2_X1 u_majority7_module_91__or_module_8_U1 ( .A1(
        n_majority7_module_91__or_module_4_res), .A2(
        n_majority7_module_91__or_module_3_res), .ZN(
        n_majority7_module_91__or_module_8_res) );
  AND2_X1 u_majority7_module_91__and_module_8_U1 ( .A1(
        n_majority7_module_91__or_module_5_res), .A2(
        n_majority7_module_91__and_module_6_res), .ZN(
        n_majority7_module_91__and_module_8_res) );
  OR2_X1 u_majority7_module_91__or_module_9_U1 ( .A1(
        n_majority7_module_91__and_module_6_res), .A2(
        n_majority7_module_91__or_module_5_res), .ZN(
        n_majority7_module_91__or_module_9_res) );
  OR2_X1 u_majority7_module_91__or_module_10_U1 ( .A1(
        n_majority7_module_91__or_module_7_res), .A2(
        n_majority7_module_91__and_module_7_res), .ZN(
        n_majority7_module_91__or_module_10_res) );
  AND2_X1 u_majority7_module_91__and_module_9_U1 ( .A1(
        n_majority7_module_91__or_module_6_res), .A2(
        n_majority7_module_91__or_module_9_res), .ZN(
        n_majority7_module_91__and_module_9_res) );
  OR2_X1 u_majority7_module_91__or_module_11_U1 ( .A1(
        n_majority7_module_91__or_module_10_res), .A2(
        n_majority7_module_91__and_module_8_res), .ZN(
        n_majority7_module_91__or_module_11_res) );
  AND2_X1 u_majority7_module_91__and_module_10_U1 ( .A1(
        n_majority7_module_91__or_module_8_res), .A2(
        n_majority7_module_91__and_module_9_res), .ZN(
        n_majority7_module_91__and_module_10_res) );
  AND2_X1 u_majority7_module_91__and_module_11_U1 ( .A1(
        n_majority7_module_91__and_module_10_res), .A2(
        n_majority7_module_91__or_module_11_res), .ZN(
        n_majority7_module_91_res) );
  DFF_X1 u_reg_module_113__cini_mul_v00_reg ( .D(n_majority7_module_91_res), 
        .CK(clock_5), .Q(n_reg_module_113_res), .QN() );
  DFF_X1 u_reg_module_114__cini_mul_v00_reg ( .D(n_and_module_86_res), .CK(
        clock_5), .Q(n_reg_module_114_res), .QN() );
  AND2_X1 u_majority7_module_92__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_92__and_module_1_res)
         );
  OR2_X1 u_majority7_module_92__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_92__or_module_1_res)
         );
  AND2_X1 u_majority7_module_92__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(n_majority7_module_92__and_module_2_res) );
  OR2_X1 u_majority7_module_92__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_92__or_module_2_res)
         );
  AND2_X1 u_majority7_module_92__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(n_majority7_module_92__and_module_3_res) );
  OR2_X1 u_majority7_module_92__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_92__or_module_3_res)
         );
  AND2_X1 u_majority7_module_92__and_module_4_U1 ( .A1(
        n_majority7_module_92__and_module_2_res), .A2(
        n_majority7_module_92__and_module_1_res), .ZN(
        n_majority7_module_92__and_module_4_res) );
  OR2_X1 u_majority7_module_92__or_module_4_U1 ( .A1(
        n_majority7_module_92__and_module_1_res), .A2(
        n_majority7_module_92__and_module_2_res), .ZN(
        n_majority7_module_92__or_module_4_res) );
  AND2_X1 u_majority7_module_92__and_module_5_U1 ( .A1(
        n_majority7_module_92__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_92__and_module_5_res) );
  OR2_X1 u_majority7_module_92__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_92__and_module_3_res), .ZN(
        n_majority7_module_92__or_module_5_res) );
  AND2_X1 u_majority7_module_92__and_module_6_U1 ( .A1(
        n_majority7_module_92__or_module_1_res), .A2(
        n_majority7_module_92__or_module_2_res), .ZN(
        n_majority7_module_92__and_module_6_res) );
  OR2_X1 u_majority7_module_92__or_module_6_U1 ( .A1(
        n_majority7_module_92__or_module_2_res), .A2(
        n_majority7_module_92__or_module_1_res), .ZN(
        n_majority7_module_92__or_module_6_res) );
  OR2_X1 u_majority7_module_92__or_module_7_U1 ( .A1(
        n_majority7_module_92__and_module_4_res), .A2(
        n_majority7_module_92__and_module_5_res), .ZN(
        n_majority7_module_92__or_module_7_res) );
  AND2_X1 u_majority7_module_92__and_module_7_U1 ( .A1(
        n_majority7_module_92__or_module_3_res), .A2(
        n_majority7_module_92__or_module_4_res), .ZN(
        n_majority7_module_92__and_module_7_res) );
  OR2_X1 u_majority7_module_92__or_module_8_U1 ( .A1(
        n_majority7_module_92__or_module_4_res), .A2(
        n_majority7_module_92__or_module_3_res), .ZN(
        n_majority7_module_92__or_module_8_res) );
  AND2_X1 u_majority7_module_92__and_module_8_U1 ( .A1(
        n_majority7_module_92__or_module_5_res), .A2(
        n_majority7_module_92__and_module_6_res), .ZN(
        n_majority7_module_92__and_module_8_res) );
  OR2_X1 u_majority7_module_92__or_module_9_U1 ( .A1(
        n_majority7_module_92__and_module_6_res), .A2(
        n_majority7_module_92__or_module_5_res), .ZN(
        n_majority7_module_92__or_module_9_res) );
  OR2_X1 u_majority7_module_92__or_module_10_U1 ( .A1(
        n_majority7_module_92__or_module_7_res), .A2(
        n_majority7_module_92__and_module_7_res), .ZN(
        n_majority7_module_92__or_module_10_res) );
  AND2_X1 u_majority7_module_92__and_module_9_U1 ( .A1(
        n_majority7_module_92__or_module_6_res), .A2(
        n_majority7_module_92__or_module_9_res), .ZN(
        n_majority7_module_92__and_module_9_res) );
  OR2_X1 u_majority7_module_92__or_module_11_U1 ( .A1(
        n_majority7_module_92__or_module_10_res), .A2(
        n_majority7_module_92__and_module_8_res), .ZN(
        n_majority7_module_92__or_module_11_res) );
  AND2_X1 u_majority7_module_92__and_module_10_U1 ( .A1(
        n_majority7_module_92__or_module_8_res), .A2(
        n_majority7_module_92__and_module_9_res), .ZN(
        n_majority7_module_92__and_module_10_res) );
  AND2_X1 u_majority7_module_92__and_module_11_U1 ( .A1(
        n_majority7_module_92__and_module_10_res), .A2(
        n_majority7_module_92__or_module_11_res), .ZN(
        n_majority7_module_92_res) );
  DFF_X1 u_reg_module_115__cini_mul_v00_reg ( .D(n_majority7_module_92_res), 
        .CK(clock_5), .Q(n_reg_module_115_res), .QN() );
  AND2_X1 u_majority7_module_93__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_93__and_module_1_res)
         );
  OR2_X1 u_majority7_module_93__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_93__or_module_1_res)
         );
  AND2_X1 u_majority7_module_93__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(n_majority7_module_93__and_module_2_res) );
  OR2_X1 u_majority7_module_93__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_93__or_module_2_res)
         );
  AND2_X1 u_majority7_module_93__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(n_majority7_module_93__and_module_3_res) );
  OR2_X1 u_majority7_module_93__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_93__or_module_3_res)
         );
  AND2_X1 u_majority7_module_93__and_module_4_U1 ( .A1(
        n_majority7_module_93__and_module_2_res), .A2(
        n_majority7_module_93__and_module_1_res), .ZN(
        n_majority7_module_93__and_module_4_res) );
  OR2_X1 u_majority7_module_93__or_module_4_U1 ( .A1(
        n_majority7_module_93__and_module_1_res), .A2(
        n_majority7_module_93__and_module_2_res), .ZN(
        n_majority7_module_93__or_module_4_res) );
  AND2_X1 u_majority7_module_93__and_module_5_U1 ( .A1(
        n_majority7_module_93__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_93__and_module_5_res) );
  OR2_X1 u_majority7_module_93__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_93__and_module_3_res), .ZN(
        n_majority7_module_93__or_module_5_res) );
  AND2_X1 u_majority7_module_93__and_module_6_U1 ( .A1(
        n_majority7_module_93__or_module_1_res), .A2(
        n_majority7_module_93__or_module_2_res), .ZN(
        n_majority7_module_93__and_module_6_res) );
  OR2_X1 u_majority7_module_93__or_module_6_U1 ( .A1(
        n_majority7_module_93__or_module_2_res), .A2(
        n_majority7_module_93__or_module_1_res), .ZN(
        n_majority7_module_93__or_module_6_res) );
  OR2_X1 u_majority7_module_93__or_module_7_U1 ( .A1(
        n_majority7_module_93__and_module_4_res), .A2(
        n_majority7_module_93__and_module_5_res), .ZN(
        n_majority7_module_93__or_module_7_res) );
  AND2_X1 u_majority7_module_93__and_module_7_U1 ( .A1(
        n_majority7_module_93__or_module_3_res), .A2(
        n_majority7_module_93__or_module_4_res), .ZN(
        n_majority7_module_93__and_module_7_res) );
  OR2_X1 u_majority7_module_93__or_module_8_U1 ( .A1(
        n_majority7_module_93__or_module_4_res), .A2(
        n_majority7_module_93__or_module_3_res), .ZN(
        n_majority7_module_93__or_module_8_res) );
  AND2_X1 u_majority7_module_93__and_module_8_U1 ( .A1(
        n_majority7_module_93__or_module_5_res), .A2(
        n_majority7_module_93__and_module_6_res), .ZN(
        n_majority7_module_93__and_module_8_res) );
  OR2_X1 u_majority7_module_93__or_module_9_U1 ( .A1(
        n_majority7_module_93__and_module_6_res), .A2(
        n_majority7_module_93__or_module_5_res), .ZN(
        n_majority7_module_93__or_module_9_res) );
  OR2_X1 u_majority7_module_93__or_module_10_U1 ( .A1(
        n_majority7_module_93__or_module_7_res), .A2(
        n_majority7_module_93__and_module_7_res), .ZN(
        n_majority7_module_93__or_module_10_res) );
  AND2_X1 u_majority7_module_93__and_module_9_U1 ( .A1(
        n_majority7_module_93__or_module_6_res), .A2(
        n_majority7_module_93__or_module_9_res), .ZN(
        n_majority7_module_93__and_module_9_res) );
  OR2_X1 u_majority7_module_93__or_module_11_U1 ( .A1(
        n_majority7_module_93__or_module_10_res), .A2(
        n_majority7_module_93__and_module_8_res), .ZN(
        n_majority7_module_93__or_module_11_res) );
  AND2_X1 u_majority7_module_93__and_module_10_U1 ( .A1(
        n_majority7_module_93__or_module_8_res), .A2(
        n_majority7_module_93__and_module_9_res), .ZN(
        n_majority7_module_93__and_module_10_res) );
  AND2_X1 u_majority7_module_93__and_module_11_U1 ( .A1(
        n_majority7_module_93__and_module_10_res), .A2(
        n_majority7_module_93__or_module_11_res), .ZN(
        n_majority7_module_93_res) );
  DFF_X1 u_reg_module_116__cini_mul_v00_reg ( .D(n_majority7_module_93_res), 
        .CK(clock_5), .Q(n_reg_module_116_res), .QN() );
  AND2_X1 u_majority7_module_94__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_94__and_module_1_res)
         );
  OR2_X1 u_majority7_module_94__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_94__or_module_1_res)
         );
  AND2_X1 u_majority7_module_94__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(n_majority7_module_94__and_module_2_res) );
  OR2_X1 u_majority7_module_94__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_94__or_module_2_res)
         );
  AND2_X1 u_majority7_module_94__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(n_majority7_module_94__and_module_3_res) );
  OR2_X1 u_majority7_module_94__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_94__or_module_3_res)
         );
  AND2_X1 u_majority7_module_94__and_module_4_U1 ( .A1(
        n_majority7_module_94__and_module_2_res), .A2(
        n_majority7_module_94__and_module_1_res), .ZN(
        n_majority7_module_94__and_module_4_res) );
  OR2_X1 u_majority7_module_94__or_module_4_U1 ( .A1(
        n_majority7_module_94__and_module_1_res), .A2(
        n_majority7_module_94__and_module_2_res), .ZN(
        n_majority7_module_94__or_module_4_res) );
  AND2_X1 u_majority7_module_94__and_module_5_U1 ( .A1(
        n_majority7_module_94__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_94__and_module_5_res) );
  OR2_X1 u_majority7_module_94__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_94__and_module_3_res), .ZN(
        n_majority7_module_94__or_module_5_res) );
  AND2_X1 u_majority7_module_94__and_module_6_U1 ( .A1(
        n_majority7_module_94__or_module_1_res), .A2(
        n_majority7_module_94__or_module_2_res), .ZN(
        n_majority7_module_94__and_module_6_res) );
  OR2_X1 u_majority7_module_94__or_module_6_U1 ( .A1(
        n_majority7_module_94__or_module_2_res), .A2(
        n_majority7_module_94__or_module_1_res), .ZN(
        n_majority7_module_94__or_module_6_res) );
  OR2_X1 u_majority7_module_94__or_module_7_U1 ( .A1(
        n_majority7_module_94__and_module_4_res), .A2(
        n_majority7_module_94__and_module_5_res), .ZN(
        n_majority7_module_94__or_module_7_res) );
  AND2_X1 u_majority7_module_94__and_module_7_U1 ( .A1(
        n_majority7_module_94__or_module_3_res), .A2(
        n_majority7_module_94__or_module_4_res), .ZN(
        n_majority7_module_94__and_module_7_res) );
  OR2_X1 u_majority7_module_94__or_module_8_U1 ( .A1(
        n_majority7_module_94__or_module_4_res), .A2(
        n_majority7_module_94__or_module_3_res), .ZN(
        n_majority7_module_94__or_module_8_res) );
  AND2_X1 u_majority7_module_94__and_module_8_U1 ( .A1(
        n_majority7_module_94__or_module_5_res), .A2(
        n_majority7_module_94__and_module_6_res), .ZN(
        n_majority7_module_94__and_module_8_res) );
  OR2_X1 u_majority7_module_94__or_module_9_U1 ( .A1(
        n_majority7_module_94__and_module_6_res), .A2(
        n_majority7_module_94__or_module_5_res), .ZN(
        n_majority7_module_94__or_module_9_res) );
  OR2_X1 u_majority7_module_94__or_module_10_U1 ( .A1(
        n_majority7_module_94__or_module_7_res), .A2(
        n_majority7_module_94__and_module_7_res), .ZN(
        n_majority7_module_94__or_module_10_res) );
  AND2_X1 u_majority7_module_94__and_module_9_U1 ( .A1(
        n_majority7_module_94__or_module_6_res), .A2(
        n_majority7_module_94__or_module_9_res), .ZN(
        n_majority7_module_94__and_module_9_res) );
  OR2_X1 u_majority7_module_94__or_module_11_U1 ( .A1(
        n_majority7_module_94__or_module_10_res), .A2(
        n_majority7_module_94__and_module_8_res), .ZN(
        n_majority7_module_94__or_module_11_res) );
  AND2_X1 u_majority7_module_94__and_module_10_U1 ( .A1(
        n_majority7_module_94__or_module_8_res), .A2(
        n_majority7_module_94__and_module_9_res), .ZN(
        n_majority7_module_94__and_module_10_res) );
  AND2_X1 u_majority7_module_94__and_module_11_U1 ( .A1(
        n_majority7_module_94__and_module_10_res), .A2(
        n_majority7_module_94__or_module_11_res), .ZN(
        n_majority7_module_94_res) );
  DFF_X1 u_reg_module_117__cini_mul_v00_reg ( .D(n_majority7_module_94_res), 
        .CK(clock_5), .Q(n_reg_module_117_res), .QN() );
  AND2_X1 u_majority7_module_95__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_95__and_module_1_res)
         );
  OR2_X1 u_majority7_module_95__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_95__or_module_1_res)
         );
  AND2_X1 u_majority7_module_95__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(n_majority7_module_95__and_module_2_res) );
  OR2_X1 u_majority7_module_95__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_95__or_module_2_res)
         );
  AND2_X1 u_majority7_module_95__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(n_majority7_module_95__and_module_3_res) );
  OR2_X1 u_majority7_module_95__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_95__or_module_3_res)
         );
  AND2_X1 u_majority7_module_95__and_module_4_U1 ( .A1(
        n_majority7_module_95__and_module_2_res), .A2(
        n_majority7_module_95__and_module_1_res), .ZN(
        n_majority7_module_95__and_module_4_res) );
  OR2_X1 u_majority7_module_95__or_module_4_U1 ( .A1(
        n_majority7_module_95__and_module_1_res), .A2(
        n_majority7_module_95__and_module_2_res), .ZN(
        n_majority7_module_95__or_module_4_res) );
  AND2_X1 u_majority7_module_95__and_module_5_U1 ( .A1(
        n_majority7_module_95__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_95__and_module_5_res) );
  OR2_X1 u_majority7_module_95__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_95__and_module_3_res), .ZN(
        n_majority7_module_95__or_module_5_res) );
  AND2_X1 u_majority7_module_95__and_module_6_U1 ( .A1(
        n_majority7_module_95__or_module_1_res), .A2(
        n_majority7_module_95__or_module_2_res), .ZN(
        n_majority7_module_95__and_module_6_res) );
  OR2_X1 u_majority7_module_95__or_module_6_U1 ( .A1(
        n_majority7_module_95__or_module_2_res), .A2(
        n_majority7_module_95__or_module_1_res), .ZN(
        n_majority7_module_95__or_module_6_res) );
  OR2_X1 u_majority7_module_95__or_module_7_U1 ( .A1(
        n_majority7_module_95__and_module_4_res), .A2(
        n_majority7_module_95__and_module_5_res), .ZN(
        n_majority7_module_95__or_module_7_res) );
  AND2_X1 u_majority7_module_95__and_module_7_U1 ( .A1(
        n_majority7_module_95__or_module_3_res), .A2(
        n_majority7_module_95__or_module_4_res), .ZN(
        n_majority7_module_95__and_module_7_res) );
  OR2_X1 u_majority7_module_95__or_module_8_U1 ( .A1(
        n_majority7_module_95__or_module_4_res), .A2(
        n_majority7_module_95__or_module_3_res), .ZN(
        n_majority7_module_95__or_module_8_res) );
  AND2_X1 u_majority7_module_95__and_module_8_U1 ( .A1(
        n_majority7_module_95__or_module_5_res), .A2(
        n_majority7_module_95__and_module_6_res), .ZN(
        n_majority7_module_95__and_module_8_res) );
  OR2_X1 u_majority7_module_95__or_module_9_U1 ( .A1(
        n_majority7_module_95__and_module_6_res), .A2(
        n_majority7_module_95__or_module_5_res), .ZN(
        n_majority7_module_95__or_module_9_res) );
  OR2_X1 u_majority7_module_95__or_module_10_U1 ( .A1(
        n_majority7_module_95__or_module_7_res), .A2(
        n_majority7_module_95__and_module_7_res), .ZN(
        n_majority7_module_95__or_module_10_res) );
  AND2_X1 u_majority7_module_95__and_module_9_U1 ( .A1(
        n_majority7_module_95__or_module_6_res), .A2(
        n_majority7_module_95__or_module_9_res), .ZN(
        n_majority7_module_95__and_module_9_res) );
  OR2_X1 u_majority7_module_95__or_module_11_U1 ( .A1(
        n_majority7_module_95__or_module_10_res), .A2(
        n_majority7_module_95__and_module_8_res), .ZN(
        n_majority7_module_95__or_module_11_res) );
  AND2_X1 u_majority7_module_95__and_module_10_U1 ( .A1(
        n_majority7_module_95__or_module_8_res), .A2(
        n_majority7_module_95__and_module_9_res), .ZN(
        n_majority7_module_95__and_module_10_res) );
  AND2_X1 u_majority7_module_95__and_module_11_U1 ( .A1(
        n_majority7_module_95__and_module_10_res), .A2(
        n_majority7_module_95__or_module_11_res), .ZN(
        n_majority7_module_95_res) );
  DFF_X1 u_reg_module_118__cini_mul_v00_reg ( .D(n_majority7_module_95_res), 
        .CK(clock_5), .Q(n_reg_module_118_res), .QN() );
  DFF_X1 u_reg_module_119__cini_mul_v00_reg ( .D(n_and_module_91_res), .CK(
        clock_5), .Q(n_reg_module_119_res), .QN() );
  AND2_X1 u_majority7_module_96__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_96__and_module_1_res)
         );
  OR2_X1 u_majority7_module_96__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_96__or_module_1_res)
         );
  AND2_X1 u_majority7_module_96__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(n_majority7_module_96__and_module_2_res) );
  OR2_X1 u_majority7_module_96__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_96__or_module_2_res)
         );
  AND2_X1 u_majority7_module_96__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(n_majority7_module_96__and_module_3_res) );
  OR2_X1 u_majority7_module_96__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_96__or_module_3_res)
         );
  AND2_X1 u_majority7_module_96__and_module_4_U1 ( .A1(
        n_majority7_module_96__and_module_2_res), .A2(
        n_majority7_module_96__and_module_1_res), .ZN(
        n_majority7_module_96__and_module_4_res) );
  OR2_X1 u_majority7_module_96__or_module_4_U1 ( .A1(
        n_majority7_module_96__and_module_1_res), .A2(
        n_majority7_module_96__and_module_2_res), .ZN(
        n_majority7_module_96__or_module_4_res) );
  AND2_X1 u_majority7_module_96__and_module_5_U1 ( .A1(
        n_majority7_module_96__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_96__and_module_5_res) );
  OR2_X1 u_majority7_module_96__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_96__and_module_3_res), .ZN(
        n_majority7_module_96__or_module_5_res) );
  AND2_X1 u_majority7_module_96__and_module_6_U1 ( .A1(
        n_majority7_module_96__or_module_1_res), .A2(
        n_majority7_module_96__or_module_2_res), .ZN(
        n_majority7_module_96__and_module_6_res) );
  OR2_X1 u_majority7_module_96__or_module_6_U1 ( .A1(
        n_majority7_module_96__or_module_2_res), .A2(
        n_majority7_module_96__or_module_1_res), .ZN(
        n_majority7_module_96__or_module_6_res) );
  OR2_X1 u_majority7_module_96__or_module_7_U1 ( .A1(
        n_majority7_module_96__and_module_4_res), .A2(
        n_majority7_module_96__and_module_5_res), .ZN(
        n_majority7_module_96__or_module_7_res) );
  AND2_X1 u_majority7_module_96__and_module_7_U1 ( .A1(
        n_majority7_module_96__or_module_3_res), .A2(
        n_majority7_module_96__or_module_4_res), .ZN(
        n_majority7_module_96__and_module_7_res) );
  OR2_X1 u_majority7_module_96__or_module_8_U1 ( .A1(
        n_majority7_module_96__or_module_4_res), .A2(
        n_majority7_module_96__or_module_3_res), .ZN(
        n_majority7_module_96__or_module_8_res) );
  AND2_X1 u_majority7_module_96__and_module_8_U1 ( .A1(
        n_majority7_module_96__or_module_5_res), .A2(
        n_majority7_module_96__and_module_6_res), .ZN(
        n_majority7_module_96__and_module_8_res) );
  OR2_X1 u_majority7_module_96__or_module_9_U1 ( .A1(
        n_majority7_module_96__and_module_6_res), .A2(
        n_majority7_module_96__or_module_5_res), .ZN(
        n_majority7_module_96__or_module_9_res) );
  OR2_X1 u_majority7_module_96__or_module_10_U1 ( .A1(
        n_majority7_module_96__or_module_7_res), .A2(
        n_majority7_module_96__and_module_7_res), .ZN(
        n_majority7_module_96__or_module_10_res) );
  AND2_X1 u_majority7_module_96__and_module_9_U1 ( .A1(
        n_majority7_module_96__or_module_6_res), .A2(
        n_majority7_module_96__or_module_9_res), .ZN(
        n_majority7_module_96__and_module_9_res) );
  OR2_X1 u_majority7_module_96__or_module_11_U1 ( .A1(
        n_majority7_module_96__or_module_10_res), .A2(
        n_majority7_module_96__and_module_8_res), .ZN(
        n_majority7_module_96__or_module_11_res) );
  AND2_X1 u_majority7_module_96__and_module_10_U1 ( .A1(
        n_majority7_module_96__or_module_8_res), .A2(
        n_majority7_module_96__and_module_9_res), .ZN(
        n_majority7_module_96__and_module_10_res) );
  AND2_X1 u_majority7_module_96__and_module_11_U1 ( .A1(
        n_majority7_module_96__and_module_10_res), .A2(
        n_majority7_module_96__or_module_11_res), .ZN(
        n_majority7_module_96_res) );
  DFF_X1 u_reg_module_120__cini_mul_v00_reg ( .D(n_majority7_module_96_res), 
        .CK(clock_5), .Q(n_reg_module_120_res), .QN() );
  AND2_X1 u_majority7_module_97__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_97__and_module_1_res)
         );
  OR2_X1 u_majority7_module_97__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_97__or_module_1_res)
         );
  AND2_X1 u_majority7_module_97__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(n_majority7_module_97__and_module_2_res) );
  OR2_X1 u_majority7_module_97__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_97__or_module_2_res)
         );
  AND2_X1 u_majority7_module_97__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(n_majority7_module_97__and_module_3_res) );
  OR2_X1 u_majority7_module_97__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_97__or_module_3_res)
         );
  AND2_X1 u_majority7_module_97__and_module_4_U1 ( .A1(
        n_majority7_module_97__and_module_2_res), .A2(
        n_majority7_module_97__and_module_1_res), .ZN(
        n_majority7_module_97__and_module_4_res) );
  OR2_X1 u_majority7_module_97__or_module_4_U1 ( .A1(
        n_majority7_module_97__and_module_1_res), .A2(
        n_majority7_module_97__and_module_2_res), .ZN(
        n_majority7_module_97__or_module_4_res) );
  AND2_X1 u_majority7_module_97__and_module_5_U1 ( .A1(
        n_majority7_module_97__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_97__and_module_5_res) );
  OR2_X1 u_majority7_module_97__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_97__and_module_3_res), .ZN(
        n_majority7_module_97__or_module_5_res) );
  AND2_X1 u_majority7_module_97__and_module_6_U1 ( .A1(
        n_majority7_module_97__or_module_1_res), .A2(
        n_majority7_module_97__or_module_2_res), .ZN(
        n_majority7_module_97__and_module_6_res) );
  OR2_X1 u_majority7_module_97__or_module_6_U1 ( .A1(
        n_majority7_module_97__or_module_2_res), .A2(
        n_majority7_module_97__or_module_1_res), .ZN(
        n_majority7_module_97__or_module_6_res) );
  OR2_X1 u_majority7_module_97__or_module_7_U1 ( .A1(
        n_majority7_module_97__and_module_4_res), .A2(
        n_majority7_module_97__and_module_5_res), .ZN(
        n_majority7_module_97__or_module_7_res) );
  AND2_X1 u_majority7_module_97__and_module_7_U1 ( .A1(
        n_majority7_module_97__or_module_3_res), .A2(
        n_majority7_module_97__or_module_4_res), .ZN(
        n_majority7_module_97__and_module_7_res) );
  OR2_X1 u_majority7_module_97__or_module_8_U1 ( .A1(
        n_majority7_module_97__or_module_4_res), .A2(
        n_majority7_module_97__or_module_3_res), .ZN(
        n_majority7_module_97__or_module_8_res) );
  AND2_X1 u_majority7_module_97__and_module_8_U1 ( .A1(
        n_majority7_module_97__or_module_5_res), .A2(
        n_majority7_module_97__and_module_6_res), .ZN(
        n_majority7_module_97__and_module_8_res) );
  OR2_X1 u_majority7_module_97__or_module_9_U1 ( .A1(
        n_majority7_module_97__and_module_6_res), .A2(
        n_majority7_module_97__or_module_5_res), .ZN(
        n_majority7_module_97__or_module_9_res) );
  OR2_X1 u_majority7_module_97__or_module_10_U1 ( .A1(
        n_majority7_module_97__or_module_7_res), .A2(
        n_majority7_module_97__and_module_7_res), .ZN(
        n_majority7_module_97__or_module_10_res) );
  AND2_X1 u_majority7_module_97__and_module_9_U1 ( .A1(
        n_majority7_module_97__or_module_6_res), .A2(
        n_majority7_module_97__or_module_9_res), .ZN(
        n_majority7_module_97__and_module_9_res) );
  OR2_X1 u_majority7_module_97__or_module_11_U1 ( .A1(
        n_majority7_module_97__or_module_10_res), .A2(
        n_majority7_module_97__and_module_8_res), .ZN(
        n_majority7_module_97__or_module_11_res) );
  AND2_X1 u_majority7_module_97__and_module_10_U1 ( .A1(
        n_majority7_module_97__or_module_8_res), .A2(
        n_majority7_module_97__and_module_9_res), .ZN(
        n_majority7_module_97__and_module_10_res) );
  AND2_X1 u_majority7_module_97__and_module_11_U1 ( .A1(
        n_majority7_module_97__and_module_10_res), .A2(
        n_majority7_module_97__or_module_11_res), .ZN(
        n_majority7_module_97_res) );
  DFF_X1 u_reg_module_121__cini_mul_v00_reg ( .D(n_majority7_module_97_res), 
        .CK(clock_5), .Q(n_reg_module_121_res), .QN() );
  AND2_X1 u_majority7_module_98__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_98__and_module_1_res)
         );
  OR2_X1 u_majority7_module_98__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_98__or_module_1_res)
         );
  AND2_X1 u_majority7_module_98__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(n_majority7_module_98__and_module_2_res) );
  OR2_X1 u_majority7_module_98__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_98__or_module_2_res)
         );
  AND2_X1 u_majority7_module_98__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(n_majority7_module_98__and_module_3_res) );
  OR2_X1 u_majority7_module_98__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_98__or_module_3_res)
         );
  AND2_X1 u_majority7_module_98__and_module_4_U1 ( .A1(
        n_majority7_module_98__and_module_2_res), .A2(
        n_majority7_module_98__and_module_1_res), .ZN(
        n_majority7_module_98__and_module_4_res) );
  OR2_X1 u_majority7_module_98__or_module_4_U1 ( .A1(
        n_majority7_module_98__and_module_1_res), .A2(
        n_majority7_module_98__and_module_2_res), .ZN(
        n_majority7_module_98__or_module_4_res) );
  AND2_X1 u_majority7_module_98__and_module_5_U1 ( .A1(
        n_majority7_module_98__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_98__and_module_5_res) );
  OR2_X1 u_majority7_module_98__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_98__and_module_3_res), .ZN(
        n_majority7_module_98__or_module_5_res) );
  AND2_X1 u_majority7_module_98__and_module_6_U1 ( .A1(
        n_majority7_module_98__or_module_1_res), .A2(
        n_majority7_module_98__or_module_2_res), .ZN(
        n_majority7_module_98__and_module_6_res) );
  OR2_X1 u_majority7_module_98__or_module_6_U1 ( .A1(
        n_majority7_module_98__or_module_2_res), .A2(
        n_majority7_module_98__or_module_1_res), .ZN(
        n_majority7_module_98__or_module_6_res) );
  OR2_X1 u_majority7_module_98__or_module_7_U1 ( .A1(
        n_majority7_module_98__and_module_4_res), .A2(
        n_majority7_module_98__and_module_5_res), .ZN(
        n_majority7_module_98__or_module_7_res) );
  AND2_X1 u_majority7_module_98__and_module_7_U1 ( .A1(
        n_majority7_module_98__or_module_3_res), .A2(
        n_majority7_module_98__or_module_4_res), .ZN(
        n_majority7_module_98__and_module_7_res) );
  OR2_X1 u_majority7_module_98__or_module_8_U1 ( .A1(
        n_majority7_module_98__or_module_4_res), .A2(
        n_majority7_module_98__or_module_3_res), .ZN(
        n_majority7_module_98__or_module_8_res) );
  AND2_X1 u_majority7_module_98__and_module_8_U1 ( .A1(
        n_majority7_module_98__or_module_5_res), .A2(
        n_majority7_module_98__and_module_6_res), .ZN(
        n_majority7_module_98__and_module_8_res) );
  OR2_X1 u_majority7_module_98__or_module_9_U1 ( .A1(
        n_majority7_module_98__and_module_6_res), .A2(
        n_majority7_module_98__or_module_5_res), .ZN(
        n_majority7_module_98__or_module_9_res) );
  OR2_X1 u_majority7_module_98__or_module_10_U1 ( .A1(
        n_majority7_module_98__or_module_7_res), .A2(
        n_majority7_module_98__and_module_7_res), .ZN(
        n_majority7_module_98__or_module_10_res) );
  AND2_X1 u_majority7_module_98__and_module_9_U1 ( .A1(
        n_majority7_module_98__or_module_6_res), .A2(
        n_majority7_module_98__or_module_9_res), .ZN(
        n_majority7_module_98__and_module_9_res) );
  OR2_X1 u_majority7_module_98__or_module_11_U1 ( .A1(
        n_majority7_module_98__or_module_10_res), .A2(
        n_majority7_module_98__and_module_8_res), .ZN(
        n_majority7_module_98__or_module_11_res) );
  AND2_X1 u_majority7_module_98__and_module_10_U1 ( .A1(
        n_majority7_module_98__or_module_8_res), .A2(
        n_majority7_module_98__and_module_9_res), .ZN(
        n_majority7_module_98__and_module_10_res) );
  AND2_X1 u_majority7_module_98__and_module_11_U1 ( .A1(
        n_majority7_module_98__and_module_10_res), .A2(
        n_majority7_module_98__or_module_11_res), .ZN(
        n_majority7_module_98_res) );
  DFF_X1 u_reg_module_122__cini_mul_v00_reg ( .D(n_majority7_module_98_res), 
        .CK(clock_5), .Q(n_reg_module_122_res), .QN() );
  AND2_X1 u_majority7_module_99__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_99__and_module_1_res)
         );
  OR2_X1 u_majority7_module_99__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_99__or_module_1_res)
         );
  AND2_X1 u_majority7_module_99__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(n_majority7_module_99__and_module_2_res) );
  OR2_X1 u_majority7_module_99__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_99__or_module_2_res)
         );
  AND2_X1 u_majority7_module_99__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(n_majority7_module_99__and_module_3_res) );
  OR2_X1 u_majority7_module_99__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_99__or_module_3_res)
         );
  AND2_X1 u_majority7_module_99__and_module_4_U1 ( .A1(
        n_majority7_module_99__and_module_2_res), .A2(
        n_majority7_module_99__and_module_1_res), .ZN(
        n_majority7_module_99__and_module_4_res) );
  OR2_X1 u_majority7_module_99__or_module_4_U1 ( .A1(
        n_majority7_module_99__and_module_1_res), .A2(
        n_majority7_module_99__and_module_2_res), .ZN(
        n_majority7_module_99__or_module_4_res) );
  AND2_X1 u_majority7_module_99__and_module_5_U1 ( .A1(
        n_majority7_module_99__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_99__and_module_5_res) );
  OR2_X1 u_majority7_module_99__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_99__and_module_3_res), .ZN(
        n_majority7_module_99__or_module_5_res) );
  AND2_X1 u_majority7_module_99__and_module_6_U1 ( .A1(
        n_majority7_module_99__or_module_1_res), .A2(
        n_majority7_module_99__or_module_2_res), .ZN(
        n_majority7_module_99__and_module_6_res) );
  OR2_X1 u_majority7_module_99__or_module_6_U1 ( .A1(
        n_majority7_module_99__or_module_2_res), .A2(
        n_majority7_module_99__or_module_1_res), .ZN(
        n_majority7_module_99__or_module_6_res) );
  OR2_X1 u_majority7_module_99__or_module_7_U1 ( .A1(
        n_majority7_module_99__and_module_4_res), .A2(
        n_majority7_module_99__and_module_5_res), .ZN(
        n_majority7_module_99__or_module_7_res) );
  AND2_X1 u_majority7_module_99__and_module_7_U1 ( .A1(
        n_majority7_module_99__or_module_3_res), .A2(
        n_majority7_module_99__or_module_4_res), .ZN(
        n_majority7_module_99__and_module_7_res) );
  OR2_X1 u_majority7_module_99__or_module_8_U1 ( .A1(
        n_majority7_module_99__or_module_4_res), .A2(
        n_majority7_module_99__or_module_3_res), .ZN(
        n_majority7_module_99__or_module_8_res) );
  AND2_X1 u_majority7_module_99__and_module_8_U1 ( .A1(
        n_majority7_module_99__or_module_5_res), .A2(
        n_majority7_module_99__and_module_6_res), .ZN(
        n_majority7_module_99__and_module_8_res) );
  OR2_X1 u_majority7_module_99__or_module_9_U1 ( .A1(
        n_majority7_module_99__and_module_6_res), .A2(
        n_majority7_module_99__or_module_5_res), .ZN(
        n_majority7_module_99__or_module_9_res) );
  OR2_X1 u_majority7_module_99__or_module_10_U1 ( .A1(
        n_majority7_module_99__or_module_7_res), .A2(
        n_majority7_module_99__and_module_7_res), .ZN(
        n_majority7_module_99__or_module_10_res) );
  AND2_X1 u_majority7_module_99__and_module_9_U1 ( .A1(
        n_majority7_module_99__or_module_6_res), .A2(
        n_majority7_module_99__or_module_9_res), .ZN(
        n_majority7_module_99__and_module_9_res) );
  OR2_X1 u_majority7_module_99__or_module_11_U1 ( .A1(
        n_majority7_module_99__or_module_10_res), .A2(
        n_majority7_module_99__and_module_8_res), .ZN(
        n_majority7_module_99__or_module_11_res) );
  AND2_X1 u_majority7_module_99__and_module_10_U1 ( .A1(
        n_majority7_module_99__or_module_8_res), .A2(
        n_majority7_module_99__and_module_9_res), .ZN(
        n_majority7_module_99__and_module_10_res) );
  AND2_X1 u_majority7_module_99__and_module_11_U1 ( .A1(
        n_majority7_module_99__and_module_10_res), .A2(
        n_majority7_module_99__or_module_11_res), .ZN(
        n_majority7_module_99_res) );
  DFF_X1 u_reg_module_123__cini_mul_v00_reg ( .D(n_majority7_module_99_res), 
        .CK(clock_5), .Q(n_reg_module_123_res), .QN() );
  DFF_X1 u_reg_module_124__cini_mul_v00_reg ( .D(n_and_module_96_res), .CK(
        clock_5), .Q(n_reg_module_124_res), .QN() );
  DFF_X1 u_reg_module_125__cini_mul_v00_reg ( .D(n_and_module_97_res), .CK(
        clock_6), .Q(n_reg_module_125_res), .QN() );
  AND2_X1 u_majority7_module_100__and_module_1_U1 ( .A1(n_xor_module_157_res), 
        .A2(n_xor_module_85_res), .ZN(n_majority7_module_100__and_module_1_res) );
  OR2_X1 u_majority7_module_100__or_module_1_U1 ( .A1(n_xor_module_85_res), 
        .A2(n_xor_module_157_res), .ZN(n_majority7_module_100__or_module_1_res) );
  AND2_X1 u_majority7_module_100__and_module_2_U1 ( .A1(n_xor_module_121_res), 
        .A2(n_xor_module_109_res), .ZN(
        n_majority7_module_100__and_module_2_res) );
  OR2_X1 u_majority7_module_100__or_module_2_U1 ( .A1(n_xor_module_109_res), 
        .A2(n_xor_module_121_res), .ZN(n_majority7_module_100__or_module_2_res) );
  AND2_X1 u_majority7_module_100__and_module_3_U1 ( .A1(n_xor_module_145_res), 
        .A2(n_xor_module_133_res), .ZN(
        n_majority7_module_100__and_module_3_res) );
  OR2_X1 u_majority7_module_100__or_module_3_U1 ( .A1(n_xor_module_133_res), 
        .A2(n_xor_module_145_res), .ZN(n_majority7_module_100__or_module_3_res) );
  AND2_X1 u_majority7_module_100__and_module_4_U1 ( .A1(
        n_majority7_module_100__and_module_2_res), .A2(
        n_majority7_module_100__and_module_1_res), .ZN(
        n_majority7_module_100__and_module_4_res) );
  OR2_X1 u_majority7_module_100__or_module_4_U1 ( .A1(
        n_majority7_module_100__and_module_1_res), .A2(
        n_majority7_module_100__and_module_2_res), .ZN(
        n_majority7_module_100__or_module_4_res) );
  AND2_X1 u_majority7_module_100__and_module_5_U1 ( .A1(
        n_majority7_module_100__and_module_3_res), .A2(n_xor_module_97_res), 
        .ZN(n_majority7_module_100__and_module_5_res) );
  OR2_X1 u_majority7_module_100__or_module_5_U1 ( .A1(n_xor_module_97_res), 
        .A2(n_majority7_module_100__and_module_3_res), .ZN(
        n_majority7_module_100__or_module_5_res) );
  AND2_X1 u_majority7_module_100__and_module_6_U1 ( .A1(
        n_majority7_module_100__or_module_1_res), .A2(
        n_majority7_module_100__or_module_2_res), .ZN(
        n_majority7_module_100__and_module_6_res) );
  OR2_X1 u_majority7_module_100__or_module_6_U1 ( .A1(
        n_majority7_module_100__or_module_2_res), .A2(
        n_majority7_module_100__or_module_1_res), .ZN(
        n_majority7_module_100__or_module_6_res) );
  OR2_X1 u_majority7_module_100__or_module_7_U1 ( .A1(
        n_majority7_module_100__and_module_4_res), .A2(
        n_majority7_module_100__and_module_5_res), .ZN(
        n_majority7_module_100__or_module_7_res) );
  AND2_X1 u_majority7_module_100__and_module_7_U1 ( .A1(
        n_majority7_module_100__or_module_3_res), .A2(
        n_majority7_module_100__or_module_4_res), .ZN(
        n_majority7_module_100__and_module_7_res) );
  OR2_X1 u_majority7_module_100__or_module_8_U1 ( .A1(
        n_majority7_module_100__or_module_4_res), .A2(
        n_majority7_module_100__or_module_3_res), .ZN(
        n_majority7_module_100__or_module_8_res) );
  AND2_X1 u_majority7_module_100__and_module_8_U1 ( .A1(
        n_majority7_module_100__or_module_5_res), .A2(
        n_majority7_module_100__and_module_6_res), .ZN(
        n_majority7_module_100__and_module_8_res) );
  OR2_X1 u_majority7_module_100__or_module_9_U1 ( .A1(
        n_majority7_module_100__and_module_6_res), .A2(
        n_majority7_module_100__or_module_5_res), .ZN(
        n_majority7_module_100__or_module_9_res) );
  OR2_X1 u_majority7_module_100__or_module_10_U1 ( .A1(
        n_majority7_module_100__or_module_7_res), .A2(
        n_majority7_module_100__and_module_7_res), .ZN(
        n_majority7_module_100__or_module_10_res) );
  AND2_X1 u_majority7_module_100__and_module_9_U1 ( .A1(
        n_majority7_module_100__or_module_6_res), .A2(
        n_majority7_module_100__or_module_9_res), .ZN(
        n_majority7_module_100__and_module_9_res) );
  OR2_X1 u_majority7_module_100__or_module_11_U1 ( .A1(
        n_majority7_module_100__or_module_10_res), .A2(
        n_majority7_module_100__and_module_8_res), .ZN(
        n_majority7_module_100__or_module_11_res) );
  AND2_X1 u_majority7_module_100__and_module_10_U1 ( .A1(
        n_majority7_module_100__or_module_8_res), .A2(
        n_majority7_module_100__and_module_9_res), .ZN(
        n_majority7_module_100__and_module_10_res) );
  AND2_X1 u_majority7_module_100__and_module_11_U1 ( .A1(
        n_majority7_module_100__and_module_10_res), .A2(
        n_majority7_module_100__or_module_11_res), .ZN(
        n_majority7_module_100_res) );
  DFF_X1 u_reg_module_126__cini_mul_v00_reg ( .D(n_majority7_module_100_res), 
        .CK(clock_6), .Q(n_reg_module_126_res), .QN() );
  AND2_X1 u_majority7_module_101__and_module_1_U1 ( .A1(n_xor_module_158_res), 
        .A2(n_xor_module_86_res), .ZN(n_majority7_module_101__and_module_1_res) );
  OR2_X1 u_majority7_module_101__or_module_1_U1 ( .A1(n_xor_module_86_res), 
        .A2(n_xor_module_158_res), .ZN(n_majority7_module_101__or_module_1_res) );
  AND2_X1 u_majority7_module_101__and_module_2_U1 ( .A1(n_xor_module_122_res), 
        .A2(n_xor_module_110_res), .ZN(
        n_majority7_module_101__and_module_2_res) );
  OR2_X1 u_majority7_module_101__or_module_2_U1 ( .A1(n_xor_module_110_res), 
        .A2(n_xor_module_122_res), .ZN(n_majority7_module_101__or_module_2_res) );
  AND2_X1 u_majority7_module_101__and_module_3_U1 ( .A1(n_xor_module_146_res), 
        .A2(n_xor_module_134_res), .ZN(
        n_majority7_module_101__and_module_3_res) );
  OR2_X1 u_majority7_module_101__or_module_3_U1 ( .A1(n_xor_module_134_res), 
        .A2(n_xor_module_146_res), .ZN(n_majority7_module_101__or_module_3_res) );
  AND2_X1 u_majority7_module_101__and_module_4_U1 ( .A1(
        n_majority7_module_101__and_module_2_res), .A2(
        n_majority7_module_101__and_module_1_res), .ZN(
        n_majority7_module_101__and_module_4_res) );
  OR2_X1 u_majority7_module_101__or_module_4_U1 ( .A1(
        n_majority7_module_101__and_module_1_res), .A2(
        n_majority7_module_101__and_module_2_res), .ZN(
        n_majority7_module_101__or_module_4_res) );
  AND2_X1 u_majority7_module_101__and_module_5_U1 ( .A1(
        n_majority7_module_101__and_module_3_res), .A2(n_xor_module_98_res), 
        .ZN(n_majority7_module_101__and_module_5_res) );
  OR2_X1 u_majority7_module_101__or_module_5_U1 ( .A1(n_xor_module_98_res), 
        .A2(n_majority7_module_101__and_module_3_res), .ZN(
        n_majority7_module_101__or_module_5_res) );
  AND2_X1 u_majority7_module_101__and_module_6_U1 ( .A1(
        n_majority7_module_101__or_module_1_res), .A2(
        n_majority7_module_101__or_module_2_res), .ZN(
        n_majority7_module_101__and_module_6_res) );
  OR2_X1 u_majority7_module_101__or_module_6_U1 ( .A1(
        n_majority7_module_101__or_module_2_res), .A2(
        n_majority7_module_101__or_module_1_res), .ZN(
        n_majority7_module_101__or_module_6_res) );
  OR2_X1 u_majority7_module_101__or_module_7_U1 ( .A1(
        n_majority7_module_101__and_module_4_res), .A2(
        n_majority7_module_101__and_module_5_res), .ZN(
        n_majority7_module_101__or_module_7_res) );
  AND2_X1 u_majority7_module_101__and_module_7_U1 ( .A1(
        n_majority7_module_101__or_module_3_res), .A2(
        n_majority7_module_101__or_module_4_res), .ZN(
        n_majority7_module_101__and_module_7_res) );
  OR2_X1 u_majority7_module_101__or_module_8_U1 ( .A1(
        n_majority7_module_101__or_module_4_res), .A2(
        n_majority7_module_101__or_module_3_res), .ZN(
        n_majority7_module_101__or_module_8_res) );
  AND2_X1 u_majority7_module_101__and_module_8_U1 ( .A1(
        n_majority7_module_101__or_module_5_res), .A2(
        n_majority7_module_101__and_module_6_res), .ZN(
        n_majority7_module_101__and_module_8_res) );
  OR2_X1 u_majority7_module_101__or_module_9_U1 ( .A1(
        n_majority7_module_101__and_module_6_res), .A2(
        n_majority7_module_101__or_module_5_res), .ZN(
        n_majority7_module_101__or_module_9_res) );
  OR2_X1 u_majority7_module_101__or_module_10_U1 ( .A1(
        n_majority7_module_101__or_module_7_res), .A2(
        n_majority7_module_101__and_module_7_res), .ZN(
        n_majority7_module_101__or_module_10_res) );
  AND2_X1 u_majority7_module_101__and_module_9_U1 ( .A1(
        n_majority7_module_101__or_module_6_res), .A2(
        n_majority7_module_101__or_module_9_res), .ZN(
        n_majority7_module_101__and_module_9_res) );
  OR2_X1 u_majority7_module_101__or_module_11_U1 ( .A1(
        n_majority7_module_101__or_module_10_res), .A2(
        n_majority7_module_101__and_module_8_res), .ZN(
        n_majority7_module_101__or_module_11_res) );
  AND2_X1 u_majority7_module_101__and_module_10_U1 ( .A1(
        n_majority7_module_101__or_module_8_res), .A2(
        n_majority7_module_101__and_module_9_res), .ZN(
        n_majority7_module_101__and_module_10_res) );
  AND2_X1 u_majority7_module_101__and_module_11_U1 ( .A1(
        n_majority7_module_101__and_module_10_res), .A2(
        n_majority7_module_101__or_module_11_res), .ZN(
        n_majority7_module_101_res) );
  DFF_X1 u_reg_module_127__cini_mul_v00_reg ( .D(n_majority7_module_101_res), 
        .CK(clock_6), .Q(n_reg_module_127_res), .QN() );
  AND2_X1 u_majority7_module_102__and_module_1_U1 ( .A1(n_xor_module_159_res), 
        .A2(n_xor_module_87_res), .ZN(n_majority7_module_102__and_module_1_res) );
  OR2_X1 u_majority7_module_102__or_module_1_U1 ( .A1(n_xor_module_87_res), 
        .A2(n_xor_module_159_res), .ZN(n_majority7_module_102__or_module_1_res) );
  AND2_X1 u_majority7_module_102__and_module_2_U1 ( .A1(n_xor_module_123_res), 
        .A2(n_xor_module_111_res), .ZN(
        n_majority7_module_102__and_module_2_res) );
  OR2_X1 u_majority7_module_102__or_module_2_U1 ( .A1(n_xor_module_111_res), 
        .A2(n_xor_module_123_res), .ZN(n_majority7_module_102__or_module_2_res) );
  AND2_X1 u_majority7_module_102__and_module_3_U1 ( .A1(n_xor_module_147_res), 
        .A2(n_xor_module_135_res), .ZN(
        n_majority7_module_102__and_module_3_res) );
  OR2_X1 u_majority7_module_102__or_module_3_U1 ( .A1(n_xor_module_135_res), 
        .A2(n_xor_module_147_res), .ZN(n_majority7_module_102__or_module_3_res) );
  AND2_X1 u_majority7_module_102__and_module_4_U1 ( .A1(
        n_majority7_module_102__and_module_2_res), .A2(
        n_majority7_module_102__and_module_1_res), .ZN(
        n_majority7_module_102__and_module_4_res) );
  OR2_X1 u_majority7_module_102__or_module_4_U1 ( .A1(
        n_majority7_module_102__and_module_1_res), .A2(
        n_majority7_module_102__and_module_2_res), .ZN(
        n_majority7_module_102__or_module_4_res) );
  AND2_X1 u_majority7_module_102__and_module_5_U1 ( .A1(
        n_majority7_module_102__and_module_3_res), .A2(n_xor_module_99_res), 
        .ZN(n_majority7_module_102__and_module_5_res) );
  OR2_X1 u_majority7_module_102__or_module_5_U1 ( .A1(n_xor_module_99_res), 
        .A2(n_majority7_module_102__and_module_3_res), .ZN(
        n_majority7_module_102__or_module_5_res) );
  AND2_X1 u_majority7_module_102__and_module_6_U1 ( .A1(
        n_majority7_module_102__or_module_1_res), .A2(
        n_majority7_module_102__or_module_2_res), .ZN(
        n_majority7_module_102__and_module_6_res) );
  OR2_X1 u_majority7_module_102__or_module_6_U1 ( .A1(
        n_majority7_module_102__or_module_2_res), .A2(
        n_majority7_module_102__or_module_1_res), .ZN(
        n_majority7_module_102__or_module_6_res) );
  OR2_X1 u_majority7_module_102__or_module_7_U1 ( .A1(
        n_majority7_module_102__and_module_4_res), .A2(
        n_majority7_module_102__and_module_5_res), .ZN(
        n_majority7_module_102__or_module_7_res) );
  AND2_X1 u_majority7_module_102__and_module_7_U1 ( .A1(
        n_majority7_module_102__or_module_3_res), .A2(
        n_majority7_module_102__or_module_4_res), .ZN(
        n_majority7_module_102__and_module_7_res) );
  OR2_X1 u_majority7_module_102__or_module_8_U1 ( .A1(
        n_majority7_module_102__or_module_4_res), .A2(
        n_majority7_module_102__or_module_3_res), .ZN(
        n_majority7_module_102__or_module_8_res) );
  AND2_X1 u_majority7_module_102__and_module_8_U1 ( .A1(
        n_majority7_module_102__or_module_5_res), .A2(
        n_majority7_module_102__and_module_6_res), .ZN(
        n_majority7_module_102__and_module_8_res) );
  OR2_X1 u_majority7_module_102__or_module_9_U1 ( .A1(
        n_majority7_module_102__and_module_6_res), .A2(
        n_majority7_module_102__or_module_5_res), .ZN(
        n_majority7_module_102__or_module_9_res) );
  OR2_X1 u_majority7_module_102__or_module_10_U1 ( .A1(
        n_majority7_module_102__or_module_7_res), .A2(
        n_majority7_module_102__and_module_7_res), .ZN(
        n_majority7_module_102__or_module_10_res) );
  AND2_X1 u_majority7_module_102__and_module_9_U1 ( .A1(
        n_majority7_module_102__or_module_6_res), .A2(
        n_majority7_module_102__or_module_9_res), .ZN(
        n_majority7_module_102__and_module_9_res) );
  OR2_X1 u_majority7_module_102__or_module_11_U1 ( .A1(
        n_majority7_module_102__or_module_10_res), .A2(
        n_majority7_module_102__and_module_8_res), .ZN(
        n_majority7_module_102__or_module_11_res) );
  AND2_X1 u_majority7_module_102__and_module_10_U1 ( .A1(
        n_majority7_module_102__or_module_8_res), .A2(
        n_majority7_module_102__and_module_9_res), .ZN(
        n_majority7_module_102__and_module_10_res) );
  AND2_X1 u_majority7_module_102__and_module_11_U1 ( .A1(
        n_majority7_module_102__and_module_10_res), .A2(
        n_majority7_module_102__or_module_11_res), .ZN(
        n_majority7_module_102_res) );
  DFF_X1 u_reg_module_128__cini_mul_v00_reg ( .D(n_majority7_module_102_res), 
        .CK(clock_6), .Q(n_reg_module_128_res), .QN() );
  AND2_X1 u_majority7_module_103__and_module_1_U1 ( .A1(n_xor_module_160_res), 
        .A2(n_xor_module_88_res), .ZN(n_majority7_module_103__and_module_1_res) );
  OR2_X1 u_majority7_module_103__or_module_1_U1 ( .A1(n_xor_module_88_res), 
        .A2(n_xor_module_160_res), .ZN(n_majority7_module_103__or_module_1_res) );
  AND2_X1 u_majority7_module_103__and_module_2_U1 ( .A1(n_xor_module_124_res), 
        .A2(n_xor_module_112_res), .ZN(
        n_majority7_module_103__and_module_2_res) );
  OR2_X1 u_majority7_module_103__or_module_2_U1 ( .A1(n_xor_module_112_res), 
        .A2(n_xor_module_124_res), .ZN(n_majority7_module_103__or_module_2_res) );
  AND2_X1 u_majority7_module_103__and_module_3_U1 ( .A1(n_xor_module_148_res), 
        .A2(n_xor_module_136_res), .ZN(
        n_majority7_module_103__and_module_3_res) );
  OR2_X1 u_majority7_module_103__or_module_3_U1 ( .A1(n_xor_module_136_res), 
        .A2(n_xor_module_148_res), .ZN(n_majority7_module_103__or_module_3_res) );
  AND2_X1 u_majority7_module_103__and_module_4_U1 ( .A1(
        n_majority7_module_103__and_module_2_res), .A2(
        n_majority7_module_103__and_module_1_res), .ZN(
        n_majority7_module_103__and_module_4_res) );
  OR2_X1 u_majority7_module_103__or_module_4_U1 ( .A1(
        n_majority7_module_103__and_module_1_res), .A2(
        n_majority7_module_103__and_module_2_res), .ZN(
        n_majority7_module_103__or_module_4_res) );
  AND2_X1 u_majority7_module_103__and_module_5_U1 ( .A1(
        n_majority7_module_103__and_module_3_res), .A2(n_xor_module_100_res), 
        .ZN(n_majority7_module_103__and_module_5_res) );
  OR2_X1 u_majority7_module_103__or_module_5_U1 ( .A1(n_xor_module_100_res), 
        .A2(n_majority7_module_103__and_module_3_res), .ZN(
        n_majority7_module_103__or_module_5_res) );
  AND2_X1 u_majority7_module_103__and_module_6_U1 ( .A1(
        n_majority7_module_103__or_module_1_res), .A2(
        n_majority7_module_103__or_module_2_res), .ZN(
        n_majority7_module_103__and_module_6_res) );
  OR2_X1 u_majority7_module_103__or_module_6_U1 ( .A1(
        n_majority7_module_103__or_module_2_res), .A2(
        n_majority7_module_103__or_module_1_res), .ZN(
        n_majority7_module_103__or_module_6_res) );
  OR2_X1 u_majority7_module_103__or_module_7_U1 ( .A1(
        n_majority7_module_103__and_module_4_res), .A2(
        n_majority7_module_103__and_module_5_res), .ZN(
        n_majority7_module_103__or_module_7_res) );
  AND2_X1 u_majority7_module_103__and_module_7_U1 ( .A1(
        n_majority7_module_103__or_module_3_res), .A2(
        n_majority7_module_103__or_module_4_res), .ZN(
        n_majority7_module_103__and_module_7_res) );
  OR2_X1 u_majority7_module_103__or_module_8_U1 ( .A1(
        n_majority7_module_103__or_module_4_res), .A2(
        n_majority7_module_103__or_module_3_res), .ZN(
        n_majority7_module_103__or_module_8_res) );
  AND2_X1 u_majority7_module_103__and_module_8_U1 ( .A1(
        n_majority7_module_103__or_module_5_res), .A2(
        n_majority7_module_103__and_module_6_res), .ZN(
        n_majority7_module_103__and_module_8_res) );
  OR2_X1 u_majority7_module_103__or_module_9_U1 ( .A1(
        n_majority7_module_103__and_module_6_res), .A2(
        n_majority7_module_103__or_module_5_res), .ZN(
        n_majority7_module_103__or_module_9_res) );
  OR2_X1 u_majority7_module_103__or_module_10_U1 ( .A1(
        n_majority7_module_103__or_module_7_res), .A2(
        n_majority7_module_103__and_module_7_res), .ZN(
        n_majority7_module_103__or_module_10_res) );
  AND2_X1 u_majority7_module_103__and_module_9_U1 ( .A1(
        n_majority7_module_103__or_module_6_res), .A2(
        n_majority7_module_103__or_module_9_res), .ZN(
        n_majority7_module_103__and_module_9_res) );
  OR2_X1 u_majority7_module_103__or_module_11_U1 ( .A1(
        n_majority7_module_103__or_module_10_res), .A2(
        n_majority7_module_103__and_module_8_res), .ZN(
        n_majority7_module_103__or_module_11_res) );
  AND2_X1 u_majority7_module_103__and_module_10_U1 ( .A1(
        n_majority7_module_103__or_module_8_res), .A2(
        n_majority7_module_103__and_module_9_res), .ZN(
        n_majority7_module_103__and_module_10_res) );
  AND2_X1 u_majority7_module_103__and_module_11_U1 ( .A1(
        n_majority7_module_103__and_module_10_res), .A2(
        n_majority7_module_103__or_module_11_res), .ZN(
        n_majority7_module_103_res) );
  DFF_X1 u_reg_module_129__cini_mul_v00_reg ( .D(n_majority7_module_103_res), 
        .CK(clock_6), .Q(n_reg_module_129_res), .QN() );
  DFF_X1 u_reg_module_130__cini_mul_v00_reg ( .D(n_and_module_102_res), .CK(
        clock_6), .Q(n_reg_module_130_res), .QN() );
  AND2_X1 u_majority7_module_104__and_module_1_U1 ( .A1(n_xor_module_161_res), 
        .A2(n_xor_module_89_res), .ZN(n_majority7_module_104__and_module_1_res) );
  OR2_X1 u_majority7_module_104__or_module_1_U1 ( .A1(n_xor_module_89_res), 
        .A2(n_xor_module_161_res), .ZN(n_majority7_module_104__or_module_1_res) );
  AND2_X1 u_majority7_module_104__and_module_2_U1 ( .A1(n_xor_module_125_res), 
        .A2(n_xor_module_113_res), .ZN(
        n_majority7_module_104__and_module_2_res) );
  OR2_X1 u_majority7_module_104__or_module_2_U1 ( .A1(n_xor_module_113_res), 
        .A2(n_xor_module_125_res), .ZN(n_majority7_module_104__or_module_2_res) );
  AND2_X1 u_majority7_module_104__and_module_3_U1 ( .A1(n_xor_module_149_res), 
        .A2(n_xor_module_137_res), .ZN(
        n_majority7_module_104__and_module_3_res) );
  OR2_X1 u_majority7_module_104__or_module_3_U1 ( .A1(n_xor_module_137_res), 
        .A2(n_xor_module_149_res), .ZN(n_majority7_module_104__or_module_3_res) );
  AND2_X1 u_majority7_module_104__and_module_4_U1 ( .A1(
        n_majority7_module_104__and_module_2_res), .A2(
        n_majority7_module_104__and_module_1_res), .ZN(
        n_majority7_module_104__and_module_4_res) );
  OR2_X1 u_majority7_module_104__or_module_4_U1 ( .A1(
        n_majority7_module_104__and_module_1_res), .A2(
        n_majority7_module_104__and_module_2_res), .ZN(
        n_majority7_module_104__or_module_4_res) );
  AND2_X1 u_majority7_module_104__and_module_5_U1 ( .A1(
        n_majority7_module_104__and_module_3_res), .A2(n_xor_module_101_res), 
        .ZN(n_majority7_module_104__and_module_5_res) );
  OR2_X1 u_majority7_module_104__or_module_5_U1 ( .A1(n_xor_module_101_res), 
        .A2(n_majority7_module_104__and_module_3_res), .ZN(
        n_majority7_module_104__or_module_5_res) );
  AND2_X1 u_majority7_module_104__and_module_6_U1 ( .A1(
        n_majority7_module_104__or_module_1_res), .A2(
        n_majority7_module_104__or_module_2_res), .ZN(
        n_majority7_module_104__and_module_6_res) );
  OR2_X1 u_majority7_module_104__or_module_6_U1 ( .A1(
        n_majority7_module_104__or_module_2_res), .A2(
        n_majority7_module_104__or_module_1_res), .ZN(
        n_majority7_module_104__or_module_6_res) );
  OR2_X1 u_majority7_module_104__or_module_7_U1 ( .A1(
        n_majority7_module_104__and_module_4_res), .A2(
        n_majority7_module_104__and_module_5_res), .ZN(
        n_majority7_module_104__or_module_7_res) );
  AND2_X1 u_majority7_module_104__and_module_7_U1 ( .A1(
        n_majority7_module_104__or_module_3_res), .A2(
        n_majority7_module_104__or_module_4_res), .ZN(
        n_majority7_module_104__and_module_7_res) );
  OR2_X1 u_majority7_module_104__or_module_8_U1 ( .A1(
        n_majority7_module_104__or_module_4_res), .A2(
        n_majority7_module_104__or_module_3_res), .ZN(
        n_majority7_module_104__or_module_8_res) );
  AND2_X1 u_majority7_module_104__and_module_8_U1 ( .A1(
        n_majority7_module_104__or_module_5_res), .A2(
        n_majority7_module_104__and_module_6_res), .ZN(
        n_majority7_module_104__and_module_8_res) );
  OR2_X1 u_majority7_module_104__or_module_9_U1 ( .A1(
        n_majority7_module_104__and_module_6_res), .A2(
        n_majority7_module_104__or_module_5_res), .ZN(
        n_majority7_module_104__or_module_9_res) );
  OR2_X1 u_majority7_module_104__or_module_10_U1 ( .A1(
        n_majority7_module_104__or_module_7_res), .A2(
        n_majority7_module_104__and_module_7_res), .ZN(
        n_majority7_module_104__or_module_10_res) );
  AND2_X1 u_majority7_module_104__and_module_9_U1 ( .A1(
        n_majority7_module_104__or_module_6_res), .A2(
        n_majority7_module_104__or_module_9_res), .ZN(
        n_majority7_module_104__and_module_9_res) );
  OR2_X1 u_majority7_module_104__or_module_11_U1 ( .A1(
        n_majority7_module_104__or_module_10_res), .A2(
        n_majority7_module_104__and_module_8_res), .ZN(
        n_majority7_module_104__or_module_11_res) );
  AND2_X1 u_majority7_module_104__and_module_10_U1 ( .A1(
        n_majority7_module_104__or_module_8_res), .A2(
        n_majority7_module_104__and_module_9_res), .ZN(
        n_majority7_module_104__and_module_10_res) );
  AND2_X1 u_majority7_module_104__and_module_11_U1 ( .A1(
        n_majority7_module_104__and_module_10_res), .A2(
        n_majority7_module_104__or_module_11_res), .ZN(
        n_majority7_module_104_res) );
  DFF_X1 u_reg_module_131__cini_mul_v00_reg ( .D(n_majority7_module_104_res), 
        .CK(clock_6), .Q(n_reg_module_131_res), .QN() );
  AND2_X1 u_majority7_module_105__and_module_1_U1 ( .A1(n_xor_module_162_res), 
        .A2(n_xor_module_90_res), .ZN(n_majority7_module_105__and_module_1_res) );
  OR2_X1 u_majority7_module_105__or_module_1_U1 ( .A1(n_xor_module_90_res), 
        .A2(n_xor_module_162_res), .ZN(n_majority7_module_105__or_module_1_res) );
  AND2_X1 u_majority7_module_105__and_module_2_U1 ( .A1(n_xor_module_126_res), 
        .A2(n_xor_module_114_res), .ZN(
        n_majority7_module_105__and_module_2_res) );
  OR2_X1 u_majority7_module_105__or_module_2_U1 ( .A1(n_xor_module_114_res), 
        .A2(n_xor_module_126_res), .ZN(n_majority7_module_105__or_module_2_res) );
  AND2_X1 u_majority7_module_105__and_module_3_U1 ( .A1(n_xor_module_150_res), 
        .A2(n_xor_module_138_res), .ZN(
        n_majority7_module_105__and_module_3_res) );
  OR2_X1 u_majority7_module_105__or_module_3_U1 ( .A1(n_xor_module_138_res), 
        .A2(n_xor_module_150_res), .ZN(n_majority7_module_105__or_module_3_res) );
  AND2_X1 u_majority7_module_105__and_module_4_U1 ( .A1(
        n_majority7_module_105__and_module_2_res), .A2(
        n_majority7_module_105__and_module_1_res), .ZN(
        n_majority7_module_105__and_module_4_res) );
  OR2_X1 u_majority7_module_105__or_module_4_U1 ( .A1(
        n_majority7_module_105__and_module_1_res), .A2(
        n_majority7_module_105__and_module_2_res), .ZN(
        n_majority7_module_105__or_module_4_res) );
  AND2_X1 u_majority7_module_105__and_module_5_U1 ( .A1(
        n_majority7_module_105__and_module_3_res), .A2(n_xor_module_102_res), 
        .ZN(n_majority7_module_105__and_module_5_res) );
  OR2_X1 u_majority7_module_105__or_module_5_U1 ( .A1(n_xor_module_102_res), 
        .A2(n_majority7_module_105__and_module_3_res), .ZN(
        n_majority7_module_105__or_module_5_res) );
  AND2_X1 u_majority7_module_105__and_module_6_U1 ( .A1(
        n_majority7_module_105__or_module_1_res), .A2(
        n_majority7_module_105__or_module_2_res), .ZN(
        n_majority7_module_105__and_module_6_res) );
  OR2_X1 u_majority7_module_105__or_module_6_U1 ( .A1(
        n_majority7_module_105__or_module_2_res), .A2(
        n_majority7_module_105__or_module_1_res), .ZN(
        n_majority7_module_105__or_module_6_res) );
  OR2_X1 u_majority7_module_105__or_module_7_U1 ( .A1(
        n_majority7_module_105__and_module_4_res), .A2(
        n_majority7_module_105__and_module_5_res), .ZN(
        n_majority7_module_105__or_module_7_res) );
  AND2_X1 u_majority7_module_105__and_module_7_U1 ( .A1(
        n_majority7_module_105__or_module_3_res), .A2(
        n_majority7_module_105__or_module_4_res), .ZN(
        n_majority7_module_105__and_module_7_res) );
  OR2_X1 u_majority7_module_105__or_module_8_U1 ( .A1(
        n_majority7_module_105__or_module_4_res), .A2(
        n_majority7_module_105__or_module_3_res), .ZN(
        n_majority7_module_105__or_module_8_res) );
  AND2_X1 u_majority7_module_105__and_module_8_U1 ( .A1(
        n_majority7_module_105__or_module_5_res), .A2(
        n_majority7_module_105__and_module_6_res), .ZN(
        n_majority7_module_105__and_module_8_res) );
  OR2_X1 u_majority7_module_105__or_module_9_U1 ( .A1(
        n_majority7_module_105__and_module_6_res), .A2(
        n_majority7_module_105__or_module_5_res), .ZN(
        n_majority7_module_105__or_module_9_res) );
  OR2_X1 u_majority7_module_105__or_module_10_U1 ( .A1(
        n_majority7_module_105__or_module_7_res), .A2(
        n_majority7_module_105__and_module_7_res), .ZN(
        n_majority7_module_105__or_module_10_res) );
  AND2_X1 u_majority7_module_105__and_module_9_U1 ( .A1(
        n_majority7_module_105__or_module_6_res), .A2(
        n_majority7_module_105__or_module_9_res), .ZN(
        n_majority7_module_105__and_module_9_res) );
  OR2_X1 u_majority7_module_105__or_module_11_U1 ( .A1(
        n_majority7_module_105__or_module_10_res), .A2(
        n_majority7_module_105__and_module_8_res), .ZN(
        n_majority7_module_105__or_module_11_res) );
  AND2_X1 u_majority7_module_105__and_module_10_U1 ( .A1(
        n_majority7_module_105__or_module_8_res), .A2(
        n_majority7_module_105__and_module_9_res), .ZN(
        n_majority7_module_105__and_module_10_res) );
  AND2_X1 u_majority7_module_105__and_module_11_U1 ( .A1(
        n_majority7_module_105__and_module_10_res), .A2(
        n_majority7_module_105__or_module_11_res), .ZN(
        n_majority7_module_105_res) );
  DFF_X1 u_reg_module_132__cini_mul_v00_reg ( .D(n_majority7_module_105_res), 
        .CK(clock_6), .Q(n_reg_module_132_res), .QN() );
  AND2_X1 u_majority7_module_106__and_module_1_U1 ( .A1(n_xor_module_163_res), 
        .A2(n_xor_module_91_res), .ZN(n_majority7_module_106__and_module_1_res) );
  OR2_X1 u_majority7_module_106__or_module_1_U1 ( .A1(n_xor_module_91_res), 
        .A2(n_xor_module_163_res), .ZN(n_majority7_module_106__or_module_1_res) );
  AND2_X1 u_majority7_module_106__and_module_2_U1 ( .A1(n_xor_module_127_res), 
        .A2(n_xor_module_115_res), .ZN(
        n_majority7_module_106__and_module_2_res) );
  OR2_X1 u_majority7_module_106__or_module_2_U1 ( .A1(n_xor_module_115_res), 
        .A2(n_xor_module_127_res), .ZN(n_majority7_module_106__or_module_2_res) );
  AND2_X1 u_majority7_module_106__and_module_3_U1 ( .A1(n_xor_module_151_res), 
        .A2(n_xor_module_139_res), .ZN(
        n_majority7_module_106__and_module_3_res) );
  OR2_X1 u_majority7_module_106__or_module_3_U1 ( .A1(n_xor_module_139_res), 
        .A2(n_xor_module_151_res), .ZN(n_majority7_module_106__or_module_3_res) );
  AND2_X1 u_majority7_module_106__and_module_4_U1 ( .A1(
        n_majority7_module_106__and_module_2_res), .A2(
        n_majority7_module_106__and_module_1_res), .ZN(
        n_majority7_module_106__and_module_4_res) );
  OR2_X1 u_majority7_module_106__or_module_4_U1 ( .A1(
        n_majority7_module_106__and_module_1_res), .A2(
        n_majority7_module_106__and_module_2_res), .ZN(
        n_majority7_module_106__or_module_4_res) );
  AND2_X1 u_majority7_module_106__and_module_5_U1 ( .A1(
        n_majority7_module_106__and_module_3_res), .A2(n_xor_module_103_res), 
        .ZN(n_majority7_module_106__and_module_5_res) );
  OR2_X1 u_majority7_module_106__or_module_5_U1 ( .A1(n_xor_module_103_res), 
        .A2(n_majority7_module_106__and_module_3_res), .ZN(
        n_majority7_module_106__or_module_5_res) );
  AND2_X1 u_majority7_module_106__and_module_6_U1 ( .A1(
        n_majority7_module_106__or_module_1_res), .A2(
        n_majority7_module_106__or_module_2_res), .ZN(
        n_majority7_module_106__and_module_6_res) );
  OR2_X1 u_majority7_module_106__or_module_6_U1 ( .A1(
        n_majority7_module_106__or_module_2_res), .A2(
        n_majority7_module_106__or_module_1_res), .ZN(
        n_majority7_module_106__or_module_6_res) );
  OR2_X1 u_majority7_module_106__or_module_7_U1 ( .A1(
        n_majority7_module_106__and_module_4_res), .A2(
        n_majority7_module_106__and_module_5_res), .ZN(
        n_majority7_module_106__or_module_7_res) );
  AND2_X1 u_majority7_module_106__and_module_7_U1 ( .A1(
        n_majority7_module_106__or_module_3_res), .A2(
        n_majority7_module_106__or_module_4_res), .ZN(
        n_majority7_module_106__and_module_7_res) );
  OR2_X1 u_majority7_module_106__or_module_8_U1 ( .A1(
        n_majority7_module_106__or_module_4_res), .A2(
        n_majority7_module_106__or_module_3_res), .ZN(
        n_majority7_module_106__or_module_8_res) );
  AND2_X1 u_majority7_module_106__and_module_8_U1 ( .A1(
        n_majority7_module_106__or_module_5_res), .A2(
        n_majority7_module_106__and_module_6_res), .ZN(
        n_majority7_module_106__and_module_8_res) );
  OR2_X1 u_majority7_module_106__or_module_9_U1 ( .A1(
        n_majority7_module_106__and_module_6_res), .A2(
        n_majority7_module_106__or_module_5_res), .ZN(
        n_majority7_module_106__or_module_9_res) );
  OR2_X1 u_majority7_module_106__or_module_10_U1 ( .A1(
        n_majority7_module_106__or_module_7_res), .A2(
        n_majority7_module_106__and_module_7_res), .ZN(
        n_majority7_module_106__or_module_10_res) );
  AND2_X1 u_majority7_module_106__and_module_9_U1 ( .A1(
        n_majority7_module_106__or_module_6_res), .A2(
        n_majority7_module_106__or_module_9_res), .ZN(
        n_majority7_module_106__and_module_9_res) );
  OR2_X1 u_majority7_module_106__or_module_11_U1 ( .A1(
        n_majority7_module_106__or_module_10_res), .A2(
        n_majority7_module_106__and_module_8_res), .ZN(
        n_majority7_module_106__or_module_11_res) );
  AND2_X1 u_majority7_module_106__and_module_10_U1 ( .A1(
        n_majority7_module_106__or_module_8_res), .A2(
        n_majority7_module_106__and_module_9_res), .ZN(
        n_majority7_module_106__and_module_10_res) );
  AND2_X1 u_majority7_module_106__and_module_11_U1 ( .A1(
        n_majority7_module_106__and_module_10_res), .A2(
        n_majority7_module_106__or_module_11_res), .ZN(
        n_majority7_module_106_res) );
  DFF_X1 u_reg_module_133__cini_mul_v00_reg ( .D(n_majority7_module_106_res), 
        .CK(clock_6), .Q(n_reg_module_133_res), .QN() );
  AND2_X1 u_majority7_module_107__and_module_1_U1 ( .A1(n_xor_module_164_res), 
        .A2(n_xor_module_92_res), .ZN(n_majority7_module_107__and_module_1_res) );
  OR2_X1 u_majority7_module_107__or_module_1_U1 ( .A1(n_xor_module_92_res), 
        .A2(n_xor_module_164_res), .ZN(n_majority7_module_107__or_module_1_res) );
  AND2_X1 u_majority7_module_107__and_module_2_U1 ( .A1(n_xor_module_128_res), 
        .A2(n_xor_module_116_res), .ZN(
        n_majority7_module_107__and_module_2_res) );
  OR2_X1 u_majority7_module_107__or_module_2_U1 ( .A1(n_xor_module_116_res), 
        .A2(n_xor_module_128_res), .ZN(n_majority7_module_107__or_module_2_res) );
  AND2_X1 u_majority7_module_107__and_module_3_U1 ( .A1(n_xor_module_152_res), 
        .A2(n_xor_module_140_res), .ZN(
        n_majority7_module_107__and_module_3_res) );
  OR2_X1 u_majority7_module_107__or_module_3_U1 ( .A1(n_xor_module_140_res), 
        .A2(n_xor_module_152_res), .ZN(n_majority7_module_107__or_module_3_res) );
  AND2_X1 u_majority7_module_107__and_module_4_U1 ( .A1(
        n_majority7_module_107__and_module_2_res), .A2(
        n_majority7_module_107__and_module_1_res), .ZN(
        n_majority7_module_107__and_module_4_res) );
  OR2_X1 u_majority7_module_107__or_module_4_U1 ( .A1(
        n_majority7_module_107__and_module_1_res), .A2(
        n_majority7_module_107__and_module_2_res), .ZN(
        n_majority7_module_107__or_module_4_res) );
  AND2_X1 u_majority7_module_107__and_module_5_U1 ( .A1(
        n_majority7_module_107__and_module_3_res), .A2(n_xor_module_104_res), 
        .ZN(n_majority7_module_107__and_module_5_res) );
  OR2_X1 u_majority7_module_107__or_module_5_U1 ( .A1(n_xor_module_104_res), 
        .A2(n_majority7_module_107__and_module_3_res), .ZN(
        n_majority7_module_107__or_module_5_res) );
  AND2_X1 u_majority7_module_107__and_module_6_U1 ( .A1(
        n_majority7_module_107__or_module_1_res), .A2(
        n_majority7_module_107__or_module_2_res), .ZN(
        n_majority7_module_107__and_module_6_res) );
  OR2_X1 u_majority7_module_107__or_module_6_U1 ( .A1(
        n_majority7_module_107__or_module_2_res), .A2(
        n_majority7_module_107__or_module_1_res), .ZN(
        n_majority7_module_107__or_module_6_res) );
  OR2_X1 u_majority7_module_107__or_module_7_U1 ( .A1(
        n_majority7_module_107__and_module_4_res), .A2(
        n_majority7_module_107__and_module_5_res), .ZN(
        n_majority7_module_107__or_module_7_res) );
  AND2_X1 u_majority7_module_107__and_module_7_U1 ( .A1(
        n_majority7_module_107__or_module_3_res), .A2(
        n_majority7_module_107__or_module_4_res), .ZN(
        n_majority7_module_107__and_module_7_res) );
  OR2_X1 u_majority7_module_107__or_module_8_U1 ( .A1(
        n_majority7_module_107__or_module_4_res), .A2(
        n_majority7_module_107__or_module_3_res), .ZN(
        n_majority7_module_107__or_module_8_res) );
  AND2_X1 u_majority7_module_107__and_module_8_U1 ( .A1(
        n_majority7_module_107__or_module_5_res), .A2(
        n_majority7_module_107__and_module_6_res), .ZN(
        n_majority7_module_107__and_module_8_res) );
  OR2_X1 u_majority7_module_107__or_module_9_U1 ( .A1(
        n_majority7_module_107__and_module_6_res), .A2(
        n_majority7_module_107__or_module_5_res), .ZN(
        n_majority7_module_107__or_module_9_res) );
  OR2_X1 u_majority7_module_107__or_module_10_U1 ( .A1(
        n_majority7_module_107__or_module_7_res), .A2(
        n_majority7_module_107__and_module_7_res), .ZN(
        n_majority7_module_107__or_module_10_res) );
  AND2_X1 u_majority7_module_107__and_module_9_U1 ( .A1(
        n_majority7_module_107__or_module_6_res), .A2(
        n_majority7_module_107__or_module_9_res), .ZN(
        n_majority7_module_107__and_module_9_res) );
  OR2_X1 u_majority7_module_107__or_module_11_U1 ( .A1(
        n_majority7_module_107__or_module_10_res), .A2(
        n_majority7_module_107__and_module_8_res), .ZN(
        n_majority7_module_107__or_module_11_res) );
  AND2_X1 u_majority7_module_107__and_module_10_U1 ( .A1(
        n_majority7_module_107__or_module_8_res), .A2(
        n_majority7_module_107__and_module_9_res), .ZN(
        n_majority7_module_107__and_module_10_res) );
  AND2_X1 u_majority7_module_107__and_module_11_U1 ( .A1(
        n_majority7_module_107__and_module_10_res), .A2(
        n_majority7_module_107__or_module_11_res), .ZN(
        n_majority7_module_107_res) );
  DFF_X1 u_reg_module_134__cini_mul_v00_reg ( .D(n_majority7_module_107_res), 
        .CK(clock_6), .Q(n_reg_module_134_res), .QN() );
  DFF_X1 u_reg_module_135__cini_mul_v00_reg ( .D(n_and_module_107_res), .CK(
        clock_6), .Q(n_reg_module_135_res), .QN() );
  AND2_X1 u_majority7_module_108__and_module_1_U1 ( .A1(n_xor_module_165_res), 
        .A2(n_xor_module_93_res), .ZN(n_majority7_module_108__and_module_1_res) );
  OR2_X1 u_majority7_module_108__or_module_1_U1 ( .A1(n_xor_module_93_res), 
        .A2(n_xor_module_165_res), .ZN(n_majority7_module_108__or_module_1_res) );
  AND2_X1 u_majority7_module_108__and_module_2_U1 ( .A1(n_xor_module_129_res), 
        .A2(n_xor_module_117_res), .ZN(
        n_majority7_module_108__and_module_2_res) );
  OR2_X1 u_majority7_module_108__or_module_2_U1 ( .A1(n_xor_module_117_res), 
        .A2(n_xor_module_129_res), .ZN(n_majority7_module_108__or_module_2_res) );
  AND2_X1 u_majority7_module_108__and_module_3_U1 ( .A1(n_xor_module_153_res), 
        .A2(n_xor_module_141_res), .ZN(
        n_majority7_module_108__and_module_3_res) );
  OR2_X1 u_majority7_module_108__or_module_3_U1 ( .A1(n_xor_module_141_res), 
        .A2(n_xor_module_153_res), .ZN(n_majority7_module_108__or_module_3_res) );
  AND2_X1 u_majority7_module_108__and_module_4_U1 ( .A1(
        n_majority7_module_108__and_module_2_res), .A2(
        n_majority7_module_108__and_module_1_res), .ZN(
        n_majority7_module_108__and_module_4_res) );
  OR2_X1 u_majority7_module_108__or_module_4_U1 ( .A1(
        n_majority7_module_108__and_module_1_res), .A2(
        n_majority7_module_108__and_module_2_res), .ZN(
        n_majority7_module_108__or_module_4_res) );
  AND2_X1 u_majority7_module_108__and_module_5_U1 ( .A1(
        n_majority7_module_108__and_module_3_res), .A2(n_xor_module_105_res), 
        .ZN(n_majority7_module_108__and_module_5_res) );
  OR2_X1 u_majority7_module_108__or_module_5_U1 ( .A1(n_xor_module_105_res), 
        .A2(n_majority7_module_108__and_module_3_res), .ZN(
        n_majority7_module_108__or_module_5_res) );
  AND2_X1 u_majority7_module_108__and_module_6_U1 ( .A1(
        n_majority7_module_108__or_module_1_res), .A2(
        n_majority7_module_108__or_module_2_res), .ZN(
        n_majority7_module_108__and_module_6_res) );
  OR2_X1 u_majority7_module_108__or_module_6_U1 ( .A1(
        n_majority7_module_108__or_module_2_res), .A2(
        n_majority7_module_108__or_module_1_res), .ZN(
        n_majority7_module_108__or_module_6_res) );
  OR2_X1 u_majority7_module_108__or_module_7_U1 ( .A1(
        n_majority7_module_108__and_module_4_res), .A2(
        n_majority7_module_108__and_module_5_res), .ZN(
        n_majority7_module_108__or_module_7_res) );
  AND2_X1 u_majority7_module_108__and_module_7_U1 ( .A1(
        n_majority7_module_108__or_module_3_res), .A2(
        n_majority7_module_108__or_module_4_res), .ZN(
        n_majority7_module_108__and_module_7_res) );
  OR2_X1 u_majority7_module_108__or_module_8_U1 ( .A1(
        n_majority7_module_108__or_module_4_res), .A2(
        n_majority7_module_108__or_module_3_res), .ZN(
        n_majority7_module_108__or_module_8_res) );
  AND2_X1 u_majority7_module_108__and_module_8_U1 ( .A1(
        n_majority7_module_108__or_module_5_res), .A2(
        n_majority7_module_108__and_module_6_res), .ZN(
        n_majority7_module_108__and_module_8_res) );
  OR2_X1 u_majority7_module_108__or_module_9_U1 ( .A1(
        n_majority7_module_108__and_module_6_res), .A2(
        n_majority7_module_108__or_module_5_res), .ZN(
        n_majority7_module_108__or_module_9_res) );
  OR2_X1 u_majority7_module_108__or_module_10_U1 ( .A1(
        n_majority7_module_108__or_module_7_res), .A2(
        n_majority7_module_108__and_module_7_res), .ZN(
        n_majority7_module_108__or_module_10_res) );
  AND2_X1 u_majority7_module_108__and_module_9_U1 ( .A1(
        n_majority7_module_108__or_module_6_res), .A2(
        n_majority7_module_108__or_module_9_res), .ZN(
        n_majority7_module_108__and_module_9_res) );
  OR2_X1 u_majority7_module_108__or_module_11_U1 ( .A1(
        n_majority7_module_108__or_module_10_res), .A2(
        n_majority7_module_108__and_module_8_res), .ZN(
        n_majority7_module_108__or_module_11_res) );
  AND2_X1 u_majority7_module_108__and_module_10_U1 ( .A1(
        n_majority7_module_108__or_module_8_res), .A2(
        n_majority7_module_108__and_module_9_res), .ZN(
        n_majority7_module_108__and_module_10_res) );
  AND2_X1 u_majority7_module_108__and_module_11_U1 ( .A1(
        n_majority7_module_108__and_module_10_res), .A2(
        n_majority7_module_108__or_module_11_res), .ZN(
        n_majority7_module_108_res) );
  DFF_X1 u_reg_module_136__cini_mul_v00_reg ( .D(n_majority7_module_108_res), 
        .CK(clock_6), .Q(n_reg_module_136_res), .QN() );
  AND2_X1 u_majority7_module_109__and_module_1_U1 ( .A1(n_xor_module_166_res), 
        .A2(n_xor_module_94_res), .ZN(n_majority7_module_109__and_module_1_res) );
  OR2_X1 u_majority7_module_109__or_module_1_U1 ( .A1(n_xor_module_94_res), 
        .A2(n_xor_module_166_res), .ZN(n_majority7_module_109__or_module_1_res) );
  AND2_X1 u_majority7_module_109__and_module_2_U1 ( .A1(n_xor_module_130_res), 
        .A2(n_xor_module_118_res), .ZN(
        n_majority7_module_109__and_module_2_res) );
  OR2_X1 u_majority7_module_109__or_module_2_U1 ( .A1(n_xor_module_118_res), 
        .A2(n_xor_module_130_res), .ZN(n_majority7_module_109__or_module_2_res) );
  AND2_X1 u_majority7_module_109__and_module_3_U1 ( .A1(n_xor_module_154_res), 
        .A2(n_xor_module_142_res), .ZN(
        n_majority7_module_109__and_module_3_res) );
  OR2_X1 u_majority7_module_109__or_module_3_U1 ( .A1(n_xor_module_142_res), 
        .A2(n_xor_module_154_res), .ZN(n_majority7_module_109__or_module_3_res) );
  AND2_X1 u_majority7_module_109__and_module_4_U1 ( .A1(
        n_majority7_module_109__and_module_2_res), .A2(
        n_majority7_module_109__and_module_1_res), .ZN(
        n_majority7_module_109__and_module_4_res) );
  OR2_X1 u_majority7_module_109__or_module_4_U1 ( .A1(
        n_majority7_module_109__and_module_1_res), .A2(
        n_majority7_module_109__and_module_2_res), .ZN(
        n_majority7_module_109__or_module_4_res) );
  AND2_X1 u_majority7_module_109__and_module_5_U1 ( .A1(
        n_majority7_module_109__and_module_3_res), .A2(n_xor_module_106_res), 
        .ZN(n_majority7_module_109__and_module_5_res) );
  OR2_X1 u_majority7_module_109__or_module_5_U1 ( .A1(n_xor_module_106_res), 
        .A2(n_majority7_module_109__and_module_3_res), .ZN(
        n_majority7_module_109__or_module_5_res) );
  AND2_X1 u_majority7_module_109__and_module_6_U1 ( .A1(
        n_majority7_module_109__or_module_1_res), .A2(
        n_majority7_module_109__or_module_2_res), .ZN(
        n_majority7_module_109__and_module_6_res) );
  OR2_X1 u_majority7_module_109__or_module_6_U1 ( .A1(
        n_majority7_module_109__or_module_2_res), .A2(
        n_majority7_module_109__or_module_1_res), .ZN(
        n_majority7_module_109__or_module_6_res) );
  OR2_X1 u_majority7_module_109__or_module_7_U1 ( .A1(
        n_majority7_module_109__and_module_4_res), .A2(
        n_majority7_module_109__and_module_5_res), .ZN(
        n_majority7_module_109__or_module_7_res) );
  AND2_X1 u_majority7_module_109__and_module_7_U1 ( .A1(
        n_majority7_module_109__or_module_3_res), .A2(
        n_majority7_module_109__or_module_4_res), .ZN(
        n_majority7_module_109__and_module_7_res) );
  OR2_X1 u_majority7_module_109__or_module_8_U1 ( .A1(
        n_majority7_module_109__or_module_4_res), .A2(
        n_majority7_module_109__or_module_3_res), .ZN(
        n_majority7_module_109__or_module_8_res) );
  AND2_X1 u_majority7_module_109__and_module_8_U1 ( .A1(
        n_majority7_module_109__or_module_5_res), .A2(
        n_majority7_module_109__and_module_6_res), .ZN(
        n_majority7_module_109__and_module_8_res) );
  OR2_X1 u_majority7_module_109__or_module_9_U1 ( .A1(
        n_majority7_module_109__and_module_6_res), .A2(
        n_majority7_module_109__or_module_5_res), .ZN(
        n_majority7_module_109__or_module_9_res) );
  OR2_X1 u_majority7_module_109__or_module_10_U1 ( .A1(
        n_majority7_module_109__or_module_7_res), .A2(
        n_majority7_module_109__and_module_7_res), .ZN(
        n_majority7_module_109__or_module_10_res) );
  AND2_X1 u_majority7_module_109__and_module_9_U1 ( .A1(
        n_majority7_module_109__or_module_6_res), .A2(
        n_majority7_module_109__or_module_9_res), .ZN(
        n_majority7_module_109__and_module_9_res) );
  OR2_X1 u_majority7_module_109__or_module_11_U1 ( .A1(
        n_majority7_module_109__or_module_10_res), .A2(
        n_majority7_module_109__and_module_8_res), .ZN(
        n_majority7_module_109__or_module_11_res) );
  AND2_X1 u_majority7_module_109__and_module_10_U1 ( .A1(
        n_majority7_module_109__or_module_8_res), .A2(
        n_majority7_module_109__and_module_9_res), .ZN(
        n_majority7_module_109__and_module_10_res) );
  AND2_X1 u_majority7_module_109__and_module_11_U1 ( .A1(
        n_majority7_module_109__and_module_10_res), .A2(
        n_majority7_module_109__or_module_11_res), .ZN(
        n_majority7_module_109_res) );
  DFF_X1 u_reg_module_137__cini_mul_v00_reg ( .D(n_majority7_module_109_res), 
        .CK(clock_6), .Q(n_reg_module_137_res), .QN() );
  AND2_X1 u_majority7_module_110__and_module_1_U1 ( .A1(n_xor_module_167_res), 
        .A2(n_xor_module_95_res), .ZN(n_majority7_module_110__and_module_1_res) );
  OR2_X1 u_majority7_module_110__or_module_1_U1 ( .A1(n_xor_module_95_res), 
        .A2(n_xor_module_167_res), .ZN(n_majority7_module_110__or_module_1_res) );
  AND2_X1 u_majority7_module_110__and_module_2_U1 ( .A1(n_xor_module_131_res), 
        .A2(n_xor_module_119_res), .ZN(
        n_majority7_module_110__and_module_2_res) );
  OR2_X1 u_majority7_module_110__or_module_2_U1 ( .A1(n_xor_module_119_res), 
        .A2(n_xor_module_131_res), .ZN(n_majority7_module_110__or_module_2_res) );
  AND2_X1 u_majority7_module_110__and_module_3_U1 ( .A1(n_xor_module_155_res), 
        .A2(n_xor_module_143_res), .ZN(
        n_majority7_module_110__and_module_3_res) );
  OR2_X1 u_majority7_module_110__or_module_3_U1 ( .A1(n_xor_module_143_res), 
        .A2(n_xor_module_155_res), .ZN(n_majority7_module_110__or_module_3_res) );
  AND2_X1 u_majority7_module_110__and_module_4_U1 ( .A1(
        n_majority7_module_110__and_module_2_res), .A2(
        n_majority7_module_110__and_module_1_res), .ZN(
        n_majority7_module_110__and_module_4_res) );
  OR2_X1 u_majority7_module_110__or_module_4_U1 ( .A1(
        n_majority7_module_110__and_module_1_res), .A2(
        n_majority7_module_110__and_module_2_res), .ZN(
        n_majority7_module_110__or_module_4_res) );
  AND2_X1 u_majority7_module_110__and_module_5_U1 ( .A1(
        n_majority7_module_110__and_module_3_res), .A2(n_xor_module_107_res), 
        .ZN(n_majority7_module_110__and_module_5_res) );
  OR2_X1 u_majority7_module_110__or_module_5_U1 ( .A1(n_xor_module_107_res), 
        .A2(n_majority7_module_110__and_module_3_res), .ZN(
        n_majority7_module_110__or_module_5_res) );
  AND2_X1 u_majority7_module_110__and_module_6_U1 ( .A1(
        n_majority7_module_110__or_module_1_res), .A2(
        n_majority7_module_110__or_module_2_res), .ZN(
        n_majority7_module_110__and_module_6_res) );
  OR2_X1 u_majority7_module_110__or_module_6_U1 ( .A1(
        n_majority7_module_110__or_module_2_res), .A2(
        n_majority7_module_110__or_module_1_res), .ZN(
        n_majority7_module_110__or_module_6_res) );
  OR2_X1 u_majority7_module_110__or_module_7_U1 ( .A1(
        n_majority7_module_110__and_module_4_res), .A2(
        n_majority7_module_110__and_module_5_res), .ZN(
        n_majority7_module_110__or_module_7_res) );
  AND2_X1 u_majority7_module_110__and_module_7_U1 ( .A1(
        n_majority7_module_110__or_module_3_res), .A2(
        n_majority7_module_110__or_module_4_res), .ZN(
        n_majority7_module_110__and_module_7_res) );
  OR2_X1 u_majority7_module_110__or_module_8_U1 ( .A1(
        n_majority7_module_110__or_module_4_res), .A2(
        n_majority7_module_110__or_module_3_res), .ZN(
        n_majority7_module_110__or_module_8_res) );
  AND2_X1 u_majority7_module_110__and_module_8_U1 ( .A1(
        n_majority7_module_110__or_module_5_res), .A2(
        n_majority7_module_110__and_module_6_res), .ZN(
        n_majority7_module_110__and_module_8_res) );
  OR2_X1 u_majority7_module_110__or_module_9_U1 ( .A1(
        n_majority7_module_110__and_module_6_res), .A2(
        n_majority7_module_110__or_module_5_res), .ZN(
        n_majority7_module_110__or_module_9_res) );
  OR2_X1 u_majority7_module_110__or_module_10_U1 ( .A1(
        n_majority7_module_110__or_module_7_res), .A2(
        n_majority7_module_110__and_module_7_res), .ZN(
        n_majority7_module_110__or_module_10_res) );
  AND2_X1 u_majority7_module_110__and_module_9_U1 ( .A1(
        n_majority7_module_110__or_module_6_res), .A2(
        n_majority7_module_110__or_module_9_res), .ZN(
        n_majority7_module_110__and_module_9_res) );
  OR2_X1 u_majority7_module_110__or_module_11_U1 ( .A1(
        n_majority7_module_110__or_module_10_res), .A2(
        n_majority7_module_110__and_module_8_res), .ZN(
        n_majority7_module_110__or_module_11_res) );
  AND2_X1 u_majority7_module_110__and_module_10_U1 ( .A1(
        n_majority7_module_110__or_module_8_res), .A2(
        n_majority7_module_110__and_module_9_res), .ZN(
        n_majority7_module_110__and_module_10_res) );
  AND2_X1 u_majority7_module_110__and_module_11_U1 ( .A1(
        n_majority7_module_110__and_module_10_res), .A2(
        n_majority7_module_110__or_module_11_res), .ZN(
        n_majority7_module_110_res) );
  DFF_X1 u_reg_module_138__cini_mul_v00_reg ( .D(n_majority7_module_110_res), 
        .CK(clock_6), .Q(n_reg_module_138_res), .QN() );
  AND2_X1 u_majority7_module_111__and_module_1_U1 ( .A1(n_xor_module_168_res), 
        .A2(n_xor_module_96_res), .ZN(n_majority7_module_111__and_module_1_res) );
  OR2_X1 u_majority7_module_111__or_module_1_U1 ( .A1(n_xor_module_96_res), 
        .A2(n_xor_module_168_res), .ZN(n_majority7_module_111__or_module_1_res) );
  AND2_X1 u_majority7_module_111__and_module_2_U1 ( .A1(n_xor_module_132_res), 
        .A2(n_xor_module_120_res), .ZN(
        n_majority7_module_111__and_module_2_res) );
  OR2_X1 u_majority7_module_111__or_module_2_U1 ( .A1(n_xor_module_120_res), 
        .A2(n_xor_module_132_res), .ZN(n_majority7_module_111__or_module_2_res) );
  AND2_X1 u_majority7_module_111__and_module_3_U1 ( .A1(n_xor_module_156_res), 
        .A2(n_xor_module_144_res), .ZN(
        n_majority7_module_111__and_module_3_res) );
  OR2_X1 u_majority7_module_111__or_module_3_U1 ( .A1(n_xor_module_144_res), 
        .A2(n_xor_module_156_res), .ZN(n_majority7_module_111__or_module_3_res) );
  AND2_X1 u_majority7_module_111__and_module_4_U1 ( .A1(
        n_majority7_module_111__and_module_2_res), .A2(
        n_majority7_module_111__and_module_1_res), .ZN(
        n_majority7_module_111__and_module_4_res) );
  OR2_X1 u_majority7_module_111__or_module_4_U1 ( .A1(
        n_majority7_module_111__and_module_1_res), .A2(
        n_majority7_module_111__and_module_2_res), .ZN(
        n_majority7_module_111__or_module_4_res) );
  AND2_X1 u_majority7_module_111__and_module_5_U1 ( .A1(
        n_majority7_module_111__and_module_3_res), .A2(n_xor_module_108_res), 
        .ZN(n_majority7_module_111__and_module_5_res) );
  OR2_X1 u_majority7_module_111__or_module_5_U1 ( .A1(n_xor_module_108_res), 
        .A2(n_majority7_module_111__and_module_3_res), .ZN(
        n_majority7_module_111__or_module_5_res) );
  AND2_X1 u_majority7_module_111__and_module_6_U1 ( .A1(
        n_majority7_module_111__or_module_1_res), .A2(
        n_majority7_module_111__or_module_2_res), .ZN(
        n_majority7_module_111__and_module_6_res) );
  OR2_X1 u_majority7_module_111__or_module_6_U1 ( .A1(
        n_majority7_module_111__or_module_2_res), .A2(
        n_majority7_module_111__or_module_1_res), .ZN(
        n_majority7_module_111__or_module_6_res) );
  OR2_X1 u_majority7_module_111__or_module_7_U1 ( .A1(
        n_majority7_module_111__and_module_4_res), .A2(
        n_majority7_module_111__and_module_5_res), .ZN(
        n_majority7_module_111__or_module_7_res) );
  AND2_X1 u_majority7_module_111__and_module_7_U1 ( .A1(
        n_majority7_module_111__or_module_3_res), .A2(
        n_majority7_module_111__or_module_4_res), .ZN(
        n_majority7_module_111__and_module_7_res) );
  OR2_X1 u_majority7_module_111__or_module_8_U1 ( .A1(
        n_majority7_module_111__or_module_4_res), .A2(
        n_majority7_module_111__or_module_3_res), .ZN(
        n_majority7_module_111__or_module_8_res) );
  AND2_X1 u_majority7_module_111__and_module_8_U1 ( .A1(
        n_majority7_module_111__or_module_5_res), .A2(
        n_majority7_module_111__and_module_6_res), .ZN(
        n_majority7_module_111__and_module_8_res) );
  OR2_X1 u_majority7_module_111__or_module_9_U1 ( .A1(
        n_majority7_module_111__and_module_6_res), .A2(
        n_majority7_module_111__or_module_5_res), .ZN(
        n_majority7_module_111__or_module_9_res) );
  OR2_X1 u_majority7_module_111__or_module_10_U1 ( .A1(
        n_majority7_module_111__or_module_7_res), .A2(
        n_majority7_module_111__and_module_7_res), .ZN(
        n_majority7_module_111__or_module_10_res) );
  AND2_X1 u_majority7_module_111__and_module_9_U1 ( .A1(
        n_majority7_module_111__or_module_6_res), .A2(
        n_majority7_module_111__or_module_9_res), .ZN(
        n_majority7_module_111__and_module_9_res) );
  OR2_X1 u_majority7_module_111__or_module_11_U1 ( .A1(
        n_majority7_module_111__or_module_10_res), .A2(
        n_majority7_module_111__and_module_8_res), .ZN(
        n_majority7_module_111__or_module_11_res) );
  AND2_X1 u_majority7_module_111__and_module_10_U1 ( .A1(
        n_majority7_module_111__or_module_8_res), .A2(
        n_majority7_module_111__and_module_9_res), .ZN(
        n_majority7_module_111__and_module_10_res) );
  AND2_X1 u_majority7_module_111__and_module_11_U1 ( .A1(
        n_majority7_module_111__and_module_10_res), .A2(
        n_majority7_module_111__or_module_11_res), .ZN(
        n_majority7_module_111_res) );
  DFF_X1 u_reg_module_139__cini_mul_v00_reg ( .D(n_majority7_module_111_res), 
        .CK(clock_6), .Q(n_reg_module_139_res), .QN() );
  DFF_X1 u_reg_module_140__cini_mul_v00_reg ( .D(n_and_module_112_res), .CK(
        clock_6), .Q(n_reg_module_140_res), .QN() );
  XOR2_X1 u_xor_module_169_U1 ( .A(n_reg_module_30_res), .B(
        n_reg_module_29_res), .Z(n_xor_module_169_res) );
  XOR2_X1 u_xor_module_170_U1 ( .A(n_reg_module_31_res), .B(
        n_xor_module_169_res), .Z(n_xor_module_170_res) );
  XOR2_X1 u_xor_module_171_U1 ( .A(n_reg_module_32_res), .B(
        n_xor_module_170_res), .Z(io_o0_s0_d0) );
  XOR2_X1 u_xor_module_172_U1 ( .A(n_reg_module_33_res), .B(
        n_reg_module_34_res), .Z(n_xor_module_172_res) );
  XOR2_X1 u_xor_module_173_U1 ( .A(n_reg_module_35_res), .B(
        n_xor_module_172_res), .Z(n_xor_module_173_res) );
  XOR2_X1 u_xor_module_174_U1 ( .A(n_reg_module_36_res), .B(
        n_xor_module_173_res), .Z(io_o0_s1_d0) );
  XOR2_X1 u_xor_module_175_U1 ( .A(n_reg_module_37_res), .B(
        n_reg_module_39_res), .Z(n_xor_module_175_res) );
  XOR2_X1 u_xor_module_176_U1 ( .A(n_reg_module_38_res), .B(
        n_xor_module_175_res), .Z(n_xor_module_176_res) );
  XOR2_X1 u_xor_module_177_U1 ( .A(n_reg_module_40_res), .B(
        n_xor_module_176_res), .Z(io_o0_s2_d0) );
  XOR2_X1 u_xor_module_178_U1 ( .A(n_reg_module_41_res), .B(
        n_reg_module_44_res), .Z(n_xor_module_178_res) );
  XOR2_X1 u_xor_module_179_U1 ( .A(n_reg_module_42_res), .B(
        n_xor_module_178_res), .Z(n_xor_module_179_res) );
  XOR2_X1 u_xor_module_180_U1 ( .A(n_reg_module_43_res), .B(
        n_xor_module_179_res), .Z(io_o0_s3_d0) );
  XOR2_X1 u_xor_module_181_U1 ( .A(n_reg_module_46_res), .B(
        n_reg_module_45_res), .Z(n_xor_module_181_res) );
  XOR2_X1 u_xor_module_182_U1 ( .A(n_reg_module_47_res), .B(
        n_xor_module_181_res), .Z(n_xor_module_182_res) );
  XOR2_X1 u_xor_module_183_U1 ( .A(n_reg_module_48_res), .B(
        n_xor_module_182_res), .Z(io_o0_s0_d1) );
  XOR2_X1 u_xor_module_184_U1 ( .A(n_reg_module_49_res), .B(
        n_reg_module_50_res), .Z(n_xor_module_184_res) );
  XOR2_X1 u_xor_module_185_U1 ( .A(n_reg_module_51_res), .B(
        n_xor_module_184_res), .Z(n_xor_module_185_res) );
  XOR2_X1 u_xor_module_186_U1 ( .A(n_reg_module_52_res), .B(
        n_xor_module_185_res), .Z(io_o0_s1_d1) );
  XOR2_X1 u_xor_module_187_U1 ( .A(n_reg_module_53_res), .B(
        n_reg_module_55_res), .Z(n_xor_module_187_res) );
  XOR2_X1 u_xor_module_188_U1 ( .A(n_reg_module_54_res), .B(
        n_xor_module_187_res), .Z(n_xor_module_188_res) );
  XOR2_X1 u_xor_module_189_U1 ( .A(n_reg_module_56_res), .B(
        n_xor_module_188_res), .Z(io_o0_s2_d1) );
  XOR2_X1 u_xor_module_190_U1 ( .A(n_reg_module_57_res), .B(
        n_reg_module_60_res), .Z(n_xor_module_190_res) );
  XOR2_X1 u_xor_module_191_U1 ( .A(n_reg_module_58_res), .B(
        n_xor_module_190_res), .Z(n_xor_module_191_res) );
  XOR2_X1 u_xor_module_192_U1 ( .A(n_reg_module_59_res), .B(
        n_xor_module_191_res), .Z(io_o0_s3_d1) );
  XOR2_X1 u_xor_module_193_U1 ( .A(n_reg_module_62_res), .B(
        n_reg_module_61_res), .Z(n_xor_module_193_res) );
  XOR2_X1 u_xor_module_194_U1 ( .A(n_reg_module_63_res), .B(
        n_xor_module_193_res), .Z(n_xor_module_194_res) );
  XOR2_X1 u_xor_module_195_U1 ( .A(n_reg_module_64_res), .B(
        n_xor_module_194_res), .Z(io_o0_s0_d2) );
  XOR2_X1 u_xor_module_196_U1 ( .A(n_reg_module_65_res), .B(
        n_reg_module_66_res), .Z(n_xor_module_196_res) );
  XOR2_X1 u_xor_module_197_U1 ( .A(n_reg_module_67_res), .B(
        n_xor_module_196_res), .Z(n_xor_module_197_res) );
  XOR2_X1 u_xor_module_198_U1 ( .A(n_reg_module_68_res), .B(
        n_xor_module_197_res), .Z(io_o0_s1_d2) );
  XOR2_X1 u_xor_module_199_U1 ( .A(n_reg_module_69_res), .B(
        n_reg_module_71_res), .Z(n_xor_module_199_res) );
  XOR2_X1 u_xor_module_200_U1 ( .A(n_reg_module_70_res), .B(
        n_xor_module_199_res), .Z(n_xor_module_200_res) );
  XOR2_X1 u_xor_module_201_U1 ( .A(n_reg_module_72_res), .B(
        n_xor_module_200_res), .Z(io_o0_s2_d2) );
  XOR2_X1 u_xor_module_202_U1 ( .A(n_reg_module_73_res), .B(
        n_reg_module_76_res), .Z(n_xor_module_202_res) );
  XOR2_X1 u_xor_module_203_U1 ( .A(n_reg_module_74_res), .B(
        n_xor_module_202_res), .Z(n_xor_module_203_res) );
  XOR2_X1 u_xor_module_204_U1 ( .A(n_reg_module_75_res), .B(
        n_xor_module_203_res), .Z(io_o0_s3_d2) );
  XOR2_X1 u_xor_module_205_U1 ( .A(n_reg_module_78_res), .B(
        n_reg_module_77_res), .Z(n_xor_module_205_res) );
  XOR2_X1 u_xor_module_206_U1 ( .A(n_reg_module_79_res), .B(
        n_xor_module_205_res), .Z(n_xor_module_206_res) );
  XOR2_X1 u_xor_module_207_U1 ( .A(n_reg_module_80_res), .B(
        n_xor_module_206_res), .Z(io_o0_s0_d3) );
  XOR2_X1 u_xor_module_208_U1 ( .A(n_reg_module_81_res), .B(
        n_reg_module_82_res), .Z(n_xor_module_208_res) );
  XOR2_X1 u_xor_module_209_U1 ( .A(n_reg_module_83_res), .B(
        n_xor_module_208_res), .Z(n_xor_module_209_res) );
  XOR2_X1 u_xor_module_210_U1 ( .A(n_reg_module_84_res), .B(
        n_xor_module_209_res), .Z(io_o0_s1_d3) );
  XOR2_X1 u_xor_module_211_U1 ( .A(n_reg_module_85_res), .B(
        n_reg_module_87_res), .Z(n_xor_module_211_res) );
  XOR2_X1 u_xor_module_212_U1 ( .A(n_reg_module_86_res), .B(
        n_xor_module_211_res), .Z(n_xor_module_212_res) );
  XOR2_X1 u_xor_module_213_U1 ( .A(n_reg_module_88_res), .B(
        n_xor_module_212_res), .Z(io_o0_s2_d3) );
  XOR2_X1 u_xor_module_214_U1 ( .A(n_reg_module_89_res), .B(
        n_reg_module_92_res), .Z(n_xor_module_214_res) );
  XOR2_X1 u_xor_module_215_U1 ( .A(n_reg_module_90_res), .B(
        n_xor_module_214_res), .Z(n_xor_module_215_res) );
  XOR2_X1 u_xor_module_216_U1 ( .A(n_reg_module_91_res), .B(
        n_xor_module_215_res), .Z(io_o0_s3_d3) );
  XOR2_X1 u_xor_module_217_U1 ( .A(n_reg_module_94_res), .B(
        n_reg_module_93_res), .Z(n_xor_module_217_res) );
  XOR2_X1 u_xor_module_218_U1 ( .A(n_reg_module_95_res), .B(
        n_xor_module_217_res), .Z(n_xor_module_218_res) );
  XOR2_X1 u_xor_module_219_U1 ( .A(n_reg_module_96_res), .B(
        n_xor_module_218_res), .Z(io_o0_s0_d4) );
  XOR2_X1 u_xor_module_220_U1 ( .A(n_reg_module_97_res), .B(
        n_reg_module_98_res), .Z(n_xor_module_220_res) );
  XOR2_X1 u_xor_module_221_U1 ( .A(n_reg_module_99_res), .B(
        n_xor_module_220_res), .Z(n_xor_module_221_res) );
  XOR2_X1 u_xor_module_222_U1 ( .A(n_reg_module_100_res), .B(
        n_xor_module_221_res), .Z(io_o0_s1_d4) );
  XOR2_X1 u_xor_module_223_U1 ( .A(n_reg_module_101_res), .B(
        n_reg_module_103_res), .Z(n_xor_module_223_res) );
  XOR2_X1 u_xor_module_224_U1 ( .A(n_reg_module_102_res), .B(
        n_xor_module_223_res), .Z(n_xor_module_224_res) );
  XOR2_X1 u_xor_module_225_U1 ( .A(n_reg_module_104_res), .B(
        n_xor_module_224_res), .Z(io_o0_s2_d4) );
  XOR2_X1 u_xor_module_226_U1 ( .A(n_reg_module_105_res), .B(
        n_reg_module_108_res), .Z(n_xor_module_226_res) );
  XOR2_X1 u_xor_module_227_U1 ( .A(n_reg_module_106_res), .B(
        n_xor_module_226_res), .Z(n_xor_module_227_res) );
  XOR2_X1 u_xor_module_228_U1 ( .A(n_reg_module_107_res), .B(
        n_xor_module_227_res), .Z(io_o0_s3_d4) );
  XOR2_X1 u_xor_module_229_U1 ( .A(n_reg_module_110_res), .B(
        n_reg_module_109_res), .Z(n_xor_module_229_res) );
  XOR2_X1 u_xor_module_230_U1 ( .A(n_reg_module_111_res), .B(
        n_xor_module_229_res), .Z(n_xor_module_230_res) );
  XOR2_X1 u_xor_module_231_U1 ( .A(n_reg_module_112_res), .B(
        n_xor_module_230_res), .Z(io_o0_s0_d5) );
  XOR2_X1 u_xor_module_232_U1 ( .A(n_reg_module_113_res), .B(
        n_reg_module_114_res), .Z(n_xor_module_232_res) );
  XOR2_X1 u_xor_module_233_U1 ( .A(n_reg_module_115_res), .B(
        n_xor_module_232_res), .Z(n_xor_module_233_res) );
  XOR2_X1 u_xor_module_234_U1 ( .A(n_reg_module_116_res), .B(
        n_xor_module_233_res), .Z(io_o0_s1_d5) );
  XOR2_X1 u_xor_module_235_U1 ( .A(n_reg_module_117_res), .B(
        n_reg_module_119_res), .Z(n_xor_module_235_res) );
  XOR2_X1 u_xor_module_236_U1 ( .A(n_reg_module_118_res), .B(
        n_xor_module_235_res), .Z(n_xor_module_236_res) );
  XOR2_X1 u_xor_module_237_U1 ( .A(n_reg_module_120_res), .B(
        n_xor_module_236_res), .Z(io_o0_s2_d5) );
  XOR2_X1 u_xor_module_238_U1 ( .A(n_reg_module_121_res), .B(
        n_reg_module_124_res), .Z(n_xor_module_238_res) );
  XOR2_X1 u_xor_module_239_U1 ( .A(n_reg_module_122_res), .B(
        n_xor_module_238_res), .Z(n_xor_module_239_res) );
  XOR2_X1 u_xor_module_240_U1 ( .A(n_reg_module_123_res), .B(
        n_xor_module_239_res), .Z(io_o0_s3_d5) );
  XOR2_X1 u_xor_module_241_U1 ( .A(n_reg_module_126_res), .B(
        n_reg_module_125_res), .Z(n_xor_module_241_res) );
  XOR2_X1 u_xor_module_242_U1 ( .A(n_reg_module_127_res), .B(
        n_xor_module_241_res), .Z(n_xor_module_242_res) );
  XOR2_X1 u_xor_module_243_U1 ( .A(n_reg_module_128_res), .B(
        n_xor_module_242_res), .Z(io_o0_s0_d6) );
  XOR2_X1 u_xor_module_244_U1 ( .A(n_reg_module_129_res), .B(
        n_reg_module_130_res), .Z(n_xor_module_244_res) );
  XOR2_X1 u_xor_module_245_U1 ( .A(n_reg_module_131_res), .B(
        n_xor_module_244_res), .Z(n_xor_module_245_res) );
  XOR2_X1 u_xor_module_246_U1 ( .A(n_reg_module_132_res), .B(
        n_xor_module_245_res), .Z(io_o0_s1_d6) );
  XOR2_X1 u_xor_module_247_U1 ( .A(n_reg_module_133_res), .B(
        n_reg_module_135_res), .Z(n_xor_module_247_res) );
  XOR2_X1 u_xor_module_248_U1 ( .A(n_reg_module_134_res), .B(
        n_xor_module_247_res), .Z(n_xor_module_248_res) );
  XOR2_X1 u_xor_module_249_U1 ( .A(n_reg_module_136_res), .B(
        n_xor_module_248_res), .Z(io_o0_s2_d6) );
  XOR2_X1 u_xor_module_250_U1 ( .A(n_reg_module_137_res), .B(
        n_reg_module_140_res), .Z(n_xor_module_250_res) );
  XOR2_X1 u_xor_module_251_U1 ( .A(n_reg_module_138_res), .B(
        n_xor_module_250_res), .Z(n_xor_module_251_res) );
  XOR2_X1 u_xor_module_252_U1 ( .A(n_reg_module_139_res), .B(
        n_xor_module_251_res), .Z(io_o0_s3_d6) );
endmodule

