module KeyAddition ( clock, reset, io_state, io_key, io_out );
  input [7:0] io_state;
  input [7:0] io_key;
  output [7:0] io_out;
  input clock, reset;


  XOR2_X1 U9 ( .A(io_state[7]), .B(io_key[7]), .Z(io_out[7]) );
  XOR2_X1 U10 ( .A(io_state[6]), .B(io_key[6]), .Z(io_out[6]) );
  XOR2_X1 U11 ( .A(io_state[5]), .B(io_key[5]), .Z(io_out[5]) );
  XOR2_X1 U12 ( .A(io_state[4]), .B(io_key[4]), .Z(io_out[4]) );
  XOR2_X1 U13 ( .A(io_state[3]), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 U14 ( .A(io_state[2]), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 U15 ( .A(io_state[1]), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 U16 ( .A(io_state[0]), .B(io_key[0]), .Z(io_out[0]) );
endmodule

