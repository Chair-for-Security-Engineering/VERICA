
module Shared_Chi3_SifaTest ( port_a_in, port_b_in, port_c_in, port_det_out );
  input [1:0] port_a_in;
  input [1:0] port_b_in;
  input [1:0] port_c_in;
  output [1:0] port_det_out;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, chi3_0_st0_t0_n2,
         chi3_0_st0_t0_n1, chi3_0_st0_t2_n1, chi3_0_st0_t1_n2,
         chi3_0_st0_t1_n1, chi3_0_st0_t3_n1, chi3_0_st1_t0_n2,
         chi3_0_st1_t0_n1, chi3_0_st1_t2_n1, chi3_0_st1_t1_n2,
         chi3_0_st1_t1_n1, chi3_0_st1_t3_n1, chi3_0_st2_t0_n2,
         chi3_0_st2_t0_n1, chi3_0_st2_t2_n1, chi3_0_st2_t1_n2,
         chi3_0_st2_t1_n1, chi3_0_st2_t3_n1, chi3_1_st0_t0_n2,
         chi3_1_st0_t0_n1, chi3_1_st0_t2_n1, chi3_1_st0_t1_n2,
         chi3_1_st0_t1_n1, chi3_1_st0_t3_n1, chi3_1_st1_t0_n2,
         chi3_1_st1_t0_n1, chi3_1_st1_t2_n1, chi3_1_st1_t1_n2,
         chi3_1_st1_t1_n1, chi3_1_st1_t3_n1, chi3_1_st2_t0_n2,
         chi3_1_st2_t0_n1, chi3_1_st2_t2_n1, chi3_1_st2_t1_n2,
         chi3_1_st2_t1_n1, chi3_1_st2_t3_n1;
  wire   [1:0] chi3_0_port_a_out;
  wire   [1:0] chi3_0_port_b_out;
  wire   [1:0] chi3_0_port_c_out;
  wire   [1:0] chi3_1_port_a_out;
  wire   [1:0] chi3_1_port_b_out;
  wire   [1:0] chi3_1_port_c_out;
  wire   [1:0] chi3_0_st0_a_temp;
  wire   [1:0] chi3_0_st1_a_temp;
  wire   [1:0] chi3_0_st2_a_temp;
  wire   [1:0] chi3_1_st0_a_temp;
  wire   [1:0] chi3_1_st1_a_temp;
  wire   [1:0] chi3_1_st2_a_temp;
  wire port_a_in0, port_a_in1;

  BUF_X1 B00 ( .A(port_a_in[0]), .Z(port_a_in0) );
  BUF_X1 B01 ( .A(port_a_in[1]), .Z(port_a_in1) );

  NOR2_X1 U11 ( .A1(n9), .A2(n10), .ZN(port_det_out[1]) );
  NAND2_X1 U12 ( .A1(n11), .A2(n12), .ZN(n10) );
  XNOR2_X1 U13 ( .A(chi3_1_port_c_out[1]), .B(chi3_0_port_c_out[1]), .ZN(n12)
         );
  XNOR2_X1 U14 ( .A(chi3_1_port_b_out[1]), .B(chi3_0_port_b_out[1]), .ZN(n11)
         );
  XOR2_X1 U15 ( .A(chi3_1_port_a_out[1]), .B(chi3_0_port_a_out[1]), .Z(n9) );
  NOR2_X1 U16 ( .A1(n13), .A2(n14), .ZN(port_det_out[0]) );
  NAND2_X1 U17 ( .A1(n15), .A2(n16), .ZN(n14) );
  XNOR2_X1 U18 ( .A(chi3_1_port_c_out[0]), .B(chi3_0_port_c_out[0]), .ZN(n16)
         );
  XNOR2_X1 U19 ( .A(chi3_1_port_b_out[0]), .B(chi3_0_port_b_out[0]), .ZN(n15)
         );
  XOR2_X1 U20 ( .A(chi3_1_port_a_out[0]), .B(chi3_0_port_a_out[0]), .Z(n13) );
  INV_X1 chi3_0_st0_t0_U3 ( .A(port_c_in[1]), .ZN(chi3_0_st0_t0_n2) );
  NOR2_X1 chi3_0_st0_t0_U2 ( .A1(port_b_in[0]), .A2(chi3_0_st0_t0_n2), .ZN(
        chi3_0_st0_t0_n1) );
  XOR2_X1 chi3_0_st0_t0_U1 ( .A(port_a_in0), .B(chi3_0_st0_t0_n1), .Z(
        chi3_0_st0_a_temp[0]) );
  NAND2_X1 chi3_0_st0_t2_U2 ( .A1(port_c_in[1]), .A2(port_b_in[1]), .ZN(
        chi3_0_st0_t2_n1) );
  XNOR2_X1 chi3_0_st0_t2_U1 ( .A(port_a_in1), .B(chi3_0_st0_t2_n1), .ZN(
        chi3_0_st0_a_temp[1]) );
  INV_X1 chi3_0_st0_t1_U3 ( .A(port_c_in[0]), .ZN(chi3_0_st0_t1_n2) );
  NOR2_X1 chi3_0_st0_t1_U2 ( .A1(port_b_in[0]), .A2(chi3_0_st0_t1_n2), .ZN(
        chi3_0_st0_t1_n1) );
  XOR2_X1 chi3_0_st0_t1_U1 ( .A(chi3_0_st0_a_temp[0]), .B(chi3_0_st0_t1_n1), 
        .Z(chi3_0_port_a_out[0]) );
  NAND2_X1 chi3_0_st0_t3_U2 ( .A1(port_c_in[0]), .A2(port_b_in[1]), .ZN(
        chi3_0_st0_t3_n1) );
  XNOR2_X1 chi3_0_st0_t3_U1 ( .A(chi3_0_st0_a_temp[1]), .B(chi3_0_st0_t3_n1), 
        .ZN(chi3_0_port_a_out[1]) );
  INV_X1 chi3_0_st1_t0_U3 ( .A(port_a_in1), .ZN(chi3_0_st1_t0_n2) );
  NOR2_X1 chi3_0_st1_t0_U2 ( .A1(port_c_in[0]), .A2(chi3_0_st1_t0_n2), .ZN(
        chi3_0_st1_t0_n1) );
  XOR2_X1 chi3_0_st1_t0_U1 ( .A(port_b_in[0]), .B(chi3_0_st1_t0_n1), .Z(
        chi3_0_st1_a_temp[0]) );
  NAND2_X1 chi3_0_st1_t2_U2 ( .A1(port_a_in1), .A2(port_c_in[1]), .ZN(
        chi3_0_st1_t2_n1) );
  XNOR2_X1 chi3_0_st1_t2_U1 ( .A(port_b_in[1]), .B(chi3_0_st1_t2_n1), .ZN(
        chi3_0_st1_a_temp[1]) );
  INV_X1 chi3_0_st1_t1_U3 ( .A(port_a_in0), .ZN(chi3_0_st1_t1_n2) );
  NOR2_X1 chi3_0_st1_t1_U2 ( .A1(port_c_in[0]), .A2(chi3_0_st1_t1_n2), .ZN(
        chi3_0_st1_t1_n1) );
  XOR2_X1 chi3_0_st1_t1_U1 ( .A(chi3_0_st1_a_temp[0]), .B(chi3_0_st1_t1_n1), 
        .Z(chi3_0_port_b_out[0]) );
  NAND2_X1 chi3_0_st1_t3_U2 ( .A1(port_a_in0), .A2(port_c_in[1]), .ZN(
        chi3_0_st1_t3_n1) );
  XNOR2_X1 chi3_0_st1_t3_U1 ( .A(chi3_0_st1_a_temp[1]), .B(chi3_0_st1_t3_n1), 
        .ZN(chi3_0_port_b_out[1]) );
  INV_X1 chi3_0_st2_t0_U3 ( .A(port_b_in[1]), .ZN(chi3_0_st2_t0_n2) );
  NOR2_X1 chi3_0_st2_t0_U2 ( .A1(port_a_in0), .A2(chi3_0_st2_t0_n2), .ZN(
        chi3_0_st2_t0_n1) );
  XOR2_X1 chi3_0_st2_t0_U1 ( .A(port_c_in[0]), .B(chi3_0_st2_t0_n1), .Z(
        chi3_0_st2_a_temp[0]) );
  NAND2_X1 chi3_0_st2_t2_U2 ( .A1(port_b_in[1]), .A2(port_a_in1), .ZN(
        chi3_0_st2_t2_n1) );
  XNOR2_X1 chi3_0_st2_t2_U1 ( .A(port_c_in[1]), .B(chi3_0_st2_t2_n1), .ZN(
        chi3_0_st2_a_temp[1]) );
  INV_X1 chi3_0_st2_t1_U3 ( .A(port_b_in[0]), .ZN(chi3_0_st2_t1_n2) );
  NOR2_X1 chi3_0_st2_t1_U2 ( .A1(port_a_in0), .A2(chi3_0_st2_t1_n2), .ZN(
        chi3_0_st2_t1_n1) );
  XOR2_X1 chi3_0_st2_t1_U1 ( .A(chi3_0_st2_a_temp[0]), .B(chi3_0_st2_t1_n1), 
        .Z(chi3_0_port_c_out[0]) );
  NAND2_X1 chi3_0_st2_t3_U2 ( .A1(port_b_in[0]), .A2(port_a_in1), .ZN(
        chi3_0_st2_t3_n1) );
  XNOR2_X1 chi3_0_st2_t3_U1 ( .A(chi3_0_st2_a_temp[1]), .B(chi3_0_st2_t3_n1), 
        .ZN(chi3_0_port_c_out[1]) );
  INV_X1 chi3_1_st0_t0_U3 ( .A(port_c_in[1]), .ZN(chi3_1_st0_t0_n2) );
  NOR2_X1 chi3_1_st0_t0_U2 ( .A1(port_b_in[0]), .A2(chi3_1_st0_t0_n2), .ZN(
        chi3_1_st0_t0_n1) );
  XOR2_X1 chi3_1_st0_t0_U1 ( .A(port_a_in[0]), .B(chi3_1_st0_t0_n1), .Z(
        chi3_1_st0_a_temp[0]) );
  NAND2_X1 chi3_1_st0_t2_U2 ( .A1(port_c_in[1]), .A2(port_b_in[1]), .ZN(
        chi3_1_st0_t2_n1) );
  XNOR2_X1 chi3_1_st0_t2_U1 ( .A(port_a_in[1]), .B(chi3_1_st0_t2_n1), .ZN(
        chi3_1_st0_a_temp[1]) );
  INV_X1 chi3_1_st0_t1_U3 ( .A(port_c_in[0]), .ZN(chi3_1_st0_t1_n2) );
  NOR2_X1 chi3_1_st0_t1_U2 ( .A1(port_b_in[0]), .A2(chi3_1_st0_t1_n2), .ZN(
        chi3_1_st0_t1_n1) );
  XOR2_X1 chi3_1_st0_t1_U1 ( .A(chi3_1_st0_a_temp[0]), .B(chi3_1_st0_t1_n1), 
        .Z(chi3_1_port_a_out[0]) );
  NAND2_X1 chi3_1_st0_t3_U2 ( .A1(port_c_in[0]), .A2(port_b_in[1]), .ZN(
        chi3_1_st0_t3_n1) );
  XNOR2_X1 chi3_1_st0_t3_U1 ( .A(chi3_1_st0_a_temp[1]), .B(chi3_1_st0_t3_n1), 
        .ZN(chi3_1_port_a_out[1]) );
  INV_X1 chi3_1_st1_t0_U3 ( .A(port_a_in[1]), .ZN(chi3_1_st1_t0_n2) );
  NOR2_X1 chi3_1_st1_t0_U2 ( .A1(port_c_in[0]), .A2(chi3_1_st1_t0_n2), .ZN(
        chi3_1_st1_t0_n1) );
  XOR2_X1 chi3_1_st1_t0_U1 ( .A(port_b_in[0]), .B(chi3_1_st1_t0_n1), .Z(
        chi3_1_st1_a_temp[0]) );
  NAND2_X1 chi3_1_st1_t2_U2 ( .A1(port_a_in[1]), .A2(port_c_in[1]), .ZN(
        chi3_1_st1_t2_n1) );
  XNOR2_X1 chi3_1_st1_t2_U1 ( .A(port_b_in[1]), .B(chi3_1_st1_t2_n1), .ZN(
        chi3_1_st1_a_temp[1]) );
  INV_X1 chi3_1_st1_t1_U3 ( .A(port_a_in[0]), .ZN(chi3_1_st1_t1_n2) );
  NOR2_X1 chi3_1_st1_t1_U2 ( .A1(port_c_in[0]), .A2(chi3_1_st1_t1_n2), .ZN(
        chi3_1_st1_t1_n1) );
  XOR2_X1 chi3_1_st1_t1_U1 ( .A(chi3_1_st1_a_temp[0]), .B(chi3_1_st1_t1_n1), 
        .Z(chi3_1_port_b_out[0]) );
  NAND2_X1 chi3_1_st1_t3_U2 ( .A1(port_a_in[0]), .A2(port_c_in[1]), .ZN(
        chi3_1_st1_t3_n1) );
  XNOR2_X1 chi3_1_st1_t3_U1 ( .A(chi3_1_st1_a_temp[1]), .B(chi3_1_st1_t3_n1), 
        .ZN(chi3_1_port_b_out[1]) );
  INV_X1 chi3_1_st2_t0_U3 ( .A(port_b_in[1]), .ZN(chi3_1_st2_t0_n2) );
  NOR2_X1 chi3_1_st2_t0_U2 ( .A1(port_a_in[0]), .A2(chi3_1_st2_t0_n2), .ZN(
        chi3_1_st2_t0_n1) );
  XOR2_X1 chi3_1_st2_t0_U1 ( .A(port_c_in[0]), .B(chi3_1_st2_t0_n1), .Z(
        chi3_1_st2_a_temp[0]) );
  NAND2_X1 chi3_1_st2_t2_U2 ( .A1(port_b_in[1]), .A2(port_a_in[1]), .ZN(
        chi3_1_st2_t2_n1) );
  XNOR2_X1 chi3_1_st2_t2_U1 ( .A(port_c_in[1]), .B(chi3_1_st2_t2_n1), .ZN(
        chi3_1_st2_a_temp[1]) );
  INV_X1 chi3_1_st2_t1_U3 ( .A(port_b_in[0]), .ZN(chi3_1_st2_t1_n2) );
  NOR2_X1 chi3_1_st2_t1_U2 ( .A1(port_a_in[0]), .A2(chi3_1_st2_t1_n2), .ZN(
        chi3_1_st2_t1_n1) );
  XOR2_X1 chi3_1_st2_t1_U1 ( .A(chi3_1_st2_a_temp[0]), .B(chi3_1_st2_t1_n1), 
        .Z(chi3_1_port_c_out[0]) );
  NAND2_X1 chi3_1_st2_t3_U2 ( .A1(port_b_in[0]), .A2(port_a_in[1]), .ZN(
        chi3_1_st2_t3_n1) );
  XNOR2_X1 chi3_1_st2_t3_U1 ( .A(chi3_1_st2_a_temp[1]), .B(chi3_1_st2_t3_n1), 
        .ZN(chi3_1_port_c_out[1]) );
endmodule

