module sbox_wrapper ( clk, data_in, data_out );
  input [11:0] data_in;
  input clk;
  output data_out;
  wire   sbox_s_f_out_11_, sbox_s_g_out_reg_1_, sbox_s_g_out_reg_2_,
         sbox_s_g_out_reg_3_, sbox_s_g_out_reg_5_, sbox_s_g_out_reg_7_,
         sbox_input_data_reg_2_, sbox_input_data_reg_3_,
         sbox_input_data_reg_5_, sbox_input_data_reg_6_,
         sbox_input_data_reg_7_, sbox_input_data_reg_9_,
         sbox_input_data_reg_10_, sbox_input_data_reg_11_, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;
  wire   [7:1] sbox_s_g_out;

  DFF_X1 sbox_s_f_out_reg_reg_11_ ( .D(sbox_s_f_out_11_), .CK(clk), .Q(
        data_out), .QN() );
  DFF_X1 sbox_s_g_out_reg_reg_1_ ( .D(sbox_s_g_out[1]), .CK(clk), .Q(
        sbox_s_g_out_reg_1_), .QN() );
  DFF_X1 sbox_s_g_out_reg_reg_2_ ( .D(sbox_s_g_out[2]), .CK(clk), .Q(
        sbox_s_g_out_reg_2_), .QN() );
  DFF_X1 sbox_s_g_out_reg_reg_3_ ( .D(sbox_s_g_out[3]), .CK(clk), .Q(
        sbox_s_g_out_reg_3_), .QN() );
  DFF_X1 sbox_s_g_out_reg_reg_5_ ( .D(sbox_s_g_out[5]), .CK(clk), .Q(
        sbox_s_g_out_reg_5_), .QN() );
  DFF_X1 sbox_s_g_out_reg_reg_7_ ( .D(sbox_s_g_out[7]), .CK(clk), .Q(
        sbox_s_g_out_reg_7_), .QN() );
  DFF_X1 sbox_input_data_reg_reg_1_ ( .D(data_in[1]), .CK(clk), .Q(), .QN(n43)
         );
  DFF_X1 sbox_input_data_reg_reg_2_ ( .D(data_in[2]), .CK(clk), .Q(
        sbox_input_data_reg_2_), .QN() );
  DFF_X1 sbox_input_data_reg_reg_3_ ( .D(data_in[3]), .CK(clk), .Q(
        sbox_input_data_reg_3_), .QN() );
  DFF_X1 sbox_input_data_reg_reg_4_ ( .D(data_in[4]), .CK(clk), .Q(
        sbox_s_g_out[1]), .QN() );
  DFF_X1 sbox_input_data_reg_reg_5_ ( .D(data_in[5]), .CK(clk), .Q(
        sbox_input_data_reg_5_), .QN(n45) );
  DFF_X1 sbox_input_data_reg_reg_6_ ( .D(data_in[6]), .CK(clk), .Q(
        sbox_input_data_reg_6_), .QN() );
  DFF_X1 sbox_input_data_reg_reg_7_ ( .D(data_in[7]), .CK(clk), .Q(
        sbox_input_data_reg_7_), .QN() );
  DFF_X1 sbox_input_data_reg_reg_8_ ( .D(data_in[8]), .CK(clk), .Q(
        sbox_s_g_out[5]), .QN() );
  DFF_X1 sbox_input_data_reg_reg_9_ ( .D(data_in[9]), .CK(clk), .Q(
        sbox_input_data_reg_9_), .QN(n44) );
  DFF_X1 sbox_input_data_reg_reg_10_ ( .D(data_in[10]), .CK(clk), .Q(
        sbox_input_data_reg_10_), .QN() );
  DFF_X1 sbox_input_data_reg_reg_11_ ( .D(data_in[11]), .CK(clk), .Q(
        sbox_input_data_reg_11_), .QN() );
  XOR2_X1 U47 ( .A(n17), .B(n18), .Z(sbox_s_g_out[3]) );
  XOR2_X1 U48 ( .A(n19), .B(n20), .Z(n18) );
  XOR2_X1 U49 ( .A(n26), .B(n27), .Z(n17) );
  NAND2_X1 U50 ( .A1(n23), .A2(n24), .ZN(n19) );
  XOR2_X1 U51 ( .A(sbox_input_data_reg_11_), .B(sbox_input_data_reg_10_), .Z(
        n13) );
  XOR2_X1 U52 ( .A(sbox_s_g_out[1]), .B(sbox_input_data_reg_9_), .Z(n27) );
  XOR2_X1 U53 ( .A(n7), .B(n8), .Z(n6) );
  NAND2_X1 U54 ( .A1(sbox_input_data_reg_2_), .A2(sbox_input_data_reg_11_), 
        .ZN(n8) );
  NAND2_X1 U55 ( .A1(sbox_input_data_reg_2_), .A2(n9), .ZN(n7) );
  XOR2_X1 U56 ( .A(sbox_input_data_reg_9_), .B(sbox_input_data_reg_3_), .Z(n9)
         );
  XOR2_X1 U57 ( .A(n21), .B(n22), .Z(n20) );
  NAND2_X1 U58 ( .A1(sbox_input_data_reg_6_), .A2(sbox_input_data_reg_11_), 
        .ZN(n22) );
  XNOR2_X1 U59 ( .A(sbox_input_data_reg_6_), .B(sbox_input_data_reg_10_), .ZN(
        n38) );
  XOR2_X1 U60 ( .A(n15), .B(n16), .Z(n10) );
  NAND2_X1 U61 ( .A1(sbox_input_data_reg_3_), .A2(sbox_input_data_reg_10_), 
        .ZN(n15) );
  AND2_X1 U62 ( .A1(sbox_input_data_reg_9_), .A2(sbox_input_data_reg_3_), .ZN(
        n16) );
  XOR2_X1 U63 ( .A(n3), .B(n4), .Z(sbox_s_g_out[7]) );
  XOR2_X1 U64 ( .A(n5), .B(n6), .Z(n4) );
  XOR2_X1 U65 ( .A(n10), .B(n11), .Z(n3) );
  XOR2_X1 U66 ( .A(sbox_s_g_out[5]), .B(sbox_input_data_reg_9_), .Z(n5) );
  NAND2_X1 U67 ( .A1(sbox_input_data_reg_7_), .A2(sbox_input_data_reg_10_), 
        .ZN(n21) );
  XOR2_X1 U68 ( .A(sbox_s_g_out_reg_5_), .B(sbox_s_g_out_reg_1_), .Z(n42) );
  NAND2_X1 U69 ( .A1(sbox_input_data_reg_10_), .A2(n25), .ZN(n24) );
  OR2_X1 U70 ( .A1(sbox_input_data_reg_11_), .A2(sbox_input_data_reg_5_), .ZN(
        n25) );
  XOR2_X1 U71 ( .A(n28), .B(sbox_input_data_reg_5_), .Z(n26) );
  NAND2_X1 U72 ( .A1(sbox_input_data_reg_9_), .A2(n29), .ZN(n28) );
  XOR2_X1 U73 ( .A(n13), .B(n30), .Z(n29) );
  XOR2_X1 U74 ( .A(sbox_input_data_reg_7_), .B(sbox_input_data_reg_6_), .Z(n30) );
  NOR2_X1 U75 ( .A1(n43), .A2(n12), .ZN(n11) );
  XOR2_X1 U76 ( .A(n13), .B(n14), .Z(n12) );
  XOR2_X1 U77 ( .A(sbox_input_data_reg_3_), .B(sbox_input_data_reg_2_), .Z(n14) );
  NAND2_X1 U78 ( .A1(sbox_input_data_reg_5_), .A2(sbox_input_data_reg_11_), 
        .ZN(n23) );
  NOR2_X1 U79 ( .A1(n35), .A2(n36), .ZN(n34) );
  NOR2_X1 U80 ( .A1(sbox_input_data_reg_7_), .A2(n37), .ZN(n35) );
  NOR2_X1 U81 ( .A1(n45), .A2(n21), .ZN(n36) );
  AND2_X1 U82 ( .A1(sbox_input_data_reg_10_), .A2(sbox_input_data_reg_5_), 
        .ZN(n37) );
  XOR2_X1 U83 ( .A(n39), .B(n40), .Z(sbox_s_f_out_11_) );
  NAND2_X1 U84 ( .A1(sbox_s_g_out_reg_5_), .A2(sbox_s_g_out_reg_3_), .ZN(n39)
         );
  XOR2_X1 U85 ( .A(n41), .B(sbox_s_g_out_reg_2_), .Z(n40) );
  NAND2_X1 U86 ( .A1(sbox_s_g_out_reg_7_), .A2(n42), .ZN(n41) );
  XOR2_X1 U87 ( .A(n31), .B(n32), .Z(sbox_s_g_out[2]) );
  XOR2_X1 U88 ( .A(sbox_s_g_out[1]), .B(n44), .Z(n31) );
  XOR2_X1 U89 ( .A(n33), .B(n34), .Z(n32) );
  NOR2_X1 U90 ( .A1(n38), .A2(n44), .ZN(n33) );
endmodule
