
module CINI_HPC3 ( port_a_0, port_a_1, port_a_2, port_b_0, port_b_1, port_b_2, 
        port_c_0, port_c_1, port_c_2, port_rand_ref, port_rand_mul, clk, reset
 );
  input [4:0] port_a_0;
  input [4:0] port_a_1;
  input [4:0] port_a_2;
  input [4:0] port_b_0;
  input [4:0] port_b_1;
  input [4:0] port_b_2;
  output [4:0] port_c_0;
  output [4:0] port_c_1;
  output [4:0] port_c_2;
  input [2:0] port_rand_ref;
  input [2:0] port_rand_mul;
  input clk, reset;
  wire   simpleAnd_30_port_z, simpleAnd_31_port_z, simpleAnd_32_port_z,
         simpleAnd_33_port_z, simpleAnd_34_port_z, simpleAnd_35_port_z,
         simpleAnd_36_port_z, simpleAnd_37_port_z, simpleAnd_38_port_z,
         simpleAnd_39_port_z, simpleAnd_40_port_z, simpleAnd_41_port_z,
         simpleAnd_42_port_z, simpleAnd_43_port_z, simpleAnd_44_port_z,
         simpleAnd_45_port_z, simpleAnd_46_port_z, simpleAnd_47_port_z,
         simpleAnd_48_port_z, simpleAnd_49_port_z, simpleAnd_50_port_z,
         simpleAnd_51_port_z, simpleAnd_52_port_z, simpleAnd_53_port_z,
         simpleAnd_54_port_z, simpleAnd_55_port_z, simpleAnd_56_port_z,
         simpleAnd_57_port_z, simpleAnd_58_port_z, simpleAnd_59_port_z,
         maj_60_port_o, maj_61_port_o, maj_62_port_o, maj_63_port_o,
         maj_64_port_o, maj_65_port_o, maj_66_port_o, maj_67_port_o,
         maj_68_port_o, maj_69_port_o, maj_70_port_o, maj_71_port_o,
         maj_72_port_o, maj_73_port_o, maj_74_port_o, maj_75_port_o,
         maj_76_port_o, maj_77_port_o, maj_78_port_o, maj_79_port_o,
         maj_80_port_o, maj_81_port_o, maj_82_port_o, maj_83_port_o,
         maj_84_port_o, maj_85_port_o, maj_86_port_o, maj_87_port_o,
         maj_88_port_o, maj_89_port_o, maj_90_port_o, maj_91_port_o,
         maj_92_port_o, maj_93_port_o, maj_94_port_o, maj_95_port_o,
         maj_96_port_o, maj_97_port_o, maj_98_port_o, maj_99_port_o,
         maj_100_port_o, maj_101_port_o, maj_102_port_o, maj_103_port_o,
         maj_104_port_o, maj_105_port_o, maj_106_port_o, maj_107_port_o,
         maj_108_port_o, maj_109_port_o, maj_110_port_o, maj_111_port_o,
         maj_112_port_o, maj_113_port_o, maj_114_port_o, maj_115_port_o,
         maj_116_port_o, maj_117_port_o, maj_118_port_o, maj_119_port_o, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, maj_60_n13, maj_60_n12, maj_60_n11, maj_60_n10,
         maj_60_n9, maj_60_n8, maj_60_n7, maj_60_n6, maj_60_n5, maj_60_n4,
         maj_60_n3, maj_60_n2, maj_60_n1, maj_61_n26, maj_61_n25, maj_61_n24,
         maj_61_n23, maj_61_n22, maj_61_n21, maj_61_n20, maj_61_n19,
         maj_61_n18, maj_61_n17, maj_61_n16, maj_61_n15, maj_61_n14,
         maj_62_n26, maj_62_n25, maj_62_n24, maj_62_n23, maj_62_n22,
         maj_62_n21, maj_62_n20, maj_62_n19, maj_62_n18, maj_62_n17,
         maj_62_n16, maj_62_n15, maj_62_n14, maj_63_n26, maj_63_n25,
         maj_63_n24, maj_63_n23, maj_63_n22, maj_63_n21, maj_63_n20,
         maj_63_n19, maj_63_n18, maj_63_n17, maj_63_n16, maj_63_n15,
         maj_63_n14, maj_64_n26, maj_64_n25, maj_64_n24, maj_64_n23,
         maj_64_n22, maj_64_n21, maj_64_n20, maj_64_n19, maj_64_n18,
         maj_64_n17, maj_64_n16, maj_64_n15, maj_64_n14, maj_65_n26,
         maj_65_n25, maj_65_n24, maj_65_n23, maj_65_n22, maj_65_n21,
         maj_65_n20, maj_65_n19, maj_65_n18, maj_65_n17, maj_65_n16,
         maj_65_n15, maj_65_n14, maj_66_n26, maj_66_n25, maj_66_n24,
         maj_66_n23, maj_66_n22, maj_66_n21, maj_66_n20, maj_66_n19,
         maj_66_n18, maj_66_n17, maj_66_n16, maj_66_n15, maj_66_n14,
         maj_67_n26, maj_67_n25, maj_67_n24, maj_67_n23, maj_67_n22,
         maj_67_n21, maj_67_n20, maj_67_n19, maj_67_n18, maj_67_n17,
         maj_67_n16, maj_67_n15, maj_67_n14, maj_68_n26, maj_68_n25,
         maj_68_n24, maj_68_n23, maj_68_n22, maj_68_n21, maj_68_n20,
         maj_68_n19, maj_68_n18, maj_68_n17, maj_68_n16, maj_68_n15,
         maj_68_n14, maj_69_n26, maj_69_n25, maj_69_n24, maj_69_n23,
         maj_69_n22, maj_69_n21, maj_69_n20, maj_69_n19, maj_69_n18,
         maj_69_n17, maj_69_n16, maj_69_n15, maj_69_n14, maj_70_n26,
         maj_70_n25, maj_70_n24, maj_70_n23, maj_70_n22, maj_70_n21,
         maj_70_n20, maj_70_n19, maj_70_n18, maj_70_n17, maj_70_n16,
         maj_70_n15, maj_70_n14, maj_71_n26, maj_71_n25, maj_71_n24,
         maj_71_n23, maj_71_n22, maj_71_n21, maj_71_n20, maj_71_n19,
         maj_71_n18, maj_71_n17, maj_71_n16, maj_71_n15, maj_71_n14,
         maj_72_n26, maj_72_n25, maj_72_n24, maj_72_n23, maj_72_n22,
         maj_72_n21, maj_72_n20, maj_72_n19, maj_72_n18, maj_72_n17,
         maj_72_n16, maj_72_n15, maj_72_n14, maj_73_n26, maj_73_n25,
         maj_73_n24, maj_73_n23, maj_73_n22, maj_73_n21, maj_73_n20,
         maj_73_n19, maj_73_n18, maj_73_n17, maj_73_n16, maj_73_n15,
         maj_73_n14, maj_74_n26, maj_74_n25, maj_74_n24, maj_74_n23,
         maj_74_n22, maj_74_n21, maj_74_n20, maj_74_n19, maj_74_n18,
         maj_74_n17, maj_74_n16, maj_74_n15, maj_74_n14, maj_75_n26,
         maj_75_n25, maj_75_n24, maj_75_n23, maj_75_n22, maj_75_n21,
         maj_75_n20, maj_75_n19, maj_75_n18, maj_75_n17, maj_75_n16,
         maj_75_n15, maj_75_n14, maj_76_n26, maj_76_n25, maj_76_n24,
         maj_76_n23, maj_76_n22, maj_76_n21, maj_76_n20, maj_76_n19,
         maj_76_n18, maj_76_n17, maj_76_n16, maj_76_n15, maj_76_n14,
         maj_77_n26, maj_77_n25, maj_77_n24, maj_77_n23, maj_77_n22,
         maj_77_n21, maj_77_n20, maj_77_n19, maj_77_n18, maj_77_n17,
         maj_77_n16, maj_77_n15, maj_77_n14, maj_78_n26, maj_78_n25,
         maj_78_n24, maj_78_n23, maj_78_n22, maj_78_n21, maj_78_n20,
         maj_78_n19, maj_78_n18, maj_78_n17, maj_78_n16, maj_78_n15,
         maj_78_n14, maj_79_n26, maj_79_n25, maj_79_n24, maj_79_n23,
         maj_79_n22, maj_79_n21, maj_79_n20, maj_79_n19, maj_79_n18,
         maj_79_n17, maj_79_n16, maj_79_n15, maj_79_n14, maj_80_n26,
         maj_80_n25, maj_80_n24, maj_80_n23, maj_80_n22, maj_80_n21,
         maj_80_n20, maj_80_n19, maj_80_n18, maj_80_n17, maj_80_n16,
         maj_80_n15, maj_80_n14, maj_81_n26, maj_81_n25, maj_81_n24,
         maj_81_n23, maj_81_n22, maj_81_n21, maj_81_n20, maj_81_n19,
         maj_81_n18, maj_81_n17, maj_81_n16, maj_81_n15, maj_81_n14,
         maj_82_n26, maj_82_n25, maj_82_n24, maj_82_n23, maj_82_n22,
         maj_82_n21, maj_82_n20, maj_82_n19, maj_82_n18, maj_82_n17,
         maj_82_n16, maj_82_n15, maj_82_n14, maj_83_n26, maj_83_n25,
         maj_83_n24, maj_83_n23, maj_83_n22, maj_83_n21, maj_83_n20,
         maj_83_n19, maj_83_n18, maj_83_n17, maj_83_n16, maj_83_n15,
         maj_83_n14, maj_84_n26, maj_84_n25, maj_84_n24, maj_84_n23,
         maj_84_n22, maj_84_n21, maj_84_n20, maj_84_n19, maj_84_n18,
         maj_84_n17, maj_84_n16, maj_84_n15, maj_84_n14, maj_85_n26,
         maj_85_n25, maj_85_n24, maj_85_n23, maj_85_n22, maj_85_n21,
         maj_85_n20, maj_85_n19, maj_85_n18, maj_85_n17, maj_85_n16,
         maj_85_n15, maj_85_n14, maj_86_n26, maj_86_n25, maj_86_n24,
         maj_86_n23, maj_86_n22, maj_86_n21, maj_86_n20, maj_86_n19,
         maj_86_n18, maj_86_n17, maj_86_n16, maj_86_n15, maj_86_n14,
         maj_87_n26, maj_87_n25, maj_87_n24, maj_87_n23, maj_87_n22,
         maj_87_n21, maj_87_n20, maj_87_n19, maj_87_n18, maj_87_n17,
         maj_87_n16, maj_87_n15, maj_87_n14, maj_88_n26, maj_88_n25,
         maj_88_n24, maj_88_n23, maj_88_n22, maj_88_n21, maj_88_n20,
         maj_88_n19, maj_88_n18, maj_88_n17, maj_88_n16, maj_88_n15,
         maj_88_n14, maj_89_n26, maj_89_n25, maj_89_n24, maj_89_n23,
         maj_89_n22, maj_89_n21, maj_89_n20, maj_89_n19, maj_89_n18,
         maj_89_n17, maj_89_n16, maj_89_n15, maj_89_n14, maj_90_n26,
         maj_90_n25, maj_90_n24, maj_90_n23, maj_90_n22, maj_90_n21,
         maj_90_n20, maj_90_n19, maj_90_n18, maj_90_n17, maj_90_n16,
         maj_90_n15, maj_90_n14, maj_91_n26, maj_91_n25, maj_91_n24,
         maj_91_n23, maj_91_n22, maj_91_n21, maj_91_n20, maj_91_n19,
         maj_91_n18, maj_91_n17, maj_91_n16, maj_91_n15, maj_91_n14,
         maj_92_n26, maj_92_n25, maj_92_n24, maj_92_n23, maj_92_n22,
         maj_92_n21, maj_92_n20, maj_92_n19, maj_92_n18, maj_92_n17,
         maj_92_n16, maj_92_n15, maj_92_n14, maj_93_n26, maj_93_n25,
         maj_93_n24, maj_93_n23, maj_93_n22, maj_93_n21, maj_93_n20,
         maj_93_n19, maj_93_n18, maj_93_n17, maj_93_n16, maj_93_n15,
         maj_93_n14, maj_94_n26, maj_94_n25, maj_94_n24, maj_94_n23,
         maj_94_n22, maj_94_n21, maj_94_n20, maj_94_n19, maj_94_n18,
         maj_94_n17, maj_94_n16, maj_94_n15, maj_94_n14, maj_95_n26,
         maj_95_n25, maj_95_n24, maj_95_n23, maj_95_n22, maj_95_n21,
         maj_95_n20, maj_95_n19, maj_95_n18, maj_95_n17, maj_95_n16,
         maj_95_n15, maj_95_n14, maj_96_n26, maj_96_n25, maj_96_n24,
         maj_96_n23, maj_96_n22, maj_96_n21, maj_96_n20, maj_96_n19,
         maj_96_n18, maj_96_n17, maj_96_n16, maj_96_n15, maj_96_n14,
         maj_97_n26, maj_97_n25, maj_97_n24, maj_97_n23, maj_97_n22,
         maj_97_n21, maj_97_n20, maj_97_n19, maj_97_n18, maj_97_n17,
         maj_97_n16, maj_97_n15, maj_97_n14, maj_98_n26, maj_98_n25,
         maj_98_n24, maj_98_n23, maj_98_n22, maj_98_n21, maj_98_n20,
         maj_98_n19, maj_98_n18, maj_98_n17, maj_98_n16, maj_98_n15,
         maj_98_n14, maj_99_n26, maj_99_n25, maj_99_n24, maj_99_n23,
         maj_99_n22, maj_99_n21, maj_99_n20, maj_99_n19, maj_99_n18,
         maj_99_n17, maj_99_n16, maj_99_n15, maj_99_n14, maj_100_n26,
         maj_100_n25, maj_100_n24, maj_100_n23, maj_100_n22, maj_100_n21,
         maj_100_n20, maj_100_n19, maj_100_n18, maj_100_n17, maj_100_n16,
         maj_100_n15, maj_100_n14, maj_101_n26, maj_101_n25, maj_101_n24,
         maj_101_n23, maj_101_n22, maj_101_n21, maj_101_n20, maj_101_n19,
         maj_101_n18, maj_101_n17, maj_101_n16, maj_101_n15, maj_101_n14,
         maj_102_n26, maj_102_n25, maj_102_n24, maj_102_n23, maj_102_n22,
         maj_102_n21, maj_102_n20, maj_102_n19, maj_102_n18, maj_102_n17,
         maj_102_n16, maj_102_n15, maj_102_n14, maj_103_n26, maj_103_n25,
         maj_103_n24, maj_103_n23, maj_103_n22, maj_103_n21, maj_103_n20,
         maj_103_n19, maj_103_n18, maj_103_n17, maj_103_n16, maj_103_n15,
         maj_103_n14, maj_104_n26, maj_104_n25, maj_104_n24, maj_104_n23,
         maj_104_n22, maj_104_n21, maj_104_n20, maj_104_n19, maj_104_n18,
         maj_104_n17, maj_104_n16, maj_104_n15, maj_104_n14, maj_105_n26,
         maj_105_n25, maj_105_n24, maj_105_n23, maj_105_n22, maj_105_n21,
         maj_105_n20, maj_105_n19, maj_105_n18, maj_105_n17, maj_105_n16,
         maj_105_n15, maj_105_n14, maj_106_n26, maj_106_n25, maj_106_n24,
         maj_106_n23, maj_106_n22, maj_106_n21, maj_106_n20, maj_106_n19,
         maj_106_n18, maj_106_n17, maj_106_n16, maj_106_n15, maj_106_n14,
         maj_107_n26, maj_107_n25, maj_107_n24, maj_107_n23, maj_107_n22,
         maj_107_n21, maj_107_n20, maj_107_n19, maj_107_n18, maj_107_n17,
         maj_107_n16, maj_107_n15, maj_107_n14, maj_108_n26, maj_108_n25,
         maj_108_n24, maj_108_n23, maj_108_n22, maj_108_n21, maj_108_n20,
         maj_108_n19, maj_108_n18, maj_108_n17, maj_108_n16, maj_108_n15,
         maj_108_n14, maj_109_n26, maj_109_n25, maj_109_n24, maj_109_n23,
         maj_109_n22, maj_109_n21, maj_109_n20, maj_109_n19, maj_109_n18,
         maj_109_n17, maj_109_n16, maj_109_n15, maj_109_n14, maj_110_n26,
         maj_110_n25, maj_110_n24, maj_110_n23, maj_110_n22, maj_110_n21,
         maj_110_n20, maj_110_n19, maj_110_n18, maj_110_n17, maj_110_n16,
         maj_110_n15, maj_110_n14, maj_111_n26, maj_111_n25, maj_111_n24,
         maj_111_n23, maj_111_n22, maj_111_n21, maj_111_n20, maj_111_n19,
         maj_111_n18, maj_111_n17, maj_111_n16, maj_111_n15, maj_111_n14,
         maj_112_n26, maj_112_n25, maj_112_n24, maj_112_n23, maj_112_n22,
         maj_112_n21, maj_112_n20, maj_112_n19, maj_112_n18, maj_112_n17,
         maj_112_n16, maj_112_n15, maj_112_n14, maj_113_n26, maj_113_n25,
         maj_113_n24, maj_113_n23, maj_113_n22, maj_113_n21, maj_113_n20,
         maj_113_n19, maj_113_n18, maj_113_n17, maj_113_n16, maj_113_n15,
         maj_113_n14, maj_114_n26, maj_114_n25, maj_114_n24, maj_114_n23,
         maj_114_n22, maj_114_n21, maj_114_n20, maj_114_n19, maj_114_n18,
         maj_114_n17, maj_114_n16, maj_114_n15, maj_114_n14, maj_115_n26,
         maj_115_n25, maj_115_n24, maj_115_n23, maj_115_n22, maj_115_n21,
         maj_115_n20, maj_115_n19, maj_115_n18, maj_115_n17, maj_115_n16,
         maj_115_n15, maj_115_n14, maj_116_n26, maj_116_n25, maj_116_n24,
         maj_116_n23, maj_116_n22, maj_116_n21, maj_116_n20, maj_116_n19,
         maj_116_n18, maj_116_n17, maj_116_n16, maj_116_n15, maj_116_n14,
         maj_117_n26, maj_117_n25, maj_117_n24, maj_117_n23, maj_117_n22,
         maj_117_n21, maj_117_n20, maj_117_n19, maj_117_n18, maj_117_n17,
         maj_117_n16, maj_117_n15, maj_117_n14, maj_118_n26, maj_118_n25,
         maj_118_n24, maj_118_n23, maj_118_n22, maj_118_n21, maj_118_n20,
         maj_118_n19, maj_118_n18, maj_118_n17, maj_118_n16, maj_118_n15,
         maj_118_n14, maj_119_n26, maj_119_n25, maj_119_n24, maj_119_n23,
         maj_119_n22, maj_119_n21, maj_119_n20, maj_119_n19, maj_119_n18,
         maj_119_n17, maj_119_n16, maj_119_n15, maj_119_n14;
  wire   [4:0] u_0_0;
  wire   [4:0] v_0_0;
  wire   [4:0] u_0_1;
  wire   [4:0] v_0_1;
  wire   [4:0] u_1_0;
  wire   [4:0] v_1_0;
  wire   [4:0] u_1_1;
  wire   [4:0] v_1_1;
  wire   [4:0] u_2_0;
  wire   [4:0] v_2_0;
  wire   [4:0] u_2_1;
  wire   [4:0] v_2_1;
  wire   [4:0] temp_0_0;
  wire   [4:0] a_reg_0;
  wire   [4:0] v_reg_0_0;
  wire   [4:0] u_reg_0_0;
  wire   [4:0] v_reg_0_1;
  wire   [4:0] u_reg_0_1;
  wire   [4:0] temp_0_1;
  wire   [4:0] a_reg_1;
  wire   [4:0] v_reg_1_0;
  wire   [4:0] u_reg_1_0;
  wire   [4:0] v_reg_1_1;
  wire   [4:0] u_reg_1_1;
  wire   [4:0] temp_0_2;
  wire   [4:0] a_reg_2;
  wire   [4:0] v_reg_2_0;
  wire   [4:0] u_reg_2_0;
  wire   [4:0] v_reg_2_1;
  wire   [4:0] u_reg_2_1;

  DFF_X1 u_reg_0_0_reg_4_ ( .D(maj_108_port_o), .CK(clk), .Q(u_reg_0_0[4]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_3_ ( .D(maj_96_port_o), .CK(clk), .Q(u_reg_0_0[3]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_2_ ( .D(maj_84_port_o), .CK(clk), .Q(u_reg_0_0[2]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_1_ ( .D(maj_72_port_o), .CK(clk), .Q(u_reg_0_0[1]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_0_ ( .D(maj_60_port_o), .CK(clk), .Q(u_reg_0_0[0]), 
        .QN() );
  DFF_X1 a_reg_2_reg_4_ ( .D(port_a_2[4]), .CK(clk), .Q(a_reg_2[4]), .QN() );
  DFF_X1 a_reg_2_reg_3_ ( .D(port_a_2[3]), .CK(clk), .Q(a_reg_2[3]), .QN() );
  DFF_X1 a_reg_2_reg_2_ ( .D(port_a_2[2]), .CK(clk), .Q(a_reg_2[2]), .QN() );
  DFF_X1 a_reg_2_reg_1_ ( .D(port_a_2[1]), .CK(clk), .Q(a_reg_2[1]), .QN() );
  DFF_X1 a_reg_2_reg_0_ ( .D(port_a_2[0]), .CK(clk), .Q(a_reg_2[0]), .QN() );
  DFF_X1 v_reg_1_0_reg_4_ ( .D(maj_113_port_o), .CK(clk), .Q(v_reg_1_0[4]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_3_ ( .D(maj_101_port_o), .CK(clk), .Q(v_reg_1_0[3]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_2_ ( .D(maj_89_port_o), .CK(clk), .Q(v_reg_1_0[2]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_1_ ( .D(maj_77_port_o), .CK(clk), .Q(v_reg_1_0[1]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_0_ ( .D(maj_65_port_o), .CK(clk), .Q(v_reg_1_0[0]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_4_ ( .D(maj_110_port_o), .CK(clk), .Q(u_reg_0_1[4]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_3_ ( .D(maj_98_port_o), .CK(clk), .Q(u_reg_0_1[3]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_2_ ( .D(maj_86_port_o), .CK(clk), .Q(u_reg_0_1[2]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_1_ ( .D(maj_74_port_o), .CK(clk), .Q(u_reg_0_1[1]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_0_ ( .D(maj_62_port_o), .CK(clk), .Q(u_reg_0_1[0]), 
        .QN() );
  DFF_X1 ab_reg_2_reg_4_ ( .D(N14), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 ab_reg_2_reg_3_ ( .D(N11), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 ab_reg_2_reg_2_ ( .D(N8), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 ab_reg_2_reg_1_ ( .D(N5), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 ab_reg_2_reg_0_ ( .D(N2), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 v_reg_0_1_reg_4_ ( .D(maj_111_port_o), .CK(clk), .Q(v_reg_0_1[4]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_3_ ( .D(maj_99_port_o), .CK(clk), .Q(v_reg_0_1[3]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_2_ ( .D(maj_87_port_o), .CK(clk), .Q(v_reg_0_1[2]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_1_ ( .D(maj_75_port_o), .CK(clk), .Q(v_reg_0_1[1]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_0_ ( .D(maj_63_port_o), .CK(clk), .Q(v_reg_0_1[0]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_4_ ( .D(maj_112_port_o), .CK(clk), .Q(u_reg_1_0[4]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_3_ ( .D(maj_100_port_o), .CK(clk), .Q(u_reg_1_0[3]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_2_ ( .D(maj_88_port_o), .CK(clk), .Q(u_reg_1_0[2]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_1_ ( .D(maj_76_port_o), .CK(clk), .Q(u_reg_1_0[1]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_0_ ( .D(maj_64_port_o), .CK(clk), .Q(u_reg_1_0[0]), 
        .QN() );
  DFF_X1 a_reg_1_reg_4_ ( .D(port_a_1[4]), .CK(clk), .Q(a_reg_1[4]), .QN() );
  DFF_X1 a_reg_1_reg_3_ ( .D(port_a_1[3]), .CK(clk), .Q(a_reg_1[3]), .QN() );
  DFF_X1 a_reg_1_reg_2_ ( .D(port_a_1[2]), .CK(clk), .Q(a_reg_1[2]), .QN() );
  DFF_X1 a_reg_1_reg_1_ ( .D(port_a_1[1]), .CK(clk), .Q(a_reg_1[1]), .QN() );
  DFF_X1 a_reg_1_reg_0_ ( .D(port_a_1[0]), .CK(clk), .Q(a_reg_1[0]), .QN() );
  DFF_X1 v_reg_0_0_reg_4_ ( .D(maj_109_port_o), .CK(clk), .Q(v_reg_0_0[4]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_3_ ( .D(maj_97_port_o), .CK(clk), .Q(v_reg_0_0[3]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_2_ ( .D(maj_85_port_o), .CK(clk), .Q(v_reg_0_0[2]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_1_ ( .D(maj_73_port_o), .CK(clk), .Q(v_reg_0_0[1]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_0_ ( .D(maj_61_port_o), .CK(clk), .Q(v_reg_0_0[0]), 
        .QN() );
  DFF_X1 ab_reg_1_reg_4_ ( .D(N13), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 ab_reg_1_reg_3_ ( .D(N10), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 ab_reg_1_reg_2_ ( .D(N7), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 ab_reg_1_reg_1_ ( .D(N4), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 ab_reg_1_reg_0_ ( .D(N1), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 a_reg_0_reg_4_ ( .D(port_a_0[4]), .CK(clk), .Q(a_reg_0[4]), .QN() );
  DFF_X1 a_reg_0_reg_3_ ( .D(port_a_0[3]), .CK(clk), .Q(a_reg_0[3]), .QN() );
  DFF_X1 a_reg_0_reg_2_ ( .D(port_a_0[2]), .CK(clk), .Q(a_reg_0[2]), .QN() );
  DFF_X1 a_reg_0_reg_1_ ( .D(port_a_0[1]), .CK(clk), .Q(a_reg_0[1]), .QN() );
  DFF_X1 a_reg_0_reg_0_ ( .D(port_a_0[0]), .CK(clk), .Q(a_reg_0[0]), .QN() );
  DFF_X1 ab_reg_0_reg_4_ ( .D(N12), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 ab_reg_0_reg_3_ ( .D(N9), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 ab_reg_0_reg_2_ ( .D(N6), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 ab_reg_0_reg_1_ ( .D(N3), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 ab_reg_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 v_reg_2_1_reg_4_ ( .D(maj_119_port_o), .CK(clk), .Q(v_reg_2_1[4]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_3_ ( .D(maj_107_port_o), .CK(clk), .Q(v_reg_2_1[3]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_2_ ( .D(maj_95_port_o), .CK(clk), .Q(v_reg_2_1[2]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_1_ ( .D(maj_83_port_o), .CK(clk), .Q(v_reg_2_1[1]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_0_ ( .D(maj_71_port_o), .CK(clk), .Q(v_reg_2_1[0]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_4_ ( .D(maj_118_port_o), .CK(clk), .Q(u_reg_2_1[4]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_3_ ( .D(maj_106_port_o), .CK(clk), .Q(u_reg_2_1[3]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_2_ ( .D(maj_94_port_o), .CK(clk), .Q(u_reg_2_1[2]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_1_ ( .D(maj_82_port_o), .CK(clk), .Q(u_reg_2_1[1]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_0_ ( .D(maj_70_port_o), .CK(clk), .Q(u_reg_2_1[0]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_4_ ( .D(maj_117_port_o), .CK(clk), .Q(v_reg_2_0[4]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_3_ ( .D(maj_105_port_o), .CK(clk), .Q(v_reg_2_0[3]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_2_ ( .D(maj_93_port_o), .CK(clk), .Q(v_reg_2_0[2]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_1_ ( .D(maj_81_port_o), .CK(clk), .Q(v_reg_2_0[1]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_0_ ( .D(maj_69_port_o), .CK(clk), .Q(v_reg_2_0[0]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_4_ ( .D(maj_116_port_o), .CK(clk), .Q(u_reg_2_0[4]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_3_ ( .D(maj_104_port_o), .CK(clk), .Q(u_reg_2_0[3]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_2_ ( .D(maj_92_port_o), .CK(clk), .Q(u_reg_2_0[2]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_1_ ( .D(maj_80_port_o), .CK(clk), .Q(u_reg_2_0[1]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_0_ ( .D(maj_68_port_o), .CK(clk), .Q(u_reg_2_0[0]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_4_ ( .D(maj_115_port_o), .CK(clk), .Q(v_reg_1_1[4]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_3_ ( .D(maj_103_port_o), .CK(clk), .Q(v_reg_1_1[3]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_2_ ( .D(maj_91_port_o), .CK(clk), .Q(v_reg_1_1[2]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_1_ ( .D(maj_79_port_o), .CK(clk), .Q(v_reg_1_1[1]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_0_ ( .D(maj_67_port_o), .CK(clk), .Q(v_reg_1_1[0]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_4_ ( .D(maj_114_port_o), .CK(clk), .Q(u_reg_1_1[4]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_3_ ( .D(maj_102_port_o), .CK(clk), .Q(u_reg_1_1[3]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_2_ ( .D(maj_90_port_o), .CK(clk), .Q(u_reg_1_1[2]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_1_ ( .D(maj_78_port_o), .CK(clk), .Q(u_reg_1_1[1]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_0_ ( .D(maj_66_port_o), .CK(clk), .Q(u_reg_1_1[0]), 
        .QN() );
  XNOR2_X1 U123 ( .A(u_reg_2_1[0]), .B(u_reg_2_0[0]), .ZN(n40) );
  XNOR2_X1 U124 ( .A(u_reg_2_1[1]), .B(u_reg_2_0[1]), .ZN(n35) );
  XNOR2_X1 U125 ( .A(u_reg_2_1[2]), .B(u_reg_2_0[2]), .ZN(n30) );
  XNOR2_X1 U126 ( .A(u_reg_2_1[3]), .B(u_reg_2_0[3]), .ZN(n25) );
  XNOR2_X1 U127 ( .A(u_reg_2_1[4]), .B(u_reg_2_0[4]), .ZN(n20) );
  XNOR2_X1 U128 ( .A(u_reg_1_1[0]), .B(u_reg_1_0[0]), .ZN(n65) );
  XNOR2_X1 U129 ( .A(u_reg_1_1[1]), .B(u_reg_1_0[1]), .ZN(n60) );
  XNOR2_X1 U130 ( .A(u_reg_1_1[2]), .B(u_reg_1_0[2]), .ZN(n55) );
  XNOR2_X1 U131 ( .A(u_reg_1_1[3]), .B(u_reg_1_0[3]), .ZN(n50) );
  XNOR2_X1 U132 ( .A(u_reg_1_1[4]), .B(u_reg_1_0[4]), .ZN(n45) );
  XNOR2_X1 U133 ( .A(u_reg_0_1[0]), .B(u_reg_0_0[0]), .ZN(n90) );
  XNOR2_X1 U134 ( .A(u_reg_0_1[1]), .B(u_reg_0_0[1]), .ZN(n85) );
  XNOR2_X1 U135 ( .A(u_reg_0_1[2]), .B(u_reg_0_0[2]), .ZN(n80) );
  XNOR2_X1 U136 ( .A(u_reg_0_1[3]), .B(u_reg_0_0[3]), .ZN(n75) );
  XNOR2_X1 U137 ( .A(u_reg_0_1[4]), .B(u_reg_0_0[4]), .ZN(n70) );
  XOR2_X1 U138 ( .A(n36), .B(n37), .Z(port_c_2[0]) );
  XNOR2_X1 U139 ( .A(n38), .B(n39), .ZN(n37) );
  XOR2_X1 U140 ( .A(n40), .B(temp_0_2[0]), .Z(n36) );
  NAND2_X1 U141 ( .A1(v_reg_2_1[0]), .A2(a_reg_2[0]), .ZN(n38) );
  XOR2_X1 U142 ( .A(n31), .B(n32), .Z(port_c_2[1]) );
  XNOR2_X1 U143 ( .A(n33), .B(n34), .ZN(n32) );
  XOR2_X1 U144 ( .A(n35), .B(temp_0_2[1]), .Z(n31) );
  NAND2_X1 U145 ( .A1(v_reg_2_1[1]), .A2(a_reg_2[1]), .ZN(n33) );
  XOR2_X1 U146 ( .A(n26), .B(n27), .Z(port_c_2[2]) );
  XNOR2_X1 U147 ( .A(n28), .B(n29), .ZN(n27) );
  XOR2_X1 U148 ( .A(n30), .B(temp_0_2[2]), .Z(n26) );
  NAND2_X1 U149 ( .A1(v_reg_2_1[2]), .A2(a_reg_2[2]), .ZN(n28) );
  XOR2_X1 U150 ( .A(n21), .B(n22), .Z(port_c_2[3]) );
  XNOR2_X1 U151 ( .A(n23), .B(n24), .ZN(n22) );
  XOR2_X1 U152 ( .A(n25), .B(temp_0_2[3]), .Z(n21) );
  NAND2_X1 U153 ( .A1(v_reg_2_1[3]), .A2(a_reg_2[3]), .ZN(n23) );
  XOR2_X1 U154 ( .A(n16), .B(n17), .Z(port_c_2[4]) );
  XNOR2_X1 U155 ( .A(n18), .B(n19), .ZN(n17) );
  XOR2_X1 U156 ( .A(n20), .B(temp_0_2[4]), .Z(n16) );
  NAND2_X1 U157 ( .A1(v_reg_2_1[4]), .A2(a_reg_2[4]), .ZN(n18) );
  XOR2_X1 U158 ( .A(n61), .B(n62), .Z(port_c_1[0]) );
  XNOR2_X1 U159 ( .A(n63), .B(n64), .ZN(n62) );
  XOR2_X1 U160 ( .A(n65), .B(temp_0_1[0]), .Z(n61) );
  NAND2_X1 U161 ( .A1(v_reg_1_1[0]), .A2(a_reg_1[0]), .ZN(n63) );
  XOR2_X1 U162 ( .A(n56), .B(n57), .Z(port_c_1[1]) );
  XNOR2_X1 U163 ( .A(n58), .B(n59), .ZN(n57) );
  XOR2_X1 U164 ( .A(n60), .B(temp_0_1[1]), .Z(n56) );
  NAND2_X1 U165 ( .A1(v_reg_1_1[1]), .A2(a_reg_1[1]), .ZN(n58) );
  XOR2_X1 U166 ( .A(n51), .B(n52), .Z(port_c_1[2]) );
  XNOR2_X1 U167 ( .A(n53), .B(n54), .ZN(n52) );
  XOR2_X1 U168 ( .A(n55), .B(temp_0_1[2]), .Z(n51) );
  NAND2_X1 U169 ( .A1(v_reg_1_1[2]), .A2(a_reg_1[2]), .ZN(n53) );
  XOR2_X1 U170 ( .A(n46), .B(n47), .Z(port_c_1[3]) );
  XNOR2_X1 U171 ( .A(n48), .B(n49), .ZN(n47) );
  XOR2_X1 U172 ( .A(n50), .B(temp_0_1[3]), .Z(n46) );
  NAND2_X1 U173 ( .A1(v_reg_1_1[3]), .A2(a_reg_1[3]), .ZN(n48) );
  XOR2_X1 U174 ( .A(n41), .B(n42), .Z(port_c_1[4]) );
  XNOR2_X1 U175 ( .A(n43), .B(n44), .ZN(n42) );
  XOR2_X1 U176 ( .A(n45), .B(temp_0_1[4]), .Z(n41) );
  NAND2_X1 U177 ( .A1(v_reg_1_1[4]), .A2(a_reg_1[4]), .ZN(n43) );
  XOR2_X1 U178 ( .A(n86), .B(n87), .Z(port_c_0[0]) );
  XNOR2_X1 U179 ( .A(n88), .B(n89), .ZN(n87) );
  XOR2_X1 U180 ( .A(n90), .B(temp_0_0[0]), .Z(n86) );
  NAND2_X1 U181 ( .A1(v_reg_0_1[0]), .A2(a_reg_0[0]), .ZN(n88) );
  XOR2_X1 U182 ( .A(n81), .B(n82), .Z(port_c_0[1]) );
  XNOR2_X1 U183 ( .A(n83), .B(n84), .ZN(n82) );
  XOR2_X1 U184 ( .A(n85), .B(temp_0_0[1]), .Z(n81) );
  NAND2_X1 U185 ( .A1(v_reg_0_1[1]), .A2(a_reg_0[1]), .ZN(n83) );
  XOR2_X1 U186 ( .A(n76), .B(n77), .Z(port_c_0[2]) );
  XNOR2_X1 U187 ( .A(n78), .B(n79), .ZN(n77) );
  XOR2_X1 U188 ( .A(n80), .B(temp_0_0[2]), .Z(n76) );
  NAND2_X1 U189 ( .A1(v_reg_0_1[2]), .A2(a_reg_0[2]), .ZN(n78) );
  XOR2_X1 U190 ( .A(n71), .B(n72), .Z(port_c_0[3]) );
  XNOR2_X1 U191 ( .A(n73), .B(n74), .ZN(n72) );
  XOR2_X1 U192 ( .A(n75), .B(temp_0_0[3]), .Z(n71) );
  NAND2_X1 U193 ( .A1(v_reg_0_1[3]), .A2(a_reg_0[3]), .ZN(n73) );
  XOR2_X1 U194 ( .A(n66), .B(n67), .Z(port_c_0[4]) );
  XNOR2_X1 U195 ( .A(n68), .B(n69), .ZN(n67) );
  XOR2_X1 U196 ( .A(n70), .B(temp_0_0[4]), .Z(n66) );
  NAND2_X1 U197 ( .A1(v_reg_0_1[4]), .A2(a_reg_0[4]), .ZN(n68) );
  NAND2_X1 U198 ( .A1(v_reg_2_0[0]), .A2(a_reg_2[0]), .ZN(n39) );
  NAND2_X1 U199 ( .A1(v_reg_2_0[1]), .A2(a_reg_2[1]), .ZN(n34) );
  NAND2_X1 U200 ( .A1(v_reg_2_0[2]), .A2(a_reg_2[2]), .ZN(n29) );
  NAND2_X1 U201 ( .A1(v_reg_2_0[3]), .A2(a_reg_2[3]), .ZN(n24) );
  NAND2_X1 U202 ( .A1(v_reg_2_0[4]), .A2(a_reg_2[4]), .ZN(n19) );
  NAND2_X1 U203 ( .A1(v_reg_1_0[0]), .A2(a_reg_1[0]), .ZN(n64) );
  NAND2_X1 U204 ( .A1(v_reg_1_0[1]), .A2(a_reg_1[1]), .ZN(n59) );
  NAND2_X1 U205 ( .A1(v_reg_1_0[2]), .A2(a_reg_1[2]), .ZN(n54) );
  NAND2_X1 U206 ( .A1(v_reg_1_0[3]), .A2(a_reg_1[3]), .ZN(n49) );
  NAND2_X1 U207 ( .A1(v_reg_1_0[4]), .A2(a_reg_1[4]), .ZN(n44) );
  NAND2_X1 U208 ( .A1(v_reg_0_0[0]), .A2(a_reg_0[0]), .ZN(n89) );
  NAND2_X1 U209 ( .A1(v_reg_0_0[1]), .A2(a_reg_0[1]), .ZN(n84) );
  NAND2_X1 U210 ( .A1(v_reg_0_0[2]), .A2(a_reg_0[2]), .ZN(n79) );
  NAND2_X1 U211 ( .A1(v_reg_0_0[3]), .A2(a_reg_0[3]), .ZN(n74) );
  NAND2_X1 U212 ( .A1(v_reg_0_0[4]), .A2(a_reg_0[4]), .ZN(n69) );
  INV_X1 U213 ( .A(port_a_2[2]), .ZN(n13) );
  INV_X1 U214 ( .A(port_a_2[1]), .ZN(n14) );
  INV_X1 U215 ( .A(port_a_2[0]), .ZN(n15) );
  INV_X1 U216 ( .A(port_a_2[4]), .ZN(n11) );
  INV_X1 U217 ( .A(port_a_2[3]), .ZN(n12) );
  INV_X1 U218 ( .A(port_a_1[2]), .ZN(n8) );
  INV_X1 U219 ( .A(port_a_1[1]), .ZN(n9) );
  INV_X1 U220 ( .A(port_a_1[0]), .ZN(n10) );
  INV_X1 U221 ( .A(port_a_1[4]), .ZN(n6) );
  INV_X1 U222 ( .A(port_a_1[3]), .ZN(n7) );
  INV_X1 U223 ( .A(port_a_0[2]), .ZN(n3) );
  INV_X1 U224 ( .A(port_a_0[1]), .ZN(n4) );
  INV_X1 U225 ( .A(port_a_0[0]), .ZN(n5) );
  INV_X1 U226 ( .A(port_a_0[4]), .ZN(n1) );
  INV_X1 U227 ( .A(port_a_0[3]), .ZN(n2) );
  AND2_X1 U228 ( .A1(port_b_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U229 ( .A1(port_b_0[1]), .A2(port_a_0[1]), .ZN(N3) );
  AND2_X1 U230 ( .A1(port_b_0[2]), .A2(port_a_0[2]), .ZN(N6) );
  AND2_X1 U231 ( .A1(port_b_0[3]), .A2(port_a_0[3]), .ZN(N9) );
  AND2_X1 U232 ( .A1(port_b_0[4]), .A2(port_a_0[4]), .ZN(N12) );
  AND2_X1 U233 ( .A1(port_b_1[0]), .A2(port_a_1[0]), .ZN(N1) );
  AND2_X1 U234 ( .A1(port_b_1[1]), .A2(port_a_1[1]), .ZN(N4) );
  AND2_X1 U235 ( .A1(port_b_1[2]), .A2(port_a_1[2]), .ZN(N7) );
  AND2_X1 U236 ( .A1(port_b_1[3]), .A2(port_a_1[3]), .ZN(N10) );
  AND2_X1 U237 ( .A1(port_b_1[4]), .A2(port_a_1[4]), .ZN(N13) );
  AND2_X1 U238 ( .A1(port_b_2[0]), .A2(port_a_2[0]), .ZN(N2) );
  AND2_X1 U239 ( .A1(port_b_2[1]), .A2(port_a_2[1]), .ZN(N5) );
  AND2_X1 U240 ( .A1(port_b_2[2]), .A2(port_a_2[2]), .ZN(N8) );
  AND2_X1 U241 ( .A1(port_b_2[3]), .A2(port_a_2[3]), .ZN(N11) );
  AND2_X1 U242 ( .A1(port_b_2[4]), .A2(port_a_2[4]), .ZN(N14) );
  AND2_X1 simpleAnd_30_U1 ( .A1(port_rand_mul[0]), .A2(n5), .ZN(
        simpleAnd_30_port_z) );
  XOR2_X2 simpleXor_60_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_30_port_z), .Z(
        u_0_0[0]) );
  XOR2_X2 simpleXor_61_U1 ( .A(port_rand_mul[0]), .B(port_b_1[0]), .Z(v_0_0[0]) );
  AND2_X1 simpleAnd_31_U1 ( .A1(port_rand_mul[1]), .A2(n5), .ZN(
        simpleAnd_31_port_z) );
  XOR2_X2 simpleXor_62_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_31_port_z), .Z(
        u_0_1[0]) );
  XOR2_X2 simpleXor_63_U1 ( .A(port_rand_mul[1]), .B(port_b_2[0]), .Z(v_0_1[0]) );
  AND2_X1 simpleAnd_32_U1 ( .A1(port_rand_mul[0]), .A2(n10), .ZN(
        simpleAnd_32_port_z) );
  XOR2_X2 simpleXor_64_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_32_port_z), .Z(
        u_1_0[0]) );
  XOR2_X2 simpleXor_65_U1 ( .A(port_rand_mul[0]), .B(port_b_0[0]), .Z(v_1_0[0]) );
  AND2_X1 simpleAnd_33_U1 ( .A1(port_rand_mul[2]), .A2(n10), .ZN(
        simpleAnd_33_port_z) );
  XOR2_X2 simpleXor_66_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_33_port_z), .Z(
        u_1_1[0]) );
  XOR2_X2 simpleXor_67_U1 ( .A(port_rand_mul[2]), .B(port_b_2[0]), .Z(v_1_1[0]) );
  AND2_X1 simpleAnd_34_U1 ( .A1(port_rand_mul[1]), .A2(n15), .ZN(
        simpleAnd_34_port_z) );
  XOR2_X2 simpleXor_68_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_34_port_z), .Z(
        u_2_0[0]) );
  XOR2_X2 simpleXor_69_U1 ( .A(port_rand_mul[1]), .B(port_b_0[0]), .Z(v_2_0[0]) );
  AND2_X1 simpleAnd_35_U1 ( .A1(port_rand_mul[2]), .A2(n15), .ZN(
        simpleAnd_35_port_z) );
  XOR2_X2 simpleXor_70_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_35_port_z), .Z(
        u_2_1[0]) );
  XOR2_X2 simpleXor_71_U1 ( .A(port_rand_mul[2]), .B(port_b_1[0]), .Z(v_2_1[0]) );
  AND2_X1 simpleAnd_36_U1 ( .A1(port_rand_mul[0]), .A2(n4), .ZN(
        simpleAnd_36_port_z) );
  XOR2_X2 simpleXor_72_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_36_port_z), .Z(
        u_0_0[1]) );
  XOR2_X2 simpleXor_73_U1 ( .A(port_rand_mul[0]), .B(port_b_1[1]), .Z(v_0_0[1]) );
  AND2_X1 simpleAnd_37_U1 ( .A1(port_rand_mul[1]), .A2(n4), .ZN(
        simpleAnd_37_port_z) );
  XOR2_X2 simpleXor_74_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_37_port_z), .Z(
        u_0_1[1]) );
  XOR2_X2 simpleXor_75_U1 ( .A(port_rand_mul[1]), .B(port_b_2[1]), .Z(v_0_1[1]) );
  AND2_X1 simpleAnd_38_U1 ( .A1(port_rand_mul[0]), .A2(n9), .ZN(
        simpleAnd_38_port_z) );
  XOR2_X2 simpleXor_76_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_38_port_z), .Z(
        u_1_0[1]) );
  XOR2_X2 simpleXor_77_U1 ( .A(port_rand_mul[0]), .B(port_b_0[1]), .Z(v_1_0[1]) );
  AND2_X1 simpleAnd_39_U1 ( .A1(port_rand_mul[2]), .A2(n9), .ZN(
        simpleAnd_39_port_z) );
  XOR2_X2 simpleXor_78_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_39_port_z), .Z(
        u_1_1[1]) );
  XOR2_X2 simpleXor_79_U1 ( .A(port_rand_mul[2]), .B(port_b_2[1]), .Z(v_1_1[1]) );
  AND2_X1 simpleAnd_40_U1 ( .A1(port_rand_mul[1]), .A2(n14), .ZN(
        simpleAnd_40_port_z) );
  XOR2_X2 simpleXor_80_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_40_port_z), .Z(
        u_2_0[1]) );
  XOR2_X2 simpleXor_81_U1 ( .A(port_rand_mul[1]), .B(port_b_0[1]), .Z(v_2_0[1]) );
  AND2_X1 simpleAnd_41_U1 ( .A1(port_rand_mul[2]), .A2(n14), .ZN(
        simpleAnd_41_port_z) );
  XOR2_X2 simpleXor_82_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_41_port_z), .Z(
        u_2_1[1]) );
  XOR2_X2 simpleXor_83_U1 ( .A(port_rand_mul[2]), .B(port_b_1[1]), .Z(v_2_1[1]) );
  AND2_X1 simpleAnd_42_U1 ( .A1(port_rand_mul[0]), .A2(n3), .ZN(
        simpleAnd_42_port_z) );
  XOR2_X2 simpleXor_84_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_42_port_z), .Z(
        u_0_0[2]) );
  XOR2_X2 simpleXor_85_U1 ( .A(port_rand_mul[0]), .B(port_b_1[2]), .Z(v_0_0[2]) );
  AND2_X1 simpleAnd_43_U1 ( .A1(port_rand_mul[1]), .A2(n3), .ZN(
        simpleAnd_43_port_z) );
  XOR2_X2 simpleXor_86_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_43_port_z), .Z(
        u_0_1[2]) );
  XOR2_X2 simpleXor_87_U1 ( .A(port_rand_mul[1]), .B(port_b_2[2]), .Z(v_0_1[2]) );
  AND2_X1 simpleAnd_44_U1 ( .A1(port_rand_mul[0]), .A2(n8), .ZN(
        simpleAnd_44_port_z) );
  XOR2_X2 simpleXor_88_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_44_port_z), .Z(
        u_1_0[2]) );
  XOR2_X2 simpleXor_89_U1 ( .A(port_rand_mul[0]), .B(port_b_0[2]), .Z(v_1_0[2]) );
  AND2_X1 simpleAnd_45_U1 ( .A1(port_rand_mul[2]), .A2(n8), .ZN(
        simpleAnd_45_port_z) );
  XOR2_X2 simpleXor_90_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_45_port_z), .Z(
        u_1_1[2]) );
  XOR2_X2 simpleXor_91_U1 ( .A(port_rand_mul[2]), .B(port_b_2[2]), .Z(v_1_1[2]) );
  AND2_X1 simpleAnd_46_U1 ( .A1(port_rand_mul[1]), .A2(n13), .ZN(
        simpleAnd_46_port_z) );
  XOR2_X2 simpleXor_92_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_46_port_z), .Z(
        u_2_0[2]) );
  XOR2_X2 simpleXor_93_U1 ( .A(port_rand_mul[1]), .B(port_b_0[2]), .Z(v_2_0[2]) );
  AND2_X1 simpleAnd_47_U1 ( .A1(port_rand_mul[2]), .A2(n13), .ZN(
        simpleAnd_47_port_z) );
  XOR2_X2 simpleXor_94_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_47_port_z), .Z(
        u_2_1[2]) );
  XOR2_X2 simpleXor_95_U1 ( .A(port_rand_mul[2]), .B(port_b_1[2]), .Z(v_2_1[2]) );
  AND2_X1 simpleAnd_48_U1 ( .A1(port_rand_mul[0]), .A2(n2), .ZN(
        simpleAnd_48_port_z) );
  XOR2_X2 simpleXor_96_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_48_port_z), .Z(
        u_0_0[3]) );
  XOR2_X2 simpleXor_97_U1 ( .A(port_rand_mul[0]), .B(port_b_1[3]), .Z(v_0_0[3]) );
  AND2_X1 simpleAnd_49_U1 ( .A1(port_rand_mul[1]), .A2(n2), .ZN(
        simpleAnd_49_port_z) );
  XOR2_X2 simpleXor_98_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_49_port_z), .Z(
        u_0_1[3]) );
  XOR2_X2 simpleXor_99_U1 ( .A(port_rand_mul[1]), .B(port_b_2[3]), .Z(v_0_1[3]) );
  AND2_X1 simpleAnd_50_U1 ( .A1(port_rand_mul[0]), .A2(n7), .ZN(
        simpleAnd_50_port_z) );
  XOR2_X2 simpleXor_100_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_50_port_z), 
        .Z(u_1_0[3]) );
  XOR2_X2 simpleXor_101_U1 ( .A(port_rand_mul[0]), .B(port_b_0[3]), .Z(
        v_1_0[3]) );
  AND2_X1 simpleAnd_51_U1 ( .A1(port_rand_mul[2]), .A2(n7), .ZN(
        simpleAnd_51_port_z) );
  XOR2_X2 simpleXor_102_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_51_port_z), 
        .Z(u_1_1[3]) );
  XOR2_X2 simpleXor_103_U1 ( .A(port_rand_mul[2]), .B(port_b_2[3]), .Z(
        v_1_1[3]) );
  AND2_X1 simpleAnd_52_U1 ( .A1(port_rand_mul[1]), .A2(n12), .ZN(
        simpleAnd_52_port_z) );
  XOR2_X2 simpleXor_104_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_52_port_z), 
        .Z(u_2_0[3]) );
  XOR2_X2 simpleXor_105_U1 ( .A(port_rand_mul[1]), .B(port_b_0[3]), .Z(
        v_2_0[3]) );
  AND2_X1 simpleAnd_53_U1 ( .A1(port_rand_mul[2]), .A2(n12), .ZN(
        simpleAnd_53_port_z) );
  XOR2_X2 simpleXor_106_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_53_port_z), 
        .Z(u_2_1[3]) );
  XOR2_X2 simpleXor_107_U1 ( .A(port_rand_mul[2]), .B(port_b_1[3]), .Z(
        v_2_1[3]) );
  AND2_X1 simpleAnd_54_U1 ( .A1(port_rand_mul[0]), .A2(n1), .ZN(
        simpleAnd_54_port_z) );
  XOR2_X2 simpleXor_108_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_54_port_z), 
        .Z(u_0_0[4]) );
  XOR2_X2 simpleXor_109_U1 ( .A(port_rand_mul[0]), .B(port_b_1[4]), .Z(
        v_0_0[4]) );
  AND2_X1 simpleAnd_55_U1 ( .A1(port_rand_mul[1]), .A2(n1), .ZN(
        simpleAnd_55_port_z) );
  XOR2_X2 simpleXor_110_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_55_port_z), 
        .Z(u_0_1[4]) );
  XOR2_X2 simpleXor_111_U1 ( .A(port_rand_mul[1]), .B(port_b_2[4]), .Z(
        v_0_1[4]) );
  AND2_X1 simpleAnd_56_U1 ( .A1(port_rand_mul[0]), .A2(n6), .ZN(
        simpleAnd_56_port_z) );
  XOR2_X2 simpleXor_112_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_56_port_z), 
        .Z(u_1_0[4]) );
  XOR2_X2 simpleXor_113_U1 ( .A(port_rand_mul[0]), .B(port_b_0[4]), .Z(
        v_1_0[4]) );
  AND2_X1 simpleAnd_57_U1 ( .A1(port_rand_mul[2]), .A2(n6), .ZN(
        simpleAnd_57_port_z) );
  XOR2_X2 simpleXor_114_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_57_port_z), 
        .Z(u_1_1[4]) );
  XOR2_X2 simpleXor_115_U1 ( .A(port_rand_mul[2]), .B(port_b_2[4]), .Z(
        v_1_1[4]) );
  AND2_X1 simpleAnd_58_U1 ( .A1(port_rand_mul[1]), .A2(n11), .ZN(
        simpleAnd_58_port_z) );
  XOR2_X2 simpleXor_116_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_58_port_z), 
        .Z(u_2_0[4]) );
  XOR2_X2 simpleXor_117_U1 ( .A(port_rand_mul[1]), .B(port_b_0[4]), .Z(
        v_2_0[4]) );
  AND2_X1 simpleAnd_59_U1 ( .A1(port_rand_mul[2]), .A2(n11), .ZN(
        simpleAnd_59_port_z) );
  XOR2_X2 simpleXor_118_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_59_port_z), 
        .Z(u_2_1[4]) );
  XOR2_X2 simpleXor_119_U1 ( .A(port_rand_mul[2]), .B(port_b_1[4]), .Z(
        v_2_1[4]) );
  NAND2_X1 maj_60_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_60_n9) );
  NAND2_X1 maj_60_U14 ( .A1(maj_60_n6), .A2(maj_60_n5), .ZN(maj_60_n10) );
  NAND2_X1 maj_60_U13 ( .A1(maj_60_n9), .A2(maj_60_n10), .ZN(maj_60_n8) );
  NAND2_X1 maj_60_U12 ( .A1(u_0_0[2]), .A2(maj_60_n11), .ZN(maj_60_n13) );
  NAND2_X1 maj_60_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_60_n12) );
  NAND2_X1 maj_60_U10 ( .A1(maj_60_n12), .A2(maj_60_n13), .ZN(maj_60_n7) );
  XOR2_X1 maj_60_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_60_n5) );
  XOR2_X1 maj_60_U8 ( .A(u_0_0[2]), .B(maj_60_n11), .Z(maj_60_n6) );
  XOR2_X1 maj_60_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_60_n11) );
  OR2_X1 maj_60_U6 ( .A1(maj_60_n7), .A2(maj_60_n8), .ZN(maj_60_n3) );
  NAND2_X1 maj_60_U5 ( .A1(maj_60_n3), .A2(maj_60_n4), .ZN(maj_60_n2) );
  NAND2_X1 maj_60_U4 ( .A1(maj_60_n7), .A2(maj_60_n8), .ZN(maj_60_n1) );
  NAND2_X1 maj_60_U3 ( .A1(maj_60_n1), .A2(maj_60_n2), .ZN(maj_60_port_o) );
  XOR2_X1 maj_60_U2 ( .A(maj_60_n5), .B(maj_60_n6), .Z(maj_60_n4) );
  NAND2_X1 maj_61_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_61_n18) );
  NAND2_X1 maj_61_U14 ( .A1(maj_61_n21), .A2(maj_61_n22), .ZN(maj_61_n17) );
  NAND2_X1 maj_61_U13 ( .A1(maj_61_n18), .A2(maj_61_n17), .ZN(maj_61_n19) );
  NAND2_X1 maj_61_U12 ( .A1(v_0_0[2]), .A2(maj_61_n16), .ZN(maj_61_n14) );
  NAND2_X1 maj_61_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_61_n15) );
  NAND2_X1 maj_61_U10 ( .A1(maj_61_n15), .A2(maj_61_n14), .ZN(maj_61_n20) );
  XOR2_X1 maj_61_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_61_n22) );
  XOR2_X1 maj_61_U8 ( .A(v_0_0[2]), .B(maj_61_n16), .Z(maj_61_n21) );
  XOR2_X1 maj_61_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_61_n16) );
  OR2_X1 maj_61_U6 ( .A1(maj_61_n20), .A2(maj_61_n19), .ZN(maj_61_n24) );
  NAND2_X1 maj_61_U5 ( .A1(maj_61_n24), .A2(maj_61_n23), .ZN(maj_61_n25) );
  NAND2_X1 maj_61_U4 ( .A1(maj_61_n20), .A2(maj_61_n19), .ZN(maj_61_n26) );
  NAND2_X1 maj_61_U3 ( .A1(maj_61_n26), .A2(maj_61_n25), .ZN(maj_61_port_o) );
  XOR2_X1 maj_61_U2 ( .A(maj_61_n22), .B(maj_61_n21), .Z(maj_61_n23) );
  NAND2_X1 maj_62_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_62_n18) );
  NAND2_X1 maj_62_U14 ( .A1(maj_62_n21), .A2(maj_62_n22), .ZN(maj_62_n17) );
  NAND2_X1 maj_62_U13 ( .A1(maj_62_n18), .A2(maj_62_n17), .ZN(maj_62_n19) );
  NAND2_X1 maj_62_U12 ( .A1(u_0_1[2]), .A2(maj_62_n16), .ZN(maj_62_n14) );
  NAND2_X1 maj_62_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_62_n15) );
  NAND2_X1 maj_62_U10 ( .A1(maj_62_n15), .A2(maj_62_n14), .ZN(maj_62_n20) );
  XOR2_X1 maj_62_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_62_n22) );
  XOR2_X1 maj_62_U8 ( .A(u_0_1[2]), .B(maj_62_n16), .Z(maj_62_n21) );
  XOR2_X1 maj_62_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_62_n16) );
  OR2_X1 maj_62_U6 ( .A1(maj_62_n20), .A2(maj_62_n19), .ZN(maj_62_n24) );
  NAND2_X1 maj_62_U5 ( .A1(maj_62_n24), .A2(maj_62_n23), .ZN(maj_62_n25) );
  NAND2_X1 maj_62_U4 ( .A1(maj_62_n20), .A2(maj_62_n19), .ZN(maj_62_n26) );
  NAND2_X1 maj_62_U3 ( .A1(maj_62_n26), .A2(maj_62_n25), .ZN(maj_62_port_o) );
  XOR2_X1 maj_62_U2 ( .A(maj_62_n22), .B(maj_62_n21), .Z(maj_62_n23) );
  NAND2_X1 maj_63_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_63_n18) );
  NAND2_X1 maj_63_U14 ( .A1(maj_63_n21), .A2(maj_63_n22), .ZN(maj_63_n17) );
  NAND2_X1 maj_63_U13 ( .A1(maj_63_n18), .A2(maj_63_n17), .ZN(maj_63_n19) );
  NAND2_X1 maj_63_U12 ( .A1(v_0_1[2]), .A2(maj_63_n16), .ZN(maj_63_n14) );
  NAND2_X1 maj_63_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_63_n15) );
  NAND2_X1 maj_63_U10 ( .A1(maj_63_n15), .A2(maj_63_n14), .ZN(maj_63_n20) );
  XOR2_X1 maj_63_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_63_n22) );
  XOR2_X1 maj_63_U8 ( .A(v_0_1[2]), .B(maj_63_n16), .Z(maj_63_n21) );
  XOR2_X1 maj_63_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_63_n16) );
  OR2_X1 maj_63_U6 ( .A1(maj_63_n20), .A2(maj_63_n19), .ZN(maj_63_n24) );
  NAND2_X1 maj_63_U5 ( .A1(maj_63_n24), .A2(maj_63_n23), .ZN(maj_63_n25) );
  NAND2_X1 maj_63_U4 ( .A1(maj_63_n20), .A2(maj_63_n19), .ZN(maj_63_n26) );
  NAND2_X1 maj_63_U3 ( .A1(maj_63_n26), .A2(maj_63_n25), .ZN(maj_63_port_o) );
  XOR2_X1 maj_63_U2 ( .A(maj_63_n22), .B(maj_63_n21), .Z(maj_63_n23) );
  NAND2_X1 maj_64_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_64_n18) );
  NAND2_X1 maj_64_U14 ( .A1(maj_64_n21), .A2(maj_64_n22), .ZN(maj_64_n17) );
  NAND2_X1 maj_64_U13 ( .A1(maj_64_n18), .A2(maj_64_n17), .ZN(maj_64_n19) );
  NAND2_X1 maj_64_U12 ( .A1(u_1_0[2]), .A2(maj_64_n16), .ZN(maj_64_n14) );
  NAND2_X1 maj_64_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_64_n15) );
  NAND2_X1 maj_64_U10 ( .A1(maj_64_n15), .A2(maj_64_n14), .ZN(maj_64_n20) );
  XOR2_X1 maj_64_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_64_n22) );
  XOR2_X1 maj_64_U8 ( .A(u_1_0[2]), .B(maj_64_n16), .Z(maj_64_n21) );
  XOR2_X1 maj_64_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_64_n16) );
  OR2_X1 maj_64_U6 ( .A1(maj_64_n20), .A2(maj_64_n19), .ZN(maj_64_n24) );
  NAND2_X1 maj_64_U5 ( .A1(maj_64_n24), .A2(maj_64_n23), .ZN(maj_64_n25) );
  NAND2_X1 maj_64_U4 ( .A1(maj_64_n20), .A2(maj_64_n19), .ZN(maj_64_n26) );
  NAND2_X1 maj_64_U3 ( .A1(maj_64_n26), .A2(maj_64_n25), .ZN(maj_64_port_o) );
  XOR2_X1 maj_64_U2 ( .A(maj_64_n22), .B(maj_64_n21), .Z(maj_64_n23) );
  NAND2_X1 maj_65_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_65_n18) );
  NAND2_X1 maj_65_U14 ( .A1(maj_65_n21), .A2(maj_65_n22), .ZN(maj_65_n17) );
  NAND2_X1 maj_65_U13 ( .A1(maj_65_n18), .A2(maj_65_n17), .ZN(maj_65_n19) );
  NAND2_X1 maj_65_U12 ( .A1(v_1_0[2]), .A2(maj_65_n16), .ZN(maj_65_n14) );
  NAND2_X1 maj_65_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_65_n15) );
  NAND2_X1 maj_65_U10 ( .A1(maj_65_n15), .A2(maj_65_n14), .ZN(maj_65_n20) );
  XOR2_X1 maj_65_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_65_n22) );
  XOR2_X1 maj_65_U8 ( .A(v_1_0[2]), .B(maj_65_n16), .Z(maj_65_n21) );
  XOR2_X1 maj_65_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_65_n16) );
  OR2_X1 maj_65_U6 ( .A1(maj_65_n20), .A2(maj_65_n19), .ZN(maj_65_n24) );
  NAND2_X1 maj_65_U5 ( .A1(maj_65_n24), .A2(maj_65_n23), .ZN(maj_65_n25) );
  NAND2_X1 maj_65_U4 ( .A1(maj_65_n20), .A2(maj_65_n19), .ZN(maj_65_n26) );
  NAND2_X1 maj_65_U3 ( .A1(maj_65_n26), .A2(maj_65_n25), .ZN(maj_65_port_o) );
  XOR2_X1 maj_65_U2 ( .A(maj_65_n22), .B(maj_65_n21), .Z(maj_65_n23) );
  NAND2_X1 maj_66_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_66_n18) );
  NAND2_X1 maj_66_U14 ( .A1(maj_66_n21), .A2(maj_66_n22), .ZN(maj_66_n17) );
  NAND2_X1 maj_66_U13 ( .A1(maj_66_n18), .A2(maj_66_n17), .ZN(maj_66_n19) );
  NAND2_X1 maj_66_U12 ( .A1(u_1_1[2]), .A2(maj_66_n16), .ZN(maj_66_n14) );
  NAND2_X1 maj_66_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_66_n15) );
  NAND2_X1 maj_66_U10 ( .A1(maj_66_n15), .A2(maj_66_n14), .ZN(maj_66_n20) );
  XOR2_X1 maj_66_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_66_n22) );
  XOR2_X1 maj_66_U8 ( .A(u_1_1[2]), .B(maj_66_n16), .Z(maj_66_n21) );
  XOR2_X1 maj_66_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_66_n16) );
  OR2_X1 maj_66_U6 ( .A1(maj_66_n20), .A2(maj_66_n19), .ZN(maj_66_n24) );
  NAND2_X1 maj_66_U5 ( .A1(maj_66_n24), .A2(maj_66_n23), .ZN(maj_66_n25) );
  NAND2_X1 maj_66_U4 ( .A1(maj_66_n20), .A2(maj_66_n19), .ZN(maj_66_n26) );
  NAND2_X1 maj_66_U3 ( .A1(maj_66_n26), .A2(maj_66_n25), .ZN(maj_66_port_o) );
  XOR2_X1 maj_66_U2 ( .A(maj_66_n22), .B(maj_66_n21), .Z(maj_66_n23) );
  NAND2_X1 maj_67_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_67_n18) );
  NAND2_X1 maj_67_U14 ( .A1(maj_67_n21), .A2(maj_67_n22), .ZN(maj_67_n17) );
  NAND2_X1 maj_67_U13 ( .A1(maj_67_n18), .A2(maj_67_n17), .ZN(maj_67_n19) );
  NAND2_X1 maj_67_U12 ( .A1(v_1_1[2]), .A2(maj_67_n16), .ZN(maj_67_n14) );
  NAND2_X1 maj_67_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_67_n15) );
  NAND2_X1 maj_67_U10 ( .A1(maj_67_n15), .A2(maj_67_n14), .ZN(maj_67_n20) );
  XOR2_X1 maj_67_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_67_n22) );
  XOR2_X1 maj_67_U8 ( .A(v_1_1[2]), .B(maj_67_n16), .Z(maj_67_n21) );
  XOR2_X1 maj_67_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_67_n16) );
  OR2_X1 maj_67_U6 ( .A1(maj_67_n20), .A2(maj_67_n19), .ZN(maj_67_n24) );
  NAND2_X1 maj_67_U5 ( .A1(maj_67_n24), .A2(maj_67_n23), .ZN(maj_67_n25) );
  NAND2_X1 maj_67_U4 ( .A1(maj_67_n20), .A2(maj_67_n19), .ZN(maj_67_n26) );
  NAND2_X1 maj_67_U3 ( .A1(maj_67_n26), .A2(maj_67_n25), .ZN(maj_67_port_o) );
  XOR2_X1 maj_67_U2 ( .A(maj_67_n22), .B(maj_67_n21), .Z(maj_67_n23) );
  NAND2_X1 maj_68_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_68_n18) );
  NAND2_X1 maj_68_U14 ( .A1(maj_68_n21), .A2(maj_68_n22), .ZN(maj_68_n17) );
  NAND2_X1 maj_68_U13 ( .A1(maj_68_n18), .A2(maj_68_n17), .ZN(maj_68_n19) );
  NAND2_X1 maj_68_U12 ( .A1(u_2_0[2]), .A2(maj_68_n16), .ZN(maj_68_n14) );
  NAND2_X1 maj_68_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_68_n15) );
  NAND2_X1 maj_68_U10 ( .A1(maj_68_n15), .A2(maj_68_n14), .ZN(maj_68_n20) );
  XOR2_X1 maj_68_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_68_n22) );
  XOR2_X1 maj_68_U8 ( .A(u_2_0[2]), .B(maj_68_n16), .Z(maj_68_n21) );
  XOR2_X1 maj_68_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_68_n16) );
  OR2_X1 maj_68_U6 ( .A1(maj_68_n20), .A2(maj_68_n19), .ZN(maj_68_n24) );
  NAND2_X1 maj_68_U5 ( .A1(maj_68_n24), .A2(maj_68_n23), .ZN(maj_68_n25) );
  NAND2_X1 maj_68_U4 ( .A1(maj_68_n20), .A2(maj_68_n19), .ZN(maj_68_n26) );
  NAND2_X1 maj_68_U3 ( .A1(maj_68_n26), .A2(maj_68_n25), .ZN(maj_68_port_o) );
  XOR2_X1 maj_68_U2 ( .A(maj_68_n22), .B(maj_68_n21), .Z(maj_68_n23) );
  NAND2_X1 maj_69_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_69_n18) );
  NAND2_X1 maj_69_U14 ( .A1(maj_69_n21), .A2(maj_69_n22), .ZN(maj_69_n17) );
  NAND2_X1 maj_69_U13 ( .A1(maj_69_n18), .A2(maj_69_n17), .ZN(maj_69_n19) );
  NAND2_X1 maj_69_U12 ( .A1(v_2_0[2]), .A2(maj_69_n16), .ZN(maj_69_n14) );
  NAND2_X1 maj_69_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_69_n15) );
  NAND2_X1 maj_69_U10 ( .A1(maj_69_n15), .A2(maj_69_n14), .ZN(maj_69_n20) );
  XOR2_X1 maj_69_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_69_n22) );
  XOR2_X1 maj_69_U8 ( .A(v_2_0[2]), .B(maj_69_n16), .Z(maj_69_n21) );
  XOR2_X1 maj_69_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_69_n16) );
  OR2_X1 maj_69_U6 ( .A1(maj_69_n20), .A2(maj_69_n19), .ZN(maj_69_n24) );
  NAND2_X1 maj_69_U5 ( .A1(maj_69_n24), .A2(maj_69_n23), .ZN(maj_69_n25) );
  NAND2_X1 maj_69_U4 ( .A1(maj_69_n20), .A2(maj_69_n19), .ZN(maj_69_n26) );
  NAND2_X1 maj_69_U3 ( .A1(maj_69_n26), .A2(maj_69_n25), .ZN(maj_69_port_o) );
  XOR2_X1 maj_69_U2 ( .A(maj_69_n22), .B(maj_69_n21), .Z(maj_69_n23) );
  NAND2_X1 maj_70_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_70_n18) );
  NAND2_X1 maj_70_U14 ( .A1(maj_70_n21), .A2(maj_70_n22), .ZN(maj_70_n17) );
  NAND2_X1 maj_70_U13 ( .A1(maj_70_n18), .A2(maj_70_n17), .ZN(maj_70_n19) );
  NAND2_X1 maj_70_U12 ( .A1(u_2_1[2]), .A2(maj_70_n16), .ZN(maj_70_n14) );
  NAND2_X1 maj_70_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_70_n15) );
  NAND2_X1 maj_70_U10 ( .A1(maj_70_n15), .A2(maj_70_n14), .ZN(maj_70_n20) );
  XOR2_X1 maj_70_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_70_n22) );
  XOR2_X1 maj_70_U8 ( .A(u_2_1[2]), .B(maj_70_n16), .Z(maj_70_n21) );
  XOR2_X1 maj_70_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_70_n16) );
  OR2_X1 maj_70_U6 ( .A1(maj_70_n20), .A2(maj_70_n19), .ZN(maj_70_n24) );
  NAND2_X1 maj_70_U5 ( .A1(maj_70_n24), .A2(maj_70_n23), .ZN(maj_70_n25) );
  NAND2_X1 maj_70_U4 ( .A1(maj_70_n20), .A2(maj_70_n19), .ZN(maj_70_n26) );
  NAND2_X1 maj_70_U3 ( .A1(maj_70_n26), .A2(maj_70_n25), .ZN(maj_70_port_o) );
  XOR2_X1 maj_70_U2 ( .A(maj_70_n22), .B(maj_70_n21), .Z(maj_70_n23) );
  NAND2_X1 maj_71_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_71_n18) );
  NAND2_X1 maj_71_U14 ( .A1(maj_71_n21), .A2(maj_71_n22), .ZN(maj_71_n17) );
  NAND2_X1 maj_71_U13 ( .A1(maj_71_n18), .A2(maj_71_n17), .ZN(maj_71_n19) );
  NAND2_X1 maj_71_U12 ( .A1(v_2_1[2]), .A2(maj_71_n16), .ZN(maj_71_n14) );
  NAND2_X1 maj_71_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_71_n15) );
  NAND2_X1 maj_71_U10 ( .A1(maj_71_n15), .A2(maj_71_n14), .ZN(maj_71_n20) );
  XOR2_X1 maj_71_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_71_n22) );
  XOR2_X1 maj_71_U8 ( .A(v_2_1[2]), .B(maj_71_n16), .Z(maj_71_n21) );
  XOR2_X1 maj_71_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_71_n16) );
  OR2_X1 maj_71_U6 ( .A1(maj_71_n20), .A2(maj_71_n19), .ZN(maj_71_n24) );
  NAND2_X1 maj_71_U5 ( .A1(maj_71_n24), .A2(maj_71_n23), .ZN(maj_71_n25) );
  NAND2_X1 maj_71_U4 ( .A1(maj_71_n20), .A2(maj_71_n19), .ZN(maj_71_n26) );
  NAND2_X1 maj_71_U3 ( .A1(maj_71_n26), .A2(maj_71_n25), .ZN(maj_71_port_o) );
  XOR2_X1 maj_71_U2 ( .A(maj_71_n22), .B(maj_71_n21), .Z(maj_71_n23) );
  NAND2_X1 maj_72_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_72_n18) );
  NAND2_X1 maj_72_U14 ( .A1(maj_72_n21), .A2(maj_72_n22), .ZN(maj_72_n17) );
  NAND2_X1 maj_72_U13 ( .A1(maj_72_n18), .A2(maj_72_n17), .ZN(maj_72_n19) );
  NAND2_X1 maj_72_U12 ( .A1(u_0_0[2]), .A2(maj_72_n16), .ZN(maj_72_n14) );
  NAND2_X1 maj_72_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_72_n15) );
  NAND2_X1 maj_72_U10 ( .A1(maj_72_n15), .A2(maj_72_n14), .ZN(maj_72_n20) );
  XOR2_X1 maj_72_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_72_n22) );
  XOR2_X1 maj_72_U8 ( .A(u_0_0[2]), .B(maj_72_n16), .Z(maj_72_n21) );
  XOR2_X1 maj_72_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_72_n16) );
  OR2_X1 maj_72_U6 ( .A1(maj_72_n20), .A2(maj_72_n19), .ZN(maj_72_n24) );
  NAND2_X1 maj_72_U5 ( .A1(maj_72_n24), .A2(maj_72_n23), .ZN(maj_72_n25) );
  NAND2_X1 maj_72_U4 ( .A1(maj_72_n20), .A2(maj_72_n19), .ZN(maj_72_n26) );
  NAND2_X1 maj_72_U3 ( .A1(maj_72_n26), .A2(maj_72_n25), .ZN(maj_72_port_o) );
  XOR2_X1 maj_72_U2 ( .A(maj_72_n22), .B(maj_72_n21), .Z(maj_72_n23) );
  NAND2_X1 maj_73_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_73_n18) );
  NAND2_X1 maj_73_U14 ( .A1(maj_73_n21), .A2(maj_73_n22), .ZN(maj_73_n17) );
  NAND2_X1 maj_73_U13 ( .A1(maj_73_n18), .A2(maj_73_n17), .ZN(maj_73_n19) );
  NAND2_X1 maj_73_U12 ( .A1(v_0_0[2]), .A2(maj_73_n16), .ZN(maj_73_n14) );
  NAND2_X1 maj_73_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_73_n15) );
  NAND2_X1 maj_73_U10 ( .A1(maj_73_n15), .A2(maj_73_n14), .ZN(maj_73_n20) );
  XOR2_X1 maj_73_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_73_n22) );
  XOR2_X1 maj_73_U8 ( .A(v_0_0[2]), .B(maj_73_n16), .Z(maj_73_n21) );
  XOR2_X1 maj_73_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_73_n16) );
  OR2_X1 maj_73_U6 ( .A1(maj_73_n20), .A2(maj_73_n19), .ZN(maj_73_n24) );
  NAND2_X1 maj_73_U5 ( .A1(maj_73_n24), .A2(maj_73_n23), .ZN(maj_73_n25) );
  NAND2_X1 maj_73_U4 ( .A1(maj_73_n20), .A2(maj_73_n19), .ZN(maj_73_n26) );
  NAND2_X1 maj_73_U3 ( .A1(maj_73_n26), .A2(maj_73_n25), .ZN(maj_73_port_o) );
  XOR2_X1 maj_73_U2 ( .A(maj_73_n22), .B(maj_73_n21), .Z(maj_73_n23) );
  NAND2_X1 maj_74_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_74_n18) );
  NAND2_X1 maj_74_U14 ( .A1(maj_74_n21), .A2(maj_74_n22), .ZN(maj_74_n17) );
  NAND2_X1 maj_74_U13 ( .A1(maj_74_n18), .A2(maj_74_n17), .ZN(maj_74_n19) );
  NAND2_X1 maj_74_U12 ( .A1(u_0_1[2]), .A2(maj_74_n16), .ZN(maj_74_n14) );
  NAND2_X1 maj_74_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_74_n15) );
  NAND2_X1 maj_74_U10 ( .A1(maj_74_n15), .A2(maj_74_n14), .ZN(maj_74_n20) );
  XOR2_X1 maj_74_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_74_n22) );
  XOR2_X1 maj_74_U8 ( .A(u_0_1[2]), .B(maj_74_n16), .Z(maj_74_n21) );
  XOR2_X1 maj_74_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_74_n16) );
  OR2_X1 maj_74_U6 ( .A1(maj_74_n20), .A2(maj_74_n19), .ZN(maj_74_n24) );
  NAND2_X1 maj_74_U5 ( .A1(maj_74_n24), .A2(maj_74_n23), .ZN(maj_74_n25) );
  NAND2_X1 maj_74_U4 ( .A1(maj_74_n20), .A2(maj_74_n19), .ZN(maj_74_n26) );
  NAND2_X1 maj_74_U3 ( .A1(maj_74_n26), .A2(maj_74_n25), .ZN(maj_74_port_o) );
  XOR2_X1 maj_74_U2 ( .A(maj_74_n22), .B(maj_74_n21), .Z(maj_74_n23) );
  NAND2_X1 maj_75_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_75_n18) );
  NAND2_X1 maj_75_U14 ( .A1(maj_75_n21), .A2(maj_75_n22), .ZN(maj_75_n17) );
  NAND2_X1 maj_75_U13 ( .A1(maj_75_n18), .A2(maj_75_n17), .ZN(maj_75_n19) );
  NAND2_X1 maj_75_U12 ( .A1(v_0_1[2]), .A2(maj_75_n16), .ZN(maj_75_n14) );
  NAND2_X1 maj_75_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_75_n15) );
  NAND2_X1 maj_75_U10 ( .A1(maj_75_n15), .A2(maj_75_n14), .ZN(maj_75_n20) );
  XOR2_X1 maj_75_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_75_n22) );
  XOR2_X1 maj_75_U8 ( .A(v_0_1[2]), .B(maj_75_n16), .Z(maj_75_n21) );
  XOR2_X1 maj_75_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_75_n16) );
  OR2_X1 maj_75_U6 ( .A1(maj_75_n20), .A2(maj_75_n19), .ZN(maj_75_n24) );
  NAND2_X1 maj_75_U5 ( .A1(maj_75_n24), .A2(maj_75_n23), .ZN(maj_75_n25) );
  NAND2_X1 maj_75_U4 ( .A1(maj_75_n20), .A2(maj_75_n19), .ZN(maj_75_n26) );
  NAND2_X1 maj_75_U3 ( .A1(maj_75_n26), .A2(maj_75_n25), .ZN(maj_75_port_o) );
  XOR2_X1 maj_75_U2 ( .A(maj_75_n22), .B(maj_75_n21), .Z(maj_75_n23) );
  NAND2_X1 maj_76_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_76_n18) );
  NAND2_X1 maj_76_U14 ( .A1(maj_76_n21), .A2(maj_76_n22), .ZN(maj_76_n17) );
  NAND2_X1 maj_76_U13 ( .A1(maj_76_n18), .A2(maj_76_n17), .ZN(maj_76_n19) );
  NAND2_X1 maj_76_U12 ( .A1(u_1_0[2]), .A2(maj_76_n16), .ZN(maj_76_n14) );
  NAND2_X1 maj_76_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_76_n15) );
  NAND2_X1 maj_76_U10 ( .A1(maj_76_n15), .A2(maj_76_n14), .ZN(maj_76_n20) );
  XOR2_X1 maj_76_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_76_n22) );
  XOR2_X1 maj_76_U8 ( .A(u_1_0[2]), .B(maj_76_n16), .Z(maj_76_n21) );
  XOR2_X1 maj_76_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_76_n16) );
  OR2_X1 maj_76_U6 ( .A1(maj_76_n20), .A2(maj_76_n19), .ZN(maj_76_n24) );
  NAND2_X1 maj_76_U5 ( .A1(maj_76_n24), .A2(maj_76_n23), .ZN(maj_76_n25) );
  NAND2_X1 maj_76_U4 ( .A1(maj_76_n20), .A2(maj_76_n19), .ZN(maj_76_n26) );
  NAND2_X1 maj_76_U3 ( .A1(maj_76_n26), .A2(maj_76_n25), .ZN(maj_76_port_o) );
  XOR2_X1 maj_76_U2 ( .A(maj_76_n22), .B(maj_76_n21), .Z(maj_76_n23) );
  NAND2_X1 maj_77_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_77_n18) );
  NAND2_X1 maj_77_U14 ( .A1(maj_77_n21), .A2(maj_77_n22), .ZN(maj_77_n17) );
  NAND2_X1 maj_77_U13 ( .A1(maj_77_n18), .A2(maj_77_n17), .ZN(maj_77_n19) );
  NAND2_X1 maj_77_U12 ( .A1(v_1_0[2]), .A2(maj_77_n16), .ZN(maj_77_n14) );
  NAND2_X1 maj_77_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_77_n15) );
  NAND2_X1 maj_77_U10 ( .A1(maj_77_n15), .A2(maj_77_n14), .ZN(maj_77_n20) );
  XOR2_X1 maj_77_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_77_n22) );
  XOR2_X1 maj_77_U8 ( .A(v_1_0[2]), .B(maj_77_n16), .Z(maj_77_n21) );
  XOR2_X1 maj_77_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_77_n16) );
  OR2_X1 maj_77_U6 ( .A1(maj_77_n20), .A2(maj_77_n19), .ZN(maj_77_n24) );
  NAND2_X1 maj_77_U5 ( .A1(maj_77_n24), .A2(maj_77_n23), .ZN(maj_77_n25) );
  NAND2_X1 maj_77_U4 ( .A1(maj_77_n20), .A2(maj_77_n19), .ZN(maj_77_n26) );
  NAND2_X1 maj_77_U3 ( .A1(maj_77_n26), .A2(maj_77_n25), .ZN(maj_77_port_o) );
  XOR2_X1 maj_77_U2 ( .A(maj_77_n22), .B(maj_77_n21), .Z(maj_77_n23) );
  NAND2_X1 maj_78_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_78_n18) );
  NAND2_X1 maj_78_U14 ( .A1(maj_78_n21), .A2(maj_78_n22), .ZN(maj_78_n17) );
  NAND2_X1 maj_78_U13 ( .A1(maj_78_n18), .A2(maj_78_n17), .ZN(maj_78_n19) );
  NAND2_X1 maj_78_U12 ( .A1(u_1_1[2]), .A2(maj_78_n16), .ZN(maj_78_n14) );
  NAND2_X1 maj_78_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_78_n15) );
  NAND2_X1 maj_78_U10 ( .A1(maj_78_n15), .A2(maj_78_n14), .ZN(maj_78_n20) );
  XOR2_X1 maj_78_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_78_n22) );
  XOR2_X1 maj_78_U8 ( .A(u_1_1[2]), .B(maj_78_n16), .Z(maj_78_n21) );
  XOR2_X1 maj_78_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_78_n16) );
  OR2_X1 maj_78_U6 ( .A1(maj_78_n20), .A2(maj_78_n19), .ZN(maj_78_n24) );
  NAND2_X1 maj_78_U5 ( .A1(maj_78_n24), .A2(maj_78_n23), .ZN(maj_78_n25) );
  NAND2_X1 maj_78_U4 ( .A1(maj_78_n20), .A2(maj_78_n19), .ZN(maj_78_n26) );
  NAND2_X1 maj_78_U3 ( .A1(maj_78_n26), .A2(maj_78_n25), .ZN(maj_78_port_o) );
  XOR2_X1 maj_78_U2 ( .A(maj_78_n22), .B(maj_78_n21), .Z(maj_78_n23) );
  NAND2_X1 maj_79_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_79_n18) );
  NAND2_X1 maj_79_U14 ( .A1(maj_79_n21), .A2(maj_79_n22), .ZN(maj_79_n17) );
  NAND2_X1 maj_79_U13 ( .A1(maj_79_n18), .A2(maj_79_n17), .ZN(maj_79_n19) );
  NAND2_X1 maj_79_U12 ( .A1(v_1_1[2]), .A2(maj_79_n16), .ZN(maj_79_n14) );
  NAND2_X1 maj_79_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_79_n15) );
  NAND2_X1 maj_79_U10 ( .A1(maj_79_n15), .A2(maj_79_n14), .ZN(maj_79_n20) );
  XOR2_X1 maj_79_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_79_n22) );
  XOR2_X1 maj_79_U8 ( .A(v_1_1[2]), .B(maj_79_n16), .Z(maj_79_n21) );
  XOR2_X1 maj_79_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_79_n16) );
  OR2_X1 maj_79_U6 ( .A1(maj_79_n20), .A2(maj_79_n19), .ZN(maj_79_n24) );
  NAND2_X1 maj_79_U5 ( .A1(maj_79_n24), .A2(maj_79_n23), .ZN(maj_79_n25) );
  NAND2_X1 maj_79_U4 ( .A1(maj_79_n20), .A2(maj_79_n19), .ZN(maj_79_n26) );
  NAND2_X1 maj_79_U3 ( .A1(maj_79_n26), .A2(maj_79_n25), .ZN(maj_79_port_o) );
  XOR2_X1 maj_79_U2 ( .A(maj_79_n22), .B(maj_79_n21), .Z(maj_79_n23) );
  NAND2_X1 maj_80_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_80_n18) );
  NAND2_X1 maj_80_U14 ( .A1(maj_80_n21), .A2(maj_80_n22), .ZN(maj_80_n17) );
  NAND2_X1 maj_80_U13 ( .A1(maj_80_n18), .A2(maj_80_n17), .ZN(maj_80_n19) );
  NAND2_X1 maj_80_U12 ( .A1(u_2_0[2]), .A2(maj_80_n16), .ZN(maj_80_n14) );
  NAND2_X1 maj_80_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_80_n15) );
  NAND2_X1 maj_80_U10 ( .A1(maj_80_n15), .A2(maj_80_n14), .ZN(maj_80_n20) );
  XOR2_X1 maj_80_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_80_n22) );
  XOR2_X1 maj_80_U8 ( .A(u_2_0[2]), .B(maj_80_n16), .Z(maj_80_n21) );
  XOR2_X1 maj_80_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_80_n16) );
  OR2_X1 maj_80_U6 ( .A1(maj_80_n20), .A2(maj_80_n19), .ZN(maj_80_n24) );
  NAND2_X1 maj_80_U5 ( .A1(maj_80_n24), .A2(maj_80_n23), .ZN(maj_80_n25) );
  NAND2_X1 maj_80_U4 ( .A1(maj_80_n20), .A2(maj_80_n19), .ZN(maj_80_n26) );
  NAND2_X1 maj_80_U3 ( .A1(maj_80_n26), .A2(maj_80_n25), .ZN(maj_80_port_o) );
  XOR2_X1 maj_80_U2 ( .A(maj_80_n22), .B(maj_80_n21), .Z(maj_80_n23) );
  NAND2_X1 maj_81_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_81_n18) );
  NAND2_X1 maj_81_U14 ( .A1(maj_81_n21), .A2(maj_81_n22), .ZN(maj_81_n17) );
  NAND2_X1 maj_81_U13 ( .A1(maj_81_n18), .A2(maj_81_n17), .ZN(maj_81_n19) );
  NAND2_X1 maj_81_U12 ( .A1(v_2_0[2]), .A2(maj_81_n16), .ZN(maj_81_n14) );
  NAND2_X1 maj_81_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_81_n15) );
  NAND2_X1 maj_81_U10 ( .A1(maj_81_n15), .A2(maj_81_n14), .ZN(maj_81_n20) );
  XOR2_X1 maj_81_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_81_n22) );
  XOR2_X1 maj_81_U8 ( .A(v_2_0[2]), .B(maj_81_n16), .Z(maj_81_n21) );
  XOR2_X1 maj_81_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_81_n16) );
  OR2_X1 maj_81_U6 ( .A1(maj_81_n20), .A2(maj_81_n19), .ZN(maj_81_n24) );
  NAND2_X1 maj_81_U5 ( .A1(maj_81_n24), .A2(maj_81_n23), .ZN(maj_81_n25) );
  NAND2_X1 maj_81_U4 ( .A1(maj_81_n20), .A2(maj_81_n19), .ZN(maj_81_n26) );
  NAND2_X1 maj_81_U3 ( .A1(maj_81_n26), .A2(maj_81_n25), .ZN(maj_81_port_o) );
  XOR2_X1 maj_81_U2 ( .A(maj_81_n22), .B(maj_81_n21), .Z(maj_81_n23) );
  NAND2_X1 maj_82_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_82_n18) );
  NAND2_X1 maj_82_U14 ( .A1(maj_82_n21), .A2(maj_82_n22), .ZN(maj_82_n17) );
  NAND2_X1 maj_82_U13 ( .A1(maj_82_n18), .A2(maj_82_n17), .ZN(maj_82_n19) );
  NAND2_X1 maj_82_U12 ( .A1(u_2_1[2]), .A2(maj_82_n16), .ZN(maj_82_n14) );
  NAND2_X1 maj_82_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_82_n15) );
  NAND2_X1 maj_82_U10 ( .A1(maj_82_n15), .A2(maj_82_n14), .ZN(maj_82_n20) );
  XOR2_X1 maj_82_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_82_n22) );
  XOR2_X1 maj_82_U8 ( .A(u_2_1[2]), .B(maj_82_n16), .Z(maj_82_n21) );
  XOR2_X1 maj_82_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_82_n16) );
  OR2_X1 maj_82_U6 ( .A1(maj_82_n20), .A2(maj_82_n19), .ZN(maj_82_n24) );
  NAND2_X1 maj_82_U5 ( .A1(maj_82_n24), .A2(maj_82_n23), .ZN(maj_82_n25) );
  NAND2_X1 maj_82_U4 ( .A1(maj_82_n20), .A2(maj_82_n19), .ZN(maj_82_n26) );
  NAND2_X1 maj_82_U3 ( .A1(maj_82_n26), .A2(maj_82_n25), .ZN(maj_82_port_o) );
  XOR2_X1 maj_82_U2 ( .A(maj_82_n22), .B(maj_82_n21), .Z(maj_82_n23) );
  NAND2_X1 maj_83_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_83_n18) );
  NAND2_X1 maj_83_U14 ( .A1(maj_83_n21), .A2(maj_83_n22), .ZN(maj_83_n17) );
  NAND2_X1 maj_83_U13 ( .A1(maj_83_n18), .A2(maj_83_n17), .ZN(maj_83_n19) );
  NAND2_X1 maj_83_U12 ( .A1(v_2_1[2]), .A2(maj_83_n16), .ZN(maj_83_n14) );
  NAND2_X1 maj_83_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_83_n15) );
  NAND2_X1 maj_83_U10 ( .A1(maj_83_n15), .A2(maj_83_n14), .ZN(maj_83_n20) );
  XOR2_X1 maj_83_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_83_n22) );
  XOR2_X1 maj_83_U8 ( .A(v_2_1[2]), .B(maj_83_n16), .Z(maj_83_n21) );
  XOR2_X1 maj_83_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_83_n16) );
  OR2_X1 maj_83_U6 ( .A1(maj_83_n20), .A2(maj_83_n19), .ZN(maj_83_n24) );
  NAND2_X1 maj_83_U5 ( .A1(maj_83_n24), .A2(maj_83_n23), .ZN(maj_83_n25) );
  NAND2_X1 maj_83_U4 ( .A1(maj_83_n20), .A2(maj_83_n19), .ZN(maj_83_n26) );
  NAND2_X1 maj_83_U3 ( .A1(maj_83_n26), .A2(maj_83_n25), .ZN(maj_83_port_o) );
  XOR2_X1 maj_83_U2 ( .A(maj_83_n22), .B(maj_83_n21), .Z(maj_83_n23) );
  NAND2_X1 maj_84_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_84_n18) );
  NAND2_X1 maj_84_U14 ( .A1(maj_84_n21), .A2(maj_84_n22), .ZN(maj_84_n17) );
  NAND2_X1 maj_84_U13 ( .A1(maj_84_n18), .A2(maj_84_n17), .ZN(maj_84_n19) );
  NAND2_X1 maj_84_U12 ( .A1(u_0_0[2]), .A2(maj_84_n16), .ZN(maj_84_n14) );
  NAND2_X1 maj_84_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_84_n15) );
  NAND2_X1 maj_84_U10 ( .A1(maj_84_n15), .A2(maj_84_n14), .ZN(maj_84_n20) );
  XOR2_X1 maj_84_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_84_n22) );
  XOR2_X1 maj_84_U8 ( .A(u_0_0[2]), .B(maj_84_n16), .Z(maj_84_n21) );
  XOR2_X1 maj_84_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_84_n16) );
  OR2_X1 maj_84_U6 ( .A1(maj_84_n20), .A2(maj_84_n19), .ZN(maj_84_n24) );
  NAND2_X1 maj_84_U5 ( .A1(maj_84_n24), .A2(maj_84_n23), .ZN(maj_84_n25) );
  NAND2_X1 maj_84_U4 ( .A1(maj_84_n20), .A2(maj_84_n19), .ZN(maj_84_n26) );
  NAND2_X1 maj_84_U3 ( .A1(maj_84_n26), .A2(maj_84_n25), .ZN(maj_84_port_o) );
  XOR2_X1 maj_84_U2 ( .A(maj_84_n22), .B(maj_84_n21), .Z(maj_84_n23) );
  NAND2_X1 maj_85_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_85_n18) );
  NAND2_X1 maj_85_U14 ( .A1(maj_85_n21), .A2(maj_85_n22), .ZN(maj_85_n17) );
  NAND2_X1 maj_85_U13 ( .A1(maj_85_n18), .A2(maj_85_n17), .ZN(maj_85_n19) );
  NAND2_X1 maj_85_U12 ( .A1(v_0_0[2]), .A2(maj_85_n16), .ZN(maj_85_n14) );
  NAND2_X1 maj_85_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_85_n15) );
  NAND2_X1 maj_85_U10 ( .A1(maj_85_n15), .A2(maj_85_n14), .ZN(maj_85_n20) );
  XOR2_X1 maj_85_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_85_n22) );
  XOR2_X1 maj_85_U8 ( .A(v_0_0[2]), .B(maj_85_n16), .Z(maj_85_n21) );
  XOR2_X1 maj_85_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_85_n16) );
  OR2_X1 maj_85_U6 ( .A1(maj_85_n20), .A2(maj_85_n19), .ZN(maj_85_n24) );
  NAND2_X1 maj_85_U5 ( .A1(maj_85_n24), .A2(maj_85_n23), .ZN(maj_85_n25) );
  NAND2_X1 maj_85_U4 ( .A1(maj_85_n20), .A2(maj_85_n19), .ZN(maj_85_n26) );
  NAND2_X1 maj_85_U3 ( .A1(maj_85_n26), .A2(maj_85_n25), .ZN(maj_85_port_o) );
  XOR2_X1 maj_85_U2 ( .A(maj_85_n22), .B(maj_85_n21), .Z(maj_85_n23) );
  NAND2_X1 maj_86_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_86_n18) );
  NAND2_X1 maj_86_U14 ( .A1(maj_86_n21), .A2(maj_86_n22), .ZN(maj_86_n17) );
  NAND2_X1 maj_86_U13 ( .A1(maj_86_n18), .A2(maj_86_n17), .ZN(maj_86_n19) );
  NAND2_X1 maj_86_U12 ( .A1(u_0_1[2]), .A2(maj_86_n16), .ZN(maj_86_n14) );
  NAND2_X1 maj_86_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_86_n15) );
  NAND2_X1 maj_86_U10 ( .A1(maj_86_n15), .A2(maj_86_n14), .ZN(maj_86_n20) );
  XOR2_X1 maj_86_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_86_n22) );
  XOR2_X1 maj_86_U8 ( .A(u_0_1[2]), .B(maj_86_n16), .Z(maj_86_n21) );
  XOR2_X1 maj_86_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_86_n16) );
  OR2_X1 maj_86_U6 ( .A1(maj_86_n20), .A2(maj_86_n19), .ZN(maj_86_n24) );
  NAND2_X1 maj_86_U5 ( .A1(maj_86_n24), .A2(maj_86_n23), .ZN(maj_86_n25) );
  NAND2_X1 maj_86_U4 ( .A1(maj_86_n20), .A2(maj_86_n19), .ZN(maj_86_n26) );
  NAND2_X1 maj_86_U3 ( .A1(maj_86_n26), .A2(maj_86_n25), .ZN(maj_86_port_o) );
  XOR2_X1 maj_86_U2 ( .A(maj_86_n22), .B(maj_86_n21), .Z(maj_86_n23) );
  NAND2_X1 maj_87_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_87_n18) );
  NAND2_X1 maj_87_U14 ( .A1(maj_87_n21), .A2(maj_87_n22), .ZN(maj_87_n17) );
  NAND2_X1 maj_87_U13 ( .A1(maj_87_n18), .A2(maj_87_n17), .ZN(maj_87_n19) );
  NAND2_X1 maj_87_U12 ( .A1(v_0_1[2]), .A2(maj_87_n16), .ZN(maj_87_n14) );
  NAND2_X1 maj_87_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_87_n15) );
  NAND2_X1 maj_87_U10 ( .A1(maj_87_n15), .A2(maj_87_n14), .ZN(maj_87_n20) );
  XOR2_X1 maj_87_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_87_n22) );
  XOR2_X1 maj_87_U8 ( .A(v_0_1[2]), .B(maj_87_n16), .Z(maj_87_n21) );
  XOR2_X1 maj_87_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_87_n16) );
  OR2_X1 maj_87_U6 ( .A1(maj_87_n20), .A2(maj_87_n19), .ZN(maj_87_n24) );
  NAND2_X1 maj_87_U5 ( .A1(maj_87_n24), .A2(maj_87_n23), .ZN(maj_87_n25) );
  NAND2_X1 maj_87_U4 ( .A1(maj_87_n20), .A2(maj_87_n19), .ZN(maj_87_n26) );
  NAND2_X1 maj_87_U3 ( .A1(maj_87_n26), .A2(maj_87_n25), .ZN(maj_87_port_o) );
  XOR2_X1 maj_87_U2 ( .A(maj_87_n22), .B(maj_87_n21), .Z(maj_87_n23) );
  NAND2_X1 maj_88_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_88_n18) );
  NAND2_X1 maj_88_U14 ( .A1(maj_88_n21), .A2(maj_88_n22), .ZN(maj_88_n17) );
  NAND2_X1 maj_88_U13 ( .A1(maj_88_n18), .A2(maj_88_n17), .ZN(maj_88_n19) );
  NAND2_X1 maj_88_U12 ( .A1(u_1_0[2]), .A2(maj_88_n16), .ZN(maj_88_n14) );
  NAND2_X1 maj_88_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_88_n15) );
  NAND2_X1 maj_88_U10 ( .A1(maj_88_n15), .A2(maj_88_n14), .ZN(maj_88_n20) );
  XOR2_X1 maj_88_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_88_n22) );
  XOR2_X1 maj_88_U8 ( .A(u_1_0[2]), .B(maj_88_n16), .Z(maj_88_n21) );
  XOR2_X1 maj_88_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_88_n16) );
  OR2_X1 maj_88_U6 ( .A1(maj_88_n20), .A2(maj_88_n19), .ZN(maj_88_n24) );
  NAND2_X1 maj_88_U5 ( .A1(maj_88_n24), .A2(maj_88_n23), .ZN(maj_88_n25) );
  NAND2_X1 maj_88_U4 ( .A1(maj_88_n20), .A2(maj_88_n19), .ZN(maj_88_n26) );
  NAND2_X1 maj_88_U3 ( .A1(maj_88_n26), .A2(maj_88_n25), .ZN(maj_88_port_o) );
  XOR2_X1 maj_88_U2 ( .A(maj_88_n22), .B(maj_88_n21), .Z(maj_88_n23) );
  NAND2_X1 maj_89_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_89_n18) );
  NAND2_X1 maj_89_U14 ( .A1(maj_89_n21), .A2(maj_89_n22), .ZN(maj_89_n17) );
  NAND2_X1 maj_89_U13 ( .A1(maj_89_n18), .A2(maj_89_n17), .ZN(maj_89_n19) );
  NAND2_X1 maj_89_U12 ( .A1(v_1_0[2]), .A2(maj_89_n16), .ZN(maj_89_n14) );
  NAND2_X1 maj_89_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_89_n15) );
  NAND2_X1 maj_89_U10 ( .A1(maj_89_n15), .A2(maj_89_n14), .ZN(maj_89_n20) );
  XOR2_X1 maj_89_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_89_n22) );
  XOR2_X1 maj_89_U8 ( .A(v_1_0[2]), .B(maj_89_n16), .Z(maj_89_n21) );
  XOR2_X1 maj_89_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_89_n16) );
  OR2_X1 maj_89_U6 ( .A1(maj_89_n20), .A2(maj_89_n19), .ZN(maj_89_n24) );
  NAND2_X1 maj_89_U5 ( .A1(maj_89_n24), .A2(maj_89_n23), .ZN(maj_89_n25) );
  NAND2_X1 maj_89_U4 ( .A1(maj_89_n20), .A2(maj_89_n19), .ZN(maj_89_n26) );
  NAND2_X1 maj_89_U3 ( .A1(maj_89_n26), .A2(maj_89_n25), .ZN(maj_89_port_o) );
  XOR2_X1 maj_89_U2 ( .A(maj_89_n22), .B(maj_89_n21), .Z(maj_89_n23) );
  NAND2_X1 maj_90_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_90_n18) );
  NAND2_X1 maj_90_U14 ( .A1(maj_90_n21), .A2(maj_90_n22), .ZN(maj_90_n17) );
  NAND2_X1 maj_90_U13 ( .A1(maj_90_n18), .A2(maj_90_n17), .ZN(maj_90_n19) );
  NAND2_X1 maj_90_U12 ( .A1(u_1_1[2]), .A2(maj_90_n16), .ZN(maj_90_n14) );
  NAND2_X1 maj_90_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_90_n15) );
  NAND2_X1 maj_90_U10 ( .A1(maj_90_n15), .A2(maj_90_n14), .ZN(maj_90_n20) );
  XOR2_X1 maj_90_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_90_n22) );
  XOR2_X1 maj_90_U8 ( .A(u_1_1[2]), .B(maj_90_n16), .Z(maj_90_n21) );
  XOR2_X1 maj_90_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_90_n16) );
  OR2_X1 maj_90_U6 ( .A1(maj_90_n20), .A2(maj_90_n19), .ZN(maj_90_n24) );
  NAND2_X1 maj_90_U5 ( .A1(maj_90_n24), .A2(maj_90_n23), .ZN(maj_90_n25) );
  NAND2_X1 maj_90_U4 ( .A1(maj_90_n20), .A2(maj_90_n19), .ZN(maj_90_n26) );
  NAND2_X1 maj_90_U3 ( .A1(maj_90_n26), .A2(maj_90_n25), .ZN(maj_90_port_o) );
  XOR2_X1 maj_90_U2 ( .A(maj_90_n22), .B(maj_90_n21), .Z(maj_90_n23) );
  NAND2_X1 maj_91_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_91_n18) );
  NAND2_X1 maj_91_U14 ( .A1(maj_91_n21), .A2(maj_91_n22), .ZN(maj_91_n17) );
  NAND2_X1 maj_91_U13 ( .A1(maj_91_n18), .A2(maj_91_n17), .ZN(maj_91_n19) );
  NAND2_X1 maj_91_U12 ( .A1(v_1_1[2]), .A2(maj_91_n16), .ZN(maj_91_n14) );
  NAND2_X1 maj_91_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_91_n15) );
  NAND2_X1 maj_91_U10 ( .A1(maj_91_n15), .A2(maj_91_n14), .ZN(maj_91_n20) );
  XOR2_X1 maj_91_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_91_n22) );
  XOR2_X1 maj_91_U8 ( .A(v_1_1[2]), .B(maj_91_n16), .Z(maj_91_n21) );
  XOR2_X1 maj_91_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_91_n16) );
  OR2_X1 maj_91_U6 ( .A1(maj_91_n20), .A2(maj_91_n19), .ZN(maj_91_n24) );
  NAND2_X1 maj_91_U5 ( .A1(maj_91_n24), .A2(maj_91_n23), .ZN(maj_91_n25) );
  NAND2_X1 maj_91_U4 ( .A1(maj_91_n20), .A2(maj_91_n19), .ZN(maj_91_n26) );
  NAND2_X1 maj_91_U3 ( .A1(maj_91_n26), .A2(maj_91_n25), .ZN(maj_91_port_o) );
  XOR2_X1 maj_91_U2 ( .A(maj_91_n22), .B(maj_91_n21), .Z(maj_91_n23) );
  NAND2_X1 maj_92_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_92_n18) );
  NAND2_X1 maj_92_U14 ( .A1(maj_92_n21), .A2(maj_92_n22), .ZN(maj_92_n17) );
  NAND2_X1 maj_92_U13 ( .A1(maj_92_n18), .A2(maj_92_n17), .ZN(maj_92_n19) );
  NAND2_X1 maj_92_U12 ( .A1(u_2_0[2]), .A2(maj_92_n16), .ZN(maj_92_n14) );
  NAND2_X1 maj_92_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_92_n15) );
  NAND2_X1 maj_92_U10 ( .A1(maj_92_n15), .A2(maj_92_n14), .ZN(maj_92_n20) );
  XOR2_X1 maj_92_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_92_n22) );
  XOR2_X1 maj_92_U8 ( .A(u_2_0[2]), .B(maj_92_n16), .Z(maj_92_n21) );
  XOR2_X1 maj_92_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_92_n16) );
  OR2_X1 maj_92_U6 ( .A1(maj_92_n20), .A2(maj_92_n19), .ZN(maj_92_n24) );
  NAND2_X1 maj_92_U5 ( .A1(maj_92_n24), .A2(maj_92_n23), .ZN(maj_92_n25) );
  NAND2_X1 maj_92_U4 ( .A1(maj_92_n20), .A2(maj_92_n19), .ZN(maj_92_n26) );
  NAND2_X1 maj_92_U3 ( .A1(maj_92_n26), .A2(maj_92_n25), .ZN(maj_92_port_o) );
  XOR2_X1 maj_92_U2 ( .A(maj_92_n22), .B(maj_92_n21), .Z(maj_92_n23) );
  NAND2_X1 maj_93_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_93_n18) );
  NAND2_X1 maj_93_U14 ( .A1(maj_93_n21), .A2(maj_93_n22), .ZN(maj_93_n17) );
  NAND2_X1 maj_93_U13 ( .A1(maj_93_n18), .A2(maj_93_n17), .ZN(maj_93_n19) );
  NAND2_X1 maj_93_U12 ( .A1(v_2_0[2]), .A2(maj_93_n16), .ZN(maj_93_n14) );
  NAND2_X1 maj_93_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_93_n15) );
  NAND2_X1 maj_93_U10 ( .A1(maj_93_n15), .A2(maj_93_n14), .ZN(maj_93_n20) );
  XOR2_X1 maj_93_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_93_n22) );
  XOR2_X1 maj_93_U8 ( .A(v_2_0[2]), .B(maj_93_n16), .Z(maj_93_n21) );
  XOR2_X1 maj_93_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_93_n16) );
  OR2_X1 maj_93_U6 ( .A1(maj_93_n20), .A2(maj_93_n19), .ZN(maj_93_n24) );
  NAND2_X1 maj_93_U5 ( .A1(maj_93_n24), .A2(maj_93_n23), .ZN(maj_93_n25) );
  NAND2_X1 maj_93_U4 ( .A1(maj_93_n20), .A2(maj_93_n19), .ZN(maj_93_n26) );
  NAND2_X1 maj_93_U3 ( .A1(maj_93_n26), .A2(maj_93_n25), .ZN(maj_93_port_o) );
  XOR2_X1 maj_93_U2 ( .A(maj_93_n22), .B(maj_93_n21), .Z(maj_93_n23) );
  NAND2_X1 maj_94_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_94_n18) );
  NAND2_X1 maj_94_U14 ( .A1(maj_94_n21), .A2(maj_94_n22), .ZN(maj_94_n17) );
  NAND2_X1 maj_94_U13 ( .A1(maj_94_n18), .A2(maj_94_n17), .ZN(maj_94_n19) );
  NAND2_X1 maj_94_U12 ( .A1(u_2_1[2]), .A2(maj_94_n16), .ZN(maj_94_n14) );
  NAND2_X1 maj_94_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_94_n15) );
  NAND2_X1 maj_94_U10 ( .A1(maj_94_n15), .A2(maj_94_n14), .ZN(maj_94_n20) );
  XOR2_X1 maj_94_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_94_n22) );
  XOR2_X1 maj_94_U8 ( .A(u_2_1[2]), .B(maj_94_n16), .Z(maj_94_n21) );
  XOR2_X1 maj_94_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_94_n16) );
  OR2_X1 maj_94_U6 ( .A1(maj_94_n20), .A2(maj_94_n19), .ZN(maj_94_n24) );
  NAND2_X1 maj_94_U5 ( .A1(maj_94_n24), .A2(maj_94_n23), .ZN(maj_94_n25) );
  NAND2_X1 maj_94_U4 ( .A1(maj_94_n20), .A2(maj_94_n19), .ZN(maj_94_n26) );
  NAND2_X1 maj_94_U3 ( .A1(maj_94_n26), .A2(maj_94_n25), .ZN(maj_94_port_o) );
  XOR2_X1 maj_94_U2 ( .A(maj_94_n22), .B(maj_94_n21), .Z(maj_94_n23) );
  NAND2_X1 maj_95_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_95_n18) );
  NAND2_X1 maj_95_U14 ( .A1(maj_95_n21), .A2(maj_95_n22), .ZN(maj_95_n17) );
  NAND2_X1 maj_95_U13 ( .A1(maj_95_n18), .A2(maj_95_n17), .ZN(maj_95_n19) );
  NAND2_X1 maj_95_U12 ( .A1(v_2_1[2]), .A2(maj_95_n16), .ZN(maj_95_n14) );
  NAND2_X1 maj_95_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_95_n15) );
  NAND2_X1 maj_95_U10 ( .A1(maj_95_n15), .A2(maj_95_n14), .ZN(maj_95_n20) );
  XOR2_X1 maj_95_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_95_n22) );
  XOR2_X1 maj_95_U8 ( .A(v_2_1[2]), .B(maj_95_n16), .Z(maj_95_n21) );
  XOR2_X1 maj_95_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_95_n16) );
  OR2_X1 maj_95_U6 ( .A1(maj_95_n20), .A2(maj_95_n19), .ZN(maj_95_n24) );
  NAND2_X1 maj_95_U5 ( .A1(maj_95_n24), .A2(maj_95_n23), .ZN(maj_95_n25) );
  NAND2_X1 maj_95_U4 ( .A1(maj_95_n20), .A2(maj_95_n19), .ZN(maj_95_n26) );
  NAND2_X1 maj_95_U3 ( .A1(maj_95_n26), .A2(maj_95_n25), .ZN(maj_95_port_o) );
  XOR2_X1 maj_95_U2 ( .A(maj_95_n22), .B(maj_95_n21), .Z(maj_95_n23) );
  NAND2_X1 maj_96_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_96_n18) );
  NAND2_X1 maj_96_U14 ( .A1(maj_96_n21), .A2(maj_96_n22), .ZN(maj_96_n17) );
  NAND2_X1 maj_96_U13 ( .A1(maj_96_n18), .A2(maj_96_n17), .ZN(maj_96_n19) );
  NAND2_X1 maj_96_U12 ( .A1(u_0_0[2]), .A2(maj_96_n16), .ZN(maj_96_n14) );
  NAND2_X1 maj_96_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_96_n15) );
  NAND2_X1 maj_96_U10 ( .A1(maj_96_n15), .A2(maj_96_n14), .ZN(maj_96_n20) );
  XOR2_X1 maj_96_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_96_n22) );
  XOR2_X1 maj_96_U8 ( .A(u_0_0[2]), .B(maj_96_n16), .Z(maj_96_n21) );
  XOR2_X1 maj_96_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_96_n16) );
  OR2_X1 maj_96_U6 ( .A1(maj_96_n20), .A2(maj_96_n19), .ZN(maj_96_n24) );
  NAND2_X1 maj_96_U5 ( .A1(maj_96_n24), .A2(maj_96_n23), .ZN(maj_96_n25) );
  NAND2_X1 maj_96_U4 ( .A1(maj_96_n20), .A2(maj_96_n19), .ZN(maj_96_n26) );
  NAND2_X1 maj_96_U3 ( .A1(maj_96_n26), .A2(maj_96_n25), .ZN(maj_96_port_o) );
  XOR2_X1 maj_96_U2 ( .A(maj_96_n22), .B(maj_96_n21), .Z(maj_96_n23) );
  NAND2_X1 maj_97_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_97_n18) );
  NAND2_X1 maj_97_U14 ( .A1(maj_97_n21), .A2(maj_97_n22), .ZN(maj_97_n17) );
  NAND2_X1 maj_97_U13 ( .A1(maj_97_n18), .A2(maj_97_n17), .ZN(maj_97_n19) );
  NAND2_X1 maj_97_U12 ( .A1(v_0_0[2]), .A2(maj_97_n16), .ZN(maj_97_n14) );
  NAND2_X1 maj_97_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_97_n15) );
  NAND2_X1 maj_97_U10 ( .A1(maj_97_n15), .A2(maj_97_n14), .ZN(maj_97_n20) );
  XOR2_X1 maj_97_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_97_n22) );
  XOR2_X1 maj_97_U8 ( .A(v_0_0[2]), .B(maj_97_n16), .Z(maj_97_n21) );
  XOR2_X1 maj_97_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_97_n16) );
  OR2_X1 maj_97_U6 ( .A1(maj_97_n20), .A2(maj_97_n19), .ZN(maj_97_n24) );
  NAND2_X1 maj_97_U5 ( .A1(maj_97_n24), .A2(maj_97_n23), .ZN(maj_97_n25) );
  NAND2_X1 maj_97_U4 ( .A1(maj_97_n20), .A2(maj_97_n19), .ZN(maj_97_n26) );
  NAND2_X1 maj_97_U3 ( .A1(maj_97_n26), .A2(maj_97_n25), .ZN(maj_97_port_o) );
  XOR2_X1 maj_97_U2 ( .A(maj_97_n22), .B(maj_97_n21), .Z(maj_97_n23) );
  NAND2_X1 maj_98_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_98_n18) );
  NAND2_X1 maj_98_U14 ( .A1(maj_98_n21), .A2(maj_98_n22), .ZN(maj_98_n17) );
  NAND2_X1 maj_98_U13 ( .A1(maj_98_n18), .A2(maj_98_n17), .ZN(maj_98_n19) );
  NAND2_X1 maj_98_U12 ( .A1(u_0_1[2]), .A2(maj_98_n16), .ZN(maj_98_n14) );
  NAND2_X1 maj_98_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_98_n15) );
  NAND2_X1 maj_98_U10 ( .A1(maj_98_n15), .A2(maj_98_n14), .ZN(maj_98_n20) );
  XOR2_X1 maj_98_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_98_n22) );
  XOR2_X1 maj_98_U8 ( .A(u_0_1[2]), .B(maj_98_n16), .Z(maj_98_n21) );
  XOR2_X1 maj_98_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_98_n16) );
  OR2_X1 maj_98_U6 ( .A1(maj_98_n20), .A2(maj_98_n19), .ZN(maj_98_n24) );
  NAND2_X1 maj_98_U5 ( .A1(maj_98_n24), .A2(maj_98_n23), .ZN(maj_98_n25) );
  NAND2_X1 maj_98_U4 ( .A1(maj_98_n20), .A2(maj_98_n19), .ZN(maj_98_n26) );
  NAND2_X1 maj_98_U3 ( .A1(maj_98_n26), .A2(maj_98_n25), .ZN(maj_98_port_o) );
  XOR2_X1 maj_98_U2 ( .A(maj_98_n22), .B(maj_98_n21), .Z(maj_98_n23) );
  NAND2_X1 maj_99_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_99_n18) );
  NAND2_X1 maj_99_U14 ( .A1(maj_99_n21), .A2(maj_99_n22), .ZN(maj_99_n17) );
  NAND2_X1 maj_99_U13 ( .A1(maj_99_n18), .A2(maj_99_n17), .ZN(maj_99_n19) );
  NAND2_X1 maj_99_U12 ( .A1(v_0_1[2]), .A2(maj_99_n16), .ZN(maj_99_n14) );
  NAND2_X1 maj_99_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_99_n15) );
  NAND2_X1 maj_99_U10 ( .A1(maj_99_n15), .A2(maj_99_n14), .ZN(maj_99_n20) );
  XOR2_X1 maj_99_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_99_n22) );
  XOR2_X1 maj_99_U8 ( .A(v_0_1[2]), .B(maj_99_n16), .Z(maj_99_n21) );
  XOR2_X1 maj_99_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_99_n16) );
  OR2_X1 maj_99_U6 ( .A1(maj_99_n20), .A2(maj_99_n19), .ZN(maj_99_n24) );
  NAND2_X1 maj_99_U5 ( .A1(maj_99_n24), .A2(maj_99_n23), .ZN(maj_99_n25) );
  NAND2_X1 maj_99_U4 ( .A1(maj_99_n20), .A2(maj_99_n19), .ZN(maj_99_n26) );
  NAND2_X1 maj_99_U3 ( .A1(maj_99_n26), .A2(maj_99_n25), .ZN(maj_99_port_o) );
  XOR2_X1 maj_99_U2 ( .A(maj_99_n22), .B(maj_99_n21), .Z(maj_99_n23) );
  NAND2_X1 maj_100_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_100_n18) );
  NAND2_X1 maj_100_U14 ( .A1(maj_100_n21), .A2(maj_100_n22), .ZN(maj_100_n17)
         );
  NAND2_X1 maj_100_U13 ( .A1(maj_100_n18), .A2(maj_100_n17), .ZN(maj_100_n19)
         );
  NAND2_X1 maj_100_U12 ( .A1(u_1_0[2]), .A2(maj_100_n16), .ZN(maj_100_n14) );
  NAND2_X1 maj_100_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_100_n15) );
  NAND2_X1 maj_100_U10 ( .A1(maj_100_n15), .A2(maj_100_n14), .ZN(maj_100_n20)
         );
  XOR2_X1 maj_100_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_100_n22) );
  XOR2_X1 maj_100_U8 ( .A(u_1_0[2]), .B(maj_100_n16), .Z(maj_100_n21) );
  XOR2_X1 maj_100_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_100_n16) );
  OR2_X1 maj_100_U6 ( .A1(maj_100_n20), .A2(maj_100_n19), .ZN(maj_100_n24) );
  NAND2_X1 maj_100_U5 ( .A1(maj_100_n24), .A2(maj_100_n23), .ZN(maj_100_n25)
         );
  NAND2_X1 maj_100_U4 ( .A1(maj_100_n20), .A2(maj_100_n19), .ZN(maj_100_n26)
         );
  NAND2_X1 maj_100_U3 ( .A1(maj_100_n26), .A2(maj_100_n25), .ZN(maj_100_port_o) );
  XOR2_X1 maj_100_U2 ( .A(maj_100_n22), .B(maj_100_n21), .Z(maj_100_n23) );
  NAND2_X1 maj_101_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_101_n18) );
  NAND2_X1 maj_101_U14 ( .A1(maj_101_n21), .A2(maj_101_n22), .ZN(maj_101_n17)
         );
  NAND2_X1 maj_101_U13 ( .A1(maj_101_n18), .A2(maj_101_n17), .ZN(maj_101_n19)
         );
  NAND2_X1 maj_101_U12 ( .A1(v_1_0[2]), .A2(maj_101_n16), .ZN(maj_101_n14) );
  NAND2_X1 maj_101_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_101_n15) );
  NAND2_X1 maj_101_U10 ( .A1(maj_101_n15), .A2(maj_101_n14), .ZN(maj_101_n20)
         );
  XOR2_X1 maj_101_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_101_n22) );
  XOR2_X1 maj_101_U8 ( .A(v_1_0[2]), .B(maj_101_n16), .Z(maj_101_n21) );
  XOR2_X1 maj_101_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_101_n16) );
  OR2_X1 maj_101_U6 ( .A1(maj_101_n20), .A2(maj_101_n19), .ZN(maj_101_n24) );
  NAND2_X1 maj_101_U5 ( .A1(maj_101_n24), .A2(maj_101_n23), .ZN(maj_101_n25)
         );
  NAND2_X1 maj_101_U4 ( .A1(maj_101_n20), .A2(maj_101_n19), .ZN(maj_101_n26)
         );
  NAND2_X1 maj_101_U3 ( .A1(maj_101_n26), .A2(maj_101_n25), .ZN(maj_101_port_o) );
  XOR2_X1 maj_101_U2 ( .A(maj_101_n22), .B(maj_101_n21), .Z(maj_101_n23) );
  NAND2_X1 maj_102_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_102_n18) );
  NAND2_X1 maj_102_U14 ( .A1(maj_102_n21), .A2(maj_102_n22), .ZN(maj_102_n17)
         );
  NAND2_X1 maj_102_U13 ( .A1(maj_102_n18), .A2(maj_102_n17), .ZN(maj_102_n19)
         );
  NAND2_X1 maj_102_U12 ( .A1(u_1_1[2]), .A2(maj_102_n16), .ZN(maj_102_n14) );
  NAND2_X1 maj_102_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_102_n15) );
  NAND2_X1 maj_102_U10 ( .A1(maj_102_n15), .A2(maj_102_n14), .ZN(maj_102_n20)
         );
  XOR2_X1 maj_102_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_102_n22) );
  XOR2_X1 maj_102_U8 ( .A(u_1_1[2]), .B(maj_102_n16), .Z(maj_102_n21) );
  XOR2_X1 maj_102_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_102_n16) );
  OR2_X1 maj_102_U6 ( .A1(maj_102_n20), .A2(maj_102_n19), .ZN(maj_102_n24) );
  NAND2_X1 maj_102_U5 ( .A1(maj_102_n24), .A2(maj_102_n23), .ZN(maj_102_n25)
         );
  NAND2_X1 maj_102_U4 ( .A1(maj_102_n20), .A2(maj_102_n19), .ZN(maj_102_n26)
         );
  NAND2_X1 maj_102_U3 ( .A1(maj_102_n26), .A2(maj_102_n25), .ZN(maj_102_port_o) );
  XOR2_X1 maj_102_U2 ( .A(maj_102_n22), .B(maj_102_n21), .Z(maj_102_n23) );
  NAND2_X1 maj_103_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_103_n18) );
  NAND2_X1 maj_103_U14 ( .A1(maj_103_n21), .A2(maj_103_n22), .ZN(maj_103_n17)
         );
  NAND2_X1 maj_103_U13 ( .A1(maj_103_n18), .A2(maj_103_n17), .ZN(maj_103_n19)
         );
  NAND2_X1 maj_103_U12 ( .A1(v_1_1[2]), .A2(maj_103_n16), .ZN(maj_103_n14) );
  NAND2_X1 maj_103_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_103_n15) );
  NAND2_X1 maj_103_U10 ( .A1(maj_103_n15), .A2(maj_103_n14), .ZN(maj_103_n20)
         );
  XOR2_X1 maj_103_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_103_n22) );
  XOR2_X1 maj_103_U8 ( .A(v_1_1[2]), .B(maj_103_n16), .Z(maj_103_n21) );
  XOR2_X1 maj_103_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_103_n16) );
  OR2_X1 maj_103_U6 ( .A1(maj_103_n20), .A2(maj_103_n19), .ZN(maj_103_n24) );
  NAND2_X1 maj_103_U5 ( .A1(maj_103_n24), .A2(maj_103_n23), .ZN(maj_103_n25)
         );
  NAND2_X1 maj_103_U4 ( .A1(maj_103_n20), .A2(maj_103_n19), .ZN(maj_103_n26)
         );
  NAND2_X1 maj_103_U3 ( .A1(maj_103_n26), .A2(maj_103_n25), .ZN(maj_103_port_o) );
  XOR2_X1 maj_103_U2 ( .A(maj_103_n22), .B(maj_103_n21), .Z(maj_103_n23) );
  NAND2_X1 maj_104_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_104_n18) );
  NAND2_X1 maj_104_U14 ( .A1(maj_104_n21), .A2(maj_104_n22), .ZN(maj_104_n17)
         );
  NAND2_X1 maj_104_U13 ( .A1(maj_104_n18), .A2(maj_104_n17), .ZN(maj_104_n19)
         );
  NAND2_X1 maj_104_U12 ( .A1(u_2_0[2]), .A2(maj_104_n16), .ZN(maj_104_n14) );
  NAND2_X1 maj_104_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_104_n15) );
  NAND2_X1 maj_104_U10 ( .A1(maj_104_n15), .A2(maj_104_n14), .ZN(maj_104_n20)
         );
  XOR2_X1 maj_104_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_104_n22) );
  XOR2_X1 maj_104_U8 ( .A(u_2_0[2]), .B(maj_104_n16), .Z(maj_104_n21) );
  XOR2_X1 maj_104_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_104_n16) );
  OR2_X1 maj_104_U6 ( .A1(maj_104_n20), .A2(maj_104_n19), .ZN(maj_104_n24) );
  NAND2_X1 maj_104_U5 ( .A1(maj_104_n24), .A2(maj_104_n23), .ZN(maj_104_n25)
         );
  NAND2_X1 maj_104_U4 ( .A1(maj_104_n20), .A2(maj_104_n19), .ZN(maj_104_n26)
         );
  NAND2_X1 maj_104_U3 ( .A1(maj_104_n26), .A2(maj_104_n25), .ZN(maj_104_port_o) );
  XOR2_X1 maj_104_U2 ( .A(maj_104_n22), .B(maj_104_n21), .Z(maj_104_n23) );
  NAND2_X1 maj_105_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_105_n18) );
  NAND2_X1 maj_105_U14 ( .A1(maj_105_n21), .A2(maj_105_n22), .ZN(maj_105_n17)
         );
  NAND2_X1 maj_105_U13 ( .A1(maj_105_n18), .A2(maj_105_n17), .ZN(maj_105_n19)
         );
  NAND2_X1 maj_105_U12 ( .A1(v_2_0[2]), .A2(maj_105_n16), .ZN(maj_105_n14) );
  NAND2_X1 maj_105_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_105_n15) );
  NAND2_X1 maj_105_U10 ( .A1(maj_105_n15), .A2(maj_105_n14), .ZN(maj_105_n20)
         );
  XOR2_X1 maj_105_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_105_n22) );
  XOR2_X1 maj_105_U8 ( .A(v_2_0[2]), .B(maj_105_n16), .Z(maj_105_n21) );
  XOR2_X1 maj_105_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_105_n16) );
  OR2_X1 maj_105_U6 ( .A1(maj_105_n20), .A2(maj_105_n19), .ZN(maj_105_n24) );
  NAND2_X1 maj_105_U5 ( .A1(maj_105_n24), .A2(maj_105_n23), .ZN(maj_105_n25)
         );
  NAND2_X1 maj_105_U4 ( .A1(maj_105_n20), .A2(maj_105_n19), .ZN(maj_105_n26)
         );
  NAND2_X1 maj_105_U3 ( .A1(maj_105_n26), .A2(maj_105_n25), .ZN(maj_105_port_o) );
  XOR2_X1 maj_105_U2 ( .A(maj_105_n22), .B(maj_105_n21), .Z(maj_105_n23) );
  NAND2_X1 maj_106_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_106_n18) );
  NAND2_X1 maj_106_U14 ( .A1(maj_106_n21), .A2(maj_106_n22), .ZN(maj_106_n17)
         );
  NAND2_X1 maj_106_U13 ( .A1(maj_106_n18), .A2(maj_106_n17), .ZN(maj_106_n19)
         );
  NAND2_X1 maj_106_U12 ( .A1(u_2_1[2]), .A2(maj_106_n16), .ZN(maj_106_n14) );
  NAND2_X1 maj_106_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_106_n15) );
  NAND2_X1 maj_106_U10 ( .A1(maj_106_n15), .A2(maj_106_n14), .ZN(maj_106_n20)
         );
  XOR2_X1 maj_106_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_106_n22) );
  XOR2_X1 maj_106_U8 ( .A(u_2_1[2]), .B(maj_106_n16), .Z(maj_106_n21) );
  XOR2_X1 maj_106_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_106_n16) );
  OR2_X1 maj_106_U6 ( .A1(maj_106_n20), .A2(maj_106_n19), .ZN(maj_106_n24) );
  NAND2_X1 maj_106_U5 ( .A1(maj_106_n24), .A2(maj_106_n23), .ZN(maj_106_n25)
         );
  NAND2_X1 maj_106_U4 ( .A1(maj_106_n20), .A2(maj_106_n19), .ZN(maj_106_n26)
         );
  NAND2_X1 maj_106_U3 ( .A1(maj_106_n26), .A2(maj_106_n25), .ZN(maj_106_port_o) );
  XOR2_X1 maj_106_U2 ( .A(maj_106_n22), .B(maj_106_n21), .Z(maj_106_n23) );
  NAND2_X1 maj_107_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_107_n18) );
  NAND2_X1 maj_107_U14 ( .A1(maj_107_n21), .A2(maj_107_n22), .ZN(maj_107_n17)
         );
  NAND2_X1 maj_107_U13 ( .A1(maj_107_n18), .A2(maj_107_n17), .ZN(maj_107_n19)
         );
  NAND2_X1 maj_107_U12 ( .A1(v_2_1[2]), .A2(maj_107_n16), .ZN(maj_107_n14) );
  NAND2_X1 maj_107_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_107_n15) );
  NAND2_X1 maj_107_U10 ( .A1(maj_107_n15), .A2(maj_107_n14), .ZN(maj_107_n20)
         );
  XOR2_X1 maj_107_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_107_n22) );
  XOR2_X1 maj_107_U8 ( .A(v_2_1[2]), .B(maj_107_n16), .Z(maj_107_n21) );
  XOR2_X1 maj_107_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_107_n16) );
  OR2_X1 maj_107_U6 ( .A1(maj_107_n20), .A2(maj_107_n19), .ZN(maj_107_n24) );
  NAND2_X1 maj_107_U5 ( .A1(maj_107_n24), .A2(maj_107_n23), .ZN(maj_107_n25)
         );
  NAND2_X1 maj_107_U4 ( .A1(maj_107_n20), .A2(maj_107_n19), .ZN(maj_107_n26)
         );
  NAND2_X1 maj_107_U3 ( .A1(maj_107_n26), .A2(maj_107_n25), .ZN(maj_107_port_o) );
  XOR2_X1 maj_107_U2 ( .A(maj_107_n22), .B(maj_107_n21), .Z(maj_107_n23) );
  NAND2_X1 maj_108_U15 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_108_n18) );
  NAND2_X1 maj_108_U14 ( .A1(maj_108_n21), .A2(maj_108_n22), .ZN(maj_108_n17)
         );
  NAND2_X1 maj_108_U13 ( .A1(maj_108_n18), .A2(maj_108_n17), .ZN(maj_108_n19)
         );
  NAND2_X1 maj_108_U12 ( .A1(u_0_0[2]), .A2(maj_108_n16), .ZN(maj_108_n14) );
  NAND2_X1 maj_108_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_108_n15) );
  NAND2_X1 maj_108_U10 ( .A1(maj_108_n15), .A2(maj_108_n14), .ZN(maj_108_n20)
         );
  XOR2_X1 maj_108_U9 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_108_n22) );
  XOR2_X1 maj_108_U8 ( .A(u_0_0[2]), .B(maj_108_n16), .Z(maj_108_n21) );
  XOR2_X1 maj_108_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_108_n16) );
  OR2_X1 maj_108_U6 ( .A1(maj_108_n20), .A2(maj_108_n19), .ZN(maj_108_n24) );
  NAND2_X1 maj_108_U5 ( .A1(maj_108_n24), .A2(maj_108_n23), .ZN(maj_108_n25)
         );
  NAND2_X1 maj_108_U4 ( .A1(maj_108_n20), .A2(maj_108_n19), .ZN(maj_108_n26)
         );
  NAND2_X1 maj_108_U3 ( .A1(maj_108_n26), .A2(maj_108_n25), .ZN(maj_108_port_o) );
  XOR2_X1 maj_108_U2 ( .A(maj_108_n22), .B(maj_108_n21), .Z(maj_108_n23) );
  NAND2_X1 maj_109_U15 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_109_n18) );
  NAND2_X1 maj_109_U14 ( .A1(maj_109_n21), .A2(maj_109_n22), .ZN(maj_109_n17)
         );
  NAND2_X1 maj_109_U13 ( .A1(maj_109_n18), .A2(maj_109_n17), .ZN(maj_109_n19)
         );
  NAND2_X1 maj_109_U12 ( .A1(v_0_0[2]), .A2(maj_109_n16), .ZN(maj_109_n14) );
  NAND2_X1 maj_109_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_109_n15) );
  NAND2_X1 maj_109_U10 ( .A1(maj_109_n15), .A2(maj_109_n14), .ZN(maj_109_n20)
         );
  XOR2_X1 maj_109_U9 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_109_n22) );
  XOR2_X1 maj_109_U8 ( .A(v_0_0[2]), .B(maj_109_n16), .Z(maj_109_n21) );
  XOR2_X1 maj_109_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_109_n16) );
  OR2_X1 maj_109_U6 ( .A1(maj_109_n20), .A2(maj_109_n19), .ZN(maj_109_n24) );
  NAND2_X1 maj_109_U5 ( .A1(maj_109_n24), .A2(maj_109_n23), .ZN(maj_109_n25)
         );
  NAND2_X1 maj_109_U4 ( .A1(maj_109_n20), .A2(maj_109_n19), .ZN(maj_109_n26)
         );
  NAND2_X1 maj_109_U3 ( .A1(maj_109_n26), .A2(maj_109_n25), .ZN(maj_109_port_o) );
  XOR2_X1 maj_109_U2 ( .A(maj_109_n22), .B(maj_109_n21), .Z(maj_109_n23) );
  NAND2_X1 maj_110_U15 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_110_n18) );
  NAND2_X1 maj_110_U14 ( .A1(maj_110_n21), .A2(maj_110_n22), .ZN(maj_110_n17)
         );
  NAND2_X1 maj_110_U13 ( .A1(maj_110_n18), .A2(maj_110_n17), .ZN(maj_110_n19)
         );
  NAND2_X1 maj_110_U12 ( .A1(u_0_1[2]), .A2(maj_110_n16), .ZN(maj_110_n14) );
  NAND2_X1 maj_110_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_110_n15) );
  NAND2_X1 maj_110_U10 ( .A1(maj_110_n15), .A2(maj_110_n14), .ZN(maj_110_n20)
         );
  XOR2_X1 maj_110_U9 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_110_n22) );
  XOR2_X1 maj_110_U8 ( .A(u_0_1[2]), .B(maj_110_n16), .Z(maj_110_n21) );
  XOR2_X1 maj_110_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_110_n16) );
  OR2_X1 maj_110_U6 ( .A1(maj_110_n20), .A2(maj_110_n19), .ZN(maj_110_n24) );
  NAND2_X1 maj_110_U5 ( .A1(maj_110_n24), .A2(maj_110_n23), .ZN(maj_110_n25)
         );
  NAND2_X1 maj_110_U4 ( .A1(maj_110_n20), .A2(maj_110_n19), .ZN(maj_110_n26)
         );
  NAND2_X1 maj_110_U3 ( .A1(maj_110_n26), .A2(maj_110_n25), .ZN(maj_110_port_o) );
  XOR2_X1 maj_110_U2 ( .A(maj_110_n22), .B(maj_110_n21), .Z(maj_110_n23) );
  NAND2_X1 maj_111_U15 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_111_n18) );
  NAND2_X1 maj_111_U14 ( .A1(maj_111_n21), .A2(maj_111_n22), .ZN(maj_111_n17)
         );
  NAND2_X1 maj_111_U13 ( .A1(maj_111_n18), .A2(maj_111_n17), .ZN(maj_111_n19)
         );
  NAND2_X1 maj_111_U12 ( .A1(v_0_1[2]), .A2(maj_111_n16), .ZN(maj_111_n14) );
  NAND2_X1 maj_111_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_111_n15) );
  NAND2_X1 maj_111_U10 ( .A1(maj_111_n15), .A2(maj_111_n14), .ZN(maj_111_n20)
         );
  XOR2_X1 maj_111_U9 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_111_n22) );
  XOR2_X1 maj_111_U8 ( .A(v_0_1[2]), .B(maj_111_n16), .Z(maj_111_n21) );
  XOR2_X1 maj_111_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_111_n16) );
  OR2_X1 maj_111_U6 ( .A1(maj_111_n20), .A2(maj_111_n19), .ZN(maj_111_n24) );
  NAND2_X1 maj_111_U5 ( .A1(maj_111_n24), .A2(maj_111_n23), .ZN(maj_111_n25)
         );
  NAND2_X1 maj_111_U4 ( .A1(maj_111_n20), .A2(maj_111_n19), .ZN(maj_111_n26)
         );
  NAND2_X1 maj_111_U3 ( .A1(maj_111_n26), .A2(maj_111_n25), .ZN(maj_111_port_o) );
  XOR2_X1 maj_111_U2 ( .A(maj_111_n22), .B(maj_111_n21), .Z(maj_111_n23) );
  NAND2_X1 maj_112_U15 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_112_n18) );
  NAND2_X1 maj_112_U14 ( .A1(maj_112_n21), .A2(maj_112_n22), .ZN(maj_112_n17)
         );
  NAND2_X1 maj_112_U13 ( .A1(maj_112_n18), .A2(maj_112_n17), .ZN(maj_112_n19)
         );
  NAND2_X1 maj_112_U12 ( .A1(u_1_0[2]), .A2(maj_112_n16), .ZN(maj_112_n14) );
  NAND2_X1 maj_112_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_112_n15) );
  NAND2_X1 maj_112_U10 ( .A1(maj_112_n15), .A2(maj_112_n14), .ZN(maj_112_n20)
         );
  XOR2_X1 maj_112_U9 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_112_n22) );
  XOR2_X1 maj_112_U8 ( .A(u_1_0[2]), .B(maj_112_n16), .Z(maj_112_n21) );
  XOR2_X1 maj_112_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_112_n16) );
  OR2_X1 maj_112_U6 ( .A1(maj_112_n20), .A2(maj_112_n19), .ZN(maj_112_n24) );
  NAND2_X1 maj_112_U5 ( .A1(maj_112_n24), .A2(maj_112_n23), .ZN(maj_112_n25)
         );
  NAND2_X1 maj_112_U4 ( .A1(maj_112_n20), .A2(maj_112_n19), .ZN(maj_112_n26)
         );
  NAND2_X1 maj_112_U3 ( .A1(maj_112_n26), .A2(maj_112_n25), .ZN(maj_112_port_o) );
  XOR2_X1 maj_112_U2 ( .A(maj_112_n22), .B(maj_112_n21), .Z(maj_112_n23) );
  NAND2_X1 maj_113_U15 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_113_n18) );
  NAND2_X1 maj_113_U14 ( .A1(maj_113_n21), .A2(maj_113_n22), .ZN(maj_113_n17)
         );
  NAND2_X1 maj_113_U13 ( .A1(maj_113_n18), .A2(maj_113_n17), .ZN(maj_113_n19)
         );
  NAND2_X1 maj_113_U12 ( .A1(v_1_0[2]), .A2(maj_113_n16), .ZN(maj_113_n14) );
  NAND2_X1 maj_113_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_113_n15) );
  NAND2_X1 maj_113_U10 ( .A1(maj_113_n15), .A2(maj_113_n14), .ZN(maj_113_n20)
         );
  XOR2_X1 maj_113_U9 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_113_n22) );
  XOR2_X1 maj_113_U8 ( .A(v_1_0[2]), .B(maj_113_n16), .Z(maj_113_n21) );
  XOR2_X1 maj_113_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_113_n16) );
  OR2_X1 maj_113_U6 ( .A1(maj_113_n20), .A2(maj_113_n19), .ZN(maj_113_n24) );
  NAND2_X1 maj_113_U5 ( .A1(maj_113_n24), .A2(maj_113_n23), .ZN(maj_113_n25)
         );
  NAND2_X1 maj_113_U4 ( .A1(maj_113_n20), .A2(maj_113_n19), .ZN(maj_113_n26)
         );
  NAND2_X1 maj_113_U3 ( .A1(maj_113_n26), .A2(maj_113_n25), .ZN(maj_113_port_o) );
  XOR2_X1 maj_113_U2 ( .A(maj_113_n22), .B(maj_113_n21), .Z(maj_113_n23) );
  NAND2_X1 maj_114_U15 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_114_n18) );
  NAND2_X1 maj_114_U14 ( .A1(maj_114_n21), .A2(maj_114_n22), .ZN(maj_114_n17)
         );
  NAND2_X1 maj_114_U13 ( .A1(maj_114_n18), .A2(maj_114_n17), .ZN(maj_114_n19)
         );
  NAND2_X1 maj_114_U12 ( .A1(u_1_1[2]), .A2(maj_114_n16), .ZN(maj_114_n14) );
  NAND2_X1 maj_114_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_114_n15) );
  NAND2_X1 maj_114_U10 ( .A1(maj_114_n15), .A2(maj_114_n14), .ZN(maj_114_n20)
         );
  XOR2_X1 maj_114_U9 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_114_n22) );
  XOR2_X1 maj_114_U8 ( .A(u_1_1[2]), .B(maj_114_n16), .Z(maj_114_n21) );
  XOR2_X1 maj_114_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_114_n16) );
  OR2_X1 maj_114_U6 ( .A1(maj_114_n20), .A2(maj_114_n19), .ZN(maj_114_n24) );
  NAND2_X1 maj_114_U5 ( .A1(maj_114_n24), .A2(maj_114_n23), .ZN(maj_114_n25)
         );
  NAND2_X1 maj_114_U4 ( .A1(maj_114_n20), .A2(maj_114_n19), .ZN(maj_114_n26)
         );
  NAND2_X1 maj_114_U3 ( .A1(maj_114_n26), .A2(maj_114_n25), .ZN(maj_114_port_o) );
  XOR2_X1 maj_114_U2 ( .A(maj_114_n22), .B(maj_114_n21), .Z(maj_114_n23) );
  NAND2_X1 maj_115_U15 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_115_n18) );
  NAND2_X1 maj_115_U14 ( .A1(maj_115_n21), .A2(maj_115_n22), .ZN(maj_115_n17)
         );
  NAND2_X1 maj_115_U13 ( .A1(maj_115_n18), .A2(maj_115_n17), .ZN(maj_115_n19)
         );
  NAND2_X1 maj_115_U12 ( .A1(v_1_1[2]), .A2(maj_115_n16), .ZN(maj_115_n14) );
  NAND2_X1 maj_115_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_115_n15) );
  NAND2_X1 maj_115_U10 ( .A1(maj_115_n15), .A2(maj_115_n14), .ZN(maj_115_n20)
         );
  XOR2_X1 maj_115_U9 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_115_n22) );
  XOR2_X1 maj_115_U8 ( .A(v_1_1[2]), .B(maj_115_n16), .Z(maj_115_n21) );
  XOR2_X1 maj_115_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_115_n16) );
  OR2_X1 maj_115_U6 ( .A1(maj_115_n20), .A2(maj_115_n19), .ZN(maj_115_n24) );
  NAND2_X1 maj_115_U5 ( .A1(maj_115_n24), .A2(maj_115_n23), .ZN(maj_115_n25)
         );
  NAND2_X1 maj_115_U4 ( .A1(maj_115_n20), .A2(maj_115_n19), .ZN(maj_115_n26)
         );
  NAND2_X1 maj_115_U3 ( .A1(maj_115_n26), .A2(maj_115_n25), .ZN(maj_115_port_o) );
  XOR2_X1 maj_115_U2 ( .A(maj_115_n22), .B(maj_115_n21), .Z(maj_115_n23) );
  NAND2_X1 maj_116_U15 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_116_n18) );
  NAND2_X1 maj_116_U14 ( .A1(maj_116_n21), .A2(maj_116_n22), .ZN(maj_116_n17)
         );
  NAND2_X1 maj_116_U13 ( .A1(maj_116_n18), .A2(maj_116_n17), .ZN(maj_116_n19)
         );
  NAND2_X1 maj_116_U12 ( .A1(u_2_0[2]), .A2(maj_116_n16), .ZN(maj_116_n14) );
  NAND2_X1 maj_116_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_116_n15) );
  NAND2_X1 maj_116_U10 ( .A1(maj_116_n15), .A2(maj_116_n14), .ZN(maj_116_n20)
         );
  XOR2_X1 maj_116_U9 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_116_n22) );
  XOR2_X1 maj_116_U8 ( .A(u_2_0[2]), .B(maj_116_n16), .Z(maj_116_n21) );
  XOR2_X1 maj_116_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_116_n16) );
  OR2_X1 maj_116_U6 ( .A1(maj_116_n20), .A2(maj_116_n19), .ZN(maj_116_n24) );
  NAND2_X1 maj_116_U5 ( .A1(maj_116_n24), .A2(maj_116_n23), .ZN(maj_116_n25)
         );
  NAND2_X1 maj_116_U4 ( .A1(maj_116_n20), .A2(maj_116_n19), .ZN(maj_116_n26)
         );
  NAND2_X1 maj_116_U3 ( .A1(maj_116_n26), .A2(maj_116_n25), .ZN(maj_116_port_o) );
  XOR2_X1 maj_116_U2 ( .A(maj_116_n22), .B(maj_116_n21), .Z(maj_116_n23) );
  NAND2_X1 maj_117_U15 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_117_n18) );
  NAND2_X1 maj_117_U14 ( .A1(maj_117_n21), .A2(maj_117_n22), .ZN(maj_117_n17)
         );
  NAND2_X1 maj_117_U13 ( .A1(maj_117_n18), .A2(maj_117_n17), .ZN(maj_117_n19)
         );
  NAND2_X1 maj_117_U12 ( .A1(v_2_0[2]), .A2(maj_117_n16), .ZN(maj_117_n14) );
  NAND2_X1 maj_117_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_117_n15) );
  NAND2_X1 maj_117_U10 ( .A1(maj_117_n15), .A2(maj_117_n14), .ZN(maj_117_n20)
         );
  XOR2_X1 maj_117_U9 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_117_n22) );
  XOR2_X1 maj_117_U8 ( .A(v_2_0[2]), .B(maj_117_n16), .Z(maj_117_n21) );
  XOR2_X1 maj_117_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_117_n16) );
  OR2_X1 maj_117_U6 ( .A1(maj_117_n20), .A2(maj_117_n19), .ZN(maj_117_n24) );
  NAND2_X1 maj_117_U5 ( .A1(maj_117_n24), .A2(maj_117_n23), .ZN(maj_117_n25)
         );
  NAND2_X1 maj_117_U4 ( .A1(maj_117_n20), .A2(maj_117_n19), .ZN(maj_117_n26)
         );
  NAND2_X1 maj_117_U3 ( .A1(maj_117_n26), .A2(maj_117_n25), .ZN(maj_117_port_o) );
  XOR2_X1 maj_117_U2 ( .A(maj_117_n22), .B(maj_117_n21), .Z(maj_117_n23) );
  NAND2_X1 maj_118_U15 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_118_n18) );
  NAND2_X1 maj_118_U14 ( .A1(maj_118_n21), .A2(maj_118_n22), .ZN(maj_118_n17)
         );
  NAND2_X1 maj_118_U13 ( .A1(maj_118_n18), .A2(maj_118_n17), .ZN(maj_118_n19)
         );
  NAND2_X1 maj_118_U12 ( .A1(u_2_1[2]), .A2(maj_118_n16), .ZN(maj_118_n14) );
  NAND2_X1 maj_118_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_118_n15) );
  NAND2_X1 maj_118_U10 ( .A1(maj_118_n15), .A2(maj_118_n14), .ZN(maj_118_n20)
         );
  XOR2_X1 maj_118_U9 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_118_n22) );
  XOR2_X1 maj_118_U8 ( .A(u_2_1[2]), .B(maj_118_n16), .Z(maj_118_n21) );
  XOR2_X1 maj_118_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_118_n16) );
  OR2_X1 maj_118_U6 ( .A1(maj_118_n20), .A2(maj_118_n19), .ZN(maj_118_n24) );
  NAND2_X1 maj_118_U5 ( .A1(maj_118_n24), .A2(maj_118_n23), .ZN(maj_118_n25)
         );
  NAND2_X1 maj_118_U4 ( .A1(maj_118_n20), .A2(maj_118_n19), .ZN(maj_118_n26)
         );
  NAND2_X1 maj_118_U3 ( .A1(maj_118_n26), .A2(maj_118_n25), .ZN(maj_118_port_o) );
  XOR2_X1 maj_118_U2 ( .A(maj_118_n22), .B(maj_118_n21), .Z(maj_118_n23) );
  NAND2_X1 maj_119_U15 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_119_n18) );
  NAND2_X1 maj_119_U14 ( .A1(maj_119_n21), .A2(maj_119_n22), .ZN(maj_119_n17)
         );
  NAND2_X1 maj_119_U13 ( .A1(maj_119_n18), .A2(maj_119_n17), .ZN(maj_119_n19)
         );
  NAND2_X1 maj_119_U12 ( .A1(v_2_1[2]), .A2(maj_119_n16), .ZN(maj_119_n14) );
  NAND2_X1 maj_119_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_119_n15) );
  NAND2_X1 maj_119_U10 ( .A1(maj_119_n15), .A2(maj_119_n14), .ZN(maj_119_n20)
         );
  XOR2_X1 maj_119_U9 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_119_n22) );
  XOR2_X1 maj_119_U8 ( .A(v_2_1[2]), .B(maj_119_n16), .Z(maj_119_n21) );
  XOR2_X1 maj_119_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_119_n16) );
  OR2_X1 maj_119_U6 ( .A1(maj_119_n20), .A2(maj_119_n19), .ZN(maj_119_n24) );
  NAND2_X1 maj_119_U5 ( .A1(maj_119_n24), .A2(maj_119_n23), .ZN(maj_119_n25)
         );
  NAND2_X1 maj_119_U4 ( .A1(maj_119_n20), .A2(maj_119_n19), .ZN(maj_119_n26)
         );
  NAND2_X1 maj_119_U3 ( .A1(maj_119_n26), .A2(maj_119_n25), .ZN(maj_119_port_o) );
  XOR2_X1 maj_119_U2 ( .A(maj_119_n22), .B(maj_119_n21), .Z(maj_119_n23) );
endmodule

