
module CINI_HPC3 ( port_a_0, port_a_1, port_a_2, port_a_3, port_b_0, port_b_1, 
        port_b_2, port_b_3, port_c_0, port_c_1, port_c_2, port_c_3, 
        port_rand_ref, port_rand_mul, clk, reset );
  input [6:0] port_a_0;
  input [6:0] port_a_1;
  input [6:0] port_a_2;
  input [6:0] port_a_3;
  input [6:0] port_b_0;
  input [6:0] port_b_1;
  input [6:0] port_b_2;
  input [6:0] port_b_3;
  output [6:0] port_c_0;
  output [6:0] port_c_1;
  output [6:0] port_c_2;
  output [6:0] port_c_3;
  input [5:0] port_rand_ref;
  input [5:0] port_rand_mul;
  input clk, reset;
  wire   simpleAnd_84_port_z, simpleAnd_85_port_z, simpleAnd_86_port_z,
         simpleAnd_87_port_z, simpleAnd_88_port_z, simpleAnd_89_port_z,
         simpleAnd_90_port_z, simpleAnd_91_port_z, simpleAnd_92_port_z,
         simpleAnd_93_port_z, simpleAnd_94_port_z, simpleAnd_95_port_z,
         simpleAnd_96_port_z, simpleAnd_97_port_z, simpleAnd_98_port_z,
         simpleAnd_99_port_z, simpleAnd_100_port_z, simpleAnd_101_port_z,
         simpleAnd_102_port_z, simpleAnd_103_port_z, simpleAnd_104_port_z,
         simpleAnd_105_port_z, simpleAnd_106_port_z, simpleAnd_107_port_z,
         simpleAnd_108_port_z, simpleAnd_109_port_z, simpleAnd_110_port_z,
         simpleAnd_111_port_z, simpleAnd_112_port_z, simpleAnd_113_port_z,
         simpleAnd_114_port_z, simpleAnd_115_port_z, simpleAnd_116_port_z,
         simpleAnd_117_port_z, simpleAnd_118_port_z, simpleAnd_119_port_z,
         simpleAnd_120_port_z, simpleAnd_121_port_z, simpleAnd_122_port_z,
         simpleAnd_123_port_z, simpleAnd_124_port_z, simpleAnd_125_port_z,
         simpleAnd_126_port_z, simpleAnd_127_port_z, simpleAnd_128_port_z,
         simpleAnd_129_port_z, simpleAnd_130_port_z, simpleAnd_131_port_z,
         simpleAnd_132_port_z, simpleAnd_133_port_z, simpleAnd_134_port_z,
         simpleAnd_135_port_z, simpleAnd_136_port_z, simpleAnd_137_port_z,
         simpleAnd_138_port_z, simpleAnd_139_port_z, simpleAnd_140_port_z,
         simpleAnd_141_port_z, simpleAnd_142_port_z, simpleAnd_143_port_z,
         simpleAnd_144_port_z, simpleAnd_145_port_z, simpleAnd_146_port_z,
         simpleAnd_147_port_z, simpleAnd_148_port_z, simpleAnd_149_port_z,
         simpleAnd_150_port_z, simpleAnd_151_port_z, simpleAnd_152_port_z,
         simpleAnd_153_port_z, simpleAnd_154_port_z, simpleAnd_155_port_z,
         simpleAnd_156_port_z, simpleAnd_157_port_z, simpleAnd_158_port_z,
         simpleAnd_159_port_z, simpleAnd_160_port_z, simpleAnd_161_port_z,
         simpleAnd_162_port_z, simpleAnd_163_port_z, simpleAnd_164_port_z,
         simpleAnd_165_port_z, simpleAnd_166_port_z, simpleAnd_167_port_z,
         maj_168_port_o, maj_169_port_o, maj_170_port_o, maj_171_port_o,
         maj_172_port_o, maj_173_port_o, maj_174_port_o, maj_175_port_o,
         maj_176_port_o, maj_177_port_o, maj_178_port_o, maj_179_port_o,
         maj_180_port_o, maj_181_port_o, maj_182_port_o, maj_183_port_o,
         maj_184_port_o, maj_185_port_o, maj_186_port_o, maj_187_port_o,
         maj_188_port_o, maj_189_port_o, maj_190_port_o, maj_191_port_o,
         maj_192_port_o, maj_193_port_o, maj_194_port_o, maj_195_port_o,
         maj_196_port_o, maj_197_port_o, maj_198_port_o, maj_199_port_o,
         maj_200_port_o, maj_201_port_o, maj_202_port_o, maj_203_port_o,
         maj_204_port_o, maj_205_port_o, maj_206_port_o, maj_207_port_o,
         maj_208_port_o, maj_209_port_o, maj_210_port_o, maj_211_port_o,
         maj_212_port_o, maj_213_port_o, maj_214_port_o, maj_215_port_o,
         maj_216_port_o, maj_217_port_o, maj_218_port_o, maj_219_port_o,
         maj_220_port_o, maj_221_port_o, maj_222_port_o, maj_223_port_o,
         maj_224_port_o, maj_225_port_o, maj_226_port_o, maj_227_port_o,
         maj_228_port_o, maj_229_port_o, maj_230_port_o, maj_231_port_o,
         maj_232_port_o, maj_233_port_o, maj_234_port_o, maj_235_port_o,
         maj_236_port_o, maj_237_port_o, maj_238_port_o, maj_239_port_o,
         maj_240_port_o, maj_241_port_o, maj_242_port_o, maj_243_port_o,
         maj_244_port_o, maj_245_port_o, maj_246_port_o, maj_247_port_o,
         maj_248_port_o, maj_249_port_o, maj_250_port_o, maj_251_port_o,
         maj_252_port_o, maj_253_port_o, maj_254_port_o, maj_255_port_o,
         maj_256_port_o, maj_257_port_o, maj_258_port_o, maj_259_port_o,
         maj_260_port_o, maj_261_port_o, maj_262_port_o, maj_263_port_o,
         maj_264_port_o, maj_265_port_o, maj_266_port_o, maj_267_port_o,
         maj_268_port_o, maj_269_port_o, maj_270_port_o, maj_271_port_o,
         maj_272_port_o, maj_273_port_o, maj_274_port_o, maj_275_port_o,
         maj_276_port_o, maj_277_port_o, maj_278_port_o, maj_279_port_o,
         maj_280_port_o, maj_281_port_o, maj_282_port_o, maj_283_port_o,
         maj_284_port_o, maj_285_port_o, maj_286_port_o, maj_287_port_o,
         maj_288_port_o, maj_289_port_o, maj_290_port_o, maj_291_port_o,
         maj_292_port_o, maj_293_port_o, maj_294_port_o, maj_295_port_o,
         maj_296_port_o, maj_297_port_o, maj_298_port_o, maj_299_port_o,
         maj_300_port_o, maj_301_port_o, maj_302_port_o, maj_303_port_o,
         maj_304_port_o, maj_305_port_o, maj_306_port_o, maj_307_port_o,
         maj_308_port_o, maj_309_port_o, maj_310_port_o, maj_311_port_o,
         maj_312_port_o, maj_313_port_o, maj_314_port_o, maj_315_port_o,
         maj_316_port_o, maj_317_port_o, maj_318_port_o, maj_319_port_o,
         maj_320_port_o, maj_321_port_o, maj_322_port_o, maj_323_port_o,
         maj_324_port_o, maj_325_port_o, maj_326_port_o, maj_327_port_o,
         maj_328_port_o, maj_329_port_o, maj_330_port_o, maj_331_port_o,
         maj_332_port_o, maj_333_port_o, maj_334_port_o, maj_335_port_o, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, maj_168_n17, maj_168_n16,
         maj_168_n15, maj_168_n14, maj_168_n13, maj_168_n12, maj_168_n11,
         maj_168_n10, maj_168_n9, maj_168_n8, maj_168_n7, maj_168_n6,
         maj_168_n5, maj_168_n4, maj_168_n3, maj_168_n2, maj_168_n1,
         maj_169_n34, maj_169_n33, maj_169_n32, maj_169_n31, maj_169_n30,
         maj_169_n29, maj_169_n28, maj_169_n27, maj_169_n26, maj_169_n25,
         maj_169_n24, maj_169_n23, maj_169_n22, maj_169_n21, maj_169_n20,
         maj_169_n19, maj_169_n18, maj_170_n34, maj_170_n33, maj_170_n32,
         maj_170_n31, maj_170_n30, maj_170_n29, maj_170_n28, maj_170_n27,
         maj_170_n26, maj_170_n25, maj_170_n24, maj_170_n23, maj_170_n22,
         maj_170_n21, maj_170_n20, maj_170_n19, maj_170_n18, maj_171_n34,
         maj_171_n33, maj_171_n32, maj_171_n31, maj_171_n30, maj_171_n29,
         maj_171_n28, maj_171_n27, maj_171_n26, maj_171_n25, maj_171_n24,
         maj_171_n23, maj_171_n22, maj_171_n21, maj_171_n20, maj_171_n19,
         maj_171_n18, maj_172_n34, maj_172_n33, maj_172_n32, maj_172_n31,
         maj_172_n30, maj_172_n29, maj_172_n28, maj_172_n27, maj_172_n26,
         maj_172_n25, maj_172_n24, maj_172_n23, maj_172_n22, maj_172_n21,
         maj_172_n20, maj_172_n19, maj_172_n18, maj_173_n34, maj_173_n33,
         maj_173_n32, maj_173_n31, maj_173_n30, maj_173_n29, maj_173_n28,
         maj_173_n27, maj_173_n26, maj_173_n25, maj_173_n24, maj_173_n23,
         maj_173_n22, maj_173_n21, maj_173_n20, maj_173_n19, maj_173_n18,
         maj_174_n34, maj_174_n33, maj_174_n32, maj_174_n31, maj_174_n30,
         maj_174_n29, maj_174_n28, maj_174_n27, maj_174_n26, maj_174_n25,
         maj_174_n24, maj_174_n23, maj_174_n22, maj_174_n21, maj_174_n20,
         maj_174_n19, maj_174_n18, maj_175_n34, maj_175_n33, maj_175_n32,
         maj_175_n31, maj_175_n30, maj_175_n29, maj_175_n28, maj_175_n27,
         maj_175_n26, maj_175_n25, maj_175_n24, maj_175_n23, maj_175_n22,
         maj_175_n21, maj_175_n20, maj_175_n19, maj_175_n18, maj_176_n34,
         maj_176_n33, maj_176_n32, maj_176_n31, maj_176_n30, maj_176_n29,
         maj_176_n28, maj_176_n27, maj_176_n26, maj_176_n25, maj_176_n24,
         maj_176_n23, maj_176_n22, maj_176_n21, maj_176_n20, maj_176_n19,
         maj_176_n18, maj_177_n34, maj_177_n33, maj_177_n32, maj_177_n31,
         maj_177_n30, maj_177_n29, maj_177_n28, maj_177_n27, maj_177_n26,
         maj_177_n25, maj_177_n24, maj_177_n23, maj_177_n22, maj_177_n21,
         maj_177_n20, maj_177_n19, maj_177_n18, maj_178_n34, maj_178_n33,
         maj_178_n32, maj_178_n31, maj_178_n30, maj_178_n29, maj_178_n28,
         maj_178_n27, maj_178_n26, maj_178_n25, maj_178_n24, maj_178_n23,
         maj_178_n22, maj_178_n21, maj_178_n20, maj_178_n19, maj_178_n18,
         maj_179_n34, maj_179_n33, maj_179_n32, maj_179_n31, maj_179_n30,
         maj_179_n29, maj_179_n28, maj_179_n27, maj_179_n26, maj_179_n25,
         maj_179_n24, maj_179_n23, maj_179_n22, maj_179_n21, maj_179_n20,
         maj_179_n19, maj_179_n18, maj_180_n34, maj_180_n33, maj_180_n32,
         maj_180_n31, maj_180_n30, maj_180_n29, maj_180_n28, maj_180_n27,
         maj_180_n26, maj_180_n25, maj_180_n24, maj_180_n23, maj_180_n22,
         maj_180_n21, maj_180_n20, maj_180_n19, maj_180_n18, maj_181_n34,
         maj_181_n33, maj_181_n32, maj_181_n31, maj_181_n30, maj_181_n29,
         maj_181_n28, maj_181_n27, maj_181_n26, maj_181_n25, maj_181_n24,
         maj_181_n23, maj_181_n22, maj_181_n21, maj_181_n20, maj_181_n19,
         maj_181_n18, maj_182_n34, maj_182_n33, maj_182_n32, maj_182_n31,
         maj_182_n30, maj_182_n29, maj_182_n28, maj_182_n27, maj_182_n26,
         maj_182_n25, maj_182_n24, maj_182_n23, maj_182_n22, maj_182_n21,
         maj_182_n20, maj_182_n19, maj_182_n18, maj_183_n34, maj_183_n33,
         maj_183_n32, maj_183_n31, maj_183_n30, maj_183_n29, maj_183_n28,
         maj_183_n27, maj_183_n26, maj_183_n25, maj_183_n24, maj_183_n23,
         maj_183_n22, maj_183_n21, maj_183_n20, maj_183_n19, maj_183_n18,
         maj_184_n34, maj_184_n33, maj_184_n32, maj_184_n31, maj_184_n30,
         maj_184_n29, maj_184_n28, maj_184_n27, maj_184_n26, maj_184_n25,
         maj_184_n24, maj_184_n23, maj_184_n22, maj_184_n21, maj_184_n20,
         maj_184_n19, maj_184_n18, maj_185_n34, maj_185_n33, maj_185_n32,
         maj_185_n31, maj_185_n30, maj_185_n29, maj_185_n28, maj_185_n27,
         maj_185_n26, maj_185_n25, maj_185_n24, maj_185_n23, maj_185_n22,
         maj_185_n21, maj_185_n20, maj_185_n19, maj_185_n18, maj_186_n34,
         maj_186_n33, maj_186_n32, maj_186_n31, maj_186_n30, maj_186_n29,
         maj_186_n28, maj_186_n27, maj_186_n26, maj_186_n25, maj_186_n24,
         maj_186_n23, maj_186_n22, maj_186_n21, maj_186_n20, maj_186_n19,
         maj_186_n18, maj_187_n34, maj_187_n33, maj_187_n32, maj_187_n31,
         maj_187_n30, maj_187_n29, maj_187_n28, maj_187_n27, maj_187_n26,
         maj_187_n25, maj_187_n24, maj_187_n23, maj_187_n22, maj_187_n21,
         maj_187_n20, maj_187_n19, maj_187_n18, maj_188_n34, maj_188_n33,
         maj_188_n32, maj_188_n31, maj_188_n30, maj_188_n29, maj_188_n28,
         maj_188_n27, maj_188_n26, maj_188_n25, maj_188_n24, maj_188_n23,
         maj_188_n22, maj_188_n21, maj_188_n20, maj_188_n19, maj_188_n18,
         maj_189_n34, maj_189_n33, maj_189_n32, maj_189_n31, maj_189_n30,
         maj_189_n29, maj_189_n28, maj_189_n27, maj_189_n26, maj_189_n25,
         maj_189_n24, maj_189_n23, maj_189_n22, maj_189_n21, maj_189_n20,
         maj_189_n19, maj_189_n18, maj_190_n34, maj_190_n33, maj_190_n32,
         maj_190_n31, maj_190_n30, maj_190_n29, maj_190_n28, maj_190_n27,
         maj_190_n26, maj_190_n25, maj_190_n24, maj_190_n23, maj_190_n22,
         maj_190_n21, maj_190_n20, maj_190_n19, maj_190_n18, maj_191_n34,
         maj_191_n33, maj_191_n32, maj_191_n31, maj_191_n30, maj_191_n29,
         maj_191_n28, maj_191_n27, maj_191_n26, maj_191_n25, maj_191_n24,
         maj_191_n23, maj_191_n22, maj_191_n21, maj_191_n20, maj_191_n19,
         maj_191_n18, maj_192_n34, maj_192_n33, maj_192_n32, maj_192_n31,
         maj_192_n30, maj_192_n29, maj_192_n28, maj_192_n27, maj_192_n26,
         maj_192_n25, maj_192_n24, maj_192_n23, maj_192_n22, maj_192_n21,
         maj_192_n20, maj_192_n19, maj_192_n18, maj_193_n34, maj_193_n33,
         maj_193_n32, maj_193_n31, maj_193_n30, maj_193_n29, maj_193_n28,
         maj_193_n27, maj_193_n26, maj_193_n25, maj_193_n24, maj_193_n23,
         maj_193_n22, maj_193_n21, maj_193_n20, maj_193_n19, maj_193_n18,
         maj_194_n34, maj_194_n33, maj_194_n32, maj_194_n31, maj_194_n30,
         maj_194_n29, maj_194_n28, maj_194_n27, maj_194_n26, maj_194_n25,
         maj_194_n24, maj_194_n23, maj_194_n22, maj_194_n21, maj_194_n20,
         maj_194_n19, maj_194_n18, maj_195_n34, maj_195_n33, maj_195_n32,
         maj_195_n31, maj_195_n30, maj_195_n29, maj_195_n28, maj_195_n27,
         maj_195_n26, maj_195_n25, maj_195_n24, maj_195_n23, maj_195_n22,
         maj_195_n21, maj_195_n20, maj_195_n19, maj_195_n18, maj_196_n34,
         maj_196_n33, maj_196_n32, maj_196_n31, maj_196_n30, maj_196_n29,
         maj_196_n28, maj_196_n27, maj_196_n26, maj_196_n25, maj_196_n24,
         maj_196_n23, maj_196_n22, maj_196_n21, maj_196_n20, maj_196_n19,
         maj_196_n18, maj_197_n34, maj_197_n33, maj_197_n32, maj_197_n31,
         maj_197_n30, maj_197_n29, maj_197_n28, maj_197_n27, maj_197_n26,
         maj_197_n25, maj_197_n24, maj_197_n23, maj_197_n22, maj_197_n21,
         maj_197_n20, maj_197_n19, maj_197_n18, maj_198_n34, maj_198_n33,
         maj_198_n32, maj_198_n31, maj_198_n30, maj_198_n29, maj_198_n28,
         maj_198_n27, maj_198_n26, maj_198_n25, maj_198_n24, maj_198_n23,
         maj_198_n22, maj_198_n21, maj_198_n20, maj_198_n19, maj_198_n18,
         maj_199_n34, maj_199_n33, maj_199_n32, maj_199_n31, maj_199_n30,
         maj_199_n29, maj_199_n28, maj_199_n27, maj_199_n26, maj_199_n25,
         maj_199_n24, maj_199_n23, maj_199_n22, maj_199_n21, maj_199_n20,
         maj_199_n19, maj_199_n18, maj_200_n34, maj_200_n33, maj_200_n32,
         maj_200_n31, maj_200_n30, maj_200_n29, maj_200_n28, maj_200_n27,
         maj_200_n26, maj_200_n25, maj_200_n24, maj_200_n23, maj_200_n22,
         maj_200_n21, maj_200_n20, maj_200_n19, maj_200_n18, maj_201_n34,
         maj_201_n33, maj_201_n32, maj_201_n31, maj_201_n30, maj_201_n29,
         maj_201_n28, maj_201_n27, maj_201_n26, maj_201_n25, maj_201_n24,
         maj_201_n23, maj_201_n22, maj_201_n21, maj_201_n20, maj_201_n19,
         maj_201_n18, maj_202_n34, maj_202_n33, maj_202_n32, maj_202_n31,
         maj_202_n30, maj_202_n29, maj_202_n28, maj_202_n27, maj_202_n26,
         maj_202_n25, maj_202_n24, maj_202_n23, maj_202_n22, maj_202_n21,
         maj_202_n20, maj_202_n19, maj_202_n18, maj_203_n34, maj_203_n33,
         maj_203_n32, maj_203_n31, maj_203_n30, maj_203_n29, maj_203_n28,
         maj_203_n27, maj_203_n26, maj_203_n25, maj_203_n24, maj_203_n23,
         maj_203_n22, maj_203_n21, maj_203_n20, maj_203_n19, maj_203_n18,
         maj_204_n34, maj_204_n33, maj_204_n32, maj_204_n31, maj_204_n30,
         maj_204_n29, maj_204_n28, maj_204_n27, maj_204_n26, maj_204_n25,
         maj_204_n24, maj_204_n23, maj_204_n22, maj_204_n21, maj_204_n20,
         maj_204_n19, maj_204_n18, maj_205_n34, maj_205_n33, maj_205_n32,
         maj_205_n31, maj_205_n30, maj_205_n29, maj_205_n28, maj_205_n27,
         maj_205_n26, maj_205_n25, maj_205_n24, maj_205_n23, maj_205_n22,
         maj_205_n21, maj_205_n20, maj_205_n19, maj_205_n18, maj_206_n34,
         maj_206_n33, maj_206_n32, maj_206_n31, maj_206_n30, maj_206_n29,
         maj_206_n28, maj_206_n27, maj_206_n26, maj_206_n25, maj_206_n24,
         maj_206_n23, maj_206_n22, maj_206_n21, maj_206_n20, maj_206_n19,
         maj_206_n18, maj_207_n34, maj_207_n33, maj_207_n32, maj_207_n31,
         maj_207_n30, maj_207_n29, maj_207_n28, maj_207_n27, maj_207_n26,
         maj_207_n25, maj_207_n24, maj_207_n23, maj_207_n22, maj_207_n21,
         maj_207_n20, maj_207_n19, maj_207_n18, maj_208_n34, maj_208_n33,
         maj_208_n32, maj_208_n31, maj_208_n30, maj_208_n29, maj_208_n28,
         maj_208_n27, maj_208_n26, maj_208_n25, maj_208_n24, maj_208_n23,
         maj_208_n22, maj_208_n21, maj_208_n20, maj_208_n19, maj_208_n18,
         maj_209_n34, maj_209_n33, maj_209_n32, maj_209_n31, maj_209_n30,
         maj_209_n29, maj_209_n28, maj_209_n27, maj_209_n26, maj_209_n25,
         maj_209_n24, maj_209_n23, maj_209_n22, maj_209_n21, maj_209_n20,
         maj_209_n19, maj_209_n18, maj_210_n34, maj_210_n33, maj_210_n32,
         maj_210_n31, maj_210_n30, maj_210_n29, maj_210_n28, maj_210_n27,
         maj_210_n26, maj_210_n25, maj_210_n24, maj_210_n23, maj_210_n22,
         maj_210_n21, maj_210_n20, maj_210_n19, maj_210_n18, maj_211_n34,
         maj_211_n33, maj_211_n32, maj_211_n31, maj_211_n30, maj_211_n29,
         maj_211_n28, maj_211_n27, maj_211_n26, maj_211_n25, maj_211_n24,
         maj_211_n23, maj_211_n22, maj_211_n21, maj_211_n20, maj_211_n19,
         maj_211_n18, maj_212_n34, maj_212_n33, maj_212_n32, maj_212_n31,
         maj_212_n30, maj_212_n29, maj_212_n28, maj_212_n27, maj_212_n26,
         maj_212_n25, maj_212_n24, maj_212_n23, maj_212_n22, maj_212_n21,
         maj_212_n20, maj_212_n19, maj_212_n18, maj_213_n34, maj_213_n33,
         maj_213_n32, maj_213_n31, maj_213_n30, maj_213_n29, maj_213_n28,
         maj_213_n27, maj_213_n26, maj_213_n25, maj_213_n24, maj_213_n23,
         maj_213_n22, maj_213_n21, maj_213_n20, maj_213_n19, maj_213_n18,
         maj_214_n34, maj_214_n33, maj_214_n32, maj_214_n31, maj_214_n30,
         maj_214_n29, maj_214_n28, maj_214_n27, maj_214_n26, maj_214_n25,
         maj_214_n24, maj_214_n23, maj_214_n22, maj_214_n21, maj_214_n20,
         maj_214_n19, maj_214_n18, maj_215_n34, maj_215_n33, maj_215_n32,
         maj_215_n31, maj_215_n30, maj_215_n29, maj_215_n28, maj_215_n27,
         maj_215_n26, maj_215_n25, maj_215_n24, maj_215_n23, maj_215_n22,
         maj_215_n21, maj_215_n20, maj_215_n19, maj_215_n18, maj_216_n34,
         maj_216_n33, maj_216_n32, maj_216_n31, maj_216_n30, maj_216_n29,
         maj_216_n28, maj_216_n27, maj_216_n26, maj_216_n25, maj_216_n24,
         maj_216_n23, maj_216_n22, maj_216_n21, maj_216_n20, maj_216_n19,
         maj_216_n18, maj_217_n34, maj_217_n33, maj_217_n32, maj_217_n31,
         maj_217_n30, maj_217_n29, maj_217_n28, maj_217_n27, maj_217_n26,
         maj_217_n25, maj_217_n24, maj_217_n23, maj_217_n22, maj_217_n21,
         maj_217_n20, maj_217_n19, maj_217_n18, maj_218_n34, maj_218_n33,
         maj_218_n32, maj_218_n31, maj_218_n30, maj_218_n29, maj_218_n28,
         maj_218_n27, maj_218_n26, maj_218_n25, maj_218_n24, maj_218_n23,
         maj_218_n22, maj_218_n21, maj_218_n20, maj_218_n19, maj_218_n18,
         maj_219_n34, maj_219_n33, maj_219_n32, maj_219_n31, maj_219_n30,
         maj_219_n29, maj_219_n28, maj_219_n27, maj_219_n26, maj_219_n25,
         maj_219_n24, maj_219_n23, maj_219_n22, maj_219_n21, maj_219_n20,
         maj_219_n19, maj_219_n18, maj_220_n34, maj_220_n33, maj_220_n32,
         maj_220_n31, maj_220_n30, maj_220_n29, maj_220_n28, maj_220_n27,
         maj_220_n26, maj_220_n25, maj_220_n24, maj_220_n23, maj_220_n22,
         maj_220_n21, maj_220_n20, maj_220_n19, maj_220_n18, maj_221_n34,
         maj_221_n33, maj_221_n32, maj_221_n31, maj_221_n30, maj_221_n29,
         maj_221_n28, maj_221_n27, maj_221_n26, maj_221_n25, maj_221_n24,
         maj_221_n23, maj_221_n22, maj_221_n21, maj_221_n20, maj_221_n19,
         maj_221_n18, maj_222_n34, maj_222_n33, maj_222_n32, maj_222_n31,
         maj_222_n30, maj_222_n29, maj_222_n28, maj_222_n27, maj_222_n26,
         maj_222_n25, maj_222_n24, maj_222_n23, maj_222_n22, maj_222_n21,
         maj_222_n20, maj_222_n19, maj_222_n18, maj_223_n34, maj_223_n33,
         maj_223_n32, maj_223_n31, maj_223_n30, maj_223_n29, maj_223_n28,
         maj_223_n27, maj_223_n26, maj_223_n25, maj_223_n24, maj_223_n23,
         maj_223_n22, maj_223_n21, maj_223_n20, maj_223_n19, maj_223_n18,
         maj_224_n34, maj_224_n33, maj_224_n32, maj_224_n31, maj_224_n30,
         maj_224_n29, maj_224_n28, maj_224_n27, maj_224_n26, maj_224_n25,
         maj_224_n24, maj_224_n23, maj_224_n22, maj_224_n21, maj_224_n20,
         maj_224_n19, maj_224_n18, maj_225_n34, maj_225_n33, maj_225_n32,
         maj_225_n31, maj_225_n30, maj_225_n29, maj_225_n28, maj_225_n27,
         maj_225_n26, maj_225_n25, maj_225_n24, maj_225_n23, maj_225_n22,
         maj_225_n21, maj_225_n20, maj_225_n19, maj_225_n18, maj_226_n34,
         maj_226_n33, maj_226_n32, maj_226_n31, maj_226_n30, maj_226_n29,
         maj_226_n28, maj_226_n27, maj_226_n26, maj_226_n25, maj_226_n24,
         maj_226_n23, maj_226_n22, maj_226_n21, maj_226_n20, maj_226_n19,
         maj_226_n18, maj_227_n34, maj_227_n33, maj_227_n32, maj_227_n31,
         maj_227_n30, maj_227_n29, maj_227_n28, maj_227_n27, maj_227_n26,
         maj_227_n25, maj_227_n24, maj_227_n23, maj_227_n22, maj_227_n21,
         maj_227_n20, maj_227_n19, maj_227_n18, maj_228_n34, maj_228_n33,
         maj_228_n32, maj_228_n31, maj_228_n30, maj_228_n29, maj_228_n28,
         maj_228_n27, maj_228_n26, maj_228_n25, maj_228_n24, maj_228_n23,
         maj_228_n22, maj_228_n21, maj_228_n20, maj_228_n19, maj_228_n18,
         maj_229_n34, maj_229_n33, maj_229_n32, maj_229_n31, maj_229_n30,
         maj_229_n29, maj_229_n28, maj_229_n27, maj_229_n26, maj_229_n25,
         maj_229_n24, maj_229_n23, maj_229_n22, maj_229_n21, maj_229_n20,
         maj_229_n19, maj_229_n18, maj_230_n34, maj_230_n33, maj_230_n32,
         maj_230_n31, maj_230_n30, maj_230_n29, maj_230_n28, maj_230_n27,
         maj_230_n26, maj_230_n25, maj_230_n24, maj_230_n23, maj_230_n22,
         maj_230_n21, maj_230_n20, maj_230_n19, maj_230_n18, maj_231_n34,
         maj_231_n33, maj_231_n32, maj_231_n31, maj_231_n30, maj_231_n29,
         maj_231_n28, maj_231_n27, maj_231_n26, maj_231_n25, maj_231_n24,
         maj_231_n23, maj_231_n22, maj_231_n21, maj_231_n20, maj_231_n19,
         maj_231_n18, maj_232_n34, maj_232_n33, maj_232_n32, maj_232_n31,
         maj_232_n30, maj_232_n29, maj_232_n28, maj_232_n27, maj_232_n26,
         maj_232_n25, maj_232_n24, maj_232_n23, maj_232_n22, maj_232_n21,
         maj_232_n20, maj_232_n19, maj_232_n18, maj_233_n34, maj_233_n33,
         maj_233_n32, maj_233_n31, maj_233_n30, maj_233_n29, maj_233_n28,
         maj_233_n27, maj_233_n26, maj_233_n25, maj_233_n24, maj_233_n23,
         maj_233_n22, maj_233_n21, maj_233_n20, maj_233_n19, maj_233_n18,
         maj_234_n34, maj_234_n33, maj_234_n32, maj_234_n31, maj_234_n30,
         maj_234_n29, maj_234_n28, maj_234_n27, maj_234_n26, maj_234_n25,
         maj_234_n24, maj_234_n23, maj_234_n22, maj_234_n21, maj_234_n20,
         maj_234_n19, maj_234_n18, maj_235_n34, maj_235_n33, maj_235_n32,
         maj_235_n31, maj_235_n30, maj_235_n29, maj_235_n28, maj_235_n27,
         maj_235_n26, maj_235_n25, maj_235_n24, maj_235_n23, maj_235_n22,
         maj_235_n21, maj_235_n20, maj_235_n19, maj_235_n18, maj_236_n34,
         maj_236_n33, maj_236_n32, maj_236_n31, maj_236_n30, maj_236_n29,
         maj_236_n28, maj_236_n27, maj_236_n26, maj_236_n25, maj_236_n24,
         maj_236_n23, maj_236_n22, maj_236_n21, maj_236_n20, maj_236_n19,
         maj_236_n18, maj_237_n34, maj_237_n33, maj_237_n32, maj_237_n31,
         maj_237_n30, maj_237_n29, maj_237_n28, maj_237_n27, maj_237_n26,
         maj_237_n25, maj_237_n24, maj_237_n23, maj_237_n22, maj_237_n21,
         maj_237_n20, maj_237_n19, maj_237_n18, maj_238_n34, maj_238_n33,
         maj_238_n32, maj_238_n31, maj_238_n30, maj_238_n29, maj_238_n28,
         maj_238_n27, maj_238_n26, maj_238_n25, maj_238_n24, maj_238_n23,
         maj_238_n22, maj_238_n21, maj_238_n20, maj_238_n19, maj_238_n18,
         maj_239_n34, maj_239_n33, maj_239_n32, maj_239_n31, maj_239_n30,
         maj_239_n29, maj_239_n28, maj_239_n27, maj_239_n26, maj_239_n25,
         maj_239_n24, maj_239_n23, maj_239_n22, maj_239_n21, maj_239_n20,
         maj_239_n19, maj_239_n18, maj_240_n34, maj_240_n33, maj_240_n32,
         maj_240_n31, maj_240_n30, maj_240_n29, maj_240_n28, maj_240_n27,
         maj_240_n26, maj_240_n25, maj_240_n24, maj_240_n23, maj_240_n22,
         maj_240_n21, maj_240_n20, maj_240_n19, maj_240_n18, maj_241_n34,
         maj_241_n33, maj_241_n32, maj_241_n31, maj_241_n30, maj_241_n29,
         maj_241_n28, maj_241_n27, maj_241_n26, maj_241_n25, maj_241_n24,
         maj_241_n23, maj_241_n22, maj_241_n21, maj_241_n20, maj_241_n19,
         maj_241_n18, maj_242_n34, maj_242_n33, maj_242_n32, maj_242_n31,
         maj_242_n30, maj_242_n29, maj_242_n28, maj_242_n27, maj_242_n26,
         maj_242_n25, maj_242_n24, maj_242_n23, maj_242_n22, maj_242_n21,
         maj_242_n20, maj_242_n19, maj_242_n18, maj_243_n34, maj_243_n33,
         maj_243_n32, maj_243_n31, maj_243_n30, maj_243_n29, maj_243_n28,
         maj_243_n27, maj_243_n26, maj_243_n25, maj_243_n24, maj_243_n23,
         maj_243_n22, maj_243_n21, maj_243_n20, maj_243_n19, maj_243_n18,
         maj_244_n34, maj_244_n33, maj_244_n32, maj_244_n31, maj_244_n30,
         maj_244_n29, maj_244_n28, maj_244_n27, maj_244_n26, maj_244_n25,
         maj_244_n24, maj_244_n23, maj_244_n22, maj_244_n21, maj_244_n20,
         maj_244_n19, maj_244_n18, maj_245_n34, maj_245_n33, maj_245_n32,
         maj_245_n31, maj_245_n30, maj_245_n29, maj_245_n28, maj_245_n27,
         maj_245_n26, maj_245_n25, maj_245_n24, maj_245_n23, maj_245_n22,
         maj_245_n21, maj_245_n20, maj_245_n19, maj_245_n18, maj_246_n34,
         maj_246_n33, maj_246_n32, maj_246_n31, maj_246_n30, maj_246_n29,
         maj_246_n28, maj_246_n27, maj_246_n26, maj_246_n25, maj_246_n24,
         maj_246_n23, maj_246_n22, maj_246_n21, maj_246_n20, maj_246_n19,
         maj_246_n18, maj_247_n34, maj_247_n33, maj_247_n32, maj_247_n31,
         maj_247_n30, maj_247_n29, maj_247_n28, maj_247_n27, maj_247_n26,
         maj_247_n25, maj_247_n24, maj_247_n23, maj_247_n22, maj_247_n21,
         maj_247_n20, maj_247_n19, maj_247_n18, maj_248_n34, maj_248_n33,
         maj_248_n32, maj_248_n31, maj_248_n30, maj_248_n29, maj_248_n28,
         maj_248_n27, maj_248_n26, maj_248_n25, maj_248_n24, maj_248_n23,
         maj_248_n22, maj_248_n21, maj_248_n20, maj_248_n19, maj_248_n18,
         maj_249_n34, maj_249_n33, maj_249_n32, maj_249_n31, maj_249_n30,
         maj_249_n29, maj_249_n28, maj_249_n27, maj_249_n26, maj_249_n25,
         maj_249_n24, maj_249_n23, maj_249_n22, maj_249_n21, maj_249_n20,
         maj_249_n19, maj_249_n18, maj_250_n34, maj_250_n33, maj_250_n32,
         maj_250_n31, maj_250_n30, maj_250_n29, maj_250_n28, maj_250_n27,
         maj_250_n26, maj_250_n25, maj_250_n24, maj_250_n23, maj_250_n22,
         maj_250_n21, maj_250_n20, maj_250_n19, maj_250_n18, maj_251_n34,
         maj_251_n33, maj_251_n32, maj_251_n31, maj_251_n30, maj_251_n29,
         maj_251_n28, maj_251_n27, maj_251_n26, maj_251_n25, maj_251_n24,
         maj_251_n23, maj_251_n22, maj_251_n21, maj_251_n20, maj_251_n19,
         maj_251_n18, maj_252_n34, maj_252_n33, maj_252_n32, maj_252_n31,
         maj_252_n30, maj_252_n29, maj_252_n28, maj_252_n27, maj_252_n26,
         maj_252_n25, maj_252_n24, maj_252_n23, maj_252_n22, maj_252_n21,
         maj_252_n20, maj_252_n19, maj_252_n18, maj_253_n34, maj_253_n33,
         maj_253_n32, maj_253_n31, maj_253_n30, maj_253_n29, maj_253_n28,
         maj_253_n27, maj_253_n26, maj_253_n25, maj_253_n24, maj_253_n23,
         maj_253_n22, maj_253_n21, maj_253_n20, maj_253_n19, maj_253_n18,
         maj_254_n34, maj_254_n33, maj_254_n32, maj_254_n31, maj_254_n30,
         maj_254_n29, maj_254_n28, maj_254_n27, maj_254_n26, maj_254_n25,
         maj_254_n24, maj_254_n23, maj_254_n22, maj_254_n21, maj_254_n20,
         maj_254_n19, maj_254_n18, maj_255_n34, maj_255_n33, maj_255_n32,
         maj_255_n31, maj_255_n30, maj_255_n29, maj_255_n28, maj_255_n27,
         maj_255_n26, maj_255_n25, maj_255_n24, maj_255_n23, maj_255_n22,
         maj_255_n21, maj_255_n20, maj_255_n19, maj_255_n18, maj_256_n34,
         maj_256_n33, maj_256_n32, maj_256_n31, maj_256_n30, maj_256_n29,
         maj_256_n28, maj_256_n27, maj_256_n26, maj_256_n25, maj_256_n24,
         maj_256_n23, maj_256_n22, maj_256_n21, maj_256_n20, maj_256_n19,
         maj_256_n18, maj_257_n34, maj_257_n33, maj_257_n32, maj_257_n31,
         maj_257_n30, maj_257_n29, maj_257_n28, maj_257_n27, maj_257_n26,
         maj_257_n25, maj_257_n24, maj_257_n23, maj_257_n22, maj_257_n21,
         maj_257_n20, maj_257_n19, maj_257_n18, maj_258_n34, maj_258_n33,
         maj_258_n32, maj_258_n31, maj_258_n30, maj_258_n29, maj_258_n28,
         maj_258_n27, maj_258_n26, maj_258_n25, maj_258_n24, maj_258_n23,
         maj_258_n22, maj_258_n21, maj_258_n20, maj_258_n19, maj_258_n18,
         maj_259_n34, maj_259_n33, maj_259_n32, maj_259_n31, maj_259_n30,
         maj_259_n29, maj_259_n28, maj_259_n27, maj_259_n26, maj_259_n25,
         maj_259_n24, maj_259_n23, maj_259_n22, maj_259_n21, maj_259_n20,
         maj_259_n19, maj_259_n18, maj_260_n34, maj_260_n33, maj_260_n32,
         maj_260_n31, maj_260_n30, maj_260_n29, maj_260_n28, maj_260_n27,
         maj_260_n26, maj_260_n25, maj_260_n24, maj_260_n23, maj_260_n22,
         maj_260_n21, maj_260_n20, maj_260_n19, maj_260_n18, maj_261_n34,
         maj_261_n33, maj_261_n32, maj_261_n31, maj_261_n30, maj_261_n29,
         maj_261_n28, maj_261_n27, maj_261_n26, maj_261_n25, maj_261_n24,
         maj_261_n23, maj_261_n22, maj_261_n21, maj_261_n20, maj_261_n19,
         maj_261_n18, maj_262_n34, maj_262_n33, maj_262_n32, maj_262_n31,
         maj_262_n30, maj_262_n29, maj_262_n28, maj_262_n27, maj_262_n26,
         maj_262_n25, maj_262_n24, maj_262_n23, maj_262_n22, maj_262_n21,
         maj_262_n20, maj_262_n19, maj_262_n18, maj_263_n34, maj_263_n33,
         maj_263_n32, maj_263_n31, maj_263_n30, maj_263_n29, maj_263_n28,
         maj_263_n27, maj_263_n26, maj_263_n25, maj_263_n24, maj_263_n23,
         maj_263_n22, maj_263_n21, maj_263_n20, maj_263_n19, maj_263_n18,
         maj_264_n34, maj_264_n33, maj_264_n32, maj_264_n31, maj_264_n30,
         maj_264_n29, maj_264_n28, maj_264_n27, maj_264_n26, maj_264_n25,
         maj_264_n24, maj_264_n23, maj_264_n22, maj_264_n21, maj_264_n20,
         maj_264_n19, maj_264_n18, maj_265_n34, maj_265_n33, maj_265_n32,
         maj_265_n31, maj_265_n30, maj_265_n29, maj_265_n28, maj_265_n27,
         maj_265_n26, maj_265_n25, maj_265_n24, maj_265_n23, maj_265_n22,
         maj_265_n21, maj_265_n20, maj_265_n19, maj_265_n18, maj_266_n34,
         maj_266_n33, maj_266_n32, maj_266_n31, maj_266_n30, maj_266_n29,
         maj_266_n28, maj_266_n27, maj_266_n26, maj_266_n25, maj_266_n24,
         maj_266_n23, maj_266_n22, maj_266_n21, maj_266_n20, maj_266_n19,
         maj_266_n18, maj_267_n34, maj_267_n33, maj_267_n32, maj_267_n31,
         maj_267_n30, maj_267_n29, maj_267_n28, maj_267_n27, maj_267_n26,
         maj_267_n25, maj_267_n24, maj_267_n23, maj_267_n22, maj_267_n21,
         maj_267_n20, maj_267_n19, maj_267_n18, maj_268_n34, maj_268_n33,
         maj_268_n32, maj_268_n31, maj_268_n30, maj_268_n29, maj_268_n28,
         maj_268_n27, maj_268_n26, maj_268_n25, maj_268_n24, maj_268_n23,
         maj_268_n22, maj_268_n21, maj_268_n20, maj_268_n19, maj_268_n18,
         maj_269_n34, maj_269_n33, maj_269_n32, maj_269_n31, maj_269_n30,
         maj_269_n29, maj_269_n28, maj_269_n27, maj_269_n26, maj_269_n25,
         maj_269_n24, maj_269_n23, maj_269_n22, maj_269_n21, maj_269_n20,
         maj_269_n19, maj_269_n18, maj_270_n34, maj_270_n33, maj_270_n32,
         maj_270_n31, maj_270_n30, maj_270_n29, maj_270_n28, maj_270_n27,
         maj_270_n26, maj_270_n25, maj_270_n24, maj_270_n23, maj_270_n22,
         maj_270_n21, maj_270_n20, maj_270_n19, maj_270_n18, maj_271_n34,
         maj_271_n33, maj_271_n32, maj_271_n31, maj_271_n30, maj_271_n29,
         maj_271_n28, maj_271_n27, maj_271_n26, maj_271_n25, maj_271_n24,
         maj_271_n23, maj_271_n22, maj_271_n21, maj_271_n20, maj_271_n19,
         maj_271_n18, maj_272_n34, maj_272_n33, maj_272_n32, maj_272_n31,
         maj_272_n30, maj_272_n29, maj_272_n28, maj_272_n27, maj_272_n26,
         maj_272_n25, maj_272_n24, maj_272_n23, maj_272_n22, maj_272_n21,
         maj_272_n20, maj_272_n19, maj_272_n18, maj_273_n34, maj_273_n33,
         maj_273_n32, maj_273_n31, maj_273_n30, maj_273_n29, maj_273_n28,
         maj_273_n27, maj_273_n26, maj_273_n25, maj_273_n24, maj_273_n23,
         maj_273_n22, maj_273_n21, maj_273_n20, maj_273_n19, maj_273_n18,
         maj_274_n34, maj_274_n33, maj_274_n32, maj_274_n31, maj_274_n30,
         maj_274_n29, maj_274_n28, maj_274_n27, maj_274_n26, maj_274_n25,
         maj_274_n24, maj_274_n23, maj_274_n22, maj_274_n21, maj_274_n20,
         maj_274_n19, maj_274_n18, maj_275_n34, maj_275_n33, maj_275_n32,
         maj_275_n31, maj_275_n30, maj_275_n29, maj_275_n28, maj_275_n27,
         maj_275_n26, maj_275_n25, maj_275_n24, maj_275_n23, maj_275_n22,
         maj_275_n21, maj_275_n20, maj_275_n19, maj_275_n18, maj_276_n34,
         maj_276_n33, maj_276_n32, maj_276_n31, maj_276_n30, maj_276_n29,
         maj_276_n28, maj_276_n27, maj_276_n26, maj_276_n25, maj_276_n24,
         maj_276_n23, maj_276_n22, maj_276_n21, maj_276_n20, maj_276_n19,
         maj_276_n18, maj_277_n34, maj_277_n33, maj_277_n32, maj_277_n31,
         maj_277_n30, maj_277_n29, maj_277_n28, maj_277_n27, maj_277_n26,
         maj_277_n25, maj_277_n24, maj_277_n23, maj_277_n22, maj_277_n21,
         maj_277_n20, maj_277_n19, maj_277_n18, maj_278_n34, maj_278_n33,
         maj_278_n32, maj_278_n31, maj_278_n30, maj_278_n29, maj_278_n28,
         maj_278_n27, maj_278_n26, maj_278_n25, maj_278_n24, maj_278_n23,
         maj_278_n22, maj_278_n21, maj_278_n20, maj_278_n19, maj_278_n18,
         maj_279_n34, maj_279_n33, maj_279_n32, maj_279_n31, maj_279_n30,
         maj_279_n29, maj_279_n28, maj_279_n27, maj_279_n26, maj_279_n25,
         maj_279_n24, maj_279_n23, maj_279_n22, maj_279_n21, maj_279_n20,
         maj_279_n19, maj_279_n18, maj_280_n34, maj_280_n33, maj_280_n32,
         maj_280_n31, maj_280_n30, maj_280_n29, maj_280_n28, maj_280_n27,
         maj_280_n26, maj_280_n25, maj_280_n24, maj_280_n23, maj_280_n22,
         maj_280_n21, maj_280_n20, maj_280_n19, maj_280_n18, maj_281_n34,
         maj_281_n33, maj_281_n32, maj_281_n31, maj_281_n30, maj_281_n29,
         maj_281_n28, maj_281_n27, maj_281_n26, maj_281_n25, maj_281_n24,
         maj_281_n23, maj_281_n22, maj_281_n21, maj_281_n20, maj_281_n19,
         maj_281_n18, maj_282_n34, maj_282_n33, maj_282_n32, maj_282_n31,
         maj_282_n30, maj_282_n29, maj_282_n28, maj_282_n27, maj_282_n26,
         maj_282_n25, maj_282_n24, maj_282_n23, maj_282_n22, maj_282_n21,
         maj_282_n20, maj_282_n19, maj_282_n18, maj_283_n34, maj_283_n33,
         maj_283_n32, maj_283_n31, maj_283_n30, maj_283_n29, maj_283_n28,
         maj_283_n27, maj_283_n26, maj_283_n25, maj_283_n24, maj_283_n23,
         maj_283_n22, maj_283_n21, maj_283_n20, maj_283_n19, maj_283_n18,
         maj_284_n34, maj_284_n33, maj_284_n32, maj_284_n31, maj_284_n30,
         maj_284_n29, maj_284_n28, maj_284_n27, maj_284_n26, maj_284_n25,
         maj_284_n24, maj_284_n23, maj_284_n22, maj_284_n21, maj_284_n20,
         maj_284_n19, maj_284_n18, maj_285_n34, maj_285_n33, maj_285_n32,
         maj_285_n31, maj_285_n30, maj_285_n29, maj_285_n28, maj_285_n27,
         maj_285_n26, maj_285_n25, maj_285_n24, maj_285_n23, maj_285_n22,
         maj_285_n21, maj_285_n20, maj_285_n19, maj_285_n18, maj_286_n34,
         maj_286_n33, maj_286_n32, maj_286_n31, maj_286_n30, maj_286_n29,
         maj_286_n28, maj_286_n27, maj_286_n26, maj_286_n25, maj_286_n24,
         maj_286_n23, maj_286_n22, maj_286_n21, maj_286_n20, maj_286_n19,
         maj_286_n18, maj_287_n34, maj_287_n33, maj_287_n32, maj_287_n31,
         maj_287_n30, maj_287_n29, maj_287_n28, maj_287_n27, maj_287_n26,
         maj_287_n25, maj_287_n24, maj_287_n23, maj_287_n22, maj_287_n21,
         maj_287_n20, maj_287_n19, maj_287_n18, maj_288_n34, maj_288_n33,
         maj_288_n32, maj_288_n31, maj_288_n30, maj_288_n29, maj_288_n28,
         maj_288_n27, maj_288_n26, maj_288_n25, maj_288_n24, maj_288_n23,
         maj_288_n22, maj_288_n21, maj_288_n20, maj_288_n19, maj_288_n18,
         maj_289_n34, maj_289_n33, maj_289_n32, maj_289_n31, maj_289_n30,
         maj_289_n29, maj_289_n28, maj_289_n27, maj_289_n26, maj_289_n25,
         maj_289_n24, maj_289_n23, maj_289_n22, maj_289_n21, maj_289_n20,
         maj_289_n19, maj_289_n18, maj_290_n34, maj_290_n33, maj_290_n32,
         maj_290_n31, maj_290_n30, maj_290_n29, maj_290_n28, maj_290_n27,
         maj_290_n26, maj_290_n25, maj_290_n24, maj_290_n23, maj_290_n22,
         maj_290_n21, maj_290_n20, maj_290_n19, maj_290_n18, maj_291_n34,
         maj_291_n33, maj_291_n32, maj_291_n31, maj_291_n30, maj_291_n29,
         maj_291_n28, maj_291_n27, maj_291_n26, maj_291_n25, maj_291_n24,
         maj_291_n23, maj_291_n22, maj_291_n21, maj_291_n20, maj_291_n19,
         maj_291_n18, maj_292_n34, maj_292_n33, maj_292_n32, maj_292_n31,
         maj_292_n30, maj_292_n29, maj_292_n28, maj_292_n27, maj_292_n26,
         maj_292_n25, maj_292_n24, maj_292_n23, maj_292_n22, maj_292_n21,
         maj_292_n20, maj_292_n19, maj_292_n18, maj_293_n34, maj_293_n33,
         maj_293_n32, maj_293_n31, maj_293_n30, maj_293_n29, maj_293_n28,
         maj_293_n27, maj_293_n26, maj_293_n25, maj_293_n24, maj_293_n23,
         maj_293_n22, maj_293_n21, maj_293_n20, maj_293_n19, maj_293_n18,
         maj_294_n34, maj_294_n33, maj_294_n32, maj_294_n31, maj_294_n30,
         maj_294_n29, maj_294_n28, maj_294_n27, maj_294_n26, maj_294_n25,
         maj_294_n24, maj_294_n23, maj_294_n22, maj_294_n21, maj_294_n20,
         maj_294_n19, maj_294_n18, maj_295_n34, maj_295_n33, maj_295_n32,
         maj_295_n31, maj_295_n30, maj_295_n29, maj_295_n28, maj_295_n27,
         maj_295_n26, maj_295_n25, maj_295_n24, maj_295_n23, maj_295_n22,
         maj_295_n21, maj_295_n20, maj_295_n19, maj_295_n18, maj_296_n34,
         maj_296_n33, maj_296_n32, maj_296_n31, maj_296_n30, maj_296_n29,
         maj_296_n28, maj_296_n27, maj_296_n26, maj_296_n25, maj_296_n24,
         maj_296_n23, maj_296_n22, maj_296_n21, maj_296_n20, maj_296_n19,
         maj_296_n18, maj_297_n34, maj_297_n33, maj_297_n32, maj_297_n31,
         maj_297_n30, maj_297_n29, maj_297_n28, maj_297_n27, maj_297_n26,
         maj_297_n25, maj_297_n24, maj_297_n23, maj_297_n22, maj_297_n21,
         maj_297_n20, maj_297_n19, maj_297_n18, maj_298_n34, maj_298_n33,
         maj_298_n32, maj_298_n31, maj_298_n30, maj_298_n29, maj_298_n28,
         maj_298_n27, maj_298_n26, maj_298_n25, maj_298_n24, maj_298_n23,
         maj_298_n22, maj_298_n21, maj_298_n20, maj_298_n19, maj_298_n18,
         maj_299_n34, maj_299_n33, maj_299_n32, maj_299_n31, maj_299_n30,
         maj_299_n29, maj_299_n28, maj_299_n27, maj_299_n26, maj_299_n25,
         maj_299_n24, maj_299_n23, maj_299_n22, maj_299_n21, maj_299_n20,
         maj_299_n19, maj_299_n18, maj_300_n34, maj_300_n33, maj_300_n32,
         maj_300_n31, maj_300_n30, maj_300_n29, maj_300_n28, maj_300_n27,
         maj_300_n26, maj_300_n25, maj_300_n24, maj_300_n23, maj_300_n22,
         maj_300_n21, maj_300_n20, maj_300_n19, maj_300_n18, maj_301_n34,
         maj_301_n33, maj_301_n32, maj_301_n31, maj_301_n30, maj_301_n29,
         maj_301_n28, maj_301_n27, maj_301_n26, maj_301_n25, maj_301_n24,
         maj_301_n23, maj_301_n22, maj_301_n21, maj_301_n20, maj_301_n19,
         maj_301_n18, maj_302_n34, maj_302_n33, maj_302_n32, maj_302_n31,
         maj_302_n30, maj_302_n29, maj_302_n28, maj_302_n27, maj_302_n26,
         maj_302_n25, maj_302_n24, maj_302_n23, maj_302_n22, maj_302_n21,
         maj_302_n20, maj_302_n19, maj_302_n18, maj_303_n34, maj_303_n33,
         maj_303_n32, maj_303_n31, maj_303_n30, maj_303_n29, maj_303_n28,
         maj_303_n27, maj_303_n26, maj_303_n25, maj_303_n24, maj_303_n23,
         maj_303_n22, maj_303_n21, maj_303_n20, maj_303_n19, maj_303_n18,
         maj_304_n34, maj_304_n33, maj_304_n32, maj_304_n31, maj_304_n30,
         maj_304_n29, maj_304_n28, maj_304_n27, maj_304_n26, maj_304_n25,
         maj_304_n24, maj_304_n23, maj_304_n22, maj_304_n21, maj_304_n20,
         maj_304_n19, maj_304_n18, maj_305_n34, maj_305_n33, maj_305_n32,
         maj_305_n31, maj_305_n30, maj_305_n29, maj_305_n28, maj_305_n27,
         maj_305_n26, maj_305_n25, maj_305_n24, maj_305_n23, maj_305_n22,
         maj_305_n21, maj_305_n20, maj_305_n19, maj_305_n18, maj_306_n34,
         maj_306_n33, maj_306_n32, maj_306_n31, maj_306_n30, maj_306_n29,
         maj_306_n28, maj_306_n27, maj_306_n26, maj_306_n25, maj_306_n24,
         maj_306_n23, maj_306_n22, maj_306_n21, maj_306_n20, maj_306_n19,
         maj_306_n18, maj_307_n34, maj_307_n33, maj_307_n32, maj_307_n31,
         maj_307_n30, maj_307_n29, maj_307_n28, maj_307_n27, maj_307_n26,
         maj_307_n25, maj_307_n24, maj_307_n23, maj_307_n22, maj_307_n21,
         maj_307_n20, maj_307_n19, maj_307_n18, maj_308_n34, maj_308_n33,
         maj_308_n32, maj_308_n31, maj_308_n30, maj_308_n29, maj_308_n28,
         maj_308_n27, maj_308_n26, maj_308_n25, maj_308_n24, maj_308_n23,
         maj_308_n22, maj_308_n21, maj_308_n20, maj_308_n19, maj_308_n18,
         maj_309_n34, maj_309_n33, maj_309_n32, maj_309_n31, maj_309_n30,
         maj_309_n29, maj_309_n28, maj_309_n27, maj_309_n26, maj_309_n25,
         maj_309_n24, maj_309_n23, maj_309_n22, maj_309_n21, maj_309_n20,
         maj_309_n19, maj_309_n18, maj_310_n34, maj_310_n33, maj_310_n32,
         maj_310_n31, maj_310_n30, maj_310_n29, maj_310_n28, maj_310_n27,
         maj_310_n26, maj_310_n25, maj_310_n24, maj_310_n23, maj_310_n22,
         maj_310_n21, maj_310_n20, maj_310_n19, maj_310_n18, maj_311_n34,
         maj_311_n33, maj_311_n32, maj_311_n31, maj_311_n30, maj_311_n29,
         maj_311_n28, maj_311_n27, maj_311_n26, maj_311_n25, maj_311_n24,
         maj_311_n23, maj_311_n22, maj_311_n21, maj_311_n20, maj_311_n19,
         maj_311_n18, maj_312_n34, maj_312_n33, maj_312_n32, maj_312_n31,
         maj_312_n30, maj_312_n29, maj_312_n28, maj_312_n27, maj_312_n26,
         maj_312_n25, maj_312_n24, maj_312_n23, maj_312_n22, maj_312_n21,
         maj_312_n20, maj_312_n19, maj_312_n18, maj_313_n34, maj_313_n33,
         maj_313_n32, maj_313_n31, maj_313_n30, maj_313_n29, maj_313_n28,
         maj_313_n27, maj_313_n26, maj_313_n25, maj_313_n24, maj_313_n23,
         maj_313_n22, maj_313_n21, maj_313_n20, maj_313_n19, maj_313_n18,
         maj_314_n34, maj_314_n33, maj_314_n32, maj_314_n31, maj_314_n30,
         maj_314_n29, maj_314_n28, maj_314_n27, maj_314_n26, maj_314_n25,
         maj_314_n24, maj_314_n23, maj_314_n22, maj_314_n21, maj_314_n20,
         maj_314_n19, maj_314_n18, maj_315_n34, maj_315_n33, maj_315_n32,
         maj_315_n31, maj_315_n30, maj_315_n29, maj_315_n28, maj_315_n27,
         maj_315_n26, maj_315_n25, maj_315_n24, maj_315_n23, maj_315_n22,
         maj_315_n21, maj_315_n20, maj_315_n19, maj_315_n18, maj_316_n34,
         maj_316_n33, maj_316_n32, maj_316_n31, maj_316_n30, maj_316_n29,
         maj_316_n28, maj_316_n27, maj_316_n26, maj_316_n25, maj_316_n24,
         maj_316_n23, maj_316_n22, maj_316_n21, maj_316_n20, maj_316_n19,
         maj_316_n18, maj_317_n34, maj_317_n33, maj_317_n32, maj_317_n31,
         maj_317_n30, maj_317_n29, maj_317_n28, maj_317_n27, maj_317_n26,
         maj_317_n25, maj_317_n24, maj_317_n23, maj_317_n22, maj_317_n21,
         maj_317_n20, maj_317_n19, maj_317_n18, maj_318_n34, maj_318_n33,
         maj_318_n32, maj_318_n31, maj_318_n30, maj_318_n29, maj_318_n28,
         maj_318_n27, maj_318_n26, maj_318_n25, maj_318_n24, maj_318_n23,
         maj_318_n22, maj_318_n21, maj_318_n20, maj_318_n19, maj_318_n18,
         maj_319_n34, maj_319_n33, maj_319_n32, maj_319_n31, maj_319_n30,
         maj_319_n29, maj_319_n28, maj_319_n27, maj_319_n26, maj_319_n25,
         maj_319_n24, maj_319_n23, maj_319_n22, maj_319_n21, maj_319_n20,
         maj_319_n19, maj_319_n18, maj_320_n34, maj_320_n33, maj_320_n32,
         maj_320_n31, maj_320_n30, maj_320_n29, maj_320_n28, maj_320_n27,
         maj_320_n26, maj_320_n25, maj_320_n24, maj_320_n23, maj_320_n22,
         maj_320_n21, maj_320_n20, maj_320_n19, maj_320_n18, maj_321_n34,
         maj_321_n33, maj_321_n32, maj_321_n31, maj_321_n30, maj_321_n29,
         maj_321_n28, maj_321_n27, maj_321_n26, maj_321_n25, maj_321_n24,
         maj_321_n23, maj_321_n22, maj_321_n21, maj_321_n20, maj_321_n19,
         maj_321_n18, maj_322_n34, maj_322_n33, maj_322_n32, maj_322_n31,
         maj_322_n30, maj_322_n29, maj_322_n28, maj_322_n27, maj_322_n26,
         maj_322_n25, maj_322_n24, maj_322_n23, maj_322_n22, maj_322_n21,
         maj_322_n20, maj_322_n19, maj_322_n18, maj_323_n34, maj_323_n33,
         maj_323_n32, maj_323_n31, maj_323_n30, maj_323_n29, maj_323_n28,
         maj_323_n27, maj_323_n26, maj_323_n25, maj_323_n24, maj_323_n23,
         maj_323_n22, maj_323_n21, maj_323_n20, maj_323_n19, maj_323_n18,
         maj_324_n34, maj_324_n33, maj_324_n32, maj_324_n31, maj_324_n30,
         maj_324_n29, maj_324_n28, maj_324_n27, maj_324_n26, maj_324_n25,
         maj_324_n24, maj_324_n23, maj_324_n22, maj_324_n21, maj_324_n20,
         maj_324_n19, maj_324_n18, maj_325_n34, maj_325_n33, maj_325_n32,
         maj_325_n31, maj_325_n30, maj_325_n29, maj_325_n28, maj_325_n27,
         maj_325_n26, maj_325_n25, maj_325_n24, maj_325_n23, maj_325_n22,
         maj_325_n21, maj_325_n20, maj_325_n19, maj_325_n18, maj_326_n34,
         maj_326_n33, maj_326_n32, maj_326_n31, maj_326_n30, maj_326_n29,
         maj_326_n28, maj_326_n27, maj_326_n26, maj_326_n25, maj_326_n24,
         maj_326_n23, maj_326_n22, maj_326_n21, maj_326_n20, maj_326_n19,
         maj_326_n18, maj_327_n34, maj_327_n33, maj_327_n32, maj_327_n31,
         maj_327_n30, maj_327_n29, maj_327_n28, maj_327_n27, maj_327_n26,
         maj_327_n25, maj_327_n24, maj_327_n23, maj_327_n22, maj_327_n21,
         maj_327_n20, maj_327_n19, maj_327_n18, maj_328_n34, maj_328_n33,
         maj_328_n32, maj_328_n31, maj_328_n30, maj_328_n29, maj_328_n28,
         maj_328_n27, maj_328_n26, maj_328_n25, maj_328_n24, maj_328_n23,
         maj_328_n22, maj_328_n21, maj_328_n20, maj_328_n19, maj_328_n18,
         maj_329_n34, maj_329_n33, maj_329_n32, maj_329_n31, maj_329_n30,
         maj_329_n29, maj_329_n28, maj_329_n27, maj_329_n26, maj_329_n25,
         maj_329_n24, maj_329_n23, maj_329_n22, maj_329_n21, maj_329_n20,
         maj_329_n19, maj_329_n18, maj_330_n34, maj_330_n33, maj_330_n32,
         maj_330_n31, maj_330_n30, maj_330_n29, maj_330_n28, maj_330_n27,
         maj_330_n26, maj_330_n25, maj_330_n24, maj_330_n23, maj_330_n22,
         maj_330_n21, maj_330_n20, maj_330_n19, maj_330_n18, maj_331_n34,
         maj_331_n33, maj_331_n32, maj_331_n31, maj_331_n30, maj_331_n29,
         maj_331_n28, maj_331_n27, maj_331_n26, maj_331_n25, maj_331_n24,
         maj_331_n23, maj_331_n22, maj_331_n21, maj_331_n20, maj_331_n19,
         maj_331_n18, maj_332_n34, maj_332_n33, maj_332_n32, maj_332_n31,
         maj_332_n30, maj_332_n29, maj_332_n28, maj_332_n27, maj_332_n26,
         maj_332_n25, maj_332_n24, maj_332_n23, maj_332_n22, maj_332_n21,
         maj_332_n20, maj_332_n19, maj_332_n18, maj_333_n34, maj_333_n33,
         maj_333_n32, maj_333_n31, maj_333_n30, maj_333_n29, maj_333_n28,
         maj_333_n27, maj_333_n26, maj_333_n25, maj_333_n24, maj_333_n23,
         maj_333_n22, maj_333_n21, maj_333_n20, maj_333_n19, maj_333_n18,
         maj_334_n34, maj_334_n33, maj_334_n32, maj_334_n31, maj_334_n30,
         maj_334_n29, maj_334_n28, maj_334_n27, maj_334_n26, maj_334_n25,
         maj_334_n24, maj_334_n23, maj_334_n22, maj_334_n21, maj_334_n20,
         maj_334_n19, maj_334_n18, maj_335_n34, maj_335_n33, maj_335_n32,
         maj_335_n31, maj_335_n30, maj_335_n29, maj_335_n28, maj_335_n27,
         maj_335_n26, maj_335_n25, maj_335_n24, maj_335_n23, maj_335_n22,
         maj_335_n21, maj_335_n20, maj_335_n19, maj_335_n18;
  wire   [6:0] u_0_0;
  wire   [6:0] v_0_0;
  wire   [6:0] u_0_1;
  wire   [6:0] v_0_1;
  wire   [6:0] u_0_2;
  wire   [6:0] v_0_2;
  wire   [6:0] u_1_0;
  wire   [6:0] v_1_0;
  wire   [6:0] u_1_1;
  wire   [6:0] v_1_1;
  wire   [6:0] u_1_2;
  wire   [6:0] v_1_2;
  wire   [6:0] u_2_0;
  wire   [6:0] v_2_0;
  wire   [6:0] u_2_1;
  wire   [6:0] v_2_1;
  wire   [6:0] u_2_2;
  wire   [6:0] v_2_2;
  wire   [6:0] u_3_0;
  wire   [6:0] v_3_0;
  wire   [6:0] u_3_1;
  wire   [6:0] v_3_1;
  wire   [6:0] u_3_2;
  wire   [6:0] v_3_2;
  wire   [6:0] temp_0_0;
  wire   [6:0] a_reg_0;
  wire   [6:0] v_reg_0_0;
  wire   [6:0] u_reg_0_0;
  wire   [6:0] v_reg_0_1;
  wire   [6:0] u_reg_0_1;
  wire   [6:0] v_reg_0_2;
  wire   [6:0] u_reg_0_2;
  wire   [6:0] temp_0_1;
  wire   [6:0] a_reg_1;
  wire   [6:0] v_reg_1_0;
  wire   [6:0] u_reg_1_0;
  wire   [6:0] v_reg_1_1;
  wire   [6:0] u_reg_1_1;
  wire   [6:0] v_reg_1_2;
  wire   [6:0] u_reg_1_2;
  wire   [6:0] temp_0_2;
  wire   [6:0] a_reg_2;
  wire   [6:0] v_reg_2_0;
  wire   [6:0] u_reg_2_0;
  wire   [6:0] v_reg_2_1;
  wire   [6:0] u_reg_2_1;
  wire   [6:0] v_reg_2_2;
  wire   [6:0] u_reg_2_2;
  wire   [6:0] temp_0_3;
  wire   [6:0] a_reg_3;
  wire   [6:0] v_reg_3_0;
  wire   [6:0] u_reg_3_0;
  wire   [6:0] v_reg_3_1;
  wire   [6:0] u_reg_3_1;
  wire   [6:0] v_reg_3_2;
  wire   [6:0] u_reg_3_2;

  DFF_X1 u_reg_0_0_reg_6_ ( .D(maj_312_port_o), .CK(clk), .Q(u_reg_0_0[6]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_5_ ( .D(maj_288_port_o), .CK(clk), .Q(u_reg_0_0[5]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_4_ ( .D(maj_264_port_o), .CK(clk), .Q(u_reg_0_0[4]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_3_ ( .D(maj_240_port_o), .CK(clk), .Q(u_reg_0_0[3]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_2_ ( .D(maj_216_port_o), .CK(clk), .Q(u_reg_0_0[2]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_1_ ( .D(maj_192_port_o), .CK(clk), .Q(u_reg_0_0[1]), 
        .QN() );
  DFF_X1 u_reg_0_0_reg_0_ ( .D(maj_168_port_o), .CK(clk), .Q(u_reg_0_0[0]), 
        .QN() );
  DFF_X1 a_reg_3_reg_6_ ( .D(port_a_3[6]), .CK(clk), .Q(a_reg_3[6]), .QN() );
  DFF_X1 a_reg_3_reg_5_ ( .D(port_a_3[5]), .CK(clk), .Q(a_reg_3[5]), .QN() );
  DFF_X1 a_reg_3_reg_4_ ( .D(port_a_3[4]), .CK(clk), .Q(a_reg_3[4]), .QN() );
  DFF_X1 a_reg_3_reg_3_ ( .D(port_a_3[3]), .CK(clk), .Q(a_reg_3[3]), .QN() );
  DFF_X1 a_reg_3_reg_2_ ( .D(port_a_3[2]), .CK(clk), .Q(a_reg_3[2]), .QN() );
  DFF_X1 a_reg_3_reg_1_ ( .D(port_a_3[1]), .CK(clk), .Q(a_reg_3[1]), .QN() );
  DFF_X1 a_reg_3_reg_0_ ( .D(port_a_3[0]), .CK(clk), .Q(a_reg_3[0]), .QN() );
  DFF_X1 v_reg_1_0_reg_6_ ( .D(maj_319_port_o), .CK(clk), .Q(v_reg_1_0[6]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_5_ ( .D(maj_295_port_o), .CK(clk), .Q(v_reg_1_0[5]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_4_ ( .D(maj_271_port_o), .CK(clk), .Q(v_reg_1_0[4]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_3_ ( .D(maj_247_port_o), .CK(clk), .Q(v_reg_1_0[3]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_2_ ( .D(maj_223_port_o), .CK(clk), .Q(v_reg_1_0[2]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_1_ ( .D(maj_199_port_o), .CK(clk), .Q(v_reg_1_0[1]), 
        .QN() );
  DFF_X1 v_reg_1_0_reg_0_ ( .D(maj_175_port_o), .CK(clk), .Q(v_reg_1_0[0]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_6_ ( .D(maj_314_port_o), .CK(clk), .Q(u_reg_0_1[6]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_5_ ( .D(maj_290_port_o), .CK(clk), .Q(u_reg_0_1[5]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_4_ ( .D(maj_266_port_o), .CK(clk), .Q(u_reg_0_1[4]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_3_ ( .D(maj_242_port_o), .CK(clk), .Q(u_reg_0_1[3]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_2_ ( .D(maj_218_port_o), .CK(clk), .Q(u_reg_0_1[2]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_1_ ( .D(maj_194_port_o), .CK(clk), .Q(u_reg_0_1[1]), 
        .QN() );
  DFF_X1 u_reg_0_1_reg_0_ ( .D(maj_170_port_o), .CK(clk), .Q(u_reg_0_1[0]), 
        .QN() );
  DFF_X1 ab_reg_3_reg_6_ ( .D(N27), .CK(clk), .Q(temp_0_3[6]), .QN() );
  DFF_X1 ab_reg_3_reg_5_ ( .D(N23), .CK(clk), .Q(temp_0_3[5]), .QN() );
  DFF_X1 ab_reg_3_reg_4_ ( .D(N19), .CK(clk), .Q(temp_0_3[4]), .QN() );
  DFF_X1 ab_reg_3_reg_3_ ( .D(N15), .CK(clk), .Q(temp_0_3[3]), .QN() );
  DFF_X1 ab_reg_3_reg_2_ ( .D(N11), .CK(clk), .Q(temp_0_3[2]), .QN() );
  DFF_X1 ab_reg_3_reg_1_ ( .D(N7), .CK(clk), .Q(temp_0_3[1]), .QN() );
  DFF_X1 ab_reg_3_reg_0_ ( .D(N3), .CK(clk), .Q(temp_0_3[0]), .QN() );
  DFF_X1 v_reg_0_2_reg_6_ ( .D(maj_317_port_o), .CK(clk), .Q(v_reg_0_2[6]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_5_ ( .D(maj_293_port_o), .CK(clk), .Q(v_reg_0_2[5]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_4_ ( .D(maj_269_port_o), .CK(clk), .Q(v_reg_0_2[4]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_3_ ( .D(maj_245_port_o), .CK(clk), .Q(v_reg_0_2[3]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_2_ ( .D(maj_221_port_o), .CK(clk), .Q(v_reg_0_2[2]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_1_ ( .D(maj_197_port_o), .CK(clk), .Q(v_reg_0_2[1]), 
        .QN() );
  DFF_X1 v_reg_0_2_reg_0_ ( .D(maj_173_port_o), .CK(clk), .Q(v_reg_0_2[0]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_6_ ( .D(maj_316_port_o), .CK(clk), .Q(u_reg_0_2[6]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_5_ ( .D(maj_292_port_o), .CK(clk), .Q(u_reg_0_2[5]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_4_ ( .D(maj_268_port_o), .CK(clk), .Q(u_reg_0_2[4]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_3_ ( .D(maj_244_port_o), .CK(clk), .Q(u_reg_0_2[3]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_2_ ( .D(maj_220_port_o), .CK(clk), .Q(u_reg_0_2[2]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_1_ ( .D(maj_196_port_o), .CK(clk), .Q(u_reg_0_2[1]), 
        .QN() );
  DFF_X1 u_reg_0_2_reg_0_ ( .D(maj_172_port_o), .CK(clk), .Q(u_reg_0_2[0]), 
        .QN() );
  DFF_X1 a_reg_2_reg_6_ ( .D(port_a_2[6]), .CK(clk), .Q(a_reg_2[6]), .QN() );
  DFF_X1 a_reg_2_reg_5_ ( .D(port_a_2[5]), .CK(clk), .Q(a_reg_2[5]), .QN() );
  DFF_X1 a_reg_2_reg_4_ ( .D(port_a_2[4]), .CK(clk), .Q(a_reg_2[4]), .QN() );
  DFF_X1 a_reg_2_reg_3_ ( .D(port_a_2[3]), .CK(clk), .Q(a_reg_2[3]), .QN() );
  DFF_X1 a_reg_2_reg_2_ ( .D(port_a_2[2]), .CK(clk), .Q(a_reg_2[2]), .QN() );
  DFF_X1 a_reg_2_reg_1_ ( .D(port_a_2[1]), .CK(clk), .Q(a_reg_2[1]), .QN() );
  DFF_X1 a_reg_2_reg_0_ ( .D(port_a_2[0]), .CK(clk), .Q(a_reg_2[0]), .QN() );
  DFF_X1 v_reg_0_1_reg_6_ ( .D(maj_315_port_o), .CK(clk), .Q(v_reg_0_1[6]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_5_ ( .D(maj_291_port_o), .CK(clk), .Q(v_reg_0_1[5]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_4_ ( .D(maj_267_port_o), .CK(clk), .Q(v_reg_0_1[4]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_3_ ( .D(maj_243_port_o), .CK(clk), .Q(v_reg_0_1[3]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_2_ ( .D(maj_219_port_o), .CK(clk), .Q(v_reg_0_1[2]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_1_ ( .D(maj_195_port_o), .CK(clk), .Q(v_reg_0_1[1]), 
        .QN() );
  DFF_X1 v_reg_0_1_reg_0_ ( .D(maj_171_port_o), .CK(clk), .Q(v_reg_0_1[0]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_6_ ( .D(maj_318_port_o), .CK(clk), .Q(u_reg_1_0[6]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_5_ ( .D(maj_294_port_o), .CK(clk), .Q(u_reg_1_0[5]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_4_ ( .D(maj_270_port_o), .CK(clk), .Q(u_reg_1_0[4]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_3_ ( .D(maj_246_port_o), .CK(clk), .Q(u_reg_1_0[3]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_2_ ( .D(maj_222_port_o), .CK(clk), .Q(u_reg_1_0[2]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_1_ ( .D(maj_198_port_o), .CK(clk), .Q(u_reg_1_0[1]), 
        .QN() );
  DFF_X1 u_reg_1_0_reg_0_ ( .D(maj_174_port_o), .CK(clk), .Q(u_reg_1_0[0]), 
        .QN() );
  DFF_X1 ab_reg_2_reg_6_ ( .D(N26), .CK(clk), .Q(temp_0_2[6]), .QN() );
  DFF_X1 ab_reg_2_reg_5_ ( .D(N22), .CK(clk), .Q(temp_0_2[5]), .QN() );
  DFF_X1 ab_reg_2_reg_4_ ( .D(N18), .CK(clk), .Q(temp_0_2[4]), .QN() );
  DFF_X1 ab_reg_2_reg_3_ ( .D(N14), .CK(clk), .Q(temp_0_2[3]), .QN() );
  DFF_X1 ab_reg_2_reg_2_ ( .D(N10), .CK(clk), .Q(temp_0_2[2]), .QN() );
  DFF_X1 ab_reg_2_reg_1_ ( .D(N6), .CK(clk), .Q(temp_0_2[1]), .QN() );
  DFF_X1 ab_reg_2_reg_0_ ( .D(N2), .CK(clk), .Q(temp_0_2[0]), .QN() );
  DFF_X1 v_reg_0_0_reg_6_ ( .D(maj_313_port_o), .CK(clk), .Q(v_reg_0_0[6]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_5_ ( .D(maj_289_port_o), .CK(clk), .Q(v_reg_0_0[5]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_4_ ( .D(maj_265_port_o), .CK(clk), .Q(v_reg_0_0[4]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_3_ ( .D(maj_241_port_o), .CK(clk), .Q(v_reg_0_0[3]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_2_ ( .D(maj_217_port_o), .CK(clk), .Q(v_reg_0_0[2]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_1_ ( .D(maj_193_port_o), .CK(clk), .Q(v_reg_0_0[1]), 
        .QN() );
  DFF_X1 v_reg_0_0_reg_0_ ( .D(maj_169_port_o), .CK(clk), .Q(v_reg_0_0[0]), 
        .QN() );
  DFF_X1 a_reg_1_reg_6_ ( .D(port_a_1[6]), .CK(clk), .Q(a_reg_1[6]), .QN() );
  DFF_X1 a_reg_1_reg_5_ ( .D(port_a_1[5]), .CK(clk), .Q(a_reg_1[5]), .QN() );
  DFF_X1 a_reg_1_reg_4_ ( .D(port_a_1[4]), .CK(clk), .Q(a_reg_1[4]), .QN() );
  DFF_X1 a_reg_1_reg_3_ ( .D(port_a_1[3]), .CK(clk), .Q(a_reg_1[3]), .QN() );
  DFF_X1 a_reg_1_reg_2_ ( .D(port_a_1[2]), .CK(clk), .Q(a_reg_1[2]), .QN() );
  DFF_X1 a_reg_1_reg_1_ ( .D(port_a_1[1]), .CK(clk), .Q(a_reg_1[1]), .QN() );
  DFF_X1 a_reg_1_reg_0_ ( .D(port_a_1[0]), .CK(clk), .Q(a_reg_1[0]), .QN() );
  DFF_X1 ab_reg_1_reg_6_ ( .D(N25), .CK(clk), .Q(temp_0_1[6]), .QN() );
  DFF_X1 ab_reg_1_reg_5_ ( .D(N21), .CK(clk), .Q(temp_0_1[5]), .QN() );
  DFF_X1 ab_reg_1_reg_4_ ( .D(N17), .CK(clk), .Q(temp_0_1[4]), .QN() );
  DFF_X1 ab_reg_1_reg_3_ ( .D(N13), .CK(clk), .Q(temp_0_1[3]), .QN() );
  DFF_X1 ab_reg_1_reg_2_ ( .D(N9), .CK(clk), .Q(temp_0_1[2]), .QN() );
  DFF_X1 ab_reg_1_reg_1_ ( .D(N5), .CK(clk), .Q(temp_0_1[1]), .QN() );
  DFF_X1 ab_reg_1_reg_0_ ( .D(N1), .CK(clk), .Q(temp_0_1[0]), .QN() );
  DFF_X1 a_reg_0_reg_6_ ( .D(port_a_0[6]), .CK(clk), .Q(a_reg_0[6]), .QN() );
  DFF_X1 a_reg_0_reg_5_ ( .D(port_a_0[5]), .CK(clk), .Q(a_reg_0[5]), .QN() );
  DFF_X1 a_reg_0_reg_4_ ( .D(port_a_0[4]), .CK(clk), .Q(a_reg_0[4]), .QN() );
  DFF_X1 a_reg_0_reg_3_ ( .D(port_a_0[3]), .CK(clk), .Q(a_reg_0[3]), .QN() );
  DFF_X1 a_reg_0_reg_2_ ( .D(port_a_0[2]), .CK(clk), .Q(a_reg_0[2]), .QN() );
  DFF_X1 a_reg_0_reg_1_ ( .D(port_a_0[1]), .CK(clk), .Q(a_reg_0[1]), .QN() );
  DFF_X1 a_reg_0_reg_0_ ( .D(port_a_0[0]), .CK(clk), .Q(a_reg_0[0]), .QN() );
  DFF_X1 ab_reg_0_reg_6_ ( .D(N24), .CK(clk), .Q(temp_0_0[6]), .QN() );
  DFF_X1 ab_reg_0_reg_5_ ( .D(N20), .CK(clk), .Q(temp_0_0[5]), .QN() );
  DFF_X1 ab_reg_0_reg_4_ ( .D(N16), .CK(clk), .Q(temp_0_0[4]), .QN() );
  DFF_X1 ab_reg_0_reg_3_ ( .D(N12), .CK(clk), .Q(temp_0_0[3]), .QN() );
  DFF_X1 ab_reg_0_reg_2_ ( .D(N8), .CK(clk), .Q(temp_0_0[2]), .QN() );
  DFF_X1 ab_reg_0_reg_1_ ( .D(N4), .CK(clk), .Q(temp_0_0[1]), .QN() );
  DFF_X1 ab_reg_0_reg_0_ ( .D(N0), .CK(clk), .Q(temp_0_0[0]), .QN() );
  DFF_X1 v_reg_3_2_reg_6_ ( .D(maj_335_port_o), .CK(clk), .Q(v_reg_3_2[6]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_5_ ( .D(maj_311_port_o), .CK(clk), .Q(v_reg_3_2[5]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_4_ ( .D(maj_287_port_o), .CK(clk), .Q(v_reg_3_2[4]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_3_ ( .D(maj_263_port_o), .CK(clk), .Q(v_reg_3_2[3]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_2_ ( .D(maj_239_port_o), .CK(clk), .Q(v_reg_3_2[2]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_1_ ( .D(maj_215_port_o), .CK(clk), .Q(v_reg_3_2[1]), 
        .QN() );
  DFF_X1 v_reg_3_2_reg_0_ ( .D(maj_191_port_o), .CK(clk), .Q(v_reg_3_2[0]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_6_ ( .D(maj_334_port_o), .CK(clk), .Q(u_reg_3_2[6]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_5_ ( .D(maj_310_port_o), .CK(clk), .Q(u_reg_3_2[5]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_4_ ( .D(maj_286_port_o), .CK(clk), .Q(u_reg_3_2[4]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_3_ ( .D(maj_262_port_o), .CK(clk), .Q(u_reg_3_2[3]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_2_ ( .D(maj_238_port_o), .CK(clk), .Q(u_reg_3_2[2]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_1_ ( .D(maj_214_port_o), .CK(clk), .Q(u_reg_3_2[1]), 
        .QN() );
  DFF_X1 u_reg_3_2_reg_0_ ( .D(maj_190_port_o), .CK(clk), .Q(u_reg_3_2[0]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_6_ ( .D(maj_333_port_o), .CK(clk), .Q(v_reg_3_1[6]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_5_ ( .D(maj_309_port_o), .CK(clk), .Q(v_reg_3_1[5]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_4_ ( .D(maj_285_port_o), .CK(clk), .Q(v_reg_3_1[4]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_3_ ( .D(maj_261_port_o), .CK(clk), .Q(v_reg_3_1[3]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_2_ ( .D(maj_237_port_o), .CK(clk), .Q(v_reg_3_1[2]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_1_ ( .D(maj_213_port_o), .CK(clk), .Q(v_reg_3_1[1]), 
        .QN() );
  DFF_X1 v_reg_3_1_reg_0_ ( .D(maj_189_port_o), .CK(clk), .Q(v_reg_3_1[0]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_6_ ( .D(maj_332_port_o), .CK(clk), .Q(u_reg_3_1[6]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_5_ ( .D(maj_308_port_o), .CK(clk), .Q(u_reg_3_1[5]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_4_ ( .D(maj_284_port_o), .CK(clk), .Q(u_reg_3_1[4]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_3_ ( .D(maj_260_port_o), .CK(clk), .Q(u_reg_3_1[3]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_2_ ( .D(maj_236_port_o), .CK(clk), .Q(u_reg_3_1[2]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_1_ ( .D(maj_212_port_o), .CK(clk), .Q(u_reg_3_1[1]), 
        .QN() );
  DFF_X1 u_reg_3_1_reg_0_ ( .D(maj_188_port_o), .CK(clk), .Q(u_reg_3_1[0]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_6_ ( .D(maj_331_port_o), .CK(clk), .Q(v_reg_3_0[6]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_5_ ( .D(maj_307_port_o), .CK(clk), .Q(v_reg_3_0[5]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_4_ ( .D(maj_283_port_o), .CK(clk), .Q(v_reg_3_0[4]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_3_ ( .D(maj_259_port_o), .CK(clk), .Q(v_reg_3_0[3]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_2_ ( .D(maj_235_port_o), .CK(clk), .Q(v_reg_3_0[2]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_1_ ( .D(maj_211_port_o), .CK(clk), .Q(v_reg_3_0[1]), 
        .QN() );
  DFF_X1 v_reg_3_0_reg_0_ ( .D(maj_187_port_o), .CK(clk), .Q(v_reg_3_0[0]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_6_ ( .D(maj_330_port_o), .CK(clk), .Q(u_reg_3_0[6]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_5_ ( .D(maj_306_port_o), .CK(clk), .Q(u_reg_3_0[5]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_4_ ( .D(maj_282_port_o), .CK(clk), .Q(u_reg_3_0[4]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_3_ ( .D(maj_258_port_o), .CK(clk), .Q(u_reg_3_0[3]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_2_ ( .D(maj_234_port_o), .CK(clk), .Q(u_reg_3_0[2]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_1_ ( .D(maj_210_port_o), .CK(clk), .Q(u_reg_3_0[1]), 
        .QN() );
  DFF_X1 u_reg_3_0_reg_0_ ( .D(maj_186_port_o), .CK(clk), .Q(u_reg_3_0[0]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_6_ ( .D(maj_329_port_o), .CK(clk), .Q(v_reg_2_2[6]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_5_ ( .D(maj_305_port_o), .CK(clk), .Q(v_reg_2_2[5]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_4_ ( .D(maj_281_port_o), .CK(clk), .Q(v_reg_2_2[4]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_3_ ( .D(maj_257_port_o), .CK(clk), .Q(v_reg_2_2[3]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_2_ ( .D(maj_233_port_o), .CK(clk), .Q(v_reg_2_2[2]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_1_ ( .D(maj_209_port_o), .CK(clk), .Q(v_reg_2_2[1]), 
        .QN() );
  DFF_X1 v_reg_2_2_reg_0_ ( .D(maj_185_port_o), .CK(clk), .Q(v_reg_2_2[0]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_6_ ( .D(maj_328_port_o), .CK(clk), .Q(u_reg_2_2[6]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_5_ ( .D(maj_304_port_o), .CK(clk), .Q(u_reg_2_2[5]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_4_ ( .D(maj_280_port_o), .CK(clk), .Q(u_reg_2_2[4]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_3_ ( .D(maj_256_port_o), .CK(clk), .Q(u_reg_2_2[3]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_2_ ( .D(maj_232_port_o), .CK(clk), .Q(u_reg_2_2[2]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_1_ ( .D(maj_208_port_o), .CK(clk), .Q(u_reg_2_2[1]), 
        .QN() );
  DFF_X1 u_reg_2_2_reg_0_ ( .D(maj_184_port_o), .CK(clk), .Q(u_reg_2_2[0]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_6_ ( .D(maj_327_port_o), .CK(clk), .Q(v_reg_2_1[6]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_5_ ( .D(maj_303_port_o), .CK(clk), .Q(v_reg_2_1[5]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_4_ ( .D(maj_279_port_o), .CK(clk), .Q(v_reg_2_1[4]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_3_ ( .D(maj_255_port_o), .CK(clk), .Q(v_reg_2_1[3]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_2_ ( .D(maj_231_port_o), .CK(clk), .Q(v_reg_2_1[2]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_1_ ( .D(maj_207_port_o), .CK(clk), .Q(v_reg_2_1[1]), 
        .QN() );
  DFF_X1 v_reg_2_1_reg_0_ ( .D(maj_183_port_o), .CK(clk), .Q(v_reg_2_1[0]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_6_ ( .D(maj_326_port_o), .CK(clk), .Q(u_reg_2_1[6]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_5_ ( .D(maj_302_port_o), .CK(clk), .Q(u_reg_2_1[5]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_4_ ( .D(maj_278_port_o), .CK(clk), .Q(u_reg_2_1[4]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_3_ ( .D(maj_254_port_o), .CK(clk), .Q(u_reg_2_1[3]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_2_ ( .D(maj_230_port_o), .CK(clk), .Q(u_reg_2_1[2]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_1_ ( .D(maj_206_port_o), .CK(clk), .Q(u_reg_2_1[1]), 
        .QN() );
  DFF_X1 u_reg_2_1_reg_0_ ( .D(maj_182_port_o), .CK(clk), .Q(u_reg_2_1[0]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_6_ ( .D(maj_325_port_o), .CK(clk), .Q(v_reg_2_0[6]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_5_ ( .D(maj_301_port_o), .CK(clk), .Q(v_reg_2_0[5]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_4_ ( .D(maj_277_port_o), .CK(clk), .Q(v_reg_2_0[4]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_3_ ( .D(maj_253_port_o), .CK(clk), .Q(v_reg_2_0[3]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_2_ ( .D(maj_229_port_o), .CK(clk), .Q(v_reg_2_0[2]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_1_ ( .D(maj_205_port_o), .CK(clk), .Q(v_reg_2_0[1]), 
        .QN() );
  DFF_X1 v_reg_2_0_reg_0_ ( .D(maj_181_port_o), .CK(clk), .Q(v_reg_2_0[0]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_6_ ( .D(maj_324_port_o), .CK(clk), .Q(u_reg_2_0[6]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_5_ ( .D(maj_300_port_o), .CK(clk), .Q(u_reg_2_0[5]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_4_ ( .D(maj_276_port_o), .CK(clk), .Q(u_reg_2_0[4]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_3_ ( .D(maj_252_port_o), .CK(clk), .Q(u_reg_2_0[3]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_2_ ( .D(maj_228_port_o), .CK(clk), .Q(u_reg_2_0[2]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_1_ ( .D(maj_204_port_o), .CK(clk), .Q(u_reg_2_0[1]), 
        .QN() );
  DFF_X1 u_reg_2_0_reg_0_ ( .D(maj_180_port_o), .CK(clk), .Q(u_reg_2_0[0]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_6_ ( .D(maj_323_port_o), .CK(clk), .Q(v_reg_1_2[6]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_5_ ( .D(maj_299_port_o), .CK(clk), .Q(v_reg_1_2[5]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_4_ ( .D(maj_275_port_o), .CK(clk), .Q(v_reg_1_2[4]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_3_ ( .D(maj_251_port_o), .CK(clk), .Q(v_reg_1_2[3]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_2_ ( .D(maj_227_port_o), .CK(clk), .Q(v_reg_1_2[2]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_1_ ( .D(maj_203_port_o), .CK(clk), .Q(v_reg_1_2[1]), 
        .QN() );
  DFF_X1 v_reg_1_2_reg_0_ ( .D(maj_179_port_o), .CK(clk), .Q(v_reg_1_2[0]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_6_ ( .D(maj_322_port_o), .CK(clk), .Q(u_reg_1_2[6]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_5_ ( .D(maj_298_port_o), .CK(clk), .Q(u_reg_1_2[5]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_4_ ( .D(maj_274_port_o), .CK(clk), .Q(u_reg_1_2[4]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_3_ ( .D(maj_250_port_o), .CK(clk), .Q(u_reg_1_2[3]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_2_ ( .D(maj_226_port_o), .CK(clk), .Q(u_reg_1_2[2]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_1_ ( .D(maj_202_port_o), .CK(clk), .Q(u_reg_1_2[1]), 
        .QN() );
  DFF_X1 u_reg_1_2_reg_0_ ( .D(maj_178_port_o), .CK(clk), .Q(u_reg_1_2[0]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_6_ ( .D(maj_321_port_o), .CK(clk), .Q(v_reg_1_1[6]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_5_ ( .D(maj_297_port_o), .CK(clk), .Q(v_reg_1_1[5]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_4_ ( .D(maj_273_port_o), .CK(clk), .Q(v_reg_1_1[4]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_3_ ( .D(maj_249_port_o), .CK(clk), .Q(v_reg_1_1[3]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_2_ ( .D(maj_225_port_o), .CK(clk), .Q(v_reg_1_1[2]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_1_ ( .D(maj_201_port_o), .CK(clk), .Q(v_reg_1_1[1]), 
        .QN() );
  DFF_X1 v_reg_1_1_reg_0_ ( .D(maj_177_port_o), .CK(clk), .Q(v_reg_1_1[0]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_6_ ( .D(maj_320_port_o), .CK(clk), .Q(u_reg_1_1[6]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_5_ ( .D(maj_296_port_o), .CK(clk), .Q(u_reg_1_1[5]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_4_ ( .D(maj_272_port_o), .CK(clk), .Q(u_reg_1_1[4]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_3_ ( .D(maj_248_port_o), .CK(clk), .Q(u_reg_1_1[3]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_2_ ( .D(maj_224_port_o), .CK(clk), .Q(u_reg_1_1[2]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_1_ ( .D(maj_200_port_o), .CK(clk), .Q(u_reg_1_1[1]), 
        .QN() );
  DFF_X1 u_reg_1_1_reg_0_ ( .D(maj_176_port_o), .CK(clk), .Q(u_reg_1_1[0]), 
        .QN() );
  XNOR2_X1 U311 ( .A(n81), .B(n82), .ZN(n80) );
  NAND2_X1 U312 ( .A1(v_reg_3_1[0]), .A2(a_reg_3[0]), .ZN(n81) );
  NAND2_X1 U313 ( .A1(v_reg_3_0[0]), .A2(a_reg_3[0]), .ZN(n82) );
  XNOR2_X1 U314 ( .A(n73), .B(n74), .ZN(n72) );
  NAND2_X1 U315 ( .A1(v_reg_3_1[1]), .A2(a_reg_3[1]), .ZN(n73) );
  NAND2_X1 U316 ( .A1(v_reg_3_0[1]), .A2(a_reg_3[1]), .ZN(n74) );
  XNOR2_X1 U317 ( .A(n65), .B(n66), .ZN(n64) );
  NAND2_X1 U318 ( .A1(v_reg_3_1[2]), .A2(a_reg_3[2]), .ZN(n65) );
  NAND2_X1 U319 ( .A1(v_reg_3_0[2]), .A2(a_reg_3[2]), .ZN(n66) );
  XNOR2_X1 U320 ( .A(n57), .B(n58), .ZN(n56) );
  NAND2_X1 U321 ( .A1(v_reg_3_1[3]), .A2(a_reg_3[3]), .ZN(n57) );
  NAND2_X1 U322 ( .A1(v_reg_3_0[3]), .A2(a_reg_3[3]), .ZN(n58) );
  XNOR2_X1 U323 ( .A(n49), .B(n50), .ZN(n48) );
  NAND2_X1 U324 ( .A1(v_reg_3_1[4]), .A2(a_reg_3[4]), .ZN(n49) );
  NAND2_X1 U325 ( .A1(v_reg_3_0[4]), .A2(a_reg_3[4]), .ZN(n50) );
  XNOR2_X1 U326 ( .A(n41), .B(n42), .ZN(n40) );
  NAND2_X1 U327 ( .A1(v_reg_3_1[5]), .A2(a_reg_3[5]), .ZN(n41) );
  NAND2_X1 U328 ( .A1(v_reg_3_0[5]), .A2(a_reg_3[5]), .ZN(n42) );
  XNOR2_X1 U329 ( .A(n33), .B(n34), .ZN(n32) );
  NAND2_X1 U330 ( .A1(v_reg_3_1[6]), .A2(a_reg_3[6]), .ZN(n33) );
  NAND2_X1 U331 ( .A1(v_reg_3_0[6]), .A2(a_reg_3[6]), .ZN(n34) );
  XNOR2_X1 U332 ( .A(n137), .B(n138), .ZN(n136) );
  NAND2_X1 U333 ( .A1(v_reg_2_1[0]), .A2(a_reg_2[0]), .ZN(n137) );
  NAND2_X1 U334 ( .A1(v_reg_2_0[0]), .A2(a_reg_2[0]), .ZN(n138) );
  XNOR2_X1 U335 ( .A(n129), .B(n130), .ZN(n128) );
  NAND2_X1 U336 ( .A1(v_reg_2_1[1]), .A2(a_reg_2[1]), .ZN(n129) );
  NAND2_X1 U337 ( .A1(v_reg_2_0[1]), .A2(a_reg_2[1]), .ZN(n130) );
  XNOR2_X1 U338 ( .A(n121), .B(n122), .ZN(n120) );
  NAND2_X1 U339 ( .A1(v_reg_2_1[2]), .A2(a_reg_2[2]), .ZN(n121) );
  NAND2_X1 U340 ( .A1(v_reg_2_0[2]), .A2(a_reg_2[2]), .ZN(n122) );
  XNOR2_X1 U341 ( .A(n113), .B(n114), .ZN(n112) );
  NAND2_X1 U342 ( .A1(v_reg_2_1[3]), .A2(a_reg_2[3]), .ZN(n113) );
  NAND2_X1 U343 ( .A1(v_reg_2_0[3]), .A2(a_reg_2[3]), .ZN(n114) );
  XNOR2_X1 U344 ( .A(n105), .B(n106), .ZN(n104) );
  NAND2_X1 U345 ( .A1(v_reg_2_1[4]), .A2(a_reg_2[4]), .ZN(n105) );
  NAND2_X1 U346 ( .A1(v_reg_2_0[4]), .A2(a_reg_2[4]), .ZN(n106) );
  XNOR2_X1 U347 ( .A(n97), .B(n98), .ZN(n96) );
  NAND2_X1 U348 ( .A1(v_reg_2_1[5]), .A2(a_reg_2[5]), .ZN(n97) );
  NAND2_X1 U349 ( .A1(v_reg_2_0[5]), .A2(a_reg_2[5]), .ZN(n98) );
  XNOR2_X1 U350 ( .A(n89), .B(n90), .ZN(n88) );
  NAND2_X1 U351 ( .A1(v_reg_2_1[6]), .A2(a_reg_2[6]), .ZN(n89) );
  NAND2_X1 U352 ( .A1(v_reg_2_0[6]), .A2(a_reg_2[6]), .ZN(n90) );
  XNOR2_X1 U353 ( .A(n193), .B(n194), .ZN(n192) );
  NAND2_X1 U354 ( .A1(v_reg_1_1[0]), .A2(a_reg_1[0]), .ZN(n193) );
  NAND2_X1 U355 ( .A1(v_reg_1_0[0]), .A2(a_reg_1[0]), .ZN(n194) );
  XNOR2_X1 U356 ( .A(n185), .B(n186), .ZN(n184) );
  NAND2_X1 U357 ( .A1(v_reg_1_1[1]), .A2(a_reg_1[1]), .ZN(n185) );
  NAND2_X1 U358 ( .A1(v_reg_1_0[1]), .A2(a_reg_1[1]), .ZN(n186) );
  XNOR2_X1 U359 ( .A(n177), .B(n178), .ZN(n176) );
  NAND2_X1 U360 ( .A1(v_reg_1_1[2]), .A2(a_reg_1[2]), .ZN(n177) );
  NAND2_X1 U361 ( .A1(v_reg_1_0[2]), .A2(a_reg_1[2]), .ZN(n178) );
  XNOR2_X1 U362 ( .A(n169), .B(n170), .ZN(n168) );
  NAND2_X1 U363 ( .A1(v_reg_1_1[3]), .A2(a_reg_1[3]), .ZN(n169) );
  NAND2_X1 U364 ( .A1(v_reg_1_0[3]), .A2(a_reg_1[3]), .ZN(n170) );
  XNOR2_X1 U365 ( .A(n161), .B(n162), .ZN(n160) );
  NAND2_X1 U366 ( .A1(v_reg_1_1[4]), .A2(a_reg_1[4]), .ZN(n161) );
  NAND2_X1 U367 ( .A1(v_reg_1_0[4]), .A2(a_reg_1[4]), .ZN(n162) );
  XNOR2_X1 U368 ( .A(n153), .B(n154), .ZN(n152) );
  NAND2_X1 U369 ( .A1(v_reg_1_1[5]), .A2(a_reg_1[5]), .ZN(n153) );
  NAND2_X1 U370 ( .A1(v_reg_1_0[5]), .A2(a_reg_1[5]), .ZN(n154) );
  XNOR2_X1 U371 ( .A(n145), .B(n146), .ZN(n144) );
  NAND2_X1 U372 ( .A1(v_reg_1_1[6]), .A2(a_reg_1[6]), .ZN(n145) );
  NAND2_X1 U373 ( .A1(v_reg_1_0[6]), .A2(a_reg_1[6]), .ZN(n146) );
  XNOR2_X1 U374 ( .A(n249), .B(n250), .ZN(n248) );
  NAND2_X1 U375 ( .A1(v_reg_0_1[0]), .A2(a_reg_0[0]), .ZN(n249) );
  NAND2_X1 U376 ( .A1(v_reg_0_0[0]), .A2(a_reg_0[0]), .ZN(n250) );
  XNOR2_X1 U377 ( .A(n241), .B(n242), .ZN(n240) );
  NAND2_X1 U378 ( .A1(v_reg_0_1[1]), .A2(a_reg_0[1]), .ZN(n241) );
  NAND2_X1 U379 ( .A1(v_reg_0_0[1]), .A2(a_reg_0[1]), .ZN(n242) );
  XNOR2_X1 U380 ( .A(n233), .B(n234), .ZN(n232) );
  NAND2_X1 U381 ( .A1(v_reg_0_1[2]), .A2(a_reg_0[2]), .ZN(n233) );
  NAND2_X1 U382 ( .A1(v_reg_0_0[2]), .A2(a_reg_0[2]), .ZN(n234) );
  XNOR2_X1 U383 ( .A(n225), .B(n226), .ZN(n224) );
  NAND2_X1 U384 ( .A1(v_reg_0_1[3]), .A2(a_reg_0[3]), .ZN(n225) );
  NAND2_X1 U385 ( .A1(v_reg_0_0[3]), .A2(a_reg_0[3]), .ZN(n226) );
  XNOR2_X1 U386 ( .A(n217), .B(n218), .ZN(n216) );
  NAND2_X1 U387 ( .A1(v_reg_0_1[4]), .A2(a_reg_0[4]), .ZN(n217) );
  NAND2_X1 U388 ( .A1(v_reg_0_0[4]), .A2(a_reg_0[4]), .ZN(n218) );
  XNOR2_X1 U389 ( .A(n209), .B(n210), .ZN(n208) );
  NAND2_X1 U390 ( .A1(v_reg_0_1[5]), .A2(a_reg_0[5]), .ZN(n209) );
  NAND2_X1 U391 ( .A1(v_reg_0_0[5]), .A2(a_reg_0[5]), .ZN(n210) );
  XNOR2_X1 U392 ( .A(n201), .B(n202), .ZN(n200) );
  NAND2_X1 U393 ( .A1(v_reg_0_1[6]), .A2(a_reg_0[6]), .ZN(n201) );
  NAND2_X1 U394 ( .A1(v_reg_0_0[6]), .A2(a_reg_0[6]), .ZN(n202) );
  XNOR2_X1 U395 ( .A(u_reg_3_0[0]), .B(temp_0_3[0]), .ZN(n84) );
  XNOR2_X1 U396 ( .A(u_reg_3_0[1]), .B(temp_0_3[1]), .ZN(n76) );
  XNOR2_X1 U397 ( .A(u_reg_3_0[2]), .B(temp_0_3[2]), .ZN(n68) );
  XNOR2_X1 U398 ( .A(u_reg_3_0[3]), .B(temp_0_3[3]), .ZN(n60) );
  XNOR2_X1 U399 ( .A(u_reg_3_0[4]), .B(temp_0_3[4]), .ZN(n52) );
  XNOR2_X1 U400 ( .A(u_reg_3_0[5]), .B(temp_0_3[5]), .ZN(n44) );
  XNOR2_X1 U401 ( .A(u_reg_3_0[6]), .B(temp_0_3[6]), .ZN(n36) );
  XNOR2_X1 U402 ( .A(u_reg_2_0[0]), .B(temp_0_2[0]), .ZN(n140) );
  XNOR2_X1 U403 ( .A(u_reg_2_0[1]), .B(temp_0_2[1]), .ZN(n132) );
  XNOR2_X1 U404 ( .A(u_reg_2_0[2]), .B(temp_0_2[2]), .ZN(n124) );
  XNOR2_X1 U405 ( .A(u_reg_2_0[3]), .B(temp_0_2[3]), .ZN(n116) );
  XNOR2_X1 U406 ( .A(u_reg_2_0[4]), .B(temp_0_2[4]), .ZN(n108) );
  XNOR2_X1 U407 ( .A(u_reg_2_0[5]), .B(temp_0_2[5]), .ZN(n100) );
  XNOR2_X1 U408 ( .A(u_reg_2_0[6]), .B(temp_0_2[6]), .ZN(n92) );
  XNOR2_X1 U409 ( .A(u_reg_1_0[0]), .B(temp_0_1[0]), .ZN(n196) );
  XNOR2_X1 U410 ( .A(u_reg_1_0[1]), .B(temp_0_1[1]), .ZN(n188) );
  XNOR2_X1 U411 ( .A(u_reg_1_0[2]), .B(temp_0_1[2]), .ZN(n180) );
  XNOR2_X1 U412 ( .A(u_reg_1_0[3]), .B(temp_0_1[3]), .ZN(n172) );
  XNOR2_X1 U413 ( .A(u_reg_1_0[4]), .B(temp_0_1[4]), .ZN(n164) );
  XNOR2_X1 U414 ( .A(u_reg_1_0[5]), .B(temp_0_1[5]), .ZN(n156) );
  XNOR2_X1 U415 ( .A(u_reg_1_0[6]), .B(temp_0_1[6]), .ZN(n148) );
  XNOR2_X1 U416 ( .A(u_reg_0_0[0]), .B(temp_0_0[0]), .ZN(n252) );
  XNOR2_X1 U417 ( .A(u_reg_0_0[1]), .B(temp_0_0[1]), .ZN(n244) );
  XNOR2_X1 U418 ( .A(u_reg_0_0[2]), .B(temp_0_0[2]), .ZN(n236) );
  XNOR2_X1 U419 ( .A(u_reg_0_0[3]), .B(temp_0_0[3]), .ZN(n228) );
  XNOR2_X1 U420 ( .A(u_reg_0_0[4]), .B(temp_0_0[4]), .ZN(n220) );
  XNOR2_X1 U421 ( .A(u_reg_0_0[5]), .B(temp_0_0[5]), .ZN(n212) );
  XNOR2_X1 U422 ( .A(u_reg_0_0[6]), .B(temp_0_0[6]), .ZN(n204) );
  INV_X1 U423 ( .A(port_a_2[2]), .ZN(n19) );
  INV_X1 U424 ( .A(port_a_2[1]), .ZN(n20) );
  INV_X1 U425 ( .A(port_a_2[0]), .ZN(n21) );
  INV_X1 U426 ( .A(port_a_2[5]), .ZN(n16) );
  INV_X1 U427 ( .A(port_a_2[4]), .ZN(n17) );
  INV_X1 U428 ( .A(port_a_2[3]), .ZN(n18) );
  INV_X1 U429 ( .A(port_a_2[6]), .ZN(n15) );
  INV_X1 U430 ( .A(port_a_3[2]), .ZN(n26) );
  INV_X1 U431 ( .A(port_a_3[1]), .ZN(n27) );
  INV_X1 U432 ( .A(port_a_3[0]), .ZN(n28) );
  INV_X1 U433 ( .A(port_a_3[5]), .ZN(n23) );
  INV_X1 U434 ( .A(port_a_3[4]), .ZN(n24) );
  INV_X1 U435 ( .A(port_a_3[3]), .ZN(n25) );
  INV_X1 U436 ( .A(port_a_3[6]), .ZN(n22) );
  INV_X1 U437 ( .A(port_a_1[2]), .ZN(n12) );
  INV_X1 U438 ( .A(port_a_1[1]), .ZN(n13) );
  INV_X1 U439 ( .A(port_a_1[0]), .ZN(n14) );
  INV_X1 U440 ( .A(port_a_1[5]), .ZN(n9) );
  INV_X1 U441 ( .A(port_a_1[4]), .ZN(n10) );
  INV_X1 U442 ( .A(port_a_1[3]), .ZN(n11) );
  INV_X1 U443 ( .A(port_a_1[6]), .ZN(n8) );
  INV_X1 U444 ( .A(port_a_0[2]), .ZN(n5) );
  INV_X1 U445 ( .A(port_a_0[1]), .ZN(n6) );
  INV_X1 U446 ( .A(port_a_0[0]), .ZN(n7) );
  INV_X1 U447 ( .A(port_a_0[5]), .ZN(n2) );
  INV_X1 U448 ( .A(port_a_0[4]), .ZN(n3) );
  INV_X1 U449 ( .A(port_a_0[3]), .ZN(n4) );
  INV_X1 U450 ( .A(port_a_0[6]), .ZN(n1) );
  XOR2_X1 U451 ( .A(n77), .B(n78), .Z(port_c_3[0]) );
  XOR2_X1 U452 ( .A(n83), .B(n84), .Z(n77) );
  XOR2_X1 U453 ( .A(n79), .B(n80), .Z(n78) );
  XNOR2_X1 U454 ( .A(u_reg_3_2[0]), .B(u_reg_3_1[0]), .ZN(n83) );
  XOR2_X1 U455 ( .A(n69), .B(n70), .Z(port_c_3[1]) );
  XOR2_X1 U456 ( .A(n75), .B(n76), .Z(n69) );
  XOR2_X1 U457 ( .A(n71), .B(n72), .Z(n70) );
  XNOR2_X1 U458 ( .A(u_reg_3_2[1]), .B(u_reg_3_1[1]), .ZN(n75) );
  XOR2_X1 U459 ( .A(n61), .B(n62), .Z(port_c_3[2]) );
  XOR2_X1 U460 ( .A(n67), .B(n68), .Z(n61) );
  XOR2_X1 U461 ( .A(n63), .B(n64), .Z(n62) );
  XNOR2_X1 U462 ( .A(u_reg_3_2[2]), .B(u_reg_3_1[2]), .ZN(n67) );
  XOR2_X1 U463 ( .A(n53), .B(n54), .Z(port_c_3[3]) );
  XOR2_X1 U464 ( .A(n59), .B(n60), .Z(n53) );
  XOR2_X1 U465 ( .A(n55), .B(n56), .Z(n54) );
  XNOR2_X1 U466 ( .A(u_reg_3_2[3]), .B(u_reg_3_1[3]), .ZN(n59) );
  XOR2_X1 U467 ( .A(n45), .B(n46), .Z(port_c_3[4]) );
  XOR2_X1 U468 ( .A(n51), .B(n52), .Z(n45) );
  XOR2_X1 U469 ( .A(n47), .B(n48), .Z(n46) );
  XNOR2_X1 U470 ( .A(u_reg_3_2[4]), .B(u_reg_3_1[4]), .ZN(n51) );
  XOR2_X1 U471 ( .A(n37), .B(n38), .Z(port_c_3[5]) );
  XOR2_X1 U472 ( .A(n43), .B(n44), .Z(n37) );
  XOR2_X1 U473 ( .A(n39), .B(n40), .Z(n38) );
  XNOR2_X1 U474 ( .A(u_reg_3_2[5]), .B(u_reg_3_1[5]), .ZN(n43) );
  XOR2_X1 U475 ( .A(n29), .B(n30), .Z(port_c_3[6]) );
  XOR2_X1 U476 ( .A(n35), .B(n36), .Z(n29) );
  XOR2_X1 U477 ( .A(n31), .B(n32), .Z(n30) );
  XNOR2_X1 U478 ( .A(u_reg_3_2[6]), .B(u_reg_3_1[6]), .ZN(n35) );
  XOR2_X1 U479 ( .A(n133), .B(n134), .Z(port_c_2[0]) );
  XOR2_X1 U480 ( .A(n139), .B(n140), .Z(n133) );
  XOR2_X1 U481 ( .A(n135), .B(n136), .Z(n134) );
  XNOR2_X1 U482 ( .A(u_reg_2_2[0]), .B(u_reg_2_1[0]), .ZN(n139) );
  XOR2_X1 U483 ( .A(n125), .B(n126), .Z(port_c_2[1]) );
  XOR2_X1 U484 ( .A(n131), .B(n132), .Z(n125) );
  XOR2_X1 U485 ( .A(n127), .B(n128), .Z(n126) );
  XNOR2_X1 U486 ( .A(u_reg_2_2[1]), .B(u_reg_2_1[1]), .ZN(n131) );
  XOR2_X1 U487 ( .A(n117), .B(n118), .Z(port_c_2[2]) );
  XOR2_X1 U488 ( .A(n123), .B(n124), .Z(n117) );
  XOR2_X1 U489 ( .A(n119), .B(n120), .Z(n118) );
  XNOR2_X1 U490 ( .A(u_reg_2_2[2]), .B(u_reg_2_1[2]), .ZN(n123) );
  XOR2_X1 U491 ( .A(n109), .B(n110), .Z(port_c_2[3]) );
  XOR2_X1 U492 ( .A(n115), .B(n116), .Z(n109) );
  XOR2_X1 U493 ( .A(n111), .B(n112), .Z(n110) );
  XNOR2_X1 U494 ( .A(u_reg_2_2[3]), .B(u_reg_2_1[3]), .ZN(n115) );
  XOR2_X1 U495 ( .A(n101), .B(n102), .Z(port_c_2[4]) );
  XOR2_X1 U496 ( .A(n107), .B(n108), .Z(n101) );
  XOR2_X1 U497 ( .A(n103), .B(n104), .Z(n102) );
  XNOR2_X1 U498 ( .A(u_reg_2_2[4]), .B(u_reg_2_1[4]), .ZN(n107) );
  XOR2_X1 U499 ( .A(n93), .B(n94), .Z(port_c_2[5]) );
  XOR2_X1 U500 ( .A(n99), .B(n100), .Z(n93) );
  XOR2_X1 U501 ( .A(n95), .B(n96), .Z(n94) );
  XNOR2_X1 U502 ( .A(u_reg_2_2[5]), .B(u_reg_2_1[5]), .ZN(n99) );
  XOR2_X1 U503 ( .A(n85), .B(n86), .Z(port_c_2[6]) );
  XOR2_X1 U504 ( .A(n91), .B(n92), .Z(n85) );
  XOR2_X1 U505 ( .A(n87), .B(n88), .Z(n86) );
  XNOR2_X1 U506 ( .A(u_reg_2_2[6]), .B(u_reg_2_1[6]), .ZN(n91) );
  XOR2_X1 U507 ( .A(n189), .B(n190), .Z(port_c_1[0]) );
  XOR2_X1 U508 ( .A(n195), .B(n196), .Z(n189) );
  XOR2_X1 U509 ( .A(n191), .B(n192), .Z(n190) );
  XNOR2_X1 U510 ( .A(u_reg_1_2[0]), .B(u_reg_1_1[0]), .ZN(n195) );
  XOR2_X1 U511 ( .A(n181), .B(n182), .Z(port_c_1[1]) );
  XOR2_X1 U512 ( .A(n187), .B(n188), .Z(n181) );
  XOR2_X1 U513 ( .A(n183), .B(n184), .Z(n182) );
  XNOR2_X1 U514 ( .A(u_reg_1_2[1]), .B(u_reg_1_1[1]), .ZN(n187) );
  XOR2_X1 U515 ( .A(n173), .B(n174), .Z(port_c_1[2]) );
  XOR2_X1 U516 ( .A(n179), .B(n180), .Z(n173) );
  XOR2_X1 U517 ( .A(n175), .B(n176), .Z(n174) );
  XNOR2_X1 U518 ( .A(u_reg_1_2[2]), .B(u_reg_1_1[2]), .ZN(n179) );
  XOR2_X1 U519 ( .A(n165), .B(n166), .Z(port_c_1[3]) );
  XOR2_X1 U520 ( .A(n171), .B(n172), .Z(n165) );
  XOR2_X1 U521 ( .A(n167), .B(n168), .Z(n166) );
  XNOR2_X1 U522 ( .A(u_reg_1_2[3]), .B(u_reg_1_1[3]), .ZN(n171) );
  XOR2_X1 U523 ( .A(n157), .B(n158), .Z(port_c_1[4]) );
  XOR2_X1 U524 ( .A(n163), .B(n164), .Z(n157) );
  XOR2_X1 U525 ( .A(n159), .B(n160), .Z(n158) );
  XNOR2_X1 U526 ( .A(u_reg_1_2[4]), .B(u_reg_1_1[4]), .ZN(n163) );
  XOR2_X1 U527 ( .A(n149), .B(n150), .Z(port_c_1[5]) );
  XOR2_X1 U528 ( .A(n155), .B(n156), .Z(n149) );
  XOR2_X1 U529 ( .A(n151), .B(n152), .Z(n150) );
  XNOR2_X1 U530 ( .A(u_reg_1_2[5]), .B(u_reg_1_1[5]), .ZN(n155) );
  XOR2_X1 U531 ( .A(n141), .B(n142), .Z(port_c_1[6]) );
  XOR2_X1 U532 ( .A(n147), .B(n148), .Z(n141) );
  XOR2_X1 U533 ( .A(n143), .B(n144), .Z(n142) );
  XNOR2_X1 U534 ( .A(u_reg_1_2[6]), .B(u_reg_1_1[6]), .ZN(n147) );
  XOR2_X1 U535 ( .A(n245), .B(n246), .Z(port_c_0[0]) );
  XOR2_X1 U536 ( .A(n251), .B(n252), .Z(n245) );
  XOR2_X1 U537 ( .A(n247), .B(n248), .Z(n246) );
  XNOR2_X1 U538 ( .A(u_reg_0_2[0]), .B(u_reg_0_1[0]), .ZN(n251) );
  XOR2_X1 U539 ( .A(n237), .B(n238), .Z(port_c_0[1]) );
  XOR2_X1 U540 ( .A(n243), .B(n244), .Z(n237) );
  XOR2_X1 U541 ( .A(n239), .B(n240), .Z(n238) );
  XNOR2_X1 U542 ( .A(u_reg_0_2[1]), .B(u_reg_0_1[1]), .ZN(n243) );
  XOR2_X1 U543 ( .A(n229), .B(n230), .Z(port_c_0[2]) );
  XOR2_X1 U544 ( .A(n235), .B(n236), .Z(n229) );
  XOR2_X1 U545 ( .A(n231), .B(n232), .Z(n230) );
  XNOR2_X1 U546 ( .A(u_reg_0_2[2]), .B(u_reg_0_1[2]), .ZN(n235) );
  XOR2_X1 U547 ( .A(n221), .B(n222), .Z(port_c_0[3]) );
  XOR2_X1 U548 ( .A(n227), .B(n228), .Z(n221) );
  XOR2_X1 U549 ( .A(n223), .B(n224), .Z(n222) );
  XNOR2_X1 U550 ( .A(u_reg_0_2[3]), .B(u_reg_0_1[3]), .ZN(n227) );
  XOR2_X1 U551 ( .A(n213), .B(n214), .Z(port_c_0[4]) );
  XOR2_X1 U552 ( .A(n219), .B(n220), .Z(n213) );
  XOR2_X1 U553 ( .A(n215), .B(n216), .Z(n214) );
  XNOR2_X1 U554 ( .A(u_reg_0_2[4]), .B(u_reg_0_1[4]), .ZN(n219) );
  XOR2_X1 U555 ( .A(n205), .B(n206), .Z(port_c_0[5]) );
  XOR2_X1 U556 ( .A(n211), .B(n212), .Z(n205) );
  XOR2_X1 U557 ( .A(n207), .B(n208), .Z(n206) );
  XNOR2_X1 U558 ( .A(u_reg_0_2[5]), .B(u_reg_0_1[5]), .ZN(n211) );
  XOR2_X1 U559 ( .A(n197), .B(n198), .Z(port_c_0[6]) );
  XOR2_X1 U560 ( .A(n203), .B(n204), .Z(n197) );
  XOR2_X1 U561 ( .A(n199), .B(n200), .Z(n198) );
  XNOR2_X1 U562 ( .A(u_reg_0_2[6]), .B(u_reg_0_1[6]), .ZN(n203) );
  NAND2_X1 U563 ( .A1(v_reg_3_2[0]), .A2(a_reg_3[0]), .ZN(n79) );
  NAND2_X1 U564 ( .A1(v_reg_3_2[1]), .A2(a_reg_3[1]), .ZN(n71) );
  NAND2_X1 U565 ( .A1(v_reg_3_2[2]), .A2(a_reg_3[2]), .ZN(n63) );
  NAND2_X1 U566 ( .A1(v_reg_3_2[3]), .A2(a_reg_3[3]), .ZN(n55) );
  NAND2_X1 U567 ( .A1(v_reg_3_2[4]), .A2(a_reg_3[4]), .ZN(n47) );
  NAND2_X1 U568 ( .A1(v_reg_3_2[5]), .A2(a_reg_3[5]), .ZN(n39) );
  NAND2_X1 U569 ( .A1(v_reg_3_2[6]), .A2(a_reg_3[6]), .ZN(n31) );
  NAND2_X1 U570 ( .A1(v_reg_2_2[0]), .A2(a_reg_2[0]), .ZN(n135) );
  NAND2_X1 U571 ( .A1(v_reg_2_2[1]), .A2(a_reg_2[1]), .ZN(n127) );
  NAND2_X1 U572 ( .A1(v_reg_2_2[2]), .A2(a_reg_2[2]), .ZN(n119) );
  NAND2_X1 U573 ( .A1(v_reg_2_2[3]), .A2(a_reg_2[3]), .ZN(n111) );
  NAND2_X1 U574 ( .A1(v_reg_2_2[4]), .A2(a_reg_2[4]), .ZN(n103) );
  NAND2_X1 U575 ( .A1(v_reg_2_2[5]), .A2(a_reg_2[5]), .ZN(n95) );
  NAND2_X1 U576 ( .A1(v_reg_2_2[6]), .A2(a_reg_2[6]), .ZN(n87) );
  NAND2_X1 U577 ( .A1(v_reg_1_2[0]), .A2(a_reg_1[0]), .ZN(n191) );
  NAND2_X1 U578 ( .A1(v_reg_1_2[1]), .A2(a_reg_1[1]), .ZN(n183) );
  NAND2_X1 U579 ( .A1(v_reg_1_2[2]), .A2(a_reg_1[2]), .ZN(n175) );
  NAND2_X1 U580 ( .A1(v_reg_1_2[3]), .A2(a_reg_1[3]), .ZN(n167) );
  NAND2_X1 U581 ( .A1(v_reg_1_2[4]), .A2(a_reg_1[4]), .ZN(n159) );
  NAND2_X1 U582 ( .A1(v_reg_1_2[5]), .A2(a_reg_1[5]), .ZN(n151) );
  NAND2_X1 U583 ( .A1(v_reg_1_2[6]), .A2(a_reg_1[6]), .ZN(n143) );
  NAND2_X1 U584 ( .A1(v_reg_0_2[0]), .A2(a_reg_0[0]), .ZN(n247) );
  NAND2_X1 U585 ( .A1(v_reg_0_2[1]), .A2(a_reg_0[1]), .ZN(n239) );
  NAND2_X1 U586 ( .A1(v_reg_0_2[2]), .A2(a_reg_0[2]), .ZN(n231) );
  NAND2_X1 U587 ( .A1(v_reg_0_2[3]), .A2(a_reg_0[3]), .ZN(n223) );
  NAND2_X1 U588 ( .A1(v_reg_0_2[4]), .A2(a_reg_0[4]), .ZN(n215) );
  NAND2_X1 U589 ( .A1(v_reg_0_2[5]), .A2(a_reg_0[5]), .ZN(n207) );
  NAND2_X1 U590 ( .A1(v_reg_0_2[6]), .A2(a_reg_0[6]), .ZN(n199) );
  AND2_X1 U591 ( .A1(port_b_0[0]), .A2(port_a_0[0]), .ZN(N0) );
  AND2_X1 U592 ( .A1(port_b_0[1]), .A2(port_a_0[1]), .ZN(N4) );
  AND2_X1 U593 ( .A1(port_b_0[2]), .A2(port_a_0[2]), .ZN(N8) );
  AND2_X1 U594 ( .A1(port_b_0[3]), .A2(port_a_0[3]), .ZN(N12) );
  AND2_X1 U595 ( .A1(port_b_0[4]), .A2(port_a_0[4]), .ZN(N16) );
  AND2_X1 U596 ( .A1(port_b_0[5]), .A2(port_a_0[5]), .ZN(N20) );
  AND2_X1 U597 ( .A1(port_b_0[6]), .A2(port_a_0[6]), .ZN(N24) );
  AND2_X1 U598 ( .A1(port_b_1[0]), .A2(port_a_1[0]), .ZN(N1) );
  AND2_X1 U599 ( .A1(port_b_1[1]), .A2(port_a_1[1]), .ZN(N5) );
  AND2_X1 U600 ( .A1(port_b_1[2]), .A2(port_a_1[2]), .ZN(N9) );
  AND2_X1 U601 ( .A1(port_b_1[3]), .A2(port_a_1[3]), .ZN(N13) );
  AND2_X1 U602 ( .A1(port_b_1[4]), .A2(port_a_1[4]), .ZN(N17) );
  AND2_X1 U603 ( .A1(port_b_1[5]), .A2(port_a_1[5]), .ZN(N21) );
  AND2_X1 U604 ( .A1(port_b_1[6]), .A2(port_a_1[6]), .ZN(N25) );
  AND2_X1 U605 ( .A1(port_b_2[0]), .A2(port_a_2[0]), .ZN(N2) );
  AND2_X1 U606 ( .A1(port_b_2[1]), .A2(port_a_2[1]), .ZN(N6) );
  AND2_X1 U607 ( .A1(port_b_2[2]), .A2(port_a_2[2]), .ZN(N10) );
  AND2_X1 U608 ( .A1(port_b_2[3]), .A2(port_a_2[3]), .ZN(N14) );
  AND2_X1 U609 ( .A1(port_b_2[4]), .A2(port_a_2[4]), .ZN(N18) );
  AND2_X1 U610 ( .A1(port_b_2[5]), .A2(port_a_2[5]), .ZN(N22) );
  AND2_X1 U611 ( .A1(port_b_2[6]), .A2(port_a_2[6]), .ZN(N26) );
  AND2_X1 U612 ( .A1(port_b_3[0]), .A2(port_a_3[0]), .ZN(N3) );
  AND2_X1 U613 ( .A1(port_b_3[1]), .A2(port_a_3[1]), .ZN(N7) );
  AND2_X1 U614 ( .A1(port_b_3[2]), .A2(port_a_3[2]), .ZN(N11) );
  AND2_X1 U615 ( .A1(port_b_3[3]), .A2(port_a_3[3]), .ZN(N15) );
  AND2_X1 U616 ( .A1(port_b_3[4]), .A2(port_a_3[4]), .ZN(N19) );
  AND2_X1 U617 ( .A1(port_b_3[5]), .A2(port_a_3[5]), .ZN(N23) );
  AND2_X1 U618 ( .A1(port_b_3[6]), .A2(port_a_3[6]), .ZN(N27) );
  AND2_X1 simpleAnd_84_U1 ( .A1(port_rand_mul[0]), .A2(n7), .ZN(
        simpleAnd_84_port_z) );
  XOR2_X2 simpleXor_168_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_84_port_z), 
        .Z(u_0_0[0]) );
  XOR2_X2 simpleXor_169_U1 ( .A(port_rand_mul[0]), .B(port_b_1[0]), .Z(
        v_0_0[0]) );
  AND2_X1 simpleAnd_85_U1 ( .A1(port_rand_mul[1]), .A2(n7), .ZN(
        simpleAnd_85_port_z) );
  XOR2_X2 simpleXor_170_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_85_port_z), 
        .Z(u_0_1[0]) );
  XOR2_X2 simpleXor_171_U1 ( .A(port_rand_mul[1]), .B(port_b_2[0]), .Z(
        v_0_1[0]) );
  AND2_X1 simpleAnd_86_U1 ( .A1(port_rand_mul[2]), .A2(n7), .ZN(
        simpleAnd_86_port_z) );
  XOR2_X2 simpleXor_172_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_86_port_z), 
        .Z(u_0_2[0]) );
  XOR2_X2 simpleXor_173_U1 ( .A(port_rand_mul[2]), .B(port_b_3[0]), .Z(
        v_0_2[0]) );
  AND2_X1 simpleAnd_87_U1 ( .A1(port_rand_mul[0]), .A2(n14), .ZN(
        simpleAnd_87_port_z) );
  XOR2_X2 simpleXor_174_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_87_port_z), 
        .Z(u_1_0[0]) );
  XOR2_X2 simpleXor_175_U1 ( .A(port_rand_mul[0]), .B(port_b_0[0]), .Z(
        v_1_0[0]) );
  AND2_X1 simpleAnd_88_U1 ( .A1(port_rand_mul[3]), .A2(n14), .ZN(
        simpleAnd_88_port_z) );
  XOR2_X2 simpleXor_176_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_88_port_z), 
        .Z(u_1_1[0]) );
  XOR2_X2 simpleXor_177_U1 ( .A(port_rand_mul[3]), .B(port_b_2[0]), .Z(
        v_1_1[0]) );
  AND2_X1 simpleAnd_89_U1 ( .A1(port_rand_mul[4]), .A2(n14), .ZN(
        simpleAnd_89_port_z) );
  XOR2_X2 simpleXor_178_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_89_port_z), 
        .Z(u_1_2[0]) );
  XOR2_X2 simpleXor_179_U1 ( .A(port_rand_mul[4]), .B(port_b_3[0]), .Z(
        v_1_2[0]) );
  AND2_X1 simpleAnd_90_U1 ( .A1(port_rand_mul[1]), .A2(n21), .ZN(
        simpleAnd_90_port_z) );
  XOR2_X2 simpleXor_180_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_90_port_z), 
        .Z(u_2_0[0]) );
  XOR2_X2 simpleXor_181_U1 ( .A(port_rand_mul[1]), .B(port_b_0[0]), .Z(
        v_2_0[0]) );
  AND2_X1 simpleAnd_91_U1 ( .A1(port_rand_mul[3]), .A2(n21), .ZN(
        simpleAnd_91_port_z) );
  XOR2_X2 simpleXor_182_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_91_port_z), 
        .Z(u_2_1[0]) );
  XOR2_X2 simpleXor_183_U1 ( .A(port_rand_mul[3]), .B(port_b_1[0]), .Z(
        v_2_1[0]) );
  AND2_X1 simpleAnd_92_U1 ( .A1(port_rand_mul[5]), .A2(n21), .ZN(
        simpleAnd_92_port_z) );
  XOR2_X2 simpleXor_184_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_92_port_z), 
        .Z(u_2_2[0]) );
  XOR2_X2 simpleXor_185_U1 ( .A(port_rand_mul[5]), .B(port_b_3[0]), .Z(
        v_2_2[0]) );
  AND2_X1 simpleAnd_93_U1 ( .A1(port_rand_mul[2]), .A2(n28), .ZN(
        simpleAnd_93_port_z) );
  XOR2_X2 simpleXor_186_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_93_port_z), 
        .Z(u_3_0[0]) );
  XOR2_X2 simpleXor_187_U1 ( .A(port_rand_mul[2]), .B(port_b_0[0]), .Z(
        v_3_0[0]) );
  AND2_X1 simpleAnd_94_U1 ( .A1(port_rand_mul[4]), .A2(n28), .ZN(
        simpleAnd_94_port_z) );
  XOR2_X2 simpleXor_188_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_94_port_z), 
        .Z(u_3_1[0]) );
  XOR2_X2 simpleXor_189_U1 ( .A(port_rand_mul[4]), .B(port_b_1[0]), .Z(
        v_3_1[0]) );
  AND2_X1 simpleAnd_95_U1 ( .A1(port_rand_mul[5]), .A2(n28), .ZN(
        simpleAnd_95_port_z) );
  XOR2_X2 simpleXor_190_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_95_port_z), 
        .Z(u_3_2[0]) );
  XOR2_X2 simpleXor_191_U1 ( .A(port_rand_mul[5]), .B(port_b_2[0]), .Z(
        v_3_2[0]) );
  AND2_X1 simpleAnd_96_U1 ( .A1(port_rand_mul[0]), .A2(n6), .ZN(
        simpleAnd_96_port_z) );
  XOR2_X2 simpleXor_192_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_96_port_z), 
        .Z(u_0_0[1]) );
  XOR2_X2 simpleXor_193_U1 ( .A(port_rand_mul[0]), .B(port_b_1[1]), .Z(
        v_0_0[1]) );
  AND2_X1 simpleAnd_97_U1 ( .A1(port_rand_mul[1]), .A2(n6), .ZN(
        simpleAnd_97_port_z) );
  XOR2_X2 simpleXor_194_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_97_port_z), 
        .Z(u_0_1[1]) );
  XOR2_X2 simpleXor_195_U1 ( .A(port_rand_mul[1]), .B(port_b_2[1]), .Z(
        v_0_1[1]) );
  AND2_X1 simpleAnd_98_U1 ( .A1(port_rand_mul[2]), .A2(n6), .ZN(
        simpleAnd_98_port_z) );
  XOR2_X2 simpleXor_196_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_98_port_z), 
        .Z(u_0_2[1]) );
  XOR2_X2 simpleXor_197_U1 ( .A(port_rand_mul[2]), .B(port_b_3[1]), .Z(
        v_0_2[1]) );
  AND2_X1 simpleAnd_99_U1 ( .A1(port_rand_mul[0]), .A2(n13), .ZN(
        simpleAnd_99_port_z) );
  XOR2_X2 simpleXor_198_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_99_port_z), 
        .Z(u_1_0[1]) );
  XOR2_X2 simpleXor_199_U1 ( .A(port_rand_mul[0]), .B(port_b_0[1]), .Z(
        v_1_0[1]) );
  AND2_X1 simpleAnd_100_U1 ( .A1(port_rand_mul[3]), .A2(n13), .ZN(
        simpleAnd_100_port_z) );
  XOR2_X2 simpleXor_200_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_100_port_z), 
        .Z(u_1_1[1]) );
  XOR2_X2 simpleXor_201_U1 ( .A(port_rand_mul[3]), .B(port_b_2[1]), .Z(
        v_1_1[1]) );
  AND2_X1 simpleAnd_101_U1 ( .A1(port_rand_mul[4]), .A2(n13), .ZN(
        simpleAnd_101_port_z) );
  XOR2_X2 simpleXor_202_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_101_port_z), 
        .Z(u_1_2[1]) );
  XOR2_X2 simpleXor_203_U1 ( .A(port_rand_mul[4]), .B(port_b_3[1]), .Z(
        v_1_2[1]) );
  AND2_X1 simpleAnd_102_U1 ( .A1(port_rand_mul[1]), .A2(n20), .ZN(
        simpleAnd_102_port_z) );
  XOR2_X2 simpleXor_204_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_102_port_z), 
        .Z(u_2_0[1]) );
  XOR2_X2 simpleXor_205_U1 ( .A(port_rand_mul[1]), .B(port_b_0[1]), .Z(
        v_2_0[1]) );
  AND2_X1 simpleAnd_103_U1 ( .A1(port_rand_mul[3]), .A2(n20), .ZN(
        simpleAnd_103_port_z) );
  XOR2_X2 simpleXor_206_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_103_port_z), 
        .Z(u_2_1[1]) );
  XOR2_X2 simpleXor_207_U1 ( .A(port_rand_mul[3]), .B(port_b_1[1]), .Z(
        v_2_1[1]) );
  AND2_X1 simpleAnd_104_U1 ( .A1(port_rand_mul[5]), .A2(n20), .ZN(
        simpleAnd_104_port_z) );
  XOR2_X2 simpleXor_208_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_104_port_z), 
        .Z(u_2_2[1]) );
  XOR2_X2 simpleXor_209_U1 ( .A(port_rand_mul[5]), .B(port_b_3[1]), .Z(
        v_2_2[1]) );
  AND2_X1 simpleAnd_105_U1 ( .A1(port_rand_mul[2]), .A2(n27), .ZN(
        simpleAnd_105_port_z) );
  XOR2_X2 simpleXor_210_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_105_port_z), 
        .Z(u_3_0[1]) );
  XOR2_X2 simpleXor_211_U1 ( .A(port_rand_mul[2]), .B(port_b_0[1]), .Z(
        v_3_0[1]) );
  AND2_X1 simpleAnd_106_U1 ( .A1(port_rand_mul[4]), .A2(n27), .ZN(
        simpleAnd_106_port_z) );
  XOR2_X2 simpleXor_212_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_106_port_z), 
        .Z(u_3_1[1]) );
  XOR2_X2 simpleXor_213_U1 ( .A(port_rand_mul[4]), .B(port_b_1[1]), .Z(
        v_3_1[1]) );
  AND2_X1 simpleAnd_107_U1 ( .A1(port_rand_mul[5]), .A2(n27), .ZN(
        simpleAnd_107_port_z) );
  XOR2_X2 simpleXor_214_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_107_port_z), 
        .Z(u_3_2[1]) );
  XOR2_X2 simpleXor_215_U1 ( .A(port_rand_mul[5]), .B(port_b_2[1]), .Z(
        v_3_2[1]) );
  AND2_X1 simpleAnd_108_U1 ( .A1(port_rand_mul[0]), .A2(n5), .ZN(
        simpleAnd_108_port_z) );
  XOR2_X2 simpleXor_216_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_108_port_z), 
        .Z(u_0_0[2]) );
  XOR2_X2 simpleXor_217_U1 ( .A(port_rand_mul[0]), .B(port_b_1[2]), .Z(
        v_0_0[2]) );
  AND2_X1 simpleAnd_109_U1 ( .A1(port_rand_mul[1]), .A2(n5), .ZN(
        simpleAnd_109_port_z) );
  XOR2_X2 simpleXor_218_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_109_port_z), 
        .Z(u_0_1[2]) );
  XOR2_X2 simpleXor_219_U1 ( .A(port_rand_mul[1]), .B(port_b_2[2]), .Z(
        v_0_1[2]) );
  AND2_X1 simpleAnd_110_U1 ( .A1(port_rand_mul[2]), .A2(n5), .ZN(
        simpleAnd_110_port_z) );
  XOR2_X2 simpleXor_220_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_110_port_z), 
        .Z(u_0_2[2]) );
  XOR2_X2 simpleXor_221_U1 ( .A(port_rand_mul[2]), .B(port_b_3[2]), .Z(
        v_0_2[2]) );
  AND2_X1 simpleAnd_111_U1 ( .A1(port_rand_mul[0]), .A2(n12), .ZN(
        simpleAnd_111_port_z) );
  XOR2_X2 simpleXor_222_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_111_port_z), 
        .Z(u_1_0[2]) );
  XOR2_X2 simpleXor_223_U1 ( .A(port_rand_mul[0]), .B(port_b_0[2]), .Z(
        v_1_0[2]) );
  AND2_X1 simpleAnd_112_U1 ( .A1(port_rand_mul[3]), .A2(n12), .ZN(
        simpleAnd_112_port_z) );
  XOR2_X2 simpleXor_224_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_112_port_z), 
        .Z(u_1_1[2]) );
  XOR2_X2 simpleXor_225_U1 ( .A(port_rand_mul[3]), .B(port_b_2[2]), .Z(
        v_1_1[2]) );
  AND2_X1 simpleAnd_113_U1 ( .A1(port_rand_mul[4]), .A2(n12), .ZN(
        simpleAnd_113_port_z) );
  XOR2_X2 simpleXor_226_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_113_port_z), 
        .Z(u_1_2[2]) );
  XOR2_X2 simpleXor_227_U1 ( .A(port_rand_mul[4]), .B(port_b_3[2]), .Z(
        v_1_2[2]) );
  AND2_X1 simpleAnd_114_U1 ( .A1(port_rand_mul[1]), .A2(n19), .ZN(
        simpleAnd_114_port_z) );
  XOR2_X2 simpleXor_228_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_114_port_z), 
        .Z(u_2_0[2]) );
  XOR2_X2 simpleXor_229_U1 ( .A(port_rand_mul[1]), .B(port_b_0[2]), .Z(
        v_2_0[2]) );
  AND2_X1 simpleAnd_115_U1 ( .A1(port_rand_mul[3]), .A2(n19), .ZN(
        simpleAnd_115_port_z) );
  XOR2_X2 simpleXor_230_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_115_port_z), 
        .Z(u_2_1[2]) );
  XOR2_X2 simpleXor_231_U1 ( .A(port_rand_mul[3]), .B(port_b_1[2]), .Z(
        v_2_1[2]) );
  AND2_X1 simpleAnd_116_U1 ( .A1(port_rand_mul[5]), .A2(n19), .ZN(
        simpleAnd_116_port_z) );
  XOR2_X2 simpleXor_232_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_116_port_z), 
        .Z(u_2_2[2]) );
  XOR2_X2 simpleXor_233_U1 ( .A(port_rand_mul[5]), .B(port_b_3[2]), .Z(
        v_2_2[2]) );
  AND2_X1 simpleAnd_117_U1 ( .A1(port_rand_mul[2]), .A2(n26), .ZN(
        simpleAnd_117_port_z) );
  XOR2_X2 simpleXor_234_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_117_port_z), 
        .Z(u_3_0[2]) );
  XOR2_X2 simpleXor_235_U1 ( .A(port_rand_mul[2]), .B(port_b_0[2]), .Z(
        v_3_0[2]) );
  AND2_X1 simpleAnd_118_U1 ( .A1(port_rand_mul[4]), .A2(n26), .ZN(
        simpleAnd_118_port_z) );
  XOR2_X2 simpleXor_236_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_118_port_z), 
        .Z(u_3_1[2]) );
  XOR2_X2 simpleXor_237_U1 ( .A(port_rand_mul[4]), .B(port_b_1[2]), .Z(
        v_3_1[2]) );
  AND2_X1 simpleAnd_119_U1 ( .A1(port_rand_mul[5]), .A2(n26), .ZN(
        simpleAnd_119_port_z) );
  XOR2_X2 simpleXor_238_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_119_port_z), 
        .Z(u_3_2[2]) );
  XOR2_X2 simpleXor_239_U1 ( .A(port_rand_mul[5]), .B(port_b_2[2]), .Z(
        v_3_2[2]) );
  AND2_X1 simpleAnd_120_U1 ( .A1(port_rand_mul[0]), .A2(n4), .ZN(
        simpleAnd_120_port_z) );
  XOR2_X2 simpleXor_240_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_120_port_z), 
        .Z(u_0_0[3]) );
  XOR2_X2 simpleXor_241_U1 ( .A(port_rand_mul[0]), .B(port_b_1[3]), .Z(
        v_0_0[3]) );
  AND2_X1 simpleAnd_121_U1 ( .A1(port_rand_mul[1]), .A2(n4), .ZN(
        simpleAnd_121_port_z) );
  XOR2_X2 simpleXor_242_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_121_port_z), 
        .Z(u_0_1[3]) );
  XOR2_X2 simpleXor_243_U1 ( .A(port_rand_mul[1]), .B(port_b_2[3]), .Z(
        v_0_1[3]) );
  AND2_X1 simpleAnd_122_U1 ( .A1(port_rand_mul[2]), .A2(n4), .ZN(
        simpleAnd_122_port_z) );
  XOR2_X2 simpleXor_244_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_122_port_z), 
        .Z(u_0_2[3]) );
  XOR2_X2 simpleXor_245_U1 ( .A(port_rand_mul[2]), .B(port_b_3[3]), .Z(
        v_0_2[3]) );
  AND2_X1 simpleAnd_123_U1 ( .A1(port_rand_mul[0]), .A2(n11), .ZN(
        simpleAnd_123_port_z) );
  XOR2_X2 simpleXor_246_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_123_port_z), 
        .Z(u_1_0[3]) );
  XOR2_X2 simpleXor_247_U1 ( .A(port_rand_mul[0]), .B(port_b_0[3]), .Z(
        v_1_0[3]) );
  AND2_X1 simpleAnd_124_U1 ( .A1(port_rand_mul[3]), .A2(n11), .ZN(
        simpleAnd_124_port_z) );
  XOR2_X2 simpleXor_248_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_124_port_z), 
        .Z(u_1_1[3]) );
  XOR2_X2 simpleXor_249_U1 ( .A(port_rand_mul[3]), .B(port_b_2[3]), .Z(
        v_1_1[3]) );
  AND2_X1 simpleAnd_125_U1 ( .A1(port_rand_mul[4]), .A2(n11), .ZN(
        simpleAnd_125_port_z) );
  XOR2_X2 simpleXor_250_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_125_port_z), 
        .Z(u_1_2[3]) );
  XOR2_X2 simpleXor_251_U1 ( .A(port_rand_mul[4]), .B(port_b_3[3]), .Z(
        v_1_2[3]) );
  AND2_X1 simpleAnd_126_U1 ( .A1(port_rand_mul[1]), .A2(n18), .ZN(
        simpleAnd_126_port_z) );
  XOR2_X2 simpleXor_252_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_126_port_z), 
        .Z(u_2_0[3]) );
  XOR2_X2 simpleXor_253_U1 ( .A(port_rand_mul[1]), .B(port_b_0[3]), .Z(
        v_2_0[3]) );
  AND2_X1 simpleAnd_127_U1 ( .A1(port_rand_mul[3]), .A2(n18), .ZN(
        simpleAnd_127_port_z) );
  XOR2_X2 simpleXor_254_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_127_port_z), 
        .Z(u_2_1[3]) );
  XOR2_X2 simpleXor_255_U1 ( .A(port_rand_mul[3]), .B(port_b_1[3]), .Z(
        v_2_1[3]) );
  AND2_X1 simpleAnd_128_U1 ( .A1(port_rand_mul[5]), .A2(n18), .ZN(
        simpleAnd_128_port_z) );
  XOR2_X2 simpleXor_256_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_128_port_z), 
        .Z(u_2_2[3]) );
  XOR2_X2 simpleXor_257_U1 ( .A(port_rand_mul[5]), .B(port_b_3[3]), .Z(
        v_2_2[3]) );
  AND2_X1 simpleAnd_129_U1 ( .A1(port_rand_mul[2]), .A2(n25), .ZN(
        simpleAnd_129_port_z) );
  XOR2_X2 simpleXor_258_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_129_port_z), 
        .Z(u_3_0[3]) );
  XOR2_X2 simpleXor_259_U1 ( .A(port_rand_mul[2]), .B(port_b_0[3]), .Z(
        v_3_0[3]) );
  AND2_X1 simpleAnd_130_U1 ( .A1(port_rand_mul[4]), .A2(n25), .ZN(
        simpleAnd_130_port_z) );
  XOR2_X2 simpleXor_260_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_130_port_z), 
        .Z(u_3_1[3]) );
  XOR2_X2 simpleXor_261_U1 ( .A(port_rand_mul[4]), .B(port_b_1[3]), .Z(
        v_3_1[3]) );
  AND2_X1 simpleAnd_131_U1 ( .A1(port_rand_mul[5]), .A2(n25), .ZN(
        simpleAnd_131_port_z) );
  XOR2_X2 simpleXor_262_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_131_port_z), 
        .Z(u_3_2[3]) );
  XOR2_X2 simpleXor_263_U1 ( .A(port_rand_mul[5]), .B(port_b_2[3]), .Z(
        v_3_2[3]) );
  AND2_X1 simpleAnd_132_U1 ( .A1(port_rand_mul[0]), .A2(n3), .ZN(
        simpleAnd_132_port_z) );
  XOR2_X2 simpleXor_264_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_132_port_z), 
        .Z(u_0_0[4]) );
  XOR2_X2 simpleXor_265_U1 ( .A(port_rand_mul[0]), .B(port_b_1[4]), .Z(
        v_0_0[4]) );
  AND2_X1 simpleAnd_133_U1 ( .A1(port_rand_mul[1]), .A2(n3), .ZN(
        simpleAnd_133_port_z) );
  XOR2_X2 simpleXor_266_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_133_port_z), 
        .Z(u_0_1[4]) );
  XOR2_X2 simpleXor_267_U1 ( .A(port_rand_mul[1]), .B(port_b_2[4]), .Z(
        v_0_1[4]) );
  AND2_X1 simpleAnd_134_U1 ( .A1(port_rand_mul[2]), .A2(n3), .ZN(
        simpleAnd_134_port_z) );
  XOR2_X2 simpleXor_268_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_134_port_z), 
        .Z(u_0_2[4]) );
  XOR2_X2 simpleXor_269_U1 ( .A(port_rand_mul[2]), .B(port_b_3[4]), .Z(
        v_0_2[4]) );
  AND2_X1 simpleAnd_135_U1 ( .A1(port_rand_mul[0]), .A2(n10), .ZN(
        simpleAnd_135_port_z) );
  XOR2_X2 simpleXor_270_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_135_port_z), 
        .Z(u_1_0[4]) );
  XOR2_X2 simpleXor_271_U1 ( .A(port_rand_mul[0]), .B(port_b_0[4]), .Z(
        v_1_0[4]) );
  AND2_X1 simpleAnd_136_U1 ( .A1(port_rand_mul[3]), .A2(n10), .ZN(
        simpleAnd_136_port_z) );
  XOR2_X2 simpleXor_272_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_136_port_z), 
        .Z(u_1_1[4]) );
  XOR2_X2 simpleXor_273_U1 ( .A(port_rand_mul[3]), .B(port_b_2[4]), .Z(
        v_1_1[4]) );
  AND2_X1 simpleAnd_137_U1 ( .A1(port_rand_mul[4]), .A2(n10), .ZN(
        simpleAnd_137_port_z) );
  XOR2_X2 simpleXor_274_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_137_port_z), 
        .Z(u_1_2[4]) );
  XOR2_X2 simpleXor_275_U1 ( .A(port_rand_mul[4]), .B(port_b_3[4]), .Z(
        v_1_2[4]) );
  AND2_X1 simpleAnd_138_U1 ( .A1(port_rand_mul[1]), .A2(n17), .ZN(
        simpleAnd_138_port_z) );
  XOR2_X2 simpleXor_276_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_138_port_z), 
        .Z(u_2_0[4]) );
  XOR2_X2 simpleXor_277_U1 ( .A(port_rand_mul[1]), .B(port_b_0[4]), .Z(
        v_2_0[4]) );
  AND2_X1 simpleAnd_139_U1 ( .A1(port_rand_mul[3]), .A2(n17), .ZN(
        simpleAnd_139_port_z) );
  XOR2_X2 simpleXor_278_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_139_port_z), 
        .Z(u_2_1[4]) );
  XOR2_X2 simpleXor_279_U1 ( .A(port_rand_mul[3]), .B(port_b_1[4]), .Z(
        v_2_1[4]) );
  AND2_X1 simpleAnd_140_U1 ( .A1(port_rand_mul[5]), .A2(n17), .ZN(
        simpleAnd_140_port_z) );
  XOR2_X2 simpleXor_280_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_140_port_z), 
        .Z(u_2_2[4]) );
  XOR2_X2 simpleXor_281_U1 ( .A(port_rand_mul[5]), .B(port_b_3[4]), .Z(
        v_2_2[4]) );
  AND2_X1 simpleAnd_141_U1 ( .A1(port_rand_mul[2]), .A2(n24), .ZN(
        simpleAnd_141_port_z) );
  XOR2_X2 simpleXor_282_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_141_port_z), 
        .Z(u_3_0[4]) );
  XOR2_X2 simpleXor_283_U1 ( .A(port_rand_mul[2]), .B(port_b_0[4]), .Z(
        v_3_0[4]) );
  AND2_X1 simpleAnd_142_U1 ( .A1(port_rand_mul[4]), .A2(n24), .ZN(
        simpleAnd_142_port_z) );
  XOR2_X2 simpleXor_284_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_142_port_z), 
        .Z(u_3_1[4]) );
  XOR2_X2 simpleXor_285_U1 ( .A(port_rand_mul[4]), .B(port_b_1[4]), .Z(
        v_3_1[4]) );
  AND2_X1 simpleAnd_143_U1 ( .A1(port_rand_mul[5]), .A2(n24), .ZN(
        simpleAnd_143_port_z) );
  XOR2_X2 simpleXor_286_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_143_port_z), 
        .Z(u_3_2[4]) );
  XOR2_X2 simpleXor_287_U1 ( .A(port_rand_mul[5]), .B(port_b_2[4]), .Z(
        v_3_2[4]) );
  AND2_X1 simpleAnd_144_U1 ( .A1(port_rand_mul[0]), .A2(n2), .ZN(
        simpleAnd_144_port_z) );
  XOR2_X2 simpleXor_288_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_144_port_z), 
        .Z(u_0_0[5]) );
  XOR2_X2 simpleXor_289_U1 ( .A(port_rand_mul[0]), .B(port_b_1[5]), .Z(
        v_0_0[5]) );
  AND2_X1 simpleAnd_145_U1 ( .A1(port_rand_mul[1]), .A2(n2), .ZN(
        simpleAnd_145_port_z) );
  XOR2_X2 simpleXor_290_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_145_port_z), 
        .Z(u_0_1[5]) );
  XOR2_X2 simpleXor_291_U1 ( .A(port_rand_mul[1]), .B(port_b_2[5]), .Z(
        v_0_1[5]) );
  AND2_X1 simpleAnd_146_U1 ( .A1(port_rand_mul[2]), .A2(n2), .ZN(
        simpleAnd_146_port_z) );
  XOR2_X2 simpleXor_292_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_146_port_z), 
        .Z(u_0_2[5]) );
  XOR2_X2 simpleXor_293_U1 ( .A(port_rand_mul[2]), .B(port_b_3[5]), .Z(
        v_0_2[5]) );
  AND2_X1 simpleAnd_147_U1 ( .A1(port_rand_mul[0]), .A2(n9), .ZN(
        simpleAnd_147_port_z) );
  XOR2_X2 simpleXor_294_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_147_port_z), 
        .Z(u_1_0[5]) );
  XOR2_X2 simpleXor_295_U1 ( .A(port_rand_mul[0]), .B(port_b_0[5]), .Z(
        v_1_0[5]) );
  AND2_X1 simpleAnd_148_U1 ( .A1(port_rand_mul[3]), .A2(n9), .ZN(
        simpleAnd_148_port_z) );
  XOR2_X2 simpleXor_296_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_148_port_z), 
        .Z(u_1_1[5]) );
  XOR2_X2 simpleXor_297_U1 ( .A(port_rand_mul[3]), .B(port_b_2[5]), .Z(
        v_1_1[5]) );
  AND2_X1 simpleAnd_149_U1 ( .A1(port_rand_mul[4]), .A2(n9), .ZN(
        simpleAnd_149_port_z) );
  XOR2_X2 simpleXor_298_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_149_port_z), 
        .Z(u_1_2[5]) );
  XOR2_X2 simpleXor_299_U1 ( .A(port_rand_mul[4]), .B(port_b_3[5]), .Z(
        v_1_2[5]) );
  AND2_X1 simpleAnd_150_U1 ( .A1(port_rand_mul[1]), .A2(n16), .ZN(
        simpleAnd_150_port_z) );
  XOR2_X2 simpleXor_300_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_150_port_z), 
        .Z(u_2_0[5]) );
  XOR2_X2 simpleXor_301_U1 ( .A(port_rand_mul[1]), .B(port_b_0[5]), .Z(
        v_2_0[5]) );
  AND2_X1 simpleAnd_151_U1 ( .A1(port_rand_mul[3]), .A2(n16), .ZN(
        simpleAnd_151_port_z) );
  XOR2_X2 simpleXor_302_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_151_port_z), 
        .Z(u_2_1[5]) );
  XOR2_X2 simpleXor_303_U1 ( .A(port_rand_mul[3]), .B(port_b_1[5]), .Z(
        v_2_1[5]) );
  AND2_X1 simpleAnd_152_U1 ( .A1(port_rand_mul[5]), .A2(n16), .ZN(
        simpleAnd_152_port_z) );
  XOR2_X2 simpleXor_304_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_152_port_z), 
        .Z(u_2_2[5]) );
  XOR2_X2 simpleXor_305_U1 ( .A(port_rand_mul[5]), .B(port_b_3[5]), .Z(
        v_2_2[5]) );
  AND2_X1 simpleAnd_153_U1 ( .A1(port_rand_mul[2]), .A2(n23), .ZN(
        simpleAnd_153_port_z) );
  XOR2_X2 simpleXor_306_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_153_port_z), 
        .Z(u_3_0[5]) );
  XOR2_X2 simpleXor_307_U1 ( .A(port_rand_mul[2]), .B(port_b_0[5]), .Z(
        v_3_0[5]) );
  AND2_X1 simpleAnd_154_U1 ( .A1(port_rand_mul[4]), .A2(n23), .ZN(
        simpleAnd_154_port_z) );
  XOR2_X2 simpleXor_308_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_154_port_z), 
        .Z(u_3_1[5]) );
  XOR2_X2 simpleXor_309_U1 ( .A(port_rand_mul[4]), .B(port_b_1[5]), .Z(
        v_3_1[5]) );
  AND2_X1 simpleAnd_155_U1 ( .A1(port_rand_mul[5]), .A2(n23), .ZN(
        simpleAnd_155_port_z) );
  XOR2_X2 simpleXor_310_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_155_port_z), 
        .Z(u_3_2[5]) );
  XOR2_X2 simpleXor_311_U1 ( .A(port_rand_mul[5]), .B(port_b_2[5]), .Z(
        v_3_2[5]) );
  AND2_X1 simpleAnd_156_U1 ( .A1(port_rand_mul[0]), .A2(n1), .ZN(
        simpleAnd_156_port_z) );
  XOR2_X1 simpleXor_312_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_156_port_z), 
        .Z(u_0_0[6]) );
  XOR2_X1 simpleXor_313_U1 ( .A(port_rand_mul[0]), .B(port_b_1[6]), .Z(
        v_0_0[6]) );
  AND2_X1 simpleAnd_157_U1 ( .A1(port_rand_mul[1]), .A2(n1), .ZN(
        simpleAnd_157_port_z) );
  XOR2_X1 simpleXor_314_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_157_port_z), 
        .Z(u_0_1[6]) );
  XOR2_X1 simpleXor_315_U1 ( .A(port_rand_mul[1]), .B(port_b_2[6]), .Z(
        v_0_1[6]) );
  AND2_X1 simpleAnd_158_U1 ( .A1(port_rand_mul[2]), .A2(n1), .ZN(
        simpleAnd_158_port_z) );
  XOR2_X1 simpleXor_316_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_158_port_z), 
        .Z(u_0_2[6]) );
  XOR2_X1 simpleXor_317_U1 ( .A(port_rand_mul[2]), .B(port_b_3[6]), .Z(
        v_0_2[6]) );
  AND2_X1 simpleAnd_159_U1 ( .A1(port_rand_mul[0]), .A2(n8), .ZN(
        simpleAnd_159_port_z) );
  XOR2_X1 simpleXor_318_U1 ( .A(port_rand_ref[0]), .B(simpleAnd_159_port_z), 
        .Z(u_1_0[6]) );
  XOR2_X1 simpleXor_319_U1 ( .A(port_rand_mul[0]), .B(port_b_0[6]), .Z(
        v_1_0[6]) );
  AND2_X1 simpleAnd_160_U1 ( .A1(port_rand_mul[3]), .A2(n8), .ZN(
        simpleAnd_160_port_z) );
  XOR2_X1 simpleXor_320_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_160_port_z), 
        .Z(u_1_1[6]) );
  XOR2_X1 simpleXor_321_U1 ( .A(port_rand_mul[3]), .B(port_b_2[6]), .Z(
        v_1_1[6]) );
  AND2_X1 simpleAnd_161_U1 ( .A1(port_rand_mul[4]), .A2(n8), .ZN(
        simpleAnd_161_port_z) );
  XOR2_X1 simpleXor_322_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_161_port_z), 
        .Z(u_1_2[6]) );
  XOR2_X1 simpleXor_323_U1 ( .A(port_rand_mul[4]), .B(port_b_3[6]), .Z(
        v_1_2[6]) );
  AND2_X1 simpleAnd_162_U1 ( .A1(port_rand_mul[1]), .A2(n15), .ZN(
        simpleAnd_162_port_z) );
  XOR2_X1 simpleXor_324_U1 ( .A(port_rand_ref[1]), .B(simpleAnd_162_port_z), 
        .Z(u_2_0[6]) );
  XOR2_X1 simpleXor_325_U1 ( .A(port_rand_mul[1]), .B(port_b_0[6]), .Z(
        v_2_0[6]) );
  AND2_X1 simpleAnd_163_U1 ( .A1(port_rand_mul[3]), .A2(n15), .ZN(
        simpleAnd_163_port_z) );
  XOR2_X1 simpleXor_326_U1 ( .A(port_rand_ref[3]), .B(simpleAnd_163_port_z), 
        .Z(u_2_1[6]) );
  XOR2_X1 simpleXor_327_U1 ( .A(port_rand_mul[3]), .B(port_b_1[6]), .Z(
        v_2_1[6]) );
  AND2_X1 simpleAnd_164_U1 ( .A1(port_rand_mul[5]), .A2(n15), .ZN(
        simpleAnd_164_port_z) );
  XOR2_X1 simpleXor_328_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_164_port_z), 
        .Z(u_2_2[6]) );
  XOR2_X1 simpleXor_329_U1 ( .A(port_rand_mul[5]), .B(port_b_3[6]), .Z(
        v_2_2[6]) );
  AND2_X1 simpleAnd_165_U1 ( .A1(port_rand_mul[2]), .A2(n22), .ZN(
        simpleAnd_165_port_z) );
  XOR2_X1 simpleXor_330_U1 ( .A(port_rand_ref[2]), .B(simpleAnd_165_port_z), 
        .Z(u_3_0[6]) );
  XOR2_X1 simpleXor_331_U1 ( .A(port_rand_mul[2]), .B(port_b_0[6]), .Z(
        v_3_0[6]) );
  AND2_X1 simpleAnd_166_U1 ( .A1(port_rand_mul[4]), .A2(n22), .ZN(
        simpleAnd_166_port_z) );
  XOR2_X1 simpleXor_332_U1 ( .A(port_rand_ref[4]), .B(simpleAnd_166_port_z), 
        .Z(u_3_1[6]) );
  XOR2_X1 simpleXor_333_U1 ( .A(port_rand_mul[4]), .B(port_b_1[6]), .Z(
        v_3_1[6]) );
  AND2_X1 simpleAnd_167_U1 ( .A1(port_rand_mul[5]), .A2(n22), .ZN(
        simpleAnd_167_port_z) );
  XOR2_X1 simpleXor_334_U1 ( .A(port_rand_ref[5]), .B(simpleAnd_167_port_z), 
        .Z(u_3_2[6]) );
  XOR2_X1 simpleXor_335_U1 ( .A(port_rand_mul[5]), .B(port_b_2[6]), .Z(
        v_3_2[6]) );
  OR2_X1 maj_168_U19 ( .A1(maj_168_n8), .A2(maj_168_n9), .ZN(maj_168_n7) );
  NAND2_X1 maj_168_U18 ( .A1(u_0_0[6]), .A2(maj_168_n7), .ZN(maj_168_n6) );
  NAND2_X1 maj_168_U17 ( .A1(maj_168_n9), .A2(maj_168_n8), .ZN(maj_168_n5) );
  NAND2_X1 maj_168_U16 ( .A1(maj_168_n5), .A2(maj_168_n6), .ZN(maj_168_n4) );
  NAND2_X1 maj_168_U15 ( .A1(u_0_0[5]), .A2(maj_168_n10), .ZN(maj_168_n17) );
  NAND2_X1 maj_168_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_168_n16) );
  NAND2_X1 maj_168_U13 ( .A1(maj_168_n16), .A2(maj_168_n17), .ZN(maj_168_n13)
         );
  NAND2_X1 maj_168_U12 ( .A1(u_0_0[2]), .A2(maj_168_n11), .ZN(maj_168_n15) );
  NAND2_X1 maj_168_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_168_n14) );
  NAND2_X1 maj_168_U10 ( .A1(maj_168_n14), .A2(maj_168_n15), .ZN(maj_168_n12)
         );
  XOR2_X1 maj_168_U9 ( .A(u_0_0[2]), .B(maj_168_n11), .Z(maj_168_n9) );
  XOR2_X1 maj_168_U8 ( .A(u_0_0[5]), .B(maj_168_n10), .Z(maj_168_n8) );
  XOR2_X1 maj_168_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_168_n11) );
  XOR2_X1 maj_168_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_168_n10) );
  OR2_X1 maj_168_U5 ( .A1(maj_168_n12), .A2(maj_168_n13), .ZN(maj_168_n3) );
  NAND2_X1 maj_168_U4 ( .A1(maj_168_n13), .A2(maj_168_n12), .ZN(maj_168_n1) );
  NAND2_X1 maj_168_U3 ( .A1(maj_168_n3), .A2(maj_168_n4), .ZN(maj_168_n2) );
  NAND2_X1 maj_168_U2 ( .A1(maj_168_n1), .A2(maj_168_n2), .ZN(maj_168_port_o)
         );
  OR2_X1 maj_169_U19 ( .A1(maj_169_n27), .A2(maj_169_n26), .ZN(maj_169_n28) );
  NAND2_X1 maj_169_U18 ( .A1(v_0_0[6]), .A2(maj_169_n28), .ZN(maj_169_n29) );
  NAND2_X1 maj_169_U17 ( .A1(maj_169_n26), .A2(maj_169_n27), .ZN(maj_169_n30)
         );
  NAND2_X1 maj_169_U16 ( .A1(maj_169_n30), .A2(maj_169_n29), .ZN(maj_169_n31)
         );
  NAND2_X1 maj_169_U15 ( .A1(v_0_0[5]), .A2(maj_169_n25), .ZN(maj_169_n18) );
  NAND2_X1 maj_169_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_169_n19) );
  NAND2_X1 maj_169_U13 ( .A1(maj_169_n19), .A2(maj_169_n18), .ZN(maj_169_n22)
         );
  NAND2_X1 maj_169_U12 ( .A1(v_0_0[2]), .A2(maj_169_n24), .ZN(maj_169_n20) );
  NAND2_X1 maj_169_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_169_n21) );
  NAND2_X1 maj_169_U10 ( .A1(maj_169_n21), .A2(maj_169_n20), .ZN(maj_169_n23)
         );
  XOR2_X1 maj_169_U9 ( .A(v_0_0[2]), .B(maj_169_n24), .Z(maj_169_n26) );
  XOR2_X1 maj_169_U8 ( .A(v_0_0[5]), .B(maj_169_n25), .Z(maj_169_n27) );
  XOR2_X1 maj_169_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_169_n24) );
  XOR2_X1 maj_169_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_169_n25) );
  OR2_X1 maj_169_U5 ( .A1(maj_169_n23), .A2(maj_169_n22), .ZN(maj_169_n32) );
  NAND2_X1 maj_169_U4 ( .A1(maj_169_n22), .A2(maj_169_n23), .ZN(maj_169_n34)
         );
  NAND2_X1 maj_169_U3 ( .A1(maj_169_n32), .A2(maj_169_n31), .ZN(maj_169_n33)
         );
  NAND2_X1 maj_169_U2 ( .A1(maj_169_n34), .A2(maj_169_n33), .ZN(maj_169_port_o) );
  OR2_X1 maj_170_U19 ( .A1(maj_170_n27), .A2(maj_170_n26), .ZN(maj_170_n28) );
  NAND2_X1 maj_170_U18 ( .A1(u_0_1[6]), .A2(maj_170_n28), .ZN(maj_170_n29) );
  NAND2_X1 maj_170_U17 ( .A1(maj_170_n26), .A2(maj_170_n27), .ZN(maj_170_n30)
         );
  NAND2_X1 maj_170_U16 ( .A1(maj_170_n30), .A2(maj_170_n29), .ZN(maj_170_n31)
         );
  NAND2_X1 maj_170_U15 ( .A1(u_0_1[5]), .A2(maj_170_n25), .ZN(maj_170_n18) );
  NAND2_X1 maj_170_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_170_n19) );
  NAND2_X1 maj_170_U13 ( .A1(maj_170_n19), .A2(maj_170_n18), .ZN(maj_170_n22)
         );
  NAND2_X1 maj_170_U12 ( .A1(u_0_1[2]), .A2(maj_170_n24), .ZN(maj_170_n20) );
  NAND2_X1 maj_170_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_170_n21) );
  NAND2_X1 maj_170_U10 ( .A1(maj_170_n21), .A2(maj_170_n20), .ZN(maj_170_n23)
         );
  XOR2_X1 maj_170_U9 ( .A(u_0_1[2]), .B(maj_170_n24), .Z(maj_170_n26) );
  XOR2_X1 maj_170_U8 ( .A(u_0_1[5]), .B(maj_170_n25), .Z(maj_170_n27) );
  XOR2_X1 maj_170_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_170_n24) );
  XOR2_X1 maj_170_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_170_n25) );
  OR2_X1 maj_170_U5 ( .A1(maj_170_n23), .A2(maj_170_n22), .ZN(maj_170_n32) );
  NAND2_X1 maj_170_U4 ( .A1(maj_170_n22), .A2(maj_170_n23), .ZN(maj_170_n34)
         );
  NAND2_X1 maj_170_U3 ( .A1(maj_170_n32), .A2(maj_170_n31), .ZN(maj_170_n33)
         );
  NAND2_X1 maj_170_U2 ( .A1(maj_170_n34), .A2(maj_170_n33), .ZN(maj_170_port_o) );
  OR2_X1 maj_171_U19 ( .A1(maj_171_n27), .A2(maj_171_n26), .ZN(maj_171_n28) );
  NAND2_X1 maj_171_U18 ( .A1(v_0_1[6]), .A2(maj_171_n28), .ZN(maj_171_n29) );
  NAND2_X1 maj_171_U17 ( .A1(maj_171_n26), .A2(maj_171_n27), .ZN(maj_171_n30)
         );
  NAND2_X1 maj_171_U16 ( .A1(maj_171_n30), .A2(maj_171_n29), .ZN(maj_171_n31)
         );
  NAND2_X1 maj_171_U15 ( .A1(v_0_1[5]), .A2(maj_171_n25), .ZN(maj_171_n18) );
  NAND2_X1 maj_171_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_171_n19) );
  NAND2_X1 maj_171_U13 ( .A1(maj_171_n19), .A2(maj_171_n18), .ZN(maj_171_n22)
         );
  NAND2_X1 maj_171_U12 ( .A1(v_0_1[2]), .A2(maj_171_n24), .ZN(maj_171_n20) );
  NAND2_X1 maj_171_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_171_n21) );
  NAND2_X1 maj_171_U10 ( .A1(maj_171_n21), .A2(maj_171_n20), .ZN(maj_171_n23)
         );
  XOR2_X1 maj_171_U9 ( .A(v_0_1[2]), .B(maj_171_n24), .Z(maj_171_n26) );
  XOR2_X1 maj_171_U8 ( .A(v_0_1[5]), .B(maj_171_n25), .Z(maj_171_n27) );
  XOR2_X1 maj_171_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_171_n24) );
  XOR2_X1 maj_171_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_171_n25) );
  OR2_X1 maj_171_U5 ( .A1(maj_171_n23), .A2(maj_171_n22), .ZN(maj_171_n32) );
  NAND2_X1 maj_171_U4 ( .A1(maj_171_n22), .A2(maj_171_n23), .ZN(maj_171_n34)
         );
  NAND2_X1 maj_171_U3 ( .A1(maj_171_n32), .A2(maj_171_n31), .ZN(maj_171_n33)
         );
  NAND2_X1 maj_171_U2 ( .A1(maj_171_n34), .A2(maj_171_n33), .ZN(maj_171_port_o) );
  OR2_X1 maj_172_U19 ( .A1(maj_172_n27), .A2(maj_172_n26), .ZN(maj_172_n28) );
  NAND2_X1 maj_172_U18 ( .A1(u_0_2[6]), .A2(maj_172_n28), .ZN(maj_172_n29) );
  NAND2_X1 maj_172_U17 ( .A1(maj_172_n26), .A2(maj_172_n27), .ZN(maj_172_n30)
         );
  NAND2_X1 maj_172_U16 ( .A1(maj_172_n30), .A2(maj_172_n29), .ZN(maj_172_n31)
         );
  NAND2_X1 maj_172_U15 ( .A1(u_0_2[5]), .A2(maj_172_n25), .ZN(maj_172_n18) );
  NAND2_X1 maj_172_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_172_n19) );
  NAND2_X1 maj_172_U13 ( .A1(maj_172_n19), .A2(maj_172_n18), .ZN(maj_172_n22)
         );
  NAND2_X1 maj_172_U12 ( .A1(u_0_2[2]), .A2(maj_172_n24), .ZN(maj_172_n20) );
  NAND2_X1 maj_172_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_172_n21) );
  NAND2_X1 maj_172_U10 ( .A1(maj_172_n21), .A2(maj_172_n20), .ZN(maj_172_n23)
         );
  XOR2_X1 maj_172_U9 ( .A(u_0_2[2]), .B(maj_172_n24), .Z(maj_172_n26) );
  XOR2_X1 maj_172_U8 ( .A(u_0_2[5]), .B(maj_172_n25), .Z(maj_172_n27) );
  XOR2_X1 maj_172_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_172_n24) );
  XOR2_X1 maj_172_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_172_n25) );
  OR2_X1 maj_172_U5 ( .A1(maj_172_n23), .A2(maj_172_n22), .ZN(maj_172_n32) );
  NAND2_X1 maj_172_U4 ( .A1(maj_172_n22), .A2(maj_172_n23), .ZN(maj_172_n34)
         );
  NAND2_X1 maj_172_U3 ( .A1(maj_172_n32), .A2(maj_172_n31), .ZN(maj_172_n33)
         );
  NAND2_X1 maj_172_U2 ( .A1(maj_172_n34), .A2(maj_172_n33), .ZN(maj_172_port_o) );
  OR2_X1 maj_173_U19 ( .A1(maj_173_n27), .A2(maj_173_n26), .ZN(maj_173_n28) );
  NAND2_X1 maj_173_U18 ( .A1(v_0_2[6]), .A2(maj_173_n28), .ZN(maj_173_n29) );
  NAND2_X1 maj_173_U17 ( .A1(maj_173_n26), .A2(maj_173_n27), .ZN(maj_173_n30)
         );
  NAND2_X1 maj_173_U16 ( .A1(maj_173_n30), .A2(maj_173_n29), .ZN(maj_173_n31)
         );
  NAND2_X1 maj_173_U15 ( .A1(v_0_2[5]), .A2(maj_173_n25), .ZN(maj_173_n18) );
  NAND2_X1 maj_173_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_173_n19) );
  NAND2_X1 maj_173_U13 ( .A1(maj_173_n19), .A2(maj_173_n18), .ZN(maj_173_n22)
         );
  NAND2_X1 maj_173_U12 ( .A1(v_0_2[2]), .A2(maj_173_n24), .ZN(maj_173_n20) );
  NAND2_X1 maj_173_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_173_n21) );
  NAND2_X1 maj_173_U10 ( .A1(maj_173_n21), .A2(maj_173_n20), .ZN(maj_173_n23)
         );
  XOR2_X1 maj_173_U9 ( .A(v_0_2[2]), .B(maj_173_n24), .Z(maj_173_n26) );
  XOR2_X1 maj_173_U8 ( .A(v_0_2[5]), .B(maj_173_n25), .Z(maj_173_n27) );
  XOR2_X1 maj_173_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_173_n24) );
  XOR2_X1 maj_173_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_173_n25) );
  OR2_X1 maj_173_U5 ( .A1(maj_173_n23), .A2(maj_173_n22), .ZN(maj_173_n32) );
  NAND2_X1 maj_173_U4 ( .A1(maj_173_n22), .A2(maj_173_n23), .ZN(maj_173_n34)
         );
  NAND2_X1 maj_173_U3 ( .A1(maj_173_n32), .A2(maj_173_n31), .ZN(maj_173_n33)
         );
  NAND2_X1 maj_173_U2 ( .A1(maj_173_n34), .A2(maj_173_n33), .ZN(maj_173_port_o) );
  OR2_X1 maj_174_U19 ( .A1(maj_174_n27), .A2(maj_174_n26), .ZN(maj_174_n28) );
  NAND2_X1 maj_174_U18 ( .A1(u_1_0[6]), .A2(maj_174_n28), .ZN(maj_174_n29) );
  NAND2_X1 maj_174_U17 ( .A1(maj_174_n26), .A2(maj_174_n27), .ZN(maj_174_n30)
         );
  NAND2_X1 maj_174_U16 ( .A1(maj_174_n30), .A2(maj_174_n29), .ZN(maj_174_n31)
         );
  NAND2_X1 maj_174_U15 ( .A1(u_1_0[5]), .A2(maj_174_n25), .ZN(maj_174_n18) );
  NAND2_X1 maj_174_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_174_n19) );
  NAND2_X1 maj_174_U13 ( .A1(maj_174_n19), .A2(maj_174_n18), .ZN(maj_174_n22)
         );
  NAND2_X1 maj_174_U12 ( .A1(u_1_0[2]), .A2(maj_174_n24), .ZN(maj_174_n20) );
  NAND2_X1 maj_174_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_174_n21) );
  NAND2_X1 maj_174_U10 ( .A1(maj_174_n21), .A2(maj_174_n20), .ZN(maj_174_n23)
         );
  XOR2_X1 maj_174_U9 ( .A(u_1_0[2]), .B(maj_174_n24), .Z(maj_174_n26) );
  XOR2_X1 maj_174_U8 ( .A(u_1_0[5]), .B(maj_174_n25), .Z(maj_174_n27) );
  XOR2_X1 maj_174_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_174_n24) );
  XOR2_X1 maj_174_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_174_n25) );
  OR2_X1 maj_174_U5 ( .A1(maj_174_n23), .A2(maj_174_n22), .ZN(maj_174_n32) );
  NAND2_X1 maj_174_U4 ( .A1(maj_174_n22), .A2(maj_174_n23), .ZN(maj_174_n34)
         );
  NAND2_X1 maj_174_U3 ( .A1(maj_174_n32), .A2(maj_174_n31), .ZN(maj_174_n33)
         );
  NAND2_X1 maj_174_U2 ( .A1(maj_174_n34), .A2(maj_174_n33), .ZN(maj_174_port_o) );
  OR2_X1 maj_175_U19 ( .A1(maj_175_n27), .A2(maj_175_n26), .ZN(maj_175_n28) );
  NAND2_X1 maj_175_U18 ( .A1(v_1_0[6]), .A2(maj_175_n28), .ZN(maj_175_n29) );
  NAND2_X1 maj_175_U17 ( .A1(maj_175_n26), .A2(maj_175_n27), .ZN(maj_175_n30)
         );
  NAND2_X1 maj_175_U16 ( .A1(maj_175_n30), .A2(maj_175_n29), .ZN(maj_175_n31)
         );
  NAND2_X1 maj_175_U15 ( .A1(v_1_0[5]), .A2(maj_175_n25), .ZN(maj_175_n18) );
  NAND2_X1 maj_175_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_175_n19) );
  NAND2_X1 maj_175_U13 ( .A1(maj_175_n19), .A2(maj_175_n18), .ZN(maj_175_n22)
         );
  NAND2_X1 maj_175_U12 ( .A1(v_1_0[2]), .A2(maj_175_n24), .ZN(maj_175_n20) );
  NAND2_X1 maj_175_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_175_n21) );
  NAND2_X1 maj_175_U10 ( .A1(maj_175_n21), .A2(maj_175_n20), .ZN(maj_175_n23)
         );
  XOR2_X1 maj_175_U9 ( .A(v_1_0[2]), .B(maj_175_n24), .Z(maj_175_n26) );
  XOR2_X1 maj_175_U8 ( .A(v_1_0[5]), .B(maj_175_n25), .Z(maj_175_n27) );
  XOR2_X1 maj_175_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_175_n24) );
  XOR2_X1 maj_175_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_175_n25) );
  OR2_X1 maj_175_U5 ( .A1(maj_175_n23), .A2(maj_175_n22), .ZN(maj_175_n32) );
  NAND2_X1 maj_175_U4 ( .A1(maj_175_n22), .A2(maj_175_n23), .ZN(maj_175_n34)
         );
  NAND2_X1 maj_175_U3 ( .A1(maj_175_n32), .A2(maj_175_n31), .ZN(maj_175_n33)
         );
  NAND2_X1 maj_175_U2 ( .A1(maj_175_n34), .A2(maj_175_n33), .ZN(maj_175_port_o) );
  OR2_X1 maj_176_U19 ( .A1(maj_176_n27), .A2(maj_176_n26), .ZN(maj_176_n28) );
  NAND2_X1 maj_176_U18 ( .A1(u_1_1[6]), .A2(maj_176_n28), .ZN(maj_176_n29) );
  NAND2_X1 maj_176_U17 ( .A1(maj_176_n26), .A2(maj_176_n27), .ZN(maj_176_n30)
         );
  NAND2_X1 maj_176_U16 ( .A1(maj_176_n30), .A2(maj_176_n29), .ZN(maj_176_n31)
         );
  NAND2_X1 maj_176_U15 ( .A1(u_1_1[5]), .A2(maj_176_n25), .ZN(maj_176_n18) );
  NAND2_X1 maj_176_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_176_n19) );
  NAND2_X1 maj_176_U13 ( .A1(maj_176_n19), .A2(maj_176_n18), .ZN(maj_176_n22)
         );
  NAND2_X1 maj_176_U12 ( .A1(u_1_1[2]), .A2(maj_176_n24), .ZN(maj_176_n20) );
  NAND2_X1 maj_176_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_176_n21) );
  NAND2_X1 maj_176_U10 ( .A1(maj_176_n21), .A2(maj_176_n20), .ZN(maj_176_n23)
         );
  XOR2_X1 maj_176_U9 ( .A(u_1_1[2]), .B(maj_176_n24), .Z(maj_176_n26) );
  XOR2_X1 maj_176_U8 ( .A(u_1_1[5]), .B(maj_176_n25), .Z(maj_176_n27) );
  XOR2_X1 maj_176_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_176_n24) );
  XOR2_X1 maj_176_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_176_n25) );
  OR2_X1 maj_176_U5 ( .A1(maj_176_n23), .A2(maj_176_n22), .ZN(maj_176_n32) );
  NAND2_X1 maj_176_U4 ( .A1(maj_176_n22), .A2(maj_176_n23), .ZN(maj_176_n34)
         );
  NAND2_X1 maj_176_U3 ( .A1(maj_176_n32), .A2(maj_176_n31), .ZN(maj_176_n33)
         );
  NAND2_X1 maj_176_U2 ( .A1(maj_176_n34), .A2(maj_176_n33), .ZN(maj_176_port_o) );
  OR2_X1 maj_177_U19 ( .A1(maj_177_n27), .A2(maj_177_n26), .ZN(maj_177_n28) );
  NAND2_X1 maj_177_U18 ( .A1(v_1_1[6]), .A2(maj_177_n28), .ZN(maj_177_n29) );
  NAND2_X1 maj_177_U17 ( .A1(maj_177_n26), .A2(maj_177_n27), .ZN(maj_177_n30)
         );
  NAND2_X1 maj_177_U16 ( .A1(maj_177_n30), .A2(maj_177_n29), .ZN(maj_177_n31)
         );
  NAND2_X1 maj_177_U15 ( .A1(v_1_1[5]), .A2(maj_177_n25), .ZN(maj_177_n18) );
  NAND2_X1 maj_177_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_177_n19) );
  NAND2_X1 maj_177_U13 ( .A1(maj_177_n19), .A2(maj_177_n18), .ZN(maj_177_n22)
         );
  NAND2_X1 maj_177_U12 ( .A1(v_1_1[2]), .A2(maj_177_n24), .ZN(maj_177_n20) );
  NAND2_X1 maj_177_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_177_n21) );
  NAND2_X1 maj_177_U10 ( .A1(maj_177_n21), .A2(maj_177_n20), .ZN(maj_177_n23)
         );
  XOR2_X1 maj_177_U9 ( .A(v_1_1[2]), .B(maj_177_n24), .Z(maj_177_n26) );
  XOR2_X1 maj_177_U8 ( .A(v_1_1[5]), .B(maj_177_n25), .Z(maj_177_n27) );
  XOR2_X1 maj_177_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_177_n24) );
  XOR2_X1 maj_177_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_177_n25) );
  OR2_X1 maj_177_U5 ( .A1(maj_177_n23), .A2(maj_177_n22), .ZN(maj_177_n32) );
  NAND2_X1 maj_177_U4 ( .A1(maj_177_n22), .A2(maj_177_n23), .ZN(maj_177_n34)
         );
  NAND2_X1 maj_177_U3 ( .A1(maj_177_n32), .A2(maj_177_n31), .ZN(maj_177_n33)
         );
  NAND2_X1 maj_177_U2 ( .A1(maj_177_n34), .A2(maj_177_n33), .ZN(maj_177_port_o) );
  OR2_X1 maj_178_U19 ( .A1(maj_178_n27), .A2(maj_178_n26), .ZN(maj_178_n28) );
  NAND2_X1 maj_178_U18 ( .A1(u_1_2[6]), .A2(maj_178_n28), .ZN(maj_178_n29) );
  NAND2_X1 maj_178_U17 ( .A1(maj_178_n26), .A2(maj_178_n27), .ZN(maj_178_n30)
         );
  NAND2_X1 maj_178_U16 ( .A1(maj_178_n30), .A2(maj_178_n29), .ZN(maj_178_n31)
         );
  NAND2_X1 maj_178_U15 ( .A1(u_1_2[5]), .A2(maj_178_n25), .ZN(maj_178_n18) );
  NAND2_X1 maj_178_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_178_n19) );
  NAND2_X1 maj_178_U13 ( .A1(maj_178_n19), .A2(maj_178_n18), .ZN(maj_178_n22)
         );
  NAND2_X1 maj_178_U12 ( .A1(u_1_2[2]), .A2(maj_178_n24), .ZN(maj_178_n20) );
  NAND2_X1 maj_178_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_178_n21) );
  NAND2_X1 maj_178_U10 ( .A1(maj_178_n21), .A2(maj_178_n20), .ZN(maj_178_n23)
         );
  XOR2_X1 maj_178_U9 ( .A(u_1_2[2]), .B(maj_178_n24), .Z(maj_178_n26) );
  XOR2_X1 maj_178_U8 ( .A(u_1_2[5]), .B(maj_178_n25), .Z(maj_178_n27) );
  XOR2_X1 maj_178_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_178_n24) );
  XOR2_X1 maj_178_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_178_n25) );
  OR2_X1 maj_178_U5 ( .A1(maj_178_n23), .A2(maj_178_n22), .ZN(maj_178_n32) );
  NAND2_X1 maj_178_U4 ( .A1(maj_178_n22), .A2(maj_178_n23), .ZN(maj_178_n34)
         );
  NAND2_X1 maj_178_U3 ( .A1(maj_178_n32), .A2(maj_178_n31), .ZN(maj_178_n33)
         );
  NAND2_X1 maj_178_U2 ( .A1(maj_178_n34), .A2(maj_178_n33), .ZN(maj_178_port_o) );
  OR2_X1 maj_179_U19 ( .A1(maj_179_n27), .A2(maj_179_n26), .ZN(maj_179_n28) );
  NAND2_X1 maj_179_U18 ( .A1(v_1_2[6]), .A2(maj_179_n28), .ZN(maj_179_n29) );
  NAND2_X1 maj_179_U17 ( .A1(maj_179_n26), .A2(maj_179_n27), .ZN(maj_179_n30)
         );
  NAND2_X1 maj_179_U16 ( .A1(maj_179_n30), .A2(maj_179_n29), .ZN(maj_179_n31)
         );
  NAND2_X1 maj_179_U15 ( .A1(v_1_2[5]), .A2(maj_179_n25), .ZN(maj_179_n18) );
  NAND2_X1 maj_179_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_179_n19) );
  NAND2_X1 maj_179_U13 ( .A1(maj_179_n19), .A2(maj_179_n18), .ZN(maj_179_n22)
         );
  NAND2_X1 maj_179_U12 ( .A1(v_1_2[2]), .A2(maj_179_n24), .ZN(maj_179_n20) );
  NAND2_X1 maj_179_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_179_n21) );
  NAND2_X1 maj_179_U10 ( .A1(maj_179_n21), .A2(maj_179_n20), .ZN(maj_179_n23)
         );
  XOR2_X1 maj_179_U9 ( .A(v_1_2[2]), .B(maj_179_n24), .Z(maj_179_n26) );
  XOR2_X1 maj_179_U8 ( .A(v_1_2[5]), .B(maj_179_n25), .Z(maj_179_n27) );
  XOR2_X1 maj_179_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_179_n24) );
  XOR2_X1 maj_179_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_179_n25) );
  OR2_X1 maj_179_U5 ( .A1(maj_179_n23), .A2(maj_179_n22), .ZN(maj_179_n32) );
  NAND2_X1 maj_179_U4 ( .A1(maj_179_n22), .A2(maj_179_n23), .ZN(maj_179_n34)
         );
  NAND2_X1 maj_179_U3 ( .A1(maj_179_n32), .A2(maj_179_n31), .ZN(maj_179_n33)
         );
  NAND2_X1 maj_179_U2 ( .A1(maj_179_n34), .A2(maj_179_n33), .ZN(maj_179_port_o) );
  OR2_X1 maj_180_U19 ( .A1(maj_180_n27), .A2(maj_180_n26), .ZN(maj_180_n28) );
  NAND2_X1 maj_180_U18 ( .A1(u_2_0[6]), .A2(maj_180_n28), .ZN(maj_180_n29) );
  NAND2_X1 maj_180_U17 ( .A1(maj_180_n26), .A2(maj_180_n27), .ZN(maj_180_n30)
         );
  NAND2_X1 maj_180_U16 ( .A1(maj_180_n30), .A2(maj_180_n29), .ZN(maj_180_n31)
         );
  NAND2_X1 maj_180_U15 ( .A1(u_2_0[5]), .A2(maj_180_n25), .ZN(maj_180_n18) );
  NAND2_X1 maj_180_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_180_n19) );
  NAND2_X1 maj_180_U13 ( .A1(maj_180_n19), .A2(maj_180_n18), .ZN(maj_180_n22)
         );
  NAND2_X1 maj_180_U12 ( .A1(u_2_0[2]), .A2(maj_180_n24), .ZN(maj_180_n20) );
  NAND2_X1 maj_180_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_180_n21) );
  NAND2_X1 maj_180_U10 ( .A1(maj_180_n21), .A2(maj_180_n20), .ZN(maj_180_n23)
         );
  XOR2_X1 maj_180_U9 ( .A(u_2_0[2]), .B(maj_180_n24), .Z(maj_180_n26) );
  XOR2_X1 maj_180_U8 ( .A(u_2_0[5]), .B(maj_180_n25), .Z(maj_180_n27) );
  XOR2_X1 maj_180_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_180_n24) );
  XOR2_X1 maj_180_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_180_n25) );
  OR2_X1 maj_180_U5 ( .A1(maj_180_n23), .A2(maj_180_n22), .ZN(maj_180_n32) );
  NAND2_X1 maj_180_U4 ( .A1(maj_180_n22), .A2(maj_180_n23), .ZN(maj_180_n34)
         );
  NAND2_X1 maj_180_U3 ( .A1(maj_180_n32), .A2(maj_180_n31), .ZN(maj_180_n33)
         );
  NAND2_X1 maj_180_U2 ( .A1(maj_180_n34), .A2(maj_180_n33), .ZN(maj_180_port_o) );
  OR2_X1 maj_181_U19 ( .A1(maj_181_n27), .A2(maj_181_n26), .ZN(maj_181_n28) );
  NAND2_X1 maj_181_U18 ( .A1(v_2_0[6]), .A2(maj_181_n28), .ZN(maj_181_n29) );
  NAND2_X1 maj_181_U17 ( .A1(maj_181_n26), .A2(maj_181_n27), .ZN(maj_181_n30)
         );
  NAND2_X1 maj_181_U16 ( .A1(maj_181_n30), .A2(maj_181_n29), .ZN(maj_181_n31)
         );
  NAND2_X1 maj_181_U15 ( .A1(v_2_0[5]), .A2(maj_181_n25), .ZN(maj_181_n18) );
  NAND2_X1 maj_181_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_181_n19) );
  NAND2_X1 maj_181_U13 ( .A1(maj_181_n19), .A2(maj_181_n18), .ZN(maj_181_n22)
         );
  NAND2_X1 maj_181_U12 ( .A1(v_2_0[2]), .A2(maj_181_n24), .ZN(maj_181_n20) );
  NAND2_X1 maj_181_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_181_n21) );
  NAND2_X1 maj_181_U10 ( .A1(maj_181_n21), .A2(maj_181_n20), .ZN(maj_181_n23)
         );
  XOR2_X1 maj_181_U9 ( .A(v_2_0[2]), .B(maj_181_n24), .Z(maj_181_n26) );
  XOR2_X1 maj_181_U8 ( .A(v_2_0[5]), .B(maj_181_n25), .Z(maj_181_n27) );
  XOR2_X1 maj_181_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_181_n24) );
  XOR2_X1 maj_181_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_181_n25) );
  OR2_X1 maj_181_U5 ( .A1(maj_181_n23), .A2(maj_181_n22), .ZN(maj_181_n32) );
  NAND2_X1 maj_181_U4 ( .A1(maj_181_n22), .A2(maj_181_n23), .ZN(maj_181_n34)
         );
  NAND2_X1 maj_181_U3 ( .A1(maj_181_n32), .A2(maj_181_n31), .ZN(maj_181_n33)
         );
  NAND2_X1 maj_181_U2 ( .A1(maj_181_n34), .A2(maj_181_n33), .ZN(maj_181_port_o) );
  OR2_X1 maj_182_U19 ( .A1(maj_182_n27), .A2(maj_182_n26), .ZN(maj_182_n28) );
  NAND2_X1 maj_182_U18 ( .A1(u_2_1[6]), .A2(maj_182_n28), .ZN(maj_182_n29) );
  NAND2_X1 maj_182_U17 ( .A1(maj_182_n26), .A2(maj_182_n27), .ZN(maj_182_n30)
         );
  NAND2_X1 maj_182_U16 ( .A1(maj_182_n30), .A2(maj_182_n29), .ZN(maj_182_n31)
         );
  NAND2_X1 maj_182_U15 ( .A1(u_2_1[5]), .A2(maj_182_n25), .ZN(maj_182_n18) );
  NAND2_X1 maj_182_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_182_n19) );
  NAND2_X1 maj_182_U13 ( .A1(maj_182_n19), .A2(maj_182_n18), .ZN(maj_182_n22)
         );
  NAND2_X1 maj_182_U12 ( .A1(u_2_1[2]), .A2(maj_182_n24), .ZN(maj_182_n20) );
  NAND2_X1 maj_182_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_182_n21) );
  NAND2_X1 maj_182_U10 ( .A1(maj_182_n21), .A2(maj_182_n20), .ZN(maj_182_n23)
         );
  XOR2_X1 maj_182_U9 ( .A(u_2_1[2]), .B(maj_182_n24), .Z(maj_182_n26) );
  XOR2_X1 maj_182_U8 ( .A(u_2_1[5]), .B(maj_182_n25), .Z(maj_182_n27) );
  XOR2_X1 maj_182_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_182_n24) );
  XOR2_X1 maj_182_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_182_n25) );
  OR2_X1 maj_182_U5 ( .A1(maj_182_n23), .A2(maj_182_n22), .ZN(maj_182_n32) );
  NAND2_X1 maj_182_U4 ( .A1(maj_182_n22), .A2(maj_182_n23), .ZN(maj_182_n34)
         );
  NAND2_X1 maj_182_U3 ( .A1(maj_182_n32), .A2(maj_182_n31), .ZN(maj_182_n33)
         );
  NAND2_X1 maj_182_U2 ( .A1(maj_182_n34), .A2(maj_182_n33), .ZN(maj_182_port_o) );
  OR2_X1 maj_183_U19 ( .A1(maj_183_n27), .A2(maj_183_n26), .ZN(maj_183_n28) );
  NAND2_X1 maj_183_U18 ( .A1(v_2_1[6]), .A2(maj_183_n28), .ZN(maj_183_n29) );
  NAND2_X1 maj_183_U17 ( .A1(maj_183_n26), .A2(maj_183_n27), .ZN(maj_183_n30)
         );
  NAND2_X1 maj_183_U16 ( .A1(maj_183_n30), .A2(maj_183_n29), .ZN(maj_183_n31)
         );
  NAND2_X1 maj_183_U15 ( .A1(v_2_1[5]), .A2(maj_183_n25), .ZN(maj_183_n18) );
  NAND2_X1 maj_183_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_183_n19) );
  NAND2_X1 maj_183_U13 ( .A1(maj_183_n19), .A2(maj_183_n18), .ZN(maj_183_n22)
         );
  NAND2_X1 maj_183_U12 ( .A1(v_2_1[2]), .A2(maj_183_n24), .ZN(maj_183_n20) );
  NAND2_X1 maj_183_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_183_n21) );
  NAND2_X1 maj_183_U10 ( .A1(maj_183_n21), .A2(maj_183_n20), .ZN(maj_183_n23)
         );
  XOR2_X1 maj_183_U9 ( .A(v_2_1[2]), .B(maj_183_n24), .Z(maj_183_n26) );
  XOR2_X1 maj_183_U8 ( .A(v_2_1[5]), .B(maj_183_n25), .Z(maj_183_n27) );
  XOR2_X1 maj_183_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_183_n24) );
  XOR2_X1 maj_183_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_183_n25) );
  OR2_X1 maj_183_U5 ( .A1(maj_183_n23), .A2(maj_183_n22), .ZN(maj_183_n32) );
  NAND2_X1 maj_183_U4 ( .A1(maj_183_n22), .A2(maj_183_n23), .ZN(maj_183_n34)
         );
  NAND2_X1 maj_183_U3 ( .A1(maj_183_n32), .A2(maj_183_n31), .ZN(maj_183_n33)
         );
  NAND2_X1 maj_183_U2 ( .A1(maj_183_n34), .A2(maj_183_n33), .ZN(maj_183_port_o) );
  OR2_X1 maj_184_U19 ( .A1(maj_184_n27), .A2(maj_184_n26), .ZN(maj_184_n28) );
  NAND2_X1 maj_184_U18 ( .A1(u_2_2[6]), .A2(maj_184_n28), .ZN(maj_184_n29) );
  NAND2_X1 maj_184_U17 ( .A1(maj_184_n26), .A2(maj_184_n27), .ZN(maj_184_n30)
         );
  NAND2_X1 maj_184_U16 ( .A1(maj_184_n30), .A2(maj_184_n29), .ZN(maj_184_n31)
         );
  NAND2_X1 maj_184_U15 ( .A1(u_2_2[5]), .A2(maj_184_n25), .ZN(maj_184_n18) );
  NAND2_X1 maj_184_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_184_n19) );
  NAND2_X1 maj_184_U13 ( .A1(maj_184_n19), .A2(maj_184_n18), .ZN(maj_184_n22)
         );
  NAND2_X1 maj_184_U12 ( .A1(u_2_2[2]), .A2(maj_184_n24), .ZN(maj_184_n20) );
  NAND2_X1 maj_184_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_184_n21) );
  NAND2_X1 maj_184_U10 ( .A1(maj_184_n21), .A2(maj_184_n20), .ZN(maj_184_n23)
         );
  XOR2_X1 maj_184_U9 ( .A(u_2_2[2]), .B(maj_184_n24), .Z(maj_184_n26) );
  XOR2_X1 maj_184_U8 ( .A(u_2_2[5]), .B(maj_184_n25), .Z(maj_184_n27) );
  XOR2_X1 maj_184_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_184_n24) );
  XOR2_X1 maj_184_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_184_n25) );
  OR2_X1 maj_184_U5 ( .A1(maj_184_n23), .A2(maj_184_n22), .ZN(maj_184_n32) );
  NAND2_X1 maj_184_U4 ( .A1(maj_184_n22), .A2(maj_184_n23), .ZN(maj_184_n34)
         );
  NAND2_X1 maj_184_U3 ( .A1(maj_184_n32), .A2(maj_184_n31), .ZN(maj_184_n33)
         );
  NAND2_X1 maj_184_U2 ( .A1(maj_184_n34), .A2(maj_184_n33), .ZN(maj_184_port_o) );
  OR2_X1 maj_185_U19 ( .A1(maj_185_n27), .A2(maj_185_n26), .ZN(maj_185_n28) );
  NAND2_X1 maj_185_U18 ( .A1(v_2_2[6]), .A2(maj_185_n28), .ZN(maj_185_n29) );
  NAND2_X1 maj_185_U17 ( .A1(maj_185_n26), .A2(maj_185_n27), .ZN(maj_185_n30)
         );
  NAND2_X1 maj_185_U16 ( .A1(maj_185_n30), .A2(maj_185_n29), .ZN(maj_185_n31)
         );
  NAND2_X1 maj_185_U15 ( .A1(v_2_2[5]), .A2(maj_185_n25), .ZN(maj_185_n18) );
  NAND2_X1 maj_185_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_185_n19) );
  NAND2_X1 maj_185_U13 ( .A1(maj_185_n19), .A2(maj_185_n18), .ZN(maj_185_n22)
         );
  NAND2_X1 maj_185_U12 ( .A1(v_2_2[2]), .A2(maj_185_n24), .ZN(maj_185_n20) );
  NAND2_X1 maj_185_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_185_n21) );
  NAND2_X1 maj_185_U10 ( .A1(maj_185_n21), .A2(maj_185_n20), .ZN(maj_185_n23)
         );
  XOR2_X1 maj_185_U9 ( .A(v_2_2[2]), .B(maj_185_n24), .Z(maj_185_n26) );
  XOR2_X1 maj_185_U8 ( .A(v_2_2[5]), .B(maj_185_n25), .Z(maj_185_n27) );
  XOR2_X1 maj_185_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_185_n24) );
  XOR2_X1 maj_185_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_185_n25) );
  OR2_X1 maj_185_U5 ( .A1(maj_185_n23), .A2(maj_185_n22), .ZN(maj_185_n32) );
  NAND2_X1 maj_185_U4 ( .A1(maj_185_n22), .A2(maj_185_n23), .ZN(maj_185_n34)
         );
  NAND2_X1 maj_185_U3 ( .A1(maj_185_n32), .A2(maj_185_n31), .ZN(maj_185_n33)
         );
  NAND2_X1 maj_185_U2 ( .A1(maj_185_n34), .A2(maj_185_n33), .ZN(maj_185_port_o) );
  OR2_X1 maj_186_U19 ( .A1(maj_186_n27), .A2(maj_186_n26), .ZN(maj_186_n28) );
  NAND2_X1 maj_186_U18 ( .A1(u_3_0[6]), .A2(maj_186_n28), .ZN(maj_186_n29) );
  NAND2_X1 maj_186_U17 ( .A1(maj_186_n26), .A2(maj_186_n27), .ZN(maj_186_n30)
         );
  NAND2_X1 maj_186_U16 ( .A1(maj_186_n30), .A2(maj_186_n29), .ZN(maj_186_n31)
         );
  NAND2_X1 maj_186_U15 ( .A1(u_3_0[5]), .A2(maj_186_n25), .ZN(maj_186_n18) );
  NAND2_X1 maj_186_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_186_n19) );
  NAND2_X1 maj_186_U13 ( .A1(maj_186_n19), .A2(maj_186_n18), .ZN(maj_186_n22)
         );
  NAND2_X1 maj_186_U12 ( .A1(u_3_0[2]), .A2(maj_186_n24), .ZN(maj_186_n20) );
  NAND2_X1 maj_186_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_186_n21) );
  NAND2_X1 maj_186_U10 ( .A1(maj_186_n21), .A2(maj_186_n20), .ZN(maj_186_n23)
         );
  XOR2_X1 maj_186_U9 ( .A(u_3_0[2]), .B(maj_186_n24), .Z(maj_186_n26) );
  XOR2_X1 maj_186_U8 ( .A(u_3_0[5]), .B(maj_186_n25), .Z(maj_186_n27) );
  XOR2_X1 maj_186_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_186_n24) );
  XOR2_X1 maj_186_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_186_n25) );
  OR2_X1 maj_186_U5 ( .A1(maj_186_n23), .A2(maj_186_n22), .ZN(maj_186_n32) );
  NAND2_X1 maj_186_U4 ( .A1(maj_186_n22), .A2(maj_186_n23), .ZN(maj_186_n34)
         );
  NAND2_X1 maj_186_U3 ( .A1(maj_186_n32), .A2(maj_186_n31), .ZN(maj_186_n33)
         );
  NAND2_X1 maj_186_U2 ( .A1(maj_186_n34), .A2(maj_186_n33), .ZN(maj_186_port_o) );
  OR2_X1 maj_187_U19 ( .A1(maj_187_n27), .A2(maj_187_n26), .ZN(maj_187_n28) );
  NAND2_X1 maj_187_U18 ( .A1(v_3_0[6]), .A2(maj_187_n28), .ZN(maj_187_n29) );
  NAND2_X1 maj_187_U17 ( .A1(maj_187_n26), .A2(maj_187_n27), .ZN(maj_187_n30)
         );
  NAND2_X1 maj_187_U16 ( .A1(maj_187_n30), .A2(maj_187_n29), .ZN(maj_187_n31)
         );
  NAND2_X1 maj_187_U15 ( .A1(v_3_0[5]), .A2(maj_187_n25), .ZN(maj_187_n18) );
  NAND2_X1 maj_187_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_187_n19) );
  NAND2_X1 maj_187_U13 ( .A1(maj_187_n19), .A2(maj_187_n18), .ZN(maj_187_n22)
         );
  NAND2_X1 maj_187_U12 ( .A1(v_3_0[2]), .A2(maj_187_n24), .ZN(maj_187_n20) );
  NAND2_X1 maj_187_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_187_n21) );
  NAND2_X1 maj_187_U10 ( .A1(maj_187_n21), .A2(maj_187_n20), .ZN(maj_187_n23)
         );
  XOR2_X1 maj_187_U9 ( .A(v_3_0[2]), .B(maj_187_n24), .Z(maj_187_n26) );
  XOR2_X1 maj_187_U8 ( .A(v_3_0[5]), .B(maj_187_n25), .Z(maj_187_n27) );
  XOR2_X1 maj_187_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_187_n24) );
  XOR2_X1 maj_187_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_187_n25) );
  OR2_X1 maj_187_U5 ( .A1(maj_187_n23), .A2(maj_187_n22), .ZN(maj_187_n32) );
  NAND2_X1 maj_187_U4 ( .A1(maj_187_n22), .A2(maj_187_n23), .ZN(maj_187_n34)
         );
  NAND2_X1 maj_187_U3 ( .A1(maj_187_n32), .A2(maj_187_n31), .ZN(maj_187_n33)
         );
  NAND2_X1 maj_187_U2 ( .A1(maj_187_n34), .A2(maj_187_n33), .ZN(maj_187_port_o) );
  OR2_X1 maj_188_U19 ( .A1(maj_188_n27), .A2(maj_188_n26), .ZN(maj_188_n28) );
  NAND2_X1 maj_188_U18 ( .A1(u_3_1[6]), .A2(maj_188_n28), .ZN(maj_188_n29) );
  NAND2_X1 maj_188_U17 ( .A1(maj_188_n26), .A2(maj_188_n27), .ZN(maj_188_n30)
         );
  NAND2_X1 maj_188_U16 ( .A1(maj_188_n30), .A2(maj_188_n29), .ZN(maj_188_n31)
         );
  NAND2_X1 maj_188_U15 ( .A1(u_3_1[5]), .A2(maj_188_n25), .ZN(maj_188_n18) );
  NAND2_X1 maj_188_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_188_n19) );
  NAND2_X1 maj_188_U13 ( .A1(maj_188_n19), .A2(maj_188_n18), .ZN(maj_188_n22)
         );
  NAND2_X1 maj_188_U12 ( .A1(u_3_1[2]), .A2(maj_188_n24), .ZN(maj_188_n20) );
  NAND2_X1 maj_188_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_188_n21) );
  NAND2_X1 maj_188_U10 ( .A1(maj_188_n21), .A2(maj_188_n20), .ZN(maj_188_n23)
         );
  XOR2_X1 maj_188_U9 ( .A(u_3_1[2]), .B(maj_188_n24), .Z(maj_188_n26) );
  XOR2_X1 maj_188_U8 ( .A(u_3_1[5]), .B(maj_188_n25), .Z(maj_188_n27) );
  XOR2_X1 maj_188_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_188_n24) );
  XOR2_X1 maj_188_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_188_n25) );
  OR2_X1 maj_188_U5 ( .A1(maj_188_n23), .A2(maj_188_n22), .ZN(maj_188_n32) );
  NAND2_X1 maj_188_U4 ( .A1(maj_188_n22), .A2(maj_188_n23), .ZN(maj_188_n34)
         );
  NAND2_X1 maj_188_U3 ( .A1(maj_188_n32), .A2(maj_188_n31), .ZN(maj_188_n33)
         );
  NAND2_X1 maj_188_U2 ( .A1(maj_188_n34), .A2(maj_188_n33), .ZN(maj_188_port_o) );
  OR2_X1 maj_189_U19 ( .A1(maj_189_n27), .A2(maj_189_n26), .ZN(maj_189_n28) );
  NAND2_X1 maj_189_U18 ( .A1(v_3_1[6]), .A2(maj_189_n28), .ZN(maj_189_n29) );
  NAND2_X1 maj_189_U17 ( .A1(maj_189_n26), .A2(maj_189_n27), .ZN(maj_189_n30)
         );
  NAND2_X1 maj_189_U16 ( .A1(maj_189_n30), .A2(maj_189_n29), .ZN(maj_189_n31)
         );
  NAND2_X1 maj_189_U15 ( .A1(v_3_1[5]), .A2(maj_189_n25), .ZN(maj_189_n18) );
  NAND2_X1 maj_189_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_189_n19) );
  NAND2_X1 maj_189_U13 ( .A1(maj_189_n19), .A2(maj_189_n18), .ZN(maj_189_n22)
         );
  NAND2_X1 maj_189_U12 ( .A1(v_3_1[2]), .A2(maj_189_n24), .ZN(maj_189_n20) );
  NAND2_X1 maj_189_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_189_n21) );
  NAND2_X1 maj_189_U10 ( .A1(maj_189_n21), .A2(maj_189_n20), .ZN(maj_189_n23)
         );
  XOR2_X1 maj_189_U9 ( .A(v_3_1[2]), .B(maj_189_n24), .Z(maj_189_n26) );
  XOR2_X1 maj_189_U8 ( .A(v_3_1[5]), .B(maj_189_n25), .Z(maj_189_n27) );
  XOR2_X1 maj_189_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_189_n24) );
  XOR2_X1 maj_189_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_189_n25) );
  OR2_X1 maj_189_U5 ( .A1(maj_189_n23), .A2(maj_189_n22), .ZN(maj_189_n32) );
  NAND2_X1 maj_189_U4 ( .A1(maj_189_n22), .A2(maj_189_n23), .ZN(maj_189_n34)
         );
  NAND2_X1 maj_189_U3 ( .A1(maj_189_n32), .A2(maj_189_n31), .ZN(maj_189_n33)
         );
  NAND2_X1 maj_189_U2 ( .A1(maj_189_n34), .A2(maj_189_n33), .ZN(maj_189_port_o) );
  OR2_X1 maj_190_U19 ( .A1(maj_190_n27), .A2(maj_190_n26), .ZN(maj_190_n28) );
  NAND2_X1 maj_190_U18 ( .A1(u_3_2[6]), .A2(maj_190_n28), .ZN(maj_190_n29) );
  NAND2_X1 maj_190_U17 ( .A1(maj_190_n26), .A2(maj_190_n27), .ZN(maj_190_n30)
         );
  NAND2_X1 maj_190_U16 ( .A1(maj_190_n30), .A2(maj_190_n29), .ZN(maj_190_n31)
         );
  NAND2_X1 maj_190_U15 ( .A1(u_3_2[5]), .A2(maj_190_n25), .ZN(maj_190_n18) );
  NAND2_X1 maj_190_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_190_n19) );
  NAND2_X1 maj_190_U13 ( .A1(maj_190_n19), .A2(maj_190_n18), .ZN(maj_190_n22)
         );
  NAND2_X1 maj_190_U12 ( .A1(u_3_2[2]), .A2(maj_190_n24), .ZN(maj_190_n20) );
  NAND2_X1 maj_190_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_190_n21) );
  NAND2_X1 maj_190_U10 ( .A1(maj_190_n21), .A2(maj_190_n20), .ZN(maj_190_n23)
         );
  XOR2_X1 maj_190_U9 ( .A(u_3_2[2]), .B(maj_190_n24), .Z(maj_190_n26) );
  XOR2_X1 maj_190_U8 ( .A(u_3_2[5]), .B(maj_190_n25), .Z(maj_190_n27) );
  XOR2_X1 maj_190_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_190_n24) );
  XOR2_X1 maj_190_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_190_n25) );
  OR2_X1 maj_190_U5 ( .A1(maj_190_n23), .A2(maj_190_n22), .ZN(maj_190_n32) );
  NAND2_X1 maj_190_U4 ( .A1(maj_190_n22), .A2(maj_190_n23), .ZN(maj_190_n34)
         );
  NAND2_X1 maj_190_U3 ( .A1(maj_190_n32), .A2(maj_190_n31), .ZN(maj_190_n33)
         );
  NAND2_X1 maj_190_U2 ( .A1(maj_190_n34), .A2(maj_190_n33), .ZN(maj_190_port_o) );
  OR2_X1 maj_191_U19 ( .A1(maj_191_n27), .A2(maj_191_n26), .ZN(maj_191_n28) );
  NAND2_X1 maj_191_U18 ( .A1(v_3_2[6]), .A2(maj_191_n28), .ZN(maj_191_n29) );
  NAND2_X1 maj_191_U17 ( .A1(maj_191_n26), .A2(maj_191_n27), .ZN(maj_191_n30)
         );
  NAND2_X1 maj_191_U16 ( .A1(maj_191_n30), .A2(maj_191_n29), .ZN(maj_191_n31)
         );
  NAND2_X1 maj_191_U15 ( .A1(v_3_2[5]), .A2(maj_191_n25), .ZN(maj_191_n18) );
  NAND2_X1 maj_191_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_191_n19) );
  NAND2_X1 maj_191_U13 ( .A1(maj_191_n19), .A2(maj_191_n18), .ZN(maj_191_n22)
         );
  NAND2_X1 maj_191_U12 ( .A1(v_3_2[2]), .A2(maj_191_n24), .ZN(maj_191_n20) );
  NAND2_X1 maj_191_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_191_n21) );
  NAND2_X1 maj_191_U10 ( .A1(maj_191_n21), .A2(maj_191_n20), .ZN(maj_191_n23)
         );
  XOR2_X1 maj_191_U9 ( .A(v_3_2[2]), .B(maj_191_n24), .Z(maj_191_n26) );
  XOR2_X1 maj_191_U8 ( .A(v_3_2[5]), .B(maj_191_n25), .Z(maj_191_n27) );
  XOR2_X1 maj_191_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_191_n24) );
  XOR2_X1 maj_191_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_191_n25) );
  OR2_X1 maj_191_U5 ( .A1(maj_191_n23), .A2(maj_191_n22), .ZN(maj_191_n32) );
  NAND2_X1 maj_191_U4 ( .A1(maj_191_n22), .A2(maj_191_n23), .ZN(maj_191_n34)
         );
  NAND2_X1 maj_191_U3 ( .A1(maj_191_n32), .A2(maj_191_n31), .ZN(maj_191_n33)
         );
  NAND2_X1 maj_191_U2 ( .A1(maj_191_n34), .A2(maj_191_n33), .ZN(maj_191_port_o) );
  OR2_X1 maj_192_U19 ( .A1(maj_192_n27), .A2(maj_192_n26), .ZN(maj_192_n28) );
  NAND2_X1 maj_192_U18 ( .A1(u_0_0[6]), .A2(maj_192_n28), .ZN(maj_192_n29) );
  NAND2_X1 maj_192_U17 ( .A1(maj_192_n26), .A2(maj_192_n27), .ZN(maj_192_n30)
         );
  NAND2_X1 maj_192_U16 ( .A1(maj_192_n30), .A2(maj_192_n29), .ZN(maj_192_n31)
         );
  NAND2_X1 maj_192_U15 ( .A1(u_0_0[5]), .A2(maj_192_n25), .ZN(maj_192_n18) );
  NAND2_X1 maj_192_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_192_n19) );
  NAND2_X1 maj_192_U13 ( .A1(maj_192_n19), .A2(maj_192_n18), .ZN(maj_192_n22)
         );
  NAND2_X1 maj_192_U12 ( .A1(u_0_0[2]), .A2(maj_192_n24), .ZN(maj_192_n20) );
  NAND2_X1 maj_192_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_192_n21) );
  NAND2_X1 maj_192_U10 ( .A1(maj_192_n21), .A2(maj_192_n20), .ZN(maj_192_n23)
         );
  XOR2_X1 maj_192_U9 ( .A(u_0_0[2]), .B(maj_192_n24), .Z(maj_192_n26) );
  XOR2_X1 maj_192_U8 ( .A(u_0_0[5]), .B(maj_192_n25), .Z(maj_192_n27) );
  XOR2_X1 maj_192_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_192_n24) );
  XOR2_X1 maj_192_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_192_n25) );
  OR2_X1 maj_192_U5 ( .A1(maj_192_n23), .A2(maj_192_n22), .ZN(maj_192_n32) );
  NAND2_X1 maj_192_U4 ( .A1(maj_192_n22), .A2(maj_192_n23), .ZN(maj_192_n34)
         );
  NAND2_X1 maj_192_U3 ( .A1(maj_192_n32), .A2(maj_192_n31), .ZN(maj_192_n33)
         );
  NAND2_X1 maj_192_U2 ( .A1(maj_192_n34), .A2(maj_192_n33), .ZN(maj_192_port_o) );
  OR2_X1 maj_193_U19 ( .A1(maj_193_n27), .A2(maj_193_n26), .ZN(maj_193_n28) );
  NAND2_X1 maj_193_U18 ( .A1(v_0_0[6]), .A2(maj_193_n28), .ZN(maj_193_n29) );
  NAND2_X1 maj_193_U17 ( .A1(maj_193_n26), .A2(maj_193_n27), .ZN(maj_193_n30)
         );
  NAND2_X1 maj_193_U16 ( .A1(maj_193_n30), .A2(maj_193_n29), .ZN(maj_193_n31)
         );
  NAND2_X1 maj_193_U15 ( .A1(v_0_0[5]), .A2(maj_193_n25), .ZN(maj_193_n18) );
  NAND2_X1 maj_193_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_193_n19) );
  NAND2_X1 maj_193_U13 ( .A1(maj_193_n19), .A2(maj_193_n18), .ZN(maj_193_n22)
         );
  NAND2_X1 maj_193_U12 ( .A1(v_0_0[2]), .A2(maj_193_n24), .ZN(maj_193_n20) );
  NAND2_X1 maj_193_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_193_n21) );
  NAND2_X1 maj_193_U10 ( .A1(maj_193_n21), .A2(maj_193_n20), .ZN(maj_193_n23)
         );
  XOR2_X1 maj_193_U9 ( .A(v_0_0[2]), .B(maj_193_n24), .Z(maj_193_n26) );
  XOR2_X1 maj_193_U8 ( .A(v_0_0[5]), .B(maj_193_n25), .Z(maj_193_n27) );
  XOR2_X1 maj_193_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_193_n24) );
  XOR2_X1 maj_193_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_193_n25) );
  OR2_X1 maj_193_U5 ( .A1(maj_193_n23), .A2(maj_193_n22), .ZN(maj_193_n32) );
  NAND2_X1 maj_193_U4 ( .A1(maj_193_n22), .A2(maj_193_n23), .ZN(maj_193_n34)
         );
  NAND2_X1 maj_193_U3 ( .A1(maj_193_n32), .A2(maj_193_n31), .ZN(maj_193_n33)
         );
  NAND2_X1 maj_193_U2 ( .A1(maj_193_n34), .A2(maj_193_n33), .ZN(maj_193_port_o) );
  OR2_X1 maj_194_U19 ( .A1(maj_194_n27), .A2(maj_194_n26), .ZN(maj_194_n28) );
  NAND2_X1 maj_194_U18 ( .A1(u_0_1[6]), .A2(maj_194_n28), .ZN(maj_194_n29) );
  NAND2_X1 maj_194_U17 ( .A1(maj_194_n26), .A2(maj_194_n27), .ZN(maj_194_n30)
         );
  NAND2_X1 maj_194_U16 ( .A1(maj_194_n30), .A2(maj_194_n29), .ZN(maj_194_n31)
         );
  NAND2_X1 maj_194_U15 ( .A1(u_0_1[5]), .A2(maj_194_n25), .ZN(maj_194_n18) );
  NAND2_X1 maj_194_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_194_n19) );
  NAND2_X1 maj_194_U13 ( .A1(maj_194_n19), .A2(maj_194_n18), .ZN(maj_194_n22)
         );
  NAND2_X1 maj_194_U12 ( .A1(u_0_1[2]), .A2(maj_194_n24), .ZN(maj_194_n20) );
  NAND2_X1 maj_194_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_194_n21) );
  NAND2_X1 maj_194_U10 ( .A1(maj_194_n21), .A2(maj_194_n20), .ZN(maj_194_n23)
         );
  XOR2_X1 maj_194_U9 ( .A(u_0_1[2]), .B(maj_194_n24), .Z(maj_194_n26) );
  XOR2_X1 maj_194_U8 ( .A(u_0_1[5]), .B(maj_194_n25), .Z(maj_194_n27) );
  XOR2_X1 maj_194_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_194_n24) );
  XOR2_X1 maj_194_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_194_n25) );
  OR2_X1 maj_194_U5 ( .A1(maj_194_n23), .A2(maj_194_n22), .ZN(maj_194_n32) );
  NAND2_X1 maj_194_U4 ( .A1(maj_194_n22), .A2(maj_194_n23), .ZN(maj_194_n34)
         );
  NAND2_X1 maj_194_U3 ( .A1(maj_194_n32), .A2(maj_194_n31), .ZN(maj_194_n33)
         );
  NAND2_X1 maj_194_U2 ( .A1(maj_194_n34), .A2(maj_194_n33), .ZN(maj_194_port_o) );
  OR2_X1 maj_195_U19 ( .A1(maj_195_n27), .A2(maj_195_n26), .ZN(maj_195_n28) );
  NAND2_X1 maj_195_U18 ( .A1(v_0_1[6]), .A2(maj_195_n28), .ZN(maj_195_n29) );
  NAND2_X1 maj_195_U17 ( .A1(maj_195_n26), .A2(maj_195_n27), .ZN(maj_195_n30)
         );
  NAND2_X1 maj_195_U16 ( .A1(maj_195_n30), .A2(maj_195_n29), .ZN(maj_195_n31)
         );
  NAND2_X1 maj_195_U15 ( .A1(v_0_1[5]), .A2(maj_195_n25), .ZN(maj_195_n18) );
  NAND2_X1 maj_195_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_195_n19) );
  NAND2_X1 maj_195_U13 ( .A1(maj_195_n19), .A2(maj_195_n18), .ZN(maj_195_n22)
         );
  NAND2_X1 maj_195_U12 ( .A1(v_0_1[2]), .A2(maj_195_n24), .ZN(maj_195_n20) );
  NAND2_X1 maj_195_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_195_n21) );
  NAND2_X1 maj_195_U10 ( .A1(maj_195_n21), .A2(maj_195_n20), .ZN(maj_195_n23)
         );
  XOR2_X1 maj_195_U9 ( .A(v_0_1[2]), .B(maj_195_n24), .Z(maj_195_n26) );
  XOR2_X1 maj_195_U8 ( .A(v_0_1[5]), .B(maj_195_n25), .Z(maj_195_n27) );
  XOR2_X1 maj_195_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_195_n24) );
  XOR2_X1 maj_195_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_195_n25) );
  OR2_X1 maj_195_U5 ( .A1(maj_195_n23), .A2(maj_195_n22), .ZN(maj_195_n32) );
  NAND2_X1 maj_195_U4 ( .A1(maj_195_n22), .A2(maj_195_n23), .ZN(maj_195_n34)
         );
  NAND2_X1 maj_195_U3 ( .A1(maj_195_n32), .A2(maj_195_n31), .ZN(maj_195_n33)
         );
  NAND2_X1 maj_195_U2 ( .A1(maj_195_n34), .A2(maj_195_n33), .ZN(maj_195_port_o) );
  OR2_X1 maj_196_U19 ( .A1(maj_196_n27), .A2(maj_196_n26), .ZN(maj_196_n28) );
  NAND2_X1 maj_196_U18 ( .A1(u_0_2[6]), .A2(maj_196_n28), .ZN(maj_196_n29) );
  NAND2_X1 maj_196_U17 ( .A1(maj_196_n26), .A2(maj_196_n27), .ZN(maj_196_n30)
         );
  NAND2_X1 maj_196_U16 ( .A1(maj_196_n30), .A2(maj_196_n29), .ZN(maj_196_n31)
         );
  NAND2_X1 maj_196_U15 ( .A1(u_0_2[5]), .A2(maj_196_n25), .ZN(maj_196_n18) );
  NAND2_X1 maj_196_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_196_n19) );
  NAND2_X1 maj_196_U13 ( .A1(maj_196_n19), .A2(maj_196_n18), .ZN(maj_196_n22)
         );
  NAND2_X1 maj_196_U12 ( .A1(u_0_2[2]), .A2(maj_196_n24), .ZN(maj_196_n20) );
  NAND2_X1 maj_196_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_196_n21) );
  NAND2_X1 maj_196_U10 ( .A1(maj_196_n21), .A2(maj_196_n20), .ZN(maj_196_n23)
         );
  XOR2_X1 maj_196_U9 ( .A(u_0_2[2]), .B(maj_196_n24), .Z(maj_196_n26) );
  XOR2_X1 maj_196_U8 ( .A(u_0_2[5]), .B(maj_196_n25), .Z(maj_196_n27) );
  XOR2_X1 maj_196_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_196_n24) );
  XOR2_X1 maj_196_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_196_n25) );
  OR2_X1 maj_196_U5 ( .A1(maj_196_n23), .A2(maj_196_n22), .ZN(maj_196_n32) );
  NAND2_X1 maj_196_U4 ( .A1(maj_196_n22), .A2(maj_196_n23), .ZN(maj_196_n34)
         );
  NAND2_X1 maj_196_U3 ( .A1(maj_196_n32), .A2(maj_196_n31), .ZN(maj_196_n33)
         );
  NAND2_X1 maj_196_U2 ( .A1(maj_196_n34), .A2(maj_196_n33), .ZN(maj_196_port_o) );
  OR2_X1 maj_197_U19 ( .A1(maj_197_n27), .A2(maj_197_n26), .ZN(maj_197_n28) );
  NAND2_X1 maj_197_U18 ( .A1(v_0_2[6]), .A2(maj_197_n28), .ZN(maj_197_n29) );
  NAND2_X1 maj_197_U17 ( .A1(maj_197_n26), .A2(maj_197_n27), .ZN(maj_197_n30)
         );
  NAND2_X1 maj_197_U16 ( .A1(maj_197_n30), .A2(maj_197_n29), .ZN(maj_197_n31)
         );
  NAND2_X1 maj_197_U15 ( .A1(v_0_2[5]), .A2(maj_197_n25), .ZN(maj_197_n18) );
  NAND2_X1 maj_197_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_197_n19) );
  NAND2_X1 maj_197_U13 ( .A1(maj_197_n19), .A2(maj_197_n18), .ZN(maj_197_n22)
         );
  NAND2_X1 maj_197_U12 ( .A1(v_0_2[2]), .A2(maj_197_n24), .ZN(maj_197_n20) );
  NAND2_X1 maj_197_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_197_n21) );
  NAND2_X1 maj_197_U10 ( .A1(maj_197_n21), .A2(maj_197_n20), .ZN(maj_197_n23)
         );
  XOR2_X1 maj_197_U9 ( .A(v_0_2[2]), .B(maj_197_n24), .Z(maj_197_n26) );
  XOR2_X1 maj_197_U8 ( .A(v_0_2[5]), .B(maj_197_n25), .Z(maj_197_n27) );
  XOR2_X1 maj_197_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_197_n24) );
  XOR2_X1 maj_197_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_197_n25) );
  OR2_X1 maj_197_U5 ( .A1(maj_197_n23), .A2(maj_197_n22), .ZN(maj_197_n32) );
  NAND2_X1 maj_197_U4 ( .A1(maj_197_n22), .A2(maj_197_n23), .ZN(maj_197_n34)
         );
  NAND2_X1 maj_197_U3 ( .A1(maj_197_n32), .A2(maj_197_n31), .ZN(maj_197_n33)
         );
  NAND2_X1 maj_197_U2 ( .A1(maj_197_n34), .A2(maj_197_n33), .ZN(maj_197_port_o) );
  OR2_X1 maj_198_U19 ( .A1(maj_198_n27), .A2(maj_198_n26), .ZN(maj_198_n28) );
  NAND2_X1 maj_198_U18 ( .A1(u_1_0[6]), .A2(maj_198_n28), .ZN(maj_198_n29) );
  NAND2_X1 maj_198_U17 ( .A1(maj_198_n26), .A2(maj_198_n27), .ZN(maj_198_n30)
         );
  NAND2_X1 maj_198_U16 ( .A1(maj_198_n30), .A2(maj_198_n29), .ZN(maj_198_n31)
         );
  NAND2_X1 maj_198_U15 ( .A1(u_1_0[5]), .A2(maj_198_n25), .ZN(maj_198_n18) );
  NAND2_X1 maj_198_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_198_n19) );
  NAND2_X1 maj_198_U13 ( .A1(maj_198_n19), .A2(maj_198_n18), .ZN(maj_198_n22)
         );
  NAND2_X1 maj_198_U12 ( .A1(u_1_0[2]), .A2(maj_198_n24), .ZN(maj_198_n20) );
  NAND2_X1 maj_198_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_198_n21) );
  NAND2_X1 maj_198_U10 ( .A1(maj_198_n21), .A2(maj_198_n20), .ZN(maj_198_n23)
         );
  XOR2_X1 maj_198_U9 ( .A(u_1_0[2]), .B(maj_198_n24), .Z(maj_198_n26) );
  XOR2_X1 maj_198_U8 ( .A(u_1_0[5]), .B(maj_198_n25), .Z(maj_198_n27) );
  XOR2_X1 maj_198_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_198_n24) );
  XOR2_X1 maj_198_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_198_n25) );
  OR2_X1 maj_198_U5 ( .A1(maj_198_n23), .A2(maj_198_n22), .ZN(maj_198_n32) );
  NAND2_X1 maj_198_U4 ( .A1(maj_198_n22), .A2(maj_198_n23), .ZN(maj_198_n34)
         );
  NAND2_X1 maj_198_U3 ( .A1(maj_198_n32), .A2(maj_198_n31), .ZN(maj_198_n33)
         );
  NAND2_X1 maj_198_U2 ( .A1(maj_198_n34), .A2(maj_198_n33), .ZN(maj_198_port_o) );
  OR2_X1 maj_199_U19 ( .A1(maj_199_n27), .A2(maj_199_n26), .ZN(maj_199_n28) );
  NAND2_X1 maj_199_U18 ( .A1(v_1_0[6]), .A2(maj_199_n28), .ZN(maj_199_n29) );
  NAND2_X1 maj_199_U17 ( .A1(maj_199_n26), .A2(maj_199_n27), .ZN(maj_199_n30)
         );
  NAND2_X1 maj_199_U16 ( .A1(maj_199_n30), .A2(maj_199_n29), .ZN(maj_199_n31)
         );
  NAND2_X1 maj_199_U15 ( .A1(v_1_0[5]), .A2(maj_199_n25), .ZN(maj_199_n18) );
  NAND2_X1 maj_199_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_199_n19) );
  NAND2_X1 maj_199_U13 ( .A1(maj_199_n19), .A2(maj_199_n18), .ZN(maj_199_n22)
         );
  NAND2_X1 maj_199_U12 ( .A1(v_1_0[2]), .A2(maj_199_n24), .ZN(maj_199_n20) );
  NAND2_X1 maj_199_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_199_n21) );
  NAND2_X1 maj_199_U10 ( .A1(maj_199_n21), .A2(maj_199_n20), .ZN(maj_199_n23)
         );
  XOR2_X1 maj_199_U9 ( .A(v_1_0[2]), .B(maj_199_n24), .Z(maj_199_n26) );
  XOR2_X1 maj_199_U8 ( .A(v_1_0[5]), .B(maj_199_n25), .Z(maj_199_n27) );
  XOR2_X1 maj_199_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_199_n24) );
  XOR2_X1 maj_199_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_199_n25) );
  OR2_X1 maj_199_U5 ( .A1(maj_199_n23), .A2(maj_199_n22), .ZN(maj_199_n32) );
  NAND2_X1 maj_199_U4 ( .A1(maj_199_n22), .A2(maj_199_n23), .ZN(maj_199_n34)
         );
  NAND2_X1 maj_199_U3 ( .A1(maj_199_n32), .A2(maj_199_n31), .ZN(maj_199_n33)
         );
  NAND2_X1 maj_199_U2 ( .A1(maj_199_n34), .A2(maj_199_n33), .ZN(maj_199_port_o) );
  OR2_X1 maj_200_U19 ( .A1(maj_200_n27), .A2(maj_200_n26), .ZN(maj_200_n28) );
  NAND2_X1 maj_200_U18 ( .A1(u_1_1[6]), .A2(maj_200_n28), .ZN(maj_200_n29) );
  NAND2_X1 maj_200_U17 ( .A1(maj_200_n26), .A2(maj_200_n27), .ZN(maj_200_n30)
         );
  NAND2_X1 maj_200_U16 ( .A1(maj_200_n30), .A2(maj_200_n29), .ZN(maj_200_n31)
         );
  NAND2_X1 maj_200_U15 ( .A1(u_1_1[5]), .A2(maj_200_n25), .ZN(maj_200_n18) );
  NAND2_X1 maj_200_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_200_n19) );
  NAND2_X1 maj_200_U13 ( .A1(maj_200_n19), .A2(maj_200_n18), .ZN(maj_200_n22)
         );
  NAND2_X1 maj_200_U12 ( .A1(u_1_1[2]), .A2(maj_200_n24), .ZN(maj_200_n20) );
  NAND2_X1 maj_200_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_200_n21) );
  NAND2_X1 maj_200_U10 ( .A1(maj_200_n21), .A2(maj_200_n20), .ZN(maj_200_n23)
         );
  XOR2_X1 maj_200_U9 ( .A(u_1_1[2]), .B(maj_200_n24), .Z(maj_200_n26) );
  XOR2_X1 maj_200_U8 ( .A(u_1_1[5]), .B(maj_200_n25), .Z(maj_200_n27) );
  XOR2_X1 maj_200_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_200_n24) );
  XOR2_X1 maj_200_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_200_n25) );
  OR2_X1 maj_200_U5 ( .A1(maj_200_n23), .A2(maj_200_n22), .ZN(maj_200_n32) );
  NAND2_X1 maj_200_U4 ( .A1(maj_200_n22), .A2(maj_200_n23), .ZN(maj_200_n34)
         );
  NAND2_X1 maj_200_U3 ( .A1(maj_200_n32), .A2(maj_200_n31), .ZN(maj_200_n33)
         );
  NAND2_X1 maj_200_U2 ( .A1(maj_200_n34), .A2(maj_200_n33), .ZN(maj_200_port_o) );
  OR2_X1 maj_201_U19 ( .A1(maj_201_n27), .A2(maj_201_n26), .ZN(maj_201_n28) );
  NAND2_X1 maj_201_U18 ( .A1(v_1_1[6]), .A2(maj_201_n28), .ZN(maj_201_n29) );
  NAND2_X1 maj_201_U17 ( .A1(maj_201_n26), .A2(maj_201_n27), .ZN(maj_201_n30)
         );
  NAND2_X1 maj_201_U16 ( .A1(maj_201_n30), .A2(maj_201_n29), .ZN(maj_201_n31)
         );
  NAND2_X1 maj_201_U15 ( .A1(v_1_1[5]), .A2(maj_201_n25), .ZN(maj_201_n18) );
  NAND2_X1 maj_201_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_201_n19) );
  NAND2_X1 maj_201_U13 ( .A1(maj_201_n19), .A2(maj_201_n18), .ZN(maj_201_n22)
         );
  NAND2_X1 maj_201_U12 ( .A1(v_1_1[2]), .A2(maj_201_n24), .ZN(maj_201_n20) );
  NAND2_X1 maj_201_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_201_n21) );
  NAND2_X1 maj_201_U10 ( .A1(maj_201_n21), .A2(maj_201_n20), .ZN(maj_201_n23)
         );
  XOR2_X1 maj_201_U9 ( .A(v_1_1[2]), .B(maj_201_n24), .Z(maj_201_n26) );
  XOR2_X1 maj_201_U8 ( .A(v_1_1[5]), .B(maj_201_n25), .Z(maj_201_n27) );
  XOR2_X1 maj_201_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_201_n24) );
  XOR2_X1 maj_201_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_201_n25) );
  OR2_X1 maj_201_U5 ( .A1(maj_201_n23), .A2(maj_201_n22), .ZN(maj_201_n32) );
  NAND2_X1 maj_201_U4 ( .A1(maj_201_n22), .A2(maj_201_n23), .ZN(maj_201_n34)
         );
  NAND2_X1 maj_201_U3 ( .A1(maj_201_n32), .A2(maj_201_n31), .ZN(maj_201_n33)
         );
  NAND2_X1 maj_201_U2 ( .A1(maj_201_n34), .A2(maj_201_n33), .ZN(maj_201_port_o) );
  OR2_X1 maj_202_U19 ( .A1(maj_202_n27), .A2(maj_202_n26), .ZN(maj_202_n28) );
  NAND2_X1 maj_202_U18 ( .A1(u_1_2[6]), .A2(maj_202_n28), .ZN(maj_202_n29) );
  NAND2_X1 maj_202_U17 ( .A1(maj_202_n26), .A2(maj_202_n27), .ZN(maj_202_n30)
         );
  NAND2_X1 maj_202_U16 ( .A1(maj_202_n30), .A2(maj_202_n29), .ZN(maj_202_n31)
         );
  NAND2_X1 maj_202_U15 ( .A1(u_1_2[5]), .A2(maj_202_n25), .ZN(maj_202_n18) );
  NAND2_X1 maj_202_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_202_n19) );
  NAND2_X1 maj_202_U13 ( .A1(maj_202_n19), .A2(maj_202_n18), .ZN(maj_202_n22)
         );
  NAND2_X1 maj_202_U12 ( .A1(u_1_2[2]), .A2(maj_202_n24), .ZN(maj_202_n20) );
  NAND2_X1 maj_202_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_202_n21) );
  NAND2_X1 maj_202_U10 ( .A1(maj_202_n21), .A2(maj_202_n20), .ZN(maj_202_n23)
         );
  XOR2_X1 maj_202_U9 ( .A(u_1_2[2]), .B(maj_202_n24), .Z(maj_202_n26) );
  XOR2_X1 maj_202_U8 ( .A(u_1_2[5]), .B(maj_202_n25), .Z(maj_202_n27) );
  XOR2_X1 maj_202_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_202_n24) );
  XOR2_X1 maj_202_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_202_n25) );
  OR2_X1 maj_202_U5 ( .A1(maj_202_n23), .A2(maj_202_n22), .ZN(maj_202_n32) );
  NAND2_X1 maj_202_U4 ( .A1(maj_202_n22), .A2(maj_202_n23), .ZN(maj_202_n34)
         );
  NAND2_X1 maj_202_U3 ( .A1(maj_202_n32), .A2(maj_202_n31), .ZN(maj_202_n33)
         );
  NAND2_X1 maj_202_U2 ( .A1(maj_202_n34), .A2(maj_202_n33), .ZN(maj_202_port_o) );
  OR2_X1 maj_203_U19 ( .A1(maj_203_n27), .A2(maj_203_n26), .ZN(maj_203_n28) );
  NAND2_X1 maj_203_U18 ( .A1(v_1_2[6]), .A2(maj_203_n28), .ZN(maj_203_n29) );
  NAND2_X1 maj_203_U17 ( .A1(maj_203_n26), .A2(maj_203_n27), .ZN(maj_203_n30)
         );
  NAND2_X1 maj_203_U16 ( .A1(maj_203_n30), .A2(maj_203_n29), .ZN(maj_203_n31)
         );
  NAND2_X1 maj_203_U15 ( .A1(v_1_2[5]), .A2(maj_203_n25), .ZN(maj_203_n18) );
  NAND2_X1 maj_203_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_203_n19) );
  NAND2_X1 maj_203_U13 ( .A1(maj_203_n19), .A2(maj_203_n18), .ZN(maj_203_n22)
         );
  NAND2_X1 maj_203_U12 ( .A1(v_1_2[2]), .A2(maj_203_n24), .ZN(maj_203_n20) );
  NAND2_X1 maj_203_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_203_n21) );
  NAND2_X1 maj_203_U10 ( .A1(maj_203_n21), .A2(maj_203_n20), .ZN(maj_203_n23)
         );
  XOR2_X1 maj_203_U9 ( .A(v_1_2[2]), .B(maj_203_n24), .Z(maj_203_n26) );
  XOR2_X1 maj_203_U8 ( .A(v_1_2[5]), .B(maj_203_n25), .Z(maj_203_n27) );
  XOR2_X1 maj_203_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_203_n24) );
  XOR2_X1 maj_203_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_203_n25) );
  OR2_X1 maj_203_U5 ( .A1(maj_203_n23), .A2(maj_203_n22), .ZN(maj_203_n32) );
  NAND2_X1 maj_203_U4 ( .A1(maj_203_n22), .A2(maj_203_n23), .ZN(maj_203_n34)
         );
  NAND2_X1 maj_203_U3 ( .A1(maj_203_n32), .A2(maj_203_n31), .ZN(maj_203_n33)
         );
  NAND2_X1 maj_203_U2 ( .A1(maj_203_n34), .A2(maj_203_n33), .ZN(maj_203_port_o) );
  OR2_X1 maj_204_U19 ( .A1(maj_204_n27), .A2(maj_204_n26), .ZN(maj_204_n28) );
  NAND2_X1 maj_204_U18 ( .A1(u_2_0[6]), .A2(maj_204_n28), .ZN(maj_204_n29) );
  NAND2_X1 maj_204_U17 ( .A1(maj_204_n26), .A2(maj_204_n27), .ZN(maj_204_n30)
         );
  NAND2_X1 maj_204_U16 ( .A1(maj_204_n30), .A2(maj_204_n29), .ZN(maj_204_n31)
         );
  NAND2_X1 maj_204_U15 ( .A1(u_2_0[5]), .A2(maj_204_n25), .ZN(maj_204_n18) );
  NAND2_X1 maj_204_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_204_n19) );
  NAND2_X1 maj_204_U13 ( .A1(maj_204_n19), .A2(maj_204_n18), .ZN(maj_204_n22)
         );
  NAND2_X1 maj_204_U12 ( .A1(u_2_0[2]), .A2(maj_204_n24), .ZN(maj_204_n20) );
  NAND2_X1 maj_204_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_204_n21) );
  NAND2_X1 maj_204_U10 ( .A1(maj_204_n21), .A2(maj_204_n20), .ZN(maj_204_n23)
         );
  XOR2_X1 maj_204_U9 ( .A(u_2_0[2]), .B(maj_204_n24), .Z(maj_204_n26) );
  XOR2_X1 maj_204_U8 ( .A(u_2_0[5]), .B(maj_204_n25), .Z(maj_204_n27) );
  XOR2_X1 maj_204_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_204_n24) );
  XOR2_X1 maj_204_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_204_n25) );
  OR2_X1 maj_204_U5 ( .A1(maj_204_n23), .A2(maj_204_n22), .ZN(maj_204_n32) );
  NAND2_X1 maj_204_U4 ( .A1(maj_204_n22), .A2(maj_204_n23), .ZN(maj_204_n34)
         );
  NAND2_X1 maj_204_U3 ( .A1(maj_204_n32), .A2(maj_204_n31), .ZN(maj_204_n33)
         );
  NAND2_X1 maj_204_U2 ( .A1(maj_204_n34), .A2(maj_204_n33), .ZN(maj_204_port_o) );
  OR2_X1 maj_205_U19 ( .A1(maj_205_n27), .A2(maj_205_n26), .ZN(maj_205_n28) );
  NAND2_X1 maj_205_U18 ( .A1(v_2_0[6]), .A2(maj_205_n28), .ZN(maj_205_n29) );
  NAND2_X1 maj_205_U17 ( .A1(maj_205_n26), .A2(maj_205_n27), .ZN(maj_205_n30)
         );
  NAND2_X1 maj_205_U16 ( .A1(maj_205_n30), .A2(maj_205_n29), .ZN(maj_205_n31)
         );
  NAND2_X1 maj_205_U15 ( .A1(v_2_0[5]), .A2(maj_205_n25), .ZN(maj_205_n18) );
  NAND2_X1 maj_205_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_205_n19) );
  NAND2_X1 maj_205_U13 ( .A1(maj_205_n19), .A2(maj_205_n18), .ZN(maj_205_n22)
         );
  NAND2_X1 maj_205_U12 ( .A1(v_2_0[2]), .A2(maj_205_n24), .ZN(maj_205_n20) );
  NAND2_X1 maj_205_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_205_n21) );
  NAND2_X1 maj_205_U10 ( .A1(maj_205_n21), .A2(maj_205_n20), .ZN(maj_205_n23)
         );
  XOR2_X1 maj_205_U9 ( .A(v_2_0[2]), .B(maj_205_n24), .Z(maj_205_n26) );
  XOR2_X1 maj_205_U8 ( .A(v_2_0[5]), .B(maj_205_n25), .Z(maj_205_n27) );
  XOR2_X1 maj_205_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_205_n24) );
  XOR2_X1 maj_205_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_205_n25) );
  OR2_X1 maj_205_U5 ( .A1(maj_205_n23), .A2(maj_205_n22), .ZN(maj_205_n32) );
  NAND2_X1 maj_205_U4 ( .A1(maj_205_n22), .A2(maj_205_n23), .ZN(maj_205_n34)
         );
  NAND2_X1 maj_205_U3 ( .A1(maj_205_n32), .A2(maj_205_n31), .ZN(maj_205_n33)
         );
  NAND2_X1 maj_205_U2 ( .A1(maj_205_n34), .A2(maj_205_n33), .ZN(maj_205_port_o) );
  OR2_X1 maj_206_U19 ( .A1(maj_206_n27), .A2(maj_206_n26), .ZN(maj_206_n28) );
  NAND2_X1 maj_206_U18 ( .A1(u_2_1[6]), .A2(maj_206_n28), .ZN(maj_206_n29) );
  NAND2_X1 maj_206_U17 ( .A1(maj_206_n26), .A2(maj_206_n27), .ZN(maj_206_n30)
         );
  NAND2_X1 maj_206_U16 ( .A1(maj_206_n30), .A2(maj_206_n29), .ZN(maj_206_n31)
         );
  NAND2_X1 maj_206_U15 ( .A1(u_2_1[5]), .A2(maj_206_n25), .ZN(maj_206_n18) );
  NAND2_X1 maj_206_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_206_n19) );
  NAND2_X1 maj_206_U13 ( .A1(maj_206_n19), .A2(maj_206_n18), .ZN(maj_206_n22)
         );
  NAND2_X1 maj_206_U12 ( .A1(u_2_1[2]), .A2(maj_206_n24), .ZN(maj_206_n20) );
  NAND2_X1 maj_206_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_206_n21) );
  NAND2_X1 maj_206_U10 ( .A1(maj_206_n21), .A2(maj_206_n20), .ZN(maj_206_n23)
         );
  XOR2_X1 maj_206_U9 ( .A(u_2_1[2]), .B(maj_206_n24), .Z(maj_206_n26) );
  XOR2_X1 maj_206_U8 ( .A(u_2_1[5]), .B(maj_206_n25), .Z(maj_206_n27) );
  XOR2_X1 maj_206_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_206_n24) );
  XOR2_X1 maj_206_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_206_n25) );
  OR2_X1 maj_206_U5 ( .A1(maj_206_n23), .A2(maj_206_n22), .ZN(maj_206_n32) );
  NAND2_X1 maj_206_U4 ( .A1(maj_206_n22), .A2(maj_206_n23), .ZN(maj_206_n34)
         );
  NAND2_X1 maj_206_U3 ( .A1(maj_206_n32), .A2(maj_206_n31), .ZN(maj_206_n33)
         );
  NAND2_X1 maj_206_U2 ( .A1(maj_206_n34), .A2(maj_206_n33), .ZN(maj_206_port_o) );
  OR2_X1 maj_207_U19 ( .A1(maj_207_n27), .A2(maj_207_n26), .ZN(maj_207_n28) );
  NAND2_X1 maj_207_U18 ( .A1(v_2_1[6]), .A2(maj_207_n28), .ZN(maj_207_n29) );
  NAND2_X1 maj_207_U17 ( .A1(maj_207_n26), .A2(maj_207_n27), .ZN(maj_207_n30)
         );
  NAND2_X1 maj_207_U16 ( .A1(maj_207_n30), .A2(maj_207_n29), .ZN(maj_207_n31)
         );
  NAND2_X1 maj_207_U15 ( .A1(v_2_1[5]), .A2(maj_207_n25), .ZN(maj_207_n18) );
  NAND2_X1 maj_207_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_207_n19) );
  NAND2_X1 maj_207_U13 ( .A1(maj_207_n19), .A2(maj_207_n18), .ZN(maj_207_n22)
         );
  NAND2_X1 maj_207_U12 ( .A1(v_2_1[2]), .A2(maj_207_n24), .ZN(maj_207_n20) );
  NAND2_X1 maj_207_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_207_n21) );
  NAND2_X1 maj_207_U10 ( .A1(maj_207_n21), .A2(maj_207_n20), .ZN(maj_207_n23)
         );
  XOR2_X1 maj_207_U9 ( .A(v_2_1[2]), .B(maj_207_n24), .Z(maj_207_n26) );
  XOR2_X1 maj_207_U8 ( .A(v_2_1[5]), .B(maj_207_n25), .Z(maj_207_n27) );
  XOR2_X1 maj_207_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_207_n24) );
  XOR2_X1 maj_207_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_207_n25) );
  OR2_X1 maj_207_U5 ( .A1(maj_207_n23), .A2(maj_207_n22), .ZN(maj_207_n32) );
  NAND2_X1 maj_207_U4 ( .A1(maj_207_n22), .A2(maj_207_n23), .ZN(maj_207_n34)
         );
  NAND2_X1 maj_207_U3 ( .A1(maj_207_n32), .A2(maj_207_n31), .ZN(maj_207_n33)
         );
  NAND2_X1 maj_207_U2 ( .A1(maj_207_n34), .A2(maj_207_n33), .ZN(maj_207_port_o) );
  OR2_X1 maj_208_U19 ( .A1(maj_208_n27), .A2(maj_208_n26), .ZN(maj_208_n28) );
  NAND2_X1 maj_208_U18 ( .A1(u_2_2[6]), .A2(maj_208_n28), .ZN(maj_208_n29) );
  NAND2_X1 maj_208_U17 ( .A1(maj_208_n26), .A2(maj_208_n27), .ZN(maj_208_n30)
         );
  NAND2_X1 maj_208_U16 ( .A1(maj_208_n30), .A2(maj_208_n29), .ZN(maj_208_n31)
         );
  NAND2_X1 maj_208_U15 ( .A1(u_2_2[5]), .A2(maj_208_n25), .ZN(maj_208_n18) );
  NAND2_X1 maj_208_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_208_n19) );
  NAND2_X1 maj_208_U13 ( .A1(maj_208_n19), .A2(maj_208_n18), .ZN(maj_208_n22)
         );
  NAND2_X1 maj_208_U12 ( .A1(u_2_2[2]), .A2(maj_208_n24), .ZN(maj_208_n20) );
  NAND2_X1 maj_208_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_208_n21) );
  NAND2_X1 maj_208_U10 ( .A1(maj_208_n21), .A2(maj_208_n20), .ZN(maj_208_n23)
         );
  XOR2_X1 maj_208_U9 ( .A(u_2_2[2]), .B(maj_208_n24), .Z(maj_208_n26) );
  XOR2_X1 maj_208_U8 ( .A(u_2_2[5]), .B(maj_208_n25), .Z(maj_208_n27) );
  XOR2_X1 maj_208_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_208_n24) );
  XOR2_X1 maj_208_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_208_n25) );
  OR2_X1 maj_208_U5 ( .A1(maj_208_n23), .A2(maj_208_n22), .ZN(maj_208_n32) );
  NAND2_X1 maj_208_U4 ( .A1(maj_208_n22), .A2(maj_208_n23), .ZN(maj_208_n34)
         );
  NAND2_X1 maj_208_U3 ( .A1(maj_208_n32), .A2(maj_208_n31), .ZN(maj_208_n33)
         );
  NAND2_X1 maj_208_U2 ( .A1(maj_208_n34), .A2(maj_208_n33), .ZN(maj_208_port_o) );
  OR2_X1 maj_209_U19 ( .A1(maj_209_n27), .A2(maj_209_n26), .ZN(maj_209_n28) );
  NAND2_X1 maj_209_U18 ( .A1(v_2_2[6]), .A2(maj_209_n28), .ZN(maj_209_n29) );
  NAND2_X1 maj_209_U17 ( .A1(maj_209_n26), .A2(maj_209_n27), .ZN(maj_209_n30)
         );
  NAND2_X1 maj_209_U16 ( .A1(maj_209_n30), .A2(maj_209_n29), .ZN(maj_209_n31)
         );
  NAND2_X1 maj_209_U15 ( .A1(v_2_2[5]), .A2(maj_209_n25), .ZN(maj_209_n18) );
  NAND2_X1 maj_209_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_209_n19) );
  NAND2_X1 maj_209_U13 ( .A1(maj_209_n19), .A2(maj_209_n18), .ZN(maj_209_n22)
         );
  NAND2_X1 maj_209_U12 ( .A1(v_2_2[2]), .A2(maj_209_n24), .ZN(maj_209_n20) );
  NAND2_X1 maj_209_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_209_n21) );
  NAND2_X1 maj_209_U10 ( .A1(maj_209_n21), .A2(maj_209_n20), .ZN(maj_209_n23)
         );
  XOR2_X1 maj_209_U9 ( .A(v_2_2[2]), .B(maj_209_n24), .Z(maj_209_n26) );
  XOR2_X1 maj_209_U8 ( .A(v_2_2[5]), .B(maj_209_n25), .Z(maj_209_n27) );
  XOR2_X1 maj_209_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_209_n24) );
  XOR2_X1 maj_209_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_209_n25) );
  OR2_X1 maj_209_U5 ( .A1(maj_209_n23), .A2(maj_209_n22), .ZN(maj_209_n32) );
  NAND2_X1 maj_209_U4 ( .A1(maj_209_n22), .A2(maj_209_n23), .ZN(maj_209_n34)
         );
  NAND2_X1 maj_209_U3 ( .A1(maj_209_n32), .A2(maj_209_n31), .ZN(maj_209_n33)
         );
  NAND2_X1 maj_209_U2 ( .A1(maj_209_n34), .A2(maj_209_n33), .ZN(maj_209_port_o) );
  OR2_X1 maj_210_U19 ( .A1(maj_210_n27), .A2(maj_210_n26), .ZN(maj_210_n28) );
  NAND2_X1 maj_210_U18 ( .A1(u_3_0[6]), .A2(maj_210_n28), .ZN(maj_210_n29) );
  NAND2_X1 maj_210_U17 ( .A1(maj_210_n26), .A2(maj_210_n27), .ZN(maj_210_n30)
         );
  NAND2_X1 maj_210_U16 ( .A1(maj_210_n30), .A2(maj_210_n29), .ZN(maj_210_n31)
         );
  NAND2_X1 maj_210_U15 ( .A1(u_3_0[5]), .A2(maj_210_n25), .ZN(maj_210_n18) );
  NAND2_X1 maj_210_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_210_n19) );
  NAND2_X1 maj_210_U13 ( .A1(maj_210_n19), .A2(maj_210_n18), .ZN(maj_210_n22)
         );
  NAND2_X1 maj_210_U12 ( .A1(u_3_0[2]), .A2(maj_210_n24), .ZN(maj_210_n20) );
  NAND2_X1 maj_210_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_210_n21) );
  NAND2_X1 maj_210_U10 ( .A1(maj_210_n21), .A2(maj_210_n20), .ZN(maj_210_n23)
         );
  XOR2_X1 maj_210_U9 ( .A(u_3_0[2]), .B(maj_210_n24), .Z(maj_210_n26) );
  XOR2_X1 maj_210_U8 ( .A(u_3_0[5]), .B(maj_210_n25), .Z(maj_210_n27) );
  XOR2_X1 maj_210_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_210_n24) );
  XOR2_X1 maj_210_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_210_n25) );
  OR2_X1 maj_210_U5 ( .A1(maj_210_n23), .A2(maj_210_n22), .ZN(maj_210_n32) );
  NAND2_X1 maj_210_U4 ( .A1(maj_210_n22), .A2(maj_210_n23), .ZN(maj_210_n34)
         );
  NAND2_X1 maj_210_U3 ( .A1(maj_210_n32), .A2(maj_210_n31), .ZN(maj_210_n33)
         );
  NAND2_X1 maj_210_U2 ( .A1(maj_210_n34), .A2(maj_210_n33), .ZN(maj_210_port_o) );
  OR2_X1 maj_211_U19 ( .A1(maj_211_n27), .A2(maj_211_n26), .ZN(maj_211_n28) );
  NAND2_X1 maj_211_U18 ( .A1(v_3_0[6]), .A2(maj_211_n28), .ZN(maj_211_n29) );
  NAND2_X1 maj_211_U17 ( .A1(maj_211_n26), .A2(maj_211_n27), .ZN(maj_211_n30)
         );
  NAND2_X1 maj_211_U16 ( .A1(maj_211_n30), .A2(maj_211_n29), .ZN(maj_211_n31)
         );
  NAND2_X1 maj_211_U15 ( .A1(v_3_0[5]), .A2(maj_211_n25), .ZN(maj_211_n18) );
  NAND2_X1 maj_211_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_211_n19) );
  NAND2_X1 maj_211_U13 ( .A1(maj_211_n19), .A2(maj_211_n18), .ZN(maj_211_n22)
         );
  NAND2_X1 maj_211_U12 ( .A1(v_3_0[2]), .A2(maj_211_n24), .ZN(maj_211_n20) );
  NAND2_X1 maj_211_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_211_n21) );
  NAND2_X1 maj_211_U10 ( .A1(maj_211_n21), .A2(maj_211_n20), .ZN(maj_211_n23)
         );
  XOR2_X1 maj_211_U9 ( .A(v_3_0[2]), .B(maj_211_n24), .Z(maj_211_n26) );
  XOR2_X1 maj_211_U8 ( .A(v_3_0[5]), .B(maj_211_n25), .Z(maj_211_n27) );
  XOR2_X1 maj_211_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_211_n24) );
  XOR2_X1 maj_211_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_211_n25) );
  OR2_X1 maj_211_U5 ( .A1(maj_211_n23), .A2(maj_211_n22), .ZN(maj_211_n32) );
  NAND2_X1 maj_211_U4 ( .A1(maj_211_n22), .A2(maj_211_n23), .ZN(maj_211_n34)
         );
  NAND2_X1 maj_211_U3 ( .A1(maj_211_n32), .A2(maj_211_n31), .ZN(maj_211_n33)
         );
  NAND2_X1 maj_211_U2 ( .A1(maj_211_n34), .A2(maj_211_n33), .ZN(maj_211_port_o) );
  OR2_X1 maj_212_U19 ( .A1(maj_212_n27), .A2(maj_212_n26), .ZN(maj_212_n28) );
  NAND2_X1 maj_212_U18 ( .A1(u_3_1[6]), .A2(maj_212_n28), .ZN(maj_212_n29) );
  NAND2_X1 maj_212_U17 ( .A1(maj_212_n26), .A2(maj_212_n27), .ZN(maj_212_n30)
         );
  NAND2_X1 maj_212_U16 ( .A1(maj_212_n30), .A2(maj_212_n29), .ZN(maj_212_n31)
         );
  NAND2_X1 maj_212_U15 ( .A1(u_3_1[5]), .A2(maj_212_n25), .ZN(maj_212_n18) );
  NAND2_X1 maj_212_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_212_n19) );
  NAND2_X1 maj_212_U13 ( .A1(maj_212_n19), .A2(maj_212_n18), .ZN(maj_212_n22)
         );
  NAND2_X1 maj_212_U12 ( .A1(u_3_1[2]), .A2(maj_212_n24), .ZN(maj_212_n20) );
  NAND2_X1 maj_212_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_212_n21) );
  NAND2_X1 maj_212_U10 ( .A1(maj_212_n21), .A2(maj_212_n20), .ZN(maj_212_n23)
         );
  XOR2_X1 maj_212_U9 ( .A(u_3_1[2]), .B(maj_212_n24), .Z(maj_212_n26) );
  XOR2_X1 maj_212_U8 ( .A(u_3_1[5]), .B(maj_212_n25), .Z(maj_212_n27) );
  XOR2_X1 maj_212_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_212_n24) );
  XOR2_X1 maj_212_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_212_n25) );
  OR2_X1 maj_212_U5 ( .A1(maj_212_n23), .A2(maj_212_n22), .ZN(maj_212_n32) );
  NAND2_X1 maj_212_U4 ( .A1(maj_212_n22), .A2(maj_212_n23), .ZN(maj_212_n34)
         );
  NAND2_X1 maj_212_U3 ( .A1(maj_212_n32), .A2(maj_212_n31), .ZN(maj_212_n33)
         );
  NAND2_X1 maj_212_U2 ( .A1(maj_212_n34), .A2(maj_212_n33), .ZN(maj_212_port_o) );
  OR2_X1 maj_213_U19 ( .A1(maj_213_n27), .A2(maj_213_n26), .ZN(maj_213_n28) );
  NAND2_X1 maj_213_U18 ( .A1(v_3_1[6]), .A2(maj_213_n28), .ZN(maj_213_n29) );
  NAND2_X1 maj_213_U17 ( .A1(maj_213_n26), .A2(maj_213_n27), .ZN(maj_213_n30)
         );
  NAND2_X1 maj_213_U16 ( .A1(maj_213_n30), .A2(maj_213_n29), .ZN(maj_213_n31)
         );
  NAND2_X1 maj_213_U15 ( .A1(v_3_1[5]), .A2(maj_213_n25), .ZN(maj_213_n18) );
  NAND2_X1 maj_213_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_213_n19) );
  NAND2_X1 maj_213_U13 ( .A1(maj_213_n19), .A2(maj_213_n18), .ZN(maj_213_n22)
         );
  NAND2_X1 maj_213_U12 ( .A1(v_3_1[2]), .A2(maj_213_n24), .ZN(maj_213_n20) );
  NAND2_X1 maj_213_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_213_n21) );
  NAND2_X1 maj_213_U10 ( .A1(maj_213_n21), .A2(maj_213_n20), .ZN(maj_213_n23)
         );
  XOR2_X1 maj_213_U9 ( .A(v_3_1[2]), .B(maj_213_n24), .Z(maj_213_n26) );
  XOR2_X1 maj_213_U8 ( .A(v_3_1[5]), .B(maj_213_n25), .Z(maj_213_n27) );
  XOR2_X1 maj_213_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_213_n24) );
  XOR2_X1 maj_213_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_213_n25) );
  OR2_X1 maj_213_U5 ( .A1(maj_213_n23), .A2(maj_213_n22), .ZN(maj_213_n32) );
  NAND2_X1 maj_213_U4 ( .A1(maj_213_n22), .A2(maj_213_n23), .ZN(maj_213_n34)
         );
  NAND2_X1 maj_213_U3 ( .A1(maj_213_n32), .A2(maj_213_n31), .ZN(maj_213_n33)
         );
  NAND2_X1 maj_213_U2 ( .A1(maj_213_n34), .A2(maj_213_n33), .ZN(maj_213_port_o) );
  OR2_X1 maj_214_U19 ( .A1(maj_214_n27), .A2(maj_214_n26), .ZN(maj_214_n28) );
  NAND2_X1 maj_214_U18 ( .A1(u_3_2[6]), .A2(maj_214_n28), .ZN(maj_214_n29) );
  NAND2_X1 maj_214_U17 ( .A1(maj_214_n26), .A2(maj_214_n27), .ZN(maj_214_n30)
         );
  NAND2_X1 maj_214_U16 ( .A1(maj_214_n30), .A2(maj_214_n29), .ZN(maj_214_n31)
         );
  NAND2_X1 maj_214_U15 ( .A1(u_3_2[5]), .A2(maj_214_n25), .ZN(maj_214_n18) );
  NAND2_X1 maj_214_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_214_n19) );
  NAND2_X1 maj_214_U13 ( .A1(maj_214_n19), .A2(maj_214_n18), .ZN(maj_214_n22)
         );
  NAND2_X1 maj_214_U12 ( .A1(u_3_2[2]), .A2(maj_214_n24), .ZN(maj_214_n20) );
  NAND2_X1 maj_214_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_214_n21) );
  NAND2_X1 maj_214_U10 ( .A1(maj_214_n21), .A2(maj_214_n20), .ZN(maj_214_n23)
         );
  XOR2_X1 maj_214_U9 ( .A(u_3_2[2]), .B(maj_214_n24), .Z(maj_214_n26) );
  XOR2_X1 maj_214_U8 ( .A(u_3_2[5]), .B(maj_214_n25), .Z(maj_214_n27) );
  XOR2_X1 maj_214_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_214_n24) );
  XOR2_X1 maj_214_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_214_n25) );
  OR2_X1 maj_214_U5 ( .A1(maj_214_n23), .A2(maj_214_n22), .ZN(maj_214_n32) );
  NAND2_X1 maj_214_U4 ( .A1(maj_214_n22), .A2(maj_214_n23), .ZN(maj_214_n34)
         );
  NAND2_X1 maj_214_U3 ( .A1(maj_214_n32), .A2(maj_214_n31), .ZN(maj_214_n33)
         );
  NAND2_X1 maj_214_U2 ( .A1(maj_214_n34), .A2(maj_214_n33), .ZN(maj_214_port_o) );
  OR2_X1 maj_215_U19 ( .A1(maj_215_n27), .A2(maj_215_n26), .ZN(maj_215_n28) );
  NAND2_X1 maj_215_U18 ( .A1(v_3_2[6]), .A2(maj_215_n28), .ZN(maj_215_n29) );
  NAND2_X1 maj_215_U17 ( .A1(maj_215_n26), .A2(maj_215_n27), .ZN(maj_215_n30)
         );
  NAND2_X1 maj_215_U16 ( .A1(maj_215_n30), .A2(maj_215_n29), .ZN(maj_215_n31)
         );
  NAND2_X1 maj_215_U15 ( .A1(v_3_2[5]), .A2(maj_215_n25), .ZN(maj_215_n18) );
  NAND2_X1 maj_215_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_215_n19) );
  NAND2_X1 maj_215_U13 ( .A1(maj_215_n19), .A2(maj_215_n18), .ZN(maj_215_n22)
         );
  NAND2_X1 maj_215_U12 ( .A1(v_3_2[2]), .A2(maj_215_n24), .ZN(maj_215_n20) );
  NAND2_X1 maj_215_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_215_n21) );
  NAND2_X1 maj_215_U10 ( .A1(maj_215_n21), .A2(maj_215_n20), .ZN(maj_215_n23)
         );
  XOR2_X1 maj_215_U9 ( .A(v_3_2[2]), .B(maj_215_n24), .Z(maj_215_n26) );
  XOR2_X1 maj_215_U8 ( .A(v_3_2[5]), .B(maj_215_n25), .Z(maj_215_n27) );
  XOR2_X1 maj_215_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_215_n24) );
  XOR2_X1 maj_215_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_215_n25) );
  OR2_X1 maj_215_U5 ( .A1(maj_215_n23), .A2(maj_215_n22), .ZN(maj_215_n32) );
  NAND2_X1 maj_215_U4 ( .A1(maj_215_n22), .A2(maj_215_n23), .ZN(maj_215_n34)
         );
  NAND2_X1 maj_215_U3 ( .A1(maj_215_n32), .A2(maj_215_n31), .ZN(maj_215_n33)
         );
  NAND2_X1 maj_215_U2 ( .A1(maj_215_n34), .A2(maj_215_n33), .ZN(maj_215_port_o) );
  OR2_X1 maj_216_U19 ( .A1(maj_216_n27), .A2(maj_216_n26), .ZN(maj_216_n28) );
  NAND2_X1 maj_216_U18 ( .A1(u_0_0[6]), .A2(maj_216_n28), .ZN(maj_216_n29) );
  NAND2_X1 maj_216_U17 ( .A1(maj_216_n26), .A2(maj_216_n27), .ZN(maj_216_n30)
         );
  NAND2_X1 maj_216_U16 ( .A1(maj_216_n30), .A2(maj_216_n29), .ZN(maj_216_n31)
         );
  NAND2_X1 maj_216_U15 ( .A1(u_0_0[5]), .A2(maj_216_n25), .ZN(maj_216_n18) );
  NAND2_X1 maj_216_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_216_n19) );
  NAND2_X1 maj_216_U13 ( .A1(maj_216_n19), .A2(maj_216_n18), .ZN(maj_216_n22)
         );
  NAND2_X1 maj_216_U12 ( .A1(u_0_0[2]), .A2(maj_216_n24), .ZN(maj_216_n20) );
  NAND2_X1 maj_216_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_216_n21) );
  NAND2_X1 maj_216_U10 ( .A1(maj_216_n21), .A2(maj_216_n20), .ZN(maj_216_n23)
         );
  XOR2_X1 maj_216_U9 ( .A(u_0_0[2]), .B(maj_216_n24), .Z(maj_216_n26) );
  XOR2_X1 maj_216_U8 ( .A(u_0_0[5]), .B(maj_216_n25), .Z(maj_216_n27) );
  XOR2_X1 maj_216_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_216_n24) );
  XOR2_X1 maj_216_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_216_n25) );
  OR2_X1 maj_216_U5 ( .A1(maj_216_n23), .A2(maj_216_n22), .ZN(maj_216_n32) );
  NAND2_X1 maj_216_U4 ( .A1(maj_216_n22), .A2(maj_216_n23), .ZN(maj_216_n34)
         );
  NAND2_X1 maj_216_U3 ( .A1(maj_216_n32), .A2(maj_216_n31), .ZN(maj_216_n33)
         );
  NAND2_X1 maj_216_U2 ( .A1(maj_216_n34), .A2(maj_216_n33), .ZN(maj_216_port_o) );
  OR2_X1 maj_217_U19 ( .A1(maj_217_n27), .A2(maj_217_n26), .ZN(maj_217_n28) );
  NAND2_X1 maj_217_U18 ( .A1(v_0_0[6]), .A2(maj_217_n28), .ZN(maj_217_n29) );
  NAND2_X1 maj_217_U17 ( .A1(maj_217_n26), .A2(maj_217_n27), .ZN(maj_217_n30)
         );
  NAND2_X1 maj_217_U16 ( .A1(maj_217_n30), .A2(maj_217_n29), .ZN(maj_217_n31)
         );
  NAND2_X1 maj_217_U15 ( .A1(v_0_0[5]), .A2(maj_217_n25), .ZN(maj_217_n18) );
  NAND2_X1 maj_217_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_217_n19) );
  NAND2_X1 maj_217_U13 ( .A1(maj_217_n19), .A2(maj_217_n18), .ZN(maj_217_n22)
         );
  NAND2_X1 maj_217_U12 ( .A1(v_0_0[2]), .A2(maj_217_n24), .ZN(maj_217_n20) );
  NAND2_X1 maj_217_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_217_n21) );
  NAND2_X1 maj_217_U10 ( .A1(maj_217_n21), .A2(maj_217_n20), .ZN(maj_217_n23)
         );
  XOR2_X1 maj_217_U9 ( .A(v_0_0[2]), .B(maj_217_n24), .Z(maj_217_n26) );
  XOR2_X1 maj_217_U8 ( .A(v_0_0[5]), .B(maj_217_n25), .Z(maj_217_n27) );
  XOR2_X1 maj_217_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_217_n24) );
  XOR2_X1 maj_217_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_217_n25) );
  OR2_X1 maj_217_U5 ( .A1(maj_217_n23), .A2(maj_217_n22), .ZN(maj_217_n32) );
  NAND2_X1 maj_217_U4 ( .A1(maj_217_n22), .A2(maj_217_n23), .ZN(maj_217_n34)
         );
  NAND2_X1 maj_217_U3 ( .A1(maj_217_n32), .A2(maj_217_n31), .ZN(maj_217_n33)
         );
  NAND2_X1 maj_217_U2 ( .A1(maj_217_n34), .A2(maj_217_n33), .ZN(maj_217_port_o) );
  OR2_X1 maj_218_U19 ( .A1(maj_218_n27), .A2(maj_218_n26), .ZN(maj_218_n28) );
  NAND2_X1 maj_218_U18 ( .A1(u_0_1[6]), .A2(maj_218_n28), .ZN(maj_218_n29) );
  NAND2_X1 maj_218_U17 ( .A1(maj_218_n26), .A2(maj_218_n27), .ZN(maj_218_n30)
         );
  NAND2_X1 maj_218_U16 ( .A1(maj_218_n30), .A2(maj_218_n29), .ZN(maj_218_n31)
         );
  NAND2_X1 maj_218_U15 ( .A1(u_0_1[5]), .A2(maj_218_n25), .ZN(maj_218_n18) );
  NAND2_X1 maj_218_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_218_n19) );
  NAND2_X1 maj_218_U13 ( .A1(maj_218_n19), .A2(maj_218_n18), .ZN(maj_218_n22)
         );
  NAND2_X1 maj_218_U12 ( .A1(u_0_1[2]), .A2(maj_218_n24), .ZN(maj_218_n20) );
  NAND2_X1 maj_218_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_218_n21) );
  NAND2_X1 maj_218_U10 ( .A1(maj_218_n21), .A2(maj_218_n20), .ZN(maj_218_n23)
         );
  XOR2_X1 maj_218_U9 ( .A(u_0_1[2]), .B(maj_218_n24), .Z(maj_218_n26) );
  XOR2_X1 maj_218_U8 ( .A(u_0_1[5]), .B(maj_218_n25), .Z(maj_218_n27) );
  XOR2_X1 maj_218_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_218_n24) );
  XOR2_X1 maj_218_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_218_n25) );
  OR2_X1 maj_218_U5 ( .A1(maj_218_n23), .A2(maj_218_n22), .ZN(maj_218_n32) );
  NAND2_X1 maj_218_U4 ( .A1(maj_218_n22), .A2(maj_218_n23), .ZN(maj_218_n34)
         );
  NAND2_X1 maj_218_U3 ( .A1(maj_218_n32), .A2(maj_218_n31), .ZN(maj_218_n33)
         );
  NAND2_X1 maj_218_U2 ( .A1(maj_218_n34), .A2(maj_218_n33), .ZN(maj_218_port_o) );
  OR2_X1 maj_219_U19 ( .A1(maj_219_n27), .A2(maj_219_n26), .ZN(maj_219_n28) );
  NAND2_X1 maj_219_U18 ( .A1(v_0_1[6]), .A2(maj_219_n28), .ZN(maj_219_n29) );
  NAND2_X1 maj_219_U17 ( .A1(maj_219_n26), .A2(maj_219_n27), .ZN(maj_219_n30)
         );
  NAND2_X1 maj_219_U16 ( .A1(maj_219_n30), .A2(maj_219_n29), .ZN(maj_219_n31)
         );
  NAND2_X1 maj_219_U15 ( .A1(v_0_1[5]), .A2(maj_219_n25), .ZN(maj_219_n18) );
  NAND2_X1 maj_219_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_219_n19) );
  NAND2_X1 maj_219_U13 ( .A1(maj_219_n19), .A2(maj_219_n18), .ZN(maj_219_n22)
         );
  NAND2_X1 maj_219_U12 ( .A1(v_0_1[2]), .A2(maj_219_n24), .ZN(maj_219_n20) );
  NAND2_X1 maj_219_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_219_n21) );
  NAND2_X1 maj_219_U10 ( .A1(maj_219_n21), .A2(maj_219_n20), .ZN(maj_219_n23)
         );
  XOR2_X1 maj_219_U9 ( .A(v_0_1[2]), .B(maj_219_n24), .Z(maj_219_n26) );
  XOR2_X1 maj_219_U8 ( .A(v_0_1[5]), .B(maj_219_n25), .Z(maj_219_n27) );
  XOR2_X1 maj_219_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_219_n24) );
  XOR2_X1 maj_219_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_219_n25) );
  OR2_X1 maj_219_U5 ( .A1(maj_219_n23), .A2(maj_219_n22), .ZN(maj_219_n32) );
  NAND2_X1 maj_219_U4 ( .A1(maj_219_n22), .A2(maj_219_n23), .ZN(maj_219_n34)
         );
  NAND2_X1 maj_219_U3 ( .A1(maj_219_n32), .A2(maj_219_n31), .ZN(maj_219_n33)
         );
  NAND2_X1 maj_219_U2 ( .A1(maj_219_n34), .A2(maj_219_n33), .ZN(maj_219_port_o) );
  OR2_X1 maj_220_U19 ( .A1(maj_220_n27), .A2(maj_220_n26), .ZN(maj_220_n28) );
  NAND2_X1 maj_220_U18 ( .A1(u_0_2[6]), .A2(maj_220_n28), .ZN(maj_220_n29) );
  NAND2_X1 maj_220_U17 ( .A1(maj_220_n26), .A2(maj_220_n27), .ZN(maj_220_n30)
         );
  NAND2_X1 maj_220_U16 ( .A1(maj_220_n30), .A2(maj_220_n29), .ZN(maj_220_n31)
         );
  NAND2_X1 maj_220_U15 ( .A1(u_0_2[5]), .A2(maj_220_n25), .ZN(maj_220_n18) );
  NAND2_X1 maj_220_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_220_n19) );
  NAND2_X1 maj_220_U13 ( .A1(maj_220_n19), .A2(maj_220_n18), .ZN(maj_220_n22)
         );
  NAND2_X1 maj_220_U12 ( .A1(u_0_2[2]), .A2(maj_220_n24), .ZN(maj_220_n20) );
  NAND2_X1 maj_220_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_220_n21) );
  NAND2_X1 maj_220_U10 ( .A1(maj_220_n21), .A2(maj_220_n20), .ZN(maj_220_n23)
         );
  XOR2_X1 maj_220_U9 ( .A(u_0_2[2]), .B(maj_220_n24), .Z(maj_220_n26) );
  XOR2_X1 maj_220_U8 ( .A(u_0_2[5]), .B(maj_220_n25), .Z(maj_220_n27) );
  XOR2_X1 maj_220_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_220_n24) );
  XOR2_X1 maj_220_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_220_n25) );
  OR2_X1 maj_220_U5 ( .A1(maj_220_n23), .A2(maj_220_n22), .ZN(maj_220_n32) );
  NAND2_X1 maj_220_U4 ( .A1(maj_220_n22), .A2(maj_220_n23), .ZN(maj_220_n34)
         );
  NAND2_X1 maj_220_U3 ( .A1(maj_220_n32), .A2(maj_220_n31), .ZN(maj_220_n33)
         );
  NAND2_X1 maj_220_U2 ( .A1(maj_220_n34), .A2(maj_220_n33), .ZN(maj_220_port_o) );
  OR2_X1 maj_221_U19 ( .A1(maj_221_n27), .A2(maj_221_n26), .ZN(maj_221_n28) );
  NAND2_X1 maj_221_U18 ( .A1(v_0_2[6]), .A2(maj_221_n28), .ZN(maj_221_n29) );
  NAND2_X1 maj_221_U17 ( .A1(maj_221_n26), .A2(maj_221_n27), .ZN(maj_221_n30)
         );
  NAND2_X1 maj_221_U16 ( .A1(maj_221_n30), .A2(maj_221_n29), .ZN(maj_221_n31)
         );
  NAND2_X1 maj_221_U15 ( .A1(v_0_2[5]), .A2(maj_221_n25), .ZN(maj_221_n18) );
  NAND2_X1 maj_221_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_221_n19) );
  NAND2_X1 maj_221_U13 ( .A1(maj_221_n19), .A2(maj_221_n18), .ZN(maj_221_n22)
         );
  NAND2_X1 maj_221_U12 ( .A1(v_0_2[2]), .A2(maj_221_n24), .ZN(maj_221_n20) );
  NAND2_X1 maj_221_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_221_n21) );
  NAND2_X1 maj_221_U10 ( .A1(maj_221_n21), .A2(maj_221_n20), .ZN(maj_221_n23)
         );
  XOR2_X1 maj_221_U9 ( .A(v_0_2[2]), .B(maj_221_n24), .Z(maj_221_n26) );
  XOR2_X1 maj_221_U8 ( .A(v_0_2[5]), .B(maj_221_n25), .Z(maj_221_n27) );
  XOR2_X1 maj_221_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_221_n24) );
  XOR2_X1 maj_221_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_221_n25) );
  OR2_X1 maj_221_U5 ( .A1(maj_221_n23), .A2(maj_221_n22), .ZN(maj_221_n32) );
  NAND2_X1 maj_221_U4 ( .A1(maj_221_n22), .A2(maj_221_n23), .ZN(maj_221_n34)
         );
  NAND2_X1 maj_221_U3 ( .A1(maj_221_n32), .A2(maj_221_n31), .ZN(maj_221_n33)
         );
  NAND2_X1 maj_221_U2 ( .A1(maj_221_n34), .A2(maj_221_n33), .ZN(maj_221_port_o) );
  OR2_X1 maj_222_U19 ( .A1(maj_222_n27), .A2(maj_222_n26), .ZN(maj_222_n28) );
  NAND2_X1 maj_222_U18 ( .A1(u_1_0[6]), .A2(maj_222_n28), .ZN(maj_222_n29) );
  NAND2_X1 maj_222_U17 ( .A1(maj_222_n26), .A2(maj_222_n27), .ZN(maj_222_n30)
         );
  NAND2_X1 maj_222_U16 ( .A1(maj_222_n30), .A2(maj_222_n29), .ZN(maj_222_n31)
         );
  NAND2_X1 maj_222_U15 ( .A1(u_1_0[5]), .A2(maj_222_n25), .ZN(maj_222_n18) );
  NAND2_X1 maj_222_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_222_n19) );
  NAND2_X1 maj_222_U13 ( .A1(maj_222_n19), .A2(maj_222_n18), .ZN(maj_222_n22)
         );
  NAND2_X1 maj_222_U12 ( .A1(u_1_0[2]), .A2(maj_222_n24), .ZN(maj_222_n20) );
  NAND2_X1 maj_222_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_222_n21) );
  NAND2_X1 maj_222_U10 ( .A1(maj_222_n21), .A2(maj_222_n20), .ZN(maj_222_n23)
         );
  XOR2_X1 maj_222_U9 ( .A(u_1_0[2]), .B(maj_222_n24), .Z(maj_222_n26) );
  XOR2_X1 maj_222_U8 ( .A(u_1_0[5]), .B(maj_222_n25), .Z(maj_222_n27) );
  XOR2_X1 maj_222_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_222_n24) );
  XOR2_X1 maj_222_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_222_n25) );
  OR2_X1 maj_222_U5 ( .A1(maj_222_n23), .A2(maj_222_n22), .ZN(maj_222_n32) );
  NAND2_X1 maj_222_U4 ( .A1(maj_222_n22), .A2(maj_222_n23), .ZN(maj_222_n34)
         );
  NAND2_X1 maj_222_U3 ( .A1(maj_222_n32), .A2(maj_222_n31), .ZN(maj_222_n33)
         );
  NAND2_X1 maj_222_U2 ( .A1(maj_222_n34), .A2(maj_222_n33), .ZN(maj_222_port_o) );
  OR2_X1 maj_223_U19 ( .A1(maj_223_n27), .A2(maj_223_n26), .ZN(maj_223_n28) );
  NAND2_X1 maj_223_U18 ( .A1(v_1_0[6]), .A2(maj_223_n28), .ZN(maj_223_n29) );
  NAND2_X1 maj_223_U17 ( .A1(maj_223_n26), .A2(maj_223_n27), .ZN(maj_223_n30)
         );
  NAND2_X1 maj_223_U16 ( .A1(maj_223_n30), .A2(maj_223_n29), .ZN(maj_223_n31)
         );
  NAND2_X1 maj_223_U15 ( .A1(v_1_0[5]), .A2(maj_223_n25), .ZN(maj_223_n18) );
  NAND2_X1 maj_223_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_223_n19) );
  NAND2_X1 maj_223_U13 ( .A1(maj_223_n19), .A2(maj_223_n18), .ZN(maj_223_n22)
         );
  NAND2_X1 maj_223_U12 ( .A1(v_1_0[2]), .A2(maj_223_n24), .ZN(maj_223_n20) );
  NAND2_X1 maj_223_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_223_n21) );
  NAND2_X1 maj_223_U10 ( .A1(maj_223_n21), .A2(maj_223_n20), .ZN(maj_223_n23)
         );
  XOR2_X1 maj_223_U9 ( .A(v_1_0[2]), .B(maj_223_n24), .Z(maj_223_n26) );
  XOR2_X1 maj_223_U8 ( .A(v_1_0[5]), .B(maj_223_n25), .Z(maj_223_n27) );
  XOR2_X1 maj_223_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_223_n24) );
  XOR2_X1 maj_223_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_223_n25) );
  OR2_X1 maj_223_U5 ( .A1(maj_223_n23), .A2(maj_223_n22), .ZN(maj_223_n32) );
  NAND2_X1 maj_223_U4 ( .A1(maj_223_n22), .A2(maj_223_n23), .ZN(maj_223_n34)
         );
  NAND2_X1 maj_223_U3 ( .A1(maj_223_n32), .A2(maj_223_n31), .ZN(maj_223_n33)
         );
  NAND2_X1 maj_223_U2 ( .A1(maj_223_n34), .A2(maj_223_n33), .ZN(maj_223_port_o) );
  OR2_X1 maj_224_U19 ( .A1(maj_224_n27), .A2(maj_224_n26), .ZN(maj_224_n28) );
  NAND2_X1 maj_224_U18 ( .A1(u_1_1[6]), .A2(maj_224_n28), .ZN(maj_224_n29) );
  NAND2_X1 maj_224_U17 ( .A1(maj_224_n26), .A2(maj_224_n27), .ZN(maj_224_n30)
         );
  NAND2_X1 maj_224_U16 ( .A1(maj_224_n30), .A2(maj_224_n29), .ZN(maj_224_n31)
         );
  NAND2_X1 maj_224_U15 ( .A1(u_1_1[5]), .A2(maj_224_n25), .ZN(maj_224_n18) );
  NAND2_X1 maj_224_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_224_n19) );
  NAND2_X1 maj_224_U13 ( .A1(maj_224_n19), .A2(maj_224_n18), .ZN(maj_224_n22)
         );
  NAND2_X1 maj_224_U12 ( .A1(u_1_1[2]), .A2(maj_224_n24), .ZN(maj_224_n20) );
  NAND2_X1 maj_224_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_224_n21) );
  NAND2_X1 maj_224_U10 ( .A1(maj_224_n21), .A2(maj_224_n20), .ZN(maj_224_n23)
         );
  XOR2_X1 maj_224_U9 ( .A(u_1_1[2]), .B(maj_224_n24), .Z(maj_224_n26) );
  XOR2_X1 maj_224_U8 ( .A(u_1_1[5]), .B(maj_224_n25), .Z(maj_224_n27) );
  XOR2_X1 maj_224_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_224_n24) );
  XOR2_X1 maj_224_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_224_n25) );
  OR2_X1 maj_224_U5 ( .A1(maj_224_n23), .A2(maj_224_n22), .ZN(maj_224_n32) );
  NAND2_X1 maj_224_U4 ( .A1(maj_224_n22), .A2(maj_224_n23), .ZN(maj_224_n34)
         );
  NAND2_X1 maj_224_U3 ( .A1(maj_224_n32), .A2(maj_224_n31), .ZN(maj_224_n33)
         );
  NAND2_X1 maj_224_U2 ( .A1(maj_224_n34), .A2(maj_224_n33), .ZN(maj_224_port_o) );
  OR2_X1 maj_225_U19 ( .A1(maj_225_n27), .A2(maj_225_n26), .ZN(maj_225_n28) );
  NAND2_X1 maj_225_U18 ( .A1(v_1_1[6]), .A2(maj_225_n28), .ZN(maj_225_n29) );
  NAND2_X1 maj_225_U17 ( .A1(maj_225_n26), .A2(maj_225_n27), .ZN(maj_225_n30)
         );
  NAND2_X1 maj_225_U16 ( .A1(maj_225_n30), .A2(maj_225_n29), .ZN(maj_225_n31)
         );
  NAND2_X1 maj_225_U15 ( .A1(v_1_1[5]), .A2(maj_225_n25), .ZN(maj_225_n18) );
  NAND2_X1 maj_225_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_225_n19) );
  NAND2_X1 maj_225_U13 ( .A1(maj_225_n19), .A2(maj_225_n18), .ZN(maj_225_n22)
         );
  NAND2_X1 maj_225_U12 ( .A1(v_1_1[2]), .A2(maj_225_n24), .ZN(maj_225_n20) );
  NAND2_X1 maj_225_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_225_n21) );
  NAND2_X1 maj_225_U10 ( .A1(maj_225_n21), .A2(maj_225_n20), .ZN(maj_225_n23)
         );
  XOR2_X1 maj_225_U9 ( .A(v_1_1[2]), .B(maj_225_n24), .Z(maj_225_n26) );
  XOR2_X1 maj_225_U8 ( .A(v_1_1[5]), .B(maj_225_n25), .Z(maj_225_n27) );
  XOR2_X1 maj_225_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_225_n24) );
  XOR2_X1 maj_225_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_225_n25) );
  OR2_X1 maj_225_U5 ( .A1(maj_225_n23), .A2(maj_225_n22), .ZN(maj_225_n32) );
  NAND2_X1 maj_225_U4 ( .A1(maj_225_n22), .A2(maj_225_n23), .ZN(maj_225_n34)
         );
  NAND2_X1 maj_225_U3 ( .A1(maj_225_n32), .A2(maj_225_n31), .ZN(maj_225_n33)
         );
  NAND2_X1 maj_225_U2 ( .A1(maj_225_n34), .A2(maj_225_n33), .ZN(maj_225_port_o) );
  OR2_X1 maj_226_U19 ( .A1(maj_226_n27), .A2(maj_226_n26), .ZN(maj_226_n28) );
  NAND2_X1 maj_226_U18 ( .A1(u_1_2[6]), .A2(maj_226_n28), .ZN(maj_226_n29) );
  NAND2_X1 maj_226_U17 ( .A1(maj_226_n26), .A2(maj_226_n27), .ZN(maj_226_n30)
         );
  NAND2_X1 maj_226_U16 ( .A1(maj_226_n30), .A2(maj_226_n29), .ZN(maj_226_n31)
         );
  NAND2_X1 maj_226_U15 ( .A1(u_1_2[5]), .A2(maj_226_n25), .ZN(maj_226_n18) );
  NAND2_X1 maj_226_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_226_n19) );
  NAND2_X1 maj_226_U13 ( .A1(maj_226_n19), .A2(maj_226_n18), .ZN(maj_226_n22)
         );
  NAND2_X1 maj_226_U12 ( .A1(u_1_2[2]), .A2(maj_226_n24), .ZN(maj_226_n20) );
  NAND2_X1 maj_226_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_226_n21) );
  NAND2_X1 maj_226_U10 ( .A1(maj_226_n21), .A2(maj_226_n20), .ZN(maj_226_n23)
         );
  XOR2_X1 maj_226_U9 ( .A(u_1_2[2]), .B(maj_226_n24), .Z(maj_226_n26) );
  XOR2_X1 maj_226_U8 ( .A(u_1_2[5]), .B(maj_226_n25), .Z(maj_226_n27) );
  XOR2_X1 maj_226_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_226_n24) );
  XOR2_X1 maj_226_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_226_n25) );
  OR2_X1 maj_226_U5 ( .A1(maj_226_n23), .A2(maj_226_n22), .ZN(maj_226_n32) );
  NAND2_X1 maj_226_U4 ( .A1(maj_226_n22), .A2(maj_226_n23), .ZN(maj_226_n34)
         );
  NAND2_X1 maj_226_U3 ( .A1(maj_226_n32), .A2(maj_226_n31), .ZN(maj_226_n33)
         );
  NAND2_X1 maj_226_U2 ( .A1(maj_226_n34), .A2(maj_226_n33), .ZN(maj_226_port_o) );
  OR2_X1 maj_227_U19 ( .A1(maj_227_n27), .A2(maj_227_n26), .ZN(maj_227_n28) );
  NAND2_X1 maj_227_U18 ( .A1(v_1_2[6]), .A2(maj_227_n28), .ZN(maj_227_n29) );
  NAND2_X1 maj_227_U17 ( .A1(maj_227_n26), .A2(maj_227_n27), .ZN(maj_227_n30)
         );
  NAND2_X1 maj_227_U16 ( .A1(maj_227_n30), .A2(maj_227_n29), .ZN(maj_227_n31)
         );
  NAND2_X1 maj_227_U15 ( .A1(v_1_2[5]), .A2(maj_227_n25), .ZN(maj_227_n18) );
  NAND2_X1 maj_227_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_227_n19) );
  NAND2_X1 maj_227_U13 ( .A1(maj_227_n19), .A2(maj_227_n18), .ZN(maj_227_n22)
         );
  NAND2_X1 maj_227_U12 ( .A1(v_1_2[2]), .A2(maj_227_n24), .ZN(maj_227_n20) );
  NAND2_X1 maj_227_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_227_n21) );
  NAND2_X1 maj_227_U10 ( .A1(maj_227_n21), .A2(maj_227_n20), .ZN(maj_227_n23)
         );
  XOR2_X1 maj_227_U9 ( .A(v_1_2[2]), .B(maj_227_n24), .Z(maj_227_n26) );
  XOR2_X1 maj_227_U8 ( .A(v_1_2[5]), .B(maj_227_n25), .Z(maj_227_n27) );
  XOR2_X1 maj_227_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_227_n24) );
  XOR2_X1 maj_227_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_227_n25) );
  OR2_X1 maj_227_U5 ( .A1(maj_227_n23), .A2(maj_227_n22), .ZN(maj_227_n32) );
  NAND2_X1 maj_227_U4 ( .A1(maj_227_n22), .A2(maj_227_n23), .ZN(maj_227_n34)
         );
  NAND2_X1 maj_227_U3 ( .A1(maj_227_n32), .A2(maj_227_n31), .ZN(maj_227_n33)
         );
  NAND2_X1 maj_227_U2 ( .A1(maj_227_n34), .A2(maj_227_n33), .ZN(maj_227_port_o) );
  OR2_X1 maj_228_U19 ( .A1(maj_228_n27), .A2(maj_228_n26), .ZN(maj_228_n28) );
  NAND2_X1 maj_228_U18 ( .A1(u_2_0[6]), .A2(maj_228_n28), .ZN(maj_228_n29) );
  NAND2_X1 maj_228_U17 ( .A1(maj_228_n26), .A2(maj_228_n27), .ZN(maj_228_n30)
         );
  NAND2_X1 maj_228_U16 ( .A1(maj_228_n30), .A2(maj_228_n29), .ZN(maj_228_n31)
         );
  NAND2_X1 maj_228_U15 ( .A1(u_2_0[5]), .A2(maj_228_n25), .ZN(maj_228_n18) );
  NAND2_X1 maj_228_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_228_n19) );
  NAND2_X1 maj_228_U13 ( .A1(maj_228_n19), .A2(maj_228_n18), .ZN(maj_228_n22)
         );
  NAND2_X1 maj_228_U12 ( .A1(u_2_0[2]), .A2(maj_228_n24), .ZN(maj_228_n20) );
  NAND2_X1 maj_228_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_228_n21) );
  NAND2_X1 maj_228_U10 ( .A1(maj_228_n21), .A2(maj_228_n20), .ZN(maj_228_n23)
         );
  XOR2_X1 maj_228_U9 ( .A(u_2_0[2]), .B(maj_228_n24), .Z(maj_228_n26) );
  XOR2_X1 maj_228_U8 ( .A(u_2_0[5]), .B(maj_228_n25), .Z(maj_228_n27) );
  XOR2_X1 maj_228_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_228_n24) );
  XOR2_X1 maj_228_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_228_n25) );
  OR2_X1 maj_228_U5 ( .A1(maj_228_n23), .A2(maj_228_n22), .ZN(maj_228_n32) );
  NAND2_X1 maj_228_U4 ( .A1(maj_228_n22), .A2(maj_228_n23), .ZN(maj_228_n34)
         );
  NAND2_X1 maj_228_U3 ( .A1(maj_228_n32), .A2(maj_228_n31), .ZN(maj_228_n33)
         );
  NAND2_X1 maj_228_U2 ( .A1(maj_228_n34), .A2(maj_228_n33), .ZN(maj_228_port_o) );
  OR2_X1 maj_229_U19 ( .A1(maj_229_n27), .A2(maj_229_n26), .ZN(maj_229_n28) );
  NAND2_X1 maj_229_U18 ( .A1(v_2_0[6]), .A2(maj_229_n28), .ZN(maj_229_n29) );
  NAND2_X1 maj_229_U17 ( .A1(maj_229_n26), .A2(maj_229_n27), .ZN(maj_229_n30)
         );
  NAND2_X1 maj_229_U16 ( .A1(maj_229_n30), .A2(maj_229_n29), .ZN(maj_229_n31)
         );
  NAND2_X1 maj_229_U15 ( .A1(v_2_0[5]), .A2(maj_229_n25), .ZN(maj_229_n18) );
  NAND2_X1 maj_229_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_229_n19) );
  NAND2_X1 maj_229_U13 ( .A1(maj_229_n19), .A2(maj_229_n18), .ZN(maj_229_n22)
         );
  NAND2_X1 maj_229_U12 ( .A1(v_2_0[2]), .A2(maj_229_n24), .ZN(maj_229_n20) );
  NAND2_X1 maj_229_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_229_n21) );
  NAND2_X1 maj_229_U10 ( .A1(maj_229_n21), .A2(maj_229_n20), .ZN(maj_229_n23)
         );
  XOR2_X1 maj_229_U9 ( .A(v_2_0[2]), .B(maj_229_n24), .Z(maj_229_n26) );
  XOR2_X1 maj_229_U8 ( .A(v_2_0[5]), .B(maj_229_n25), .Z(maj_229_n27) );
  XOR2_X1 maj_229_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_229_n24) );
  XOR2_X1 maj_229_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_229_n25) );
  OR2_X1 maj_229_U5 ( .A1(maj_229_n23), .A2(maj_229_n22), .ZN(maj_229_n32) );
  NAND2_X1 maj_229_U4 ( .A1(maj_229_n22), .A2(maj_229_n23), .ZN(maj_229_n34)
         );
  NAND2_X1 maj_229_U3 ( .A1(maj_229_n32), .A2(maj_229_n31), .ZN(maj_229_n33)
         );
  NAND2_X1 maj_229_U2 ( .A1(maj_229_n34), .A2(maj_229_n33), .ZN(maj_229_port_o) );
  OR2_X1 maj_230_U19 ( .A1(maj_230_n27), .A2(maj_230_n26), .ZN(maj_230_n28) );
  NAND2_X1 maj_230_U18 ( .A1(u_2_1[6]), .A2(maj_230_n28), .ZN(maj_230_n29) );
  NAND2_X1 maj_230_U17 ( .A1(maj_230_n26), .A2(maj_230_n27), .ZN(maj_230_n30)
         );
  NAND2_X1 maj_230_U16 ( .A1(maj_230_n30), .A2(maj_230_n29), .ZN(maj_230_n31)
         );
  NAND2_X1 maj_230_U15 ( .A1(u_2_1[5]), .A2(maj_230_n25), .ZN(maj_230_n18) );
  NAND2_X1 maj_230_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_230_n19) );
  NAND2_X1 maj_230_U13 ( .A1(maj_230_n19), .A2(maj_230_n18), .ZN(maj_230_n22)
         );
  NAND2_X1 maj_230_U12 ( .A1(u_2_1[2]), .A2(maj_230_n24), .ZN(maj_230_n20) );
  NAND2_X1 maj_230_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_230_n21) );
  NAND2_X1 maj_230_U10 ( .A1(maj_230_n21), .A2(maj_230_n20), .ZN(maj_230_n23)
         );
  XOR2_X1 maj_230_U9 ( .A(u_2_1[2]), .B(maj_230_n24), .Z(maj_230_n26) );
  XOR2_X1 maj_230_U8 ( .A(u_2_1[5]), .B(maj_230_n25), .Z(maj_230_n27) );
  XOR2_X1 maj_230_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_230_n24) );
  XOR2_X1 maj_230_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_230_n25) );
  OR2_X1 maj_230_U5 ( .A1(maj_230_n23), .A2(maj_230_n22), .ZN(maj_230_n32) );
  NAND2_X1 maj_230_U4 ( .A1(maj_230_n22), .A2(maj_230_n23), .ZN(maj_230_n34)
         );
  NAND2_X1 maj_230_U3 ( .A1(maj_230_n32), .A2(maj_230_n31), .ZN(maj_230_n33)
         );
  NAND2_X1 maj_230_U2 ( .A1(maj_230_n34), .A2(maj_230_n33), .ZN(maj_230_port_o) );
  OR2_X1 maj_231_U19 ( .A1(maj_231_n27), .A2(maj_231_n26), .ZN(maj_231_n28) );
  NAND2_X1 maj_231_U18 ( .A1(v_2_1[6]), .A2(maj_231_n28), .ZN(maj_231_n29) );
  NAND2_X1 maj_231_U17 ( .A1(maj_231_n26), .A2(maj_231_n27), .ZN(maj_231_n30)
         );
  NAND2_X1 maj_231_U16 ( .A1(maj_231_n30), .A2(maj_231_n29), .ZN(maj_231_n31)
         );
  NAND2_X1 maj_231_U15 ( .A1(v_2_1[5]), .A2(maj_231_n25), .ZN(maj_231_n18) );
  NAND2_X1 maj_231_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_231_n19) );
  NAND2_X1 maj_231_U13 ( .A1(maj_231_n19), .A2(maj_231_n18), .ZN(maj_231_n22)
         );
  NAND2_X1 maj_231_U12 ( .A1(v_2_1[2]), .A2(maj_231_n24), .ZN(maj_231_n20) );
  NAND2_X1 maj_231_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_231_n21) );
  NAND2_X1 maj_231_U10 ( .A1(maj_231_n21), .A2(maj_231_n20), .ZN(maj_231_n23)
         );
  XOR2_X1 maj_231_U9 ( .A(v_2_1[2]), .B(maj_231_n24), .Z(maj_231_n26) );
  XOR2_X1 maj_231_U8 ( .A(v_2_1[5]), .B(maj_231_n25), .Z(maj_231_n27) );
  XOR2_X1 maj_231_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_231_n24) );
  XOR2_X1 maj_231_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_231_n25) );
  OR2_X1 maj_231_U5 ( .A1(maj_231_n23), .A2(maj_231_n22), .ZN(maj_231_n32) );
  NAND2_X1 maj_231_U4 ( .A1(maj_231_n22), .A2(maj_231_n23), .ZN(maj_231_n34)
         );
  NAND2_X1 maj_231_U3 ( .A1(maj_231_n32), .A2(maj_231_n31), .ZN(maj_231_n33)
         );
  NAND2_X1 maj_231_U2 ( .A1(maj_231_n34), .A2(maj_231_n33), .ZN(maj_231_port_o) );
  OR2_X1 maj_232_U19 ( .A1(maj_232_n27), .A2(maj_232_n26), .ZN(maj_232_n28) );
  NAND2_X1 maj_232_U18 ( .A1(u_2_2[6]), .A2(maj_232_n28), .ZN(maj_232_n29) );
  NAND2_X1 maj_232_U17 ( .A1(maj_232_n26), .A2(maj_232_n27), .ZN(maj_232_n30)
         );
  NAND2_X1 maj_232_U16 ( .A1(maj_232_n30), .A2(maj_232_n29), .ZN(maj_232_n31)
         );
  NAND2_X1 maj_232_U15 ( .A1(u_2_2[5]), .A2(maj_232_n25), .ZN(maj_232_n18) );
  NAND2_X1 maj_232_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_232_n19) );
  NAND2_X1 maj_232_U13 ( .A1(maj_232_n19), .A2(maj_232_n18), .ZN(maj_232_n22)
         );
  NAND2_X1 maj_232_U12 ( .A1(u_2_2[2]), .A2(maj_232_n24), .ZN(maj_232_n20) );
  NAND2_X1 maj_232_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_232_n21) );
  NAND2_X1 maj_232_U10 ( .A1(maj_232_n21), .A2(maj_232_n20), .ZN(maj_232_n23)
         );
  XOR2_X1 maj_232_U9 ( .A(u_2_2[2]), .B(maj_232_n24), .Z(maj_232_n26) );
  XOR2_X1 maj_232_U8 ( .A(u_2_2[5]), .B(maj_232_n25), .Z(maj_232_n27) );
  XOR2_X1 maj_232_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_232_n24) );
  XOR2_X1 maj_232_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_232_n25) );
  OR2_X1 maj_232_U5 ( .A1(maj_232_n23), .A2(maj_232_n22), .ZN(maj_232_n32) );
  NAND2_X1 maj_232_U4 ( .A1(maj_232_n22), .A2(maj_232_n23), .ZN(maj_232_n34)
         );
  NAND2_X1 maj_232_U3 ( .A1(maj_232_n32), .A2(maj_232_n31), .ZN(maj_232_n33)
         );
  NAND2_X1 maj_232_U2 ( .A1(maj_232_n34), .A2(maj_232_n33), .ZN(maj_232_port_o) );
  OR2_X1 maj_233_U19 ( .A1(maj_233_n27), .A2(maj_233_n26), .ZN(maj_233_n28) );
  NAND2_X1 maj_233_U18 ( .A1(v_2_2[6]), .A2(maj_233_n28), .ZN(maj_233_n29) );
  NAND2_X1 maj_233_U17 ( .A1(maj_233_n26), .A2(maj_233_n27), .ZN(maj_233_n30)
         );
  NAND2_X1 maj_233_U16 ( .A1(maj_233_n30), .A2(maj_233_n29), .ZN(maj_233_n31)
         );
  NAND2_X1 maj_233_U15 ( .A1(v_2_2[5]), .A2(maj_233_n25), .ZN(maj_233_n18) );
  NAND2_X1 maj_233_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_233_n19) );
  NAND2_X1 maj_233_U13 ( .A1(maj_233_n19), .A2(maj_233_n18), .ZN(maj_233_n22)
         );
  NAND2_X1 maj_233_U12 ( .A1(v_2_2[2]), .A2(maj_233_n24), .ZN(maj_233_n20) );
  NAND2_X1 maj_233_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_233_n21) );
  NAND2_X1 maj_233_U10 ( .A1(maj_233_n21), .A2(maj_233_n20), .ZN(maj_233_n23)
         );
  XOR2_X1 maj_233_U9 ( .A(v_2_2[2]), .B(maj_233_n24), .Z(maj_233_n26) );
  XOR2_X1 maj_233_U8 ( .A(v_2_2[5]), .B(maj_233_n25), .Z(maj_233_n27) );
  XOR2_X1 maj_233_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_233_n24) );
  XOR2_X1 maj_233_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_233_n25) );
  OR2_X1 maj_233_U5 ( .A1(maj_233_n23), .A2(maj_233_n22), .ZN(maj_233_n32) );
  NAND2_X1 maj_233_U4 ( .A1(maj_233_n22), .A2(maj_233_n23), .ZN(maj_233_n34)
         );
  NAND2_X1 maj_233_U3 ( .A1(maj_233_n32), .A2(maj_233_n31), .ZN(maj_233_n33)
         );
  NAND2_X1 maj_233_U2 ( .A1(maj_233_n34), .A2(maj_233_n33), .ZN(maj_233_port_o) );
  OR2_X1 maj_234_U19 ( .A1(maj_234_n27), .A2(maj_234_n26), .ZN(maj_234_n28) );
  NAND2_X1 maj_234_U18 ( .A1(u_3_0[6]), .A2(maj_234_n28), .ZN(maj_234_n29) );
  NAND2_X1 maj_234_U17 ( .A1(maj_234_n26), .A2(maj_234_n27), .ZN(maj_234_n30)
         );
  NAND2_X1 maj_234_U16 ( .A1(maj_234_n30), .A2(maj_234_n29), .ZN(maj_234_n31)
         );
  NAND2_X1 maj_234_U15 ( .A1(u_3_0[5]), .A2(maj_234_n25), .ZN(maj_234_n18) );
  NAND2_X1 maj_234_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_234_n19) );
  NAND2_X1 maj_234_U13 ( .A1(maj_234_n19), .A2(maj_234_n18), .ZN(maj_234_n22)
         );
  NAND2_X1 maj_234_U12 ( .A1(u_3_0[2]), .A2(maj_234_n24), .ZN(maj_234_n20) );
  NAND2_X1 maj_234_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_234_n21) );
  NAND2_X1 maj_234_U10 ( .A1(maj_234_n21), .A2(maj_234_n20), .ZN(maj_234_n23)
         );
  XOR2_X1 maj_234_U9 ( .A(u_3_0[2]), .B(maj_234_n24), .Z(maj_234_n26) );
  XOR2_X1 maj_234_U8 ( .A(u_3_0[5]), .B(maj_234_n25), .Z(maj_234_n27) );
  XOR2_X1 maj_234_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_234_n24) );
  XOR2_X1 maj_234_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_234_n25) );
  OR2_X1 maj_234_U5 ( .A1(maj_234_n23), .A2(maj_234_n22), .ZN(maj_234_n32) );
  NAND2_X1 maj_234_U4 ( .A1(maj_234_n22), .A2(maj_234_n23), .ZN(maj_234_n34)
         );
  NAND2_X1 maj_234_U3 ( .A1(maj_234_n32), .A2(maj_234_n31), .ZN(maj_234_n33)
         );
  NAND2_X1 maj_234_U2 ( .A1(maj_234_n34), .A2(maj_234_n33), .ZN(maj_234_port_o) );
  OR2_X1 maj_235_U19 ( .A1(maj_235_n27), .A2(maj_235_n26), .ZN(maj_235_n28) );
  NAND2_X1 maj_235_U18 ( .A1(v_3_0[6]), .A2(maj_235_n28), .ZN(maj_235_n29) );
  NAND2_X1 maj_235_U17 ( .A1(maj_235_n26), .A2(maj_235_n27), .ZN(maj_235_n30)
         );
  NAND2_X1 maj_235_U16 ( .A1(maj_235_n30), .A2(maj_235_n29), .ZN(maj_235_n31)
         );
  NAND2_X1 maj_235_U15 ( .A1(v_3_0[5]), .A2(maj_235_n25), .ZN(maj_235_n18) );
  NAND2_X1 maj_235_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_235_n19) );
  NAND2_X1 maj_235_U13 ( .A1(maj_235_n19), .A2(maj_235_n18), .ZN(maj_235_n22)
         );
  NAND2_X1 maj_235_U12 ( .A1(v_3_0[2]), .A2(maj_235_n24), .ZN(maj_235_n20) );
  NAND2_X1 maj_235_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_235_n21) );
  NAND2_X1 maj_235_U10 ( .A1(maj_235_n21), .A2(maj_235_n20), .ZN(maj_235_n23)
         );
  XOR2_X1 maj_235_U9 ( .A(v_3_0[2]), .B(maj_235_n24), .Z(maj_235_n26) );
  XOR2_X1 maj_235_U8 ( .A(v_3_0[5]), .B(maj_235_n25), .Z(maj_235_n27) );
  XOR2_X1 maj_235_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_235_n24) );
  XOR2_X1 maj_235_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_235_n25) );
  OR2_X1 maj_235_U5 ( .A1(maj_235_n23), .A2(maj_235_n22), .ZN(maj_235_n32) );
  NAND2_X1 maj_235_U4 ( .A1(maj_235_n22), .A2(maj_235_n23), .ZN(maj_235_n34)
         );
  NAND2_X1 maj_235_U3 ( .A1(maj_235_n32), .A2(maj_235_n31), .ZN(maj_235_n33)
         );
  NAND2_X1 maj_235_U2 ( .A1(maj_235_n34), .A2(maj_235_n33), .ZN(maj_235_port_o) );
  OR2_X1 maj_236_U19 ( .A1(maj_236_n27), .A2(maj_236_n26), .ZN(maj_236_n28) );
  NAND2_X1 maj_236_U18 ( .A1(u_3_1[6]), .A2(maj_236_n28), .ZN(maj_236_n29) );
  NAND2_X1 maj_236_U17 ( .A1(maj_236_n26), .A2(maj_236_n27), .ZN(maj_236_n30)
         );
  NAND2_X1 maj_236_U16 ( .A1(maj_236_n30), .A2(maj_236_n29), .ZN(maj_236_n31)
         );
  NAND2_X1 maj_236_U15 ( .A1(u_3_1[5]), .A2(maj_236_n25), .ZN(maj_236_n18) );
  NAND2_X1 maj_236_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_236_n19) );
  NAND2_X1 maj_236_U13 ( .A1(maj_236_n19), .A2(maj_236_n18), .ZN(maj_236_n22)
         );
  NAND2_X1 maj_236_U12 ( .A1(u_3_1[2]), .A2(maj_236_n24), .ZN(maj_236_n20) );
  NAND2_X1 maj_236_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_236_n21) );
  NAND2_X1 maj_236_U10 ( .A1(maj_236_n21), .A2(maj_236_n20), .ZN(maj_236_n23)
         );
  XOR2_X1 maj_236_U9 ( .A(u_3_1[2]), .B(maj_236_n24), .Z(maj_236_n26) );
  XOR2_X1 maj_236_U8 ( .A(u_3_1[5]), .B(maj_236_n25), .Z(maj_236_n27) );
  XOR2_X1 maj_236_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_236_n24) );
  XOR2_X1 maj_236_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_236_n25) );
  OR2_X1 maj_236_U5 ( .A1(maj_236_n23), .A2(maj_236_n22), .ZN(maj_236_n32) );
  NAND2_X1 maj_236_U4 ( .A1(maj_236_n22), .A2(maj_236_n23), .ZN(maj_236_n34)
         );
  NAND2_X1 maj_236_U3 ( .A1(maj_236_n32), .A2(maj_236_n31), .ZN(maj_236_n33)
         );
  NAND2_X1 maj_236_U2 ( .A1(maj_236_n34), .A2(maj_236_n33), .ZN(maj_236_port_o) );
  OR2_X1 maj_237_U19 ( .A1(maj_237_n27), .A2(maj_237_n26), .ZN(maj_237_n28) );
  NAND2_X1 maj_237_U18 ( .A1(v_3_1[6]), .A2(maj_237_n28), .ZN(maj_237_n29) );
  NAND2_X1 maj_237_U17 ( .A1(maj_237_n26), .A2(maj_237_n27), .ZN(maj_237_n30)
         );
  NAND2_X1 maj_237_U16 ( .A1(maj_237_n30), .A2(maj_237_n29), .ZN(maj_237_n31)
         );
  NAND2_X1 maj_237_U15 ( .A1(v_3_1[5]), .A2(maj_237_n25), .ZN(maj_237_n18) );
  NAND2_X1 maj_237_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_237_n19) );
  NAND2_X1 maj_237_U13 ( .A1(maj_237_n19), .A2(maj_237_n18), .ZN(maj_237_n22)
         );
  NAND2_X1 maj_237_U12 ( .A1(v_3_1[2]), .A2(maj_237_n24), .ZN(maj_237_n20) );
  NAND2_X1 maj_237_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_237_n21) );
  NAND2_X1 maj_237_U10 ( .A1(maj_237_n21), .A2(maj_237_n20), .ZN(maj_237_n23)
         );
  XOR2_X1 maj_237_U9 ( .A(v_3_1[2]), .B(maj_237_n24), .Z(maj_237_n26) );
  XOR2_X1 maj_237_U8 ( .A(v_3_1[5]), .B(maj_237_n25), .Z(maj_237_n27) );
  XOR2_X1 maj_237_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_237_n24) );
  XOR2_X1 maj_237_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_237_n25) );
  OR2_X1 maj_237_U5 ( .A1(maj_237_n23), .A2(maj_237_n22), .ZN(maj_237_n32) );
  NAND2_X1 maj_237_U4 ( .A1(maj_237_n22), .A2(maj_237_n23), .ZN(maj_237_n34)
         );
  NAND2_X1 maj_237_U3 ( .A1(maj_237_n32), .A2(maj_237_n31), .ZN(maj_237_n33)
         );
  NAND2_X1 maj_237_U2 ( .A1(maj_237_n34), .A2(maj_237_n33), .ZN(maj_237_port_o) );
  OR2_X1 maj_238_U19 ( .A1(maj_238_n27), .A2(maj_238_n26), .ZN(maj_238_n28) );
  NAND2_X1 maj_238_U18 ( .A1(u_3_2[6]), .A2(maj_238_n28), .ZN(maj_238_n29) );
  NAND2_X1 maj_238_U17 ( .A1(maj_238_n26), .A2(maj_238_n27), .ZN(maj_238_n30)
         );
  NAND2_X1 maj_238_U16 ( .A1(maj_238_n30), .A2(maj_238_n29), .ZN(maj_238_n31)
         );
  NAND2_X1 maj_238_U15 ( .A1(u_3_2[5]), .A2(maj_238_n25), .ZN(maj_238_n18) );
  NAND2_X1 maj_238_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_238_n19) );
  NAND2_X1 maj_238_U13 ( .A1(maj_238_n19), .A2(maj_238_n18), .ZN(maj_238_n22)
         );
  NAND2_X1 maj_238_U12 ( .A1(u_3_2[2]), .A2(maj_238_n24), .ZN(maj_238_n20) );
  NAND2_X1 maj_238_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_238_n21) );
  NAND2_X1 maj_238_U10 ( .A1(maj_238_n21), .A2(maj_238_n20), .ZN(maj_238_n23)
         );
  XOR2_X1 maj_238_U9 ( .A(u_3_2[2]), .B(maj_238_n24), .Z(maj_238_n26) );
  XOR2_X1 maj_238_U8 ( .A(u_3_2[5]), .B(maj_238_n25), .Z(maj_238_n27) );
  XOR2_X1 maj_238_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_238_n24) );
  XOR2_X1 maj_238_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_238_n25) );
  OR2_X1 maj_238_U5 ( .A1(maj_238_n23), .A2(maj_238_n22), .ZN(maj_238_n32) );
  NAND2_X1 maj_238_U4 ( .A1(maj_238_n22), .A2(maj_238_n23), .ZN(maj_238_n34)
         );
  NAND2_X1 maj_238_U3 ( .A1(maj_238_n32), .A2(maj_238_n31), .ZN(maj_238_n33)
         );
  NAND2_X1 maj_238_U2 ( .A1(maj_238_n34), .A2(maj_238_n33), .ZN(maj_238_port_o) );
  OR2_X1 maj_239_U19 ( .A1(maj_239_n27), .A2(maj_239_n26), .ZN(maj_239_n28) );
  NAND2_X1 maj_239_U18 ( .A1(v_3_2[6]), .A2(maj_239_n28), .ZN(maj_239_n29) );
  NAND2_X1 maj_239_U17 ( .A1(maj_239_n26), .A2(maj_239_n27), .ZN(maj_239_n30)
         );
  NAND2_X1 maj_239_U16 ( .A1(maj_239_n30), .A2(maj_239_n29), .ZN(maj_239_n31)
         );
  NAND2_X1 maj_239_U15 ( .A1(v_3_2[5]), .A2(maj_239_n25), .ZN(maj_239_n18) );
  NAND2_X1 maj_239_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_239_n19) );
  NAND2_X1 maj_239_U13 ( .A1(maj_239_n19), .A2(maj_239_n18), .ZN(maj_239_n22)
         );
  NAND2_X1 maj_239_U12 ( .A1(v_3_2[2]), .A2(maj_239_n24), .ZN(maj_239_n20) );
  NAND2_X1 maj_239_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_239_n21) );
  NAND2_X1 maj_239_U10 ( .A1(maj_239_n21), .A2(maj_239_n20), .ZN(maj_239_n23)
         );
  XOR2_X1 maj_239_U9 ( .A(v_3_2[2]), .B(maj_239_n24), .Z(maj_239_n26) );
  XOR2_X1 maj_239_U8 ( .A(v_3_2[5]), .B(maj_239_n25), .Z(maj_239_n27) );
  XOR2_X1 maj_239_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_239_n24) );
  XOR2_X1 maj_239_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_239_n25) );
  OR2_X1 maj_239_U5 ( .A1(maj_239_n23), .A2(maj_239_n22), .ZN(maj_239_n32) );
  NAND2_X1 maj_239_U4 ( .A1(maj_239_n22), .A2(maj_239_n23), .ZN(maj_239_n34)
         );
  NAND2_X1 maj_239_U3 ( .A1(maj_239_n32), .A2(maj_239_n31), .ZN(maj_239_n33)
         );
  NAND2_X1 maj_239_U2 ( .A1(maj_239_n34), .A2(maj_239_n33), .ZN(maj_239_port_o) );
  OR2_X1 maj_240_U19 ( .A1(maj_240_n27), .A2(maj_240_n26), .ZN(maj_240_n28) );
  NAND2_X1 maj_240_U18 ( .A1(u_0_0[6]), .A2(maj_240_n28), .ZN(maj_240_n29) );
  NAND2_X1 maj_240_U17 ( .A1(maj_240_n26), .A2(maj_240_n27), .ZN(maj_240_n30)
         );
  NAND2_X1 maj_240_U16 ( .A1(maj_240_n30), .A2(maj_240_n29), .ZN(maj_240_n31)
         );
  NAND2_X1 maj_240_U15 ( .A1(u_0_0[5]), .A2(maj_240_n25), .ZN(maj_240_n18) );
  NAND2_X1 maj_240_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_240_n19) );
  NAND2_X1 maj_240_U13 ( .A1(maj_240_n19), .A2(maj_240_n18), .ZN(maj_240_n22)
         );
  NAND2_X1 maj_240_U12 ( .A1(u_0_0[2]), .A2(maj_240_n24), .ZN(maj_240_n20) );
  NAND2_X1 maj_240_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_240_n21) );
  NAND2_X1 maj_240_U10 ( .A1(maj_240_n21), .A2(maj_240_n20), .ZN(maj_240_n23)
         );
  XOR2_X1 maj_240_U9 ( .A(u_0_0[2]), .B(maj_240_n24), .Z(maj_240_n26) );
  XOR2_X1 maj_240_U8 ( .A(u_0_0[5]), .B(maj_240_n25), .Z(maj_240_n27) );
  XOR2_X1 maj_240_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_240_n24) );
  XOR2_X1 maj_240_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_240_n25) );
  OR2_X1 maj_240_U5 ( .A1(maj_240_n23), .A2(maj_240_n22), .ZN(maj_240_n32) );
  NAND2_X1 maj_240_U4 ( .A1(maj_240_n22), .A2(maj_240_n23), .ZN(maj_240_n34)
         );
  NAND2_X1 maj_240_U3 ( .A1(maj_240_n32), .A2(maj_240_n31), .ZN(maj_240_n33)
         );
  NAND2_X1 maj_240_U2 ( .A1(maj_240_n34), .A2(maj_240_n33), .ZN(maj_240_port_o) );
  OR2_X1 maj_241_U19 ( .A1(maj_241_n27), .A2(maj_241_n26), .ZN(maj_241_n28) );
  NAND2_X1 maj_241_U18 ( .A1(v_0_0[6]), .A2(maj_241_n28), .ZN(maj_241_n29) );
  NAND2_X1 maj_241_U17 ( .A1(maj_241_n26), .A2(maj_241_n27), .ZN(maj_241_n30)
         );
  NAND2_X1 maj_241_U16 ( .A1(maj_241_n30), .A2(maj_241_n29), .ZN(maj_241_n31)
         );
  NAND2_X1 maj_241_U15 ( .A1(v_0_0[5]), .A2(maj_241_n25), .ZN(maj_241_n18) );
  NAND2_X1 maj_241_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_241_n19) );
  NAND2_X1 maj_241_U13 ( .A1(maj_241_n19), .A2(maj_241_n18), .ZN(maj_241_n22)
         );
  NAND2_X1 maj_241_U12 ( .A1(v_0_0[2]), .A2(maj_241_n24), .ZN(maj_241_n20) );
  NAND2_X1 maj_241_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_241_n21) );
  NAND2_X1 maj_241_U10 ( .A1(maj_241_n21), .A2(maj_241_n20), .ZN(maj_241_n23)
         );
  XOR2_X1 maj_241_U9 ( .A(v_0_0[2]), .B(maj_241_n24), .Z(maj_241_n26) );
  XOR2_X1 maj_241_U8 ( .A(v_0_0[5]), .B(maj_241_n25), .Z(maj_241_n27) );
  XOR2_X1 maj_241_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_241_n24) );
  XOR2_X1 maj_241_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_241_n25) );
  OR2_X1 maj_241_U5 ( .A1(maj_241_n23), .A2(maj_241_n22), .ZN(maj_241_n32) );
  NAND2_X1 maj_241_U4 ( .A1(maj_241_n22), .A2(maj_241_n23), .ZN(maj_241_n34)
         );
  NAND2_X1 maj_241_U3 ( .A1(maj_241_n32), .A2(maj_241_n31), .ZN(maj_241_n33)
         );
  NAND2_X1 maj_241_U2 ( .A1(maj_241_n34), .A2(maj_241_n33), .ZN(maj_241_port_o) );
  OR2_X1 maj_242_U19 ( .A1(maj_242_n27), .A2(maj_242_n26), .ZN(maj_242_n28) );
  NAND2_X1 maj_242_U18 ( .A1(u_0_1[6]), .A2(maj_242_n28), .ZN(maj_242_n29) );
  NAND2_X1 maj_242_U17 ( .A1(maj_242_n26), .A2(maj_242_n27), .ZN(maj_242_n30)
         );
  NAND2_X1 maj_242_U16 ( .A1(maj_242_n30), .A2(maj_242_n29), .ZN(maj_242_n31)
         );
  NAND2_X1 maj_242_U15 ( .A1(u_0_1[5]), .A2(maj_242_n25), .ZN(maj_242_n18) );
  NAND2_X1 maj_242_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_242_n19) );
  NAND2_X1 maj_242_U13 ( .A1(maj_242_n19), .A2(maj_242_n18), .ZN(maj_242_n22)
         );
  NAND2_X1 maj_242_U12 ( .A1(u_0_1[2]), .A2(maj_242_n24), .ZN(maj_242_n20) );
  NAND2_X1 maj_242_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_242_n21) );
  NAND2_X1 maj_242_U10 ( .A1(maj_242_n21), .A2(maj_242_n20), .ZN(maj_242_n23)
         );
  XOR2_X1 maj_242_U9 ( .A(u_0_1[2]), .B(maj_242_n24), .Z(maj_242_n26) );
  XOR2_X1 maj_242_U8 ( .A(u_0_1[5]), .B(maj_242_n25), .Z(maj_242_n27) );
  XOR2_X1 maj_242_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_242_n24) );
  XOR2_X1 maj_242_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_242_n25) );
  OR2_X1 maj_242_U5 ( .A1(maj_242_n23), .A2(maj_242_n22), .ZN(maj_242_n32) );
  NAND2_X1 maj_242_U4 ( .A1(maj_242_n22), .A2(maj_242_n23), .ZN(maj_242_n34)
         );
  NAND2_X1 maj_242_U3 ( .A1(maj_242_n32), .A2(maj_242_n31), .ZN(maj_242_n33)
         );
  NAND2_X1 maj_242_U2 ( .A1(maj_242_n34), .A2(maj_242_n33), .ZN(maj_242_port_o) );
  OR2_X1 maj_243_U19 ( .A1(maj_243_n27), .A2(maj_243_n26), .ZN(maj_243_n28) );
  NAND2_X1 maj_243_U18 ( .A1(v_0_1[6]), .A2(maj_243_n28), .ZN(maj_243_n29) );
  NAND2_X1 maj_243_U17 ( .A1(maj_243_n26), .A2(maj_243_n27), .ZN(maj_243_n30)
         );
  NAND2_X1 maj_243_U16 ( .A1(maj_243_n30), .A2(maj_243_n29), .ZN(maj_243_n31)
         );
  NAND2_X1 maj_243_U15 ( .A1(v_0_1[5]), .A2(maj_243_n25), .ZN(maj_243_n18) );
  NAND2_X1 maj_243_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_243_n19) );
  NAND2_X1 maj_243_U13 ( .A1(maj_243_n19), .A2(maj_243_n18), .ZN(maj_243_n22)
         );
  NAND2_X1 maj_243_U12 ( .A1(v_0_1[2]), .A2(maj_243_n24), .ZN(maj_243_n20) );
  NAND2_X1 maj_243_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_243_n21) );
  NAND2_X1 maj_243_U10 ( .A1(maj_243_n21), .A2(maj_243_n20), .ZN(maj_243_n23)
         );
  XOR2_X1 maj_243_U9 ( .A(v_0_1[2]), .B(maj_243_n24), .Z(maj_243_n26) );
  XOR2_X1 maj_243_U8 ( .A(v_0_1[5]), .B(maj_243_n25), .Z(maj_243_n27) );
  XOR2_X1 maj_243_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_243_n24) );
  XOR2_X1 maj_243_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_243_n25) );
  OR2_X1 maj_243_U5 ( .A1(maj_243_n23), .A2(maj_243_n22), .ZN(maj_243_n32) );
  NAND2_X1 maj_243_U4 ( .A1(maj_243_n22), .A2(maj_243_n23), .ZN(maj_243_n34)
         );
  NAND2_X1 maj_243_U3 ( .A1(maj_243_n32), .A2(maj_243_n31), .ZN(maj_243_n33)
         );
  NAND2_X1 maj_243_U2 ( .A1(maj_243_n34), .A2(maj_243_n33), .ZN(maj_243_port_o) );
  OR2_X1 maj_244_U19 ( .A1(maj_244_n27), .A2(maj_244_n26), .ZN(maj_244_n28) );
  NAND2_X1 maj_244_U18 ( .A1(u_0_2[6]), .A2(maj_244_n28), .ZN(maj_244_n29) );
  NAND2_X1 maj_244_U17 ( .A1(maj_244_n26), .A2(maj_244_n27), .ZN(maj_244_n30)
         );
  NAND2_X1 maj_244_U16 ( .A1(maj_244_n30), .A2(maj_244_n29), .ZN(maj_244_n31)
         );
  NAND2_X1 maj_244_U15 ( .A1(u_0_2[5]), .A2(maj_244_n25), .ZN(maj_244_n18) );
  NAND2_X1 maj_244_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_244_n19) );
  NAND2_X1 maj_244_U13 ( .A1(maj_244_n19), .A2(maj_244_n18), .ZN(maj_244_n22)
         );
  NAND2_X1 maj_244_U12 ( .A1(u_0_2[2]), .A2(maj_244_n24), .ZN(maj_244_n20) );
  NAND2_X1 maj_244_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_244_n21) );
  NAND2_X1 maj_244_U10 ( .A1(maj_244_n21), .A2(maj_244_n20), .ZN(maj_244_n23)
         );
  XOR2_X1 maj_244_U9 ( .A(u_0_2[2]), .B(maj_244_n24), .Z(maj_244_n26) );
  XOR2_X1 maj_244_U8 ( .A(u_0_2[5]), .B(maj_244_n25), .Z(maj_244_n27) );
  XOR2_X1 maj_244_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_244_n24) );
  XOR2_X1 maj_244_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_244_n25) );
  OR2_X1 maj_244_U5 ( .A1(maj_244_n23), .A2(maj_244_n22), .ZN(maj_244_n32) );
  NAND2_X1 maj_244_U4 ( .A1(maj_244_n22), .A2(maj_244_n23), .ZN(maj_244_n34)
         );
  NAND2_X1 maj_244_U3 ( .A1(maj_244_n32), .A2(maj_244_n31), .ZN(maj_244_n33)
         );
  NAND2_X1 maj_244_U2 ( .A1(maj_244_n34), .A2(maj_244_n33), .ZN(maj_244_port_o) );
  OR2_X1 maj_245_U19 ( .A1(maj_245_n27), .A2(maj_245_n26), .ZN(maj_245_n28) );
  NAND2_X1 maj_245_U18 ( .A1(v_0_2[6]), .A2(maj_245_n28), .ZN(maj_245_n29) );
  NAND2_X1 maj_245_U17 ( .A1(maj_245_n26), .A2(maj_245_n27), .ZN(maj_245_n30)
         );
  NAND2_X1 maj_245_U16 ( .A1(maj_245_n30), .A2(maj_245_n29), .ZN(maj_245_n31)
         );
  NAND2_X1 maj_245_U15 ( .A1(v_0_2[5]), .A2(maj_245_n25), .ZN(maj_245_n18) );
  NAND2_X1 maj_245_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_245_n19) );
  NAND2_X1 maj_245_U13 ( .A1(maj_245_n19), .A2(maj_245_n18), .ZN(maj_245_n22)
         );
  NAND2_X1 maj_245_U12 ( .A1(v_0_2[2]), .A2(maj_245_n24), .ZN(maj_245_n20) );
  NAND2_X1 maj_245_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_245_n21) );
  NAND2_X1 maj_245_U10 ( .A1(maj_245_n21), .A2(maj_245_n20), .ZN(maj_245_n23)
         );
  XOR2_X1 maj_245_U9 ( .A(v_0_2[2]), .B(maj_245_n24), .Z(maj_245_n26) );
  XOR2_X1 maj_245_U8 ( .A(v_0_2[5]), .B(maj_245_n25), .Z(maj_245_n27) );
  XOR2_X1 maj_245_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_245_n24) );
  XOR2_X1 maj_245_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_245_n25) );
  OR2_X1 maj_245_U5 ( .A1(maj_245_n23), .A2(maj_245_n22), .ZN(maj_245_n32) );
  NAND2_X1 maj_245_U4 ( .A1(maj_245_n22), .A2(maj_245_n23), .ZN(maj_245_n34)
         );
  NAND2_X1 maj_245_U3 ( .A1(maj_245_n32), .A2(maj_245_n31), .ZN(maj_245_n33)
         );
  NAND2_X1 maj_245_U2 ( .A1(maj_245_n34), .A2(maj_245_n33), .ZN(maj_245_port_o) );
  OR2_X1 maj_246_U19 ( .A1(maj_246_n27), .A2(maj_246_n26), .ZN(maj_246_n28) );
  NAND2_X1 maj_246_U18 ( .A1(u_1_0[6]), .A2(maj_246_n28), .ZN(maj_246_n29) );
  NAND2_X1 maj_246_U17 ( .A1(maj_246_n26), .A2(maj_246_n27), .ZN(maj_246_n30)
         );
  NAND2_X1 maj_246_U16 ( .A1(maj_246_n30), .A2(maj_246_n29), .ZN(maj_246_n31)
         );
  NAND2_X1 maj_246_U15 ( .A1(u_1_0[5]), .A2(maj_246_n25), .ZN(maj_246_n18) );
  NAND2_X1 maj_246_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_246_n19) );
  NAND2_X1 maj_246_U13 ( .A1(maj_246_n19), .A2(maj_246_n18), .ZN(maj_246_n22)
         );
  NAND2_X1 maj_246_U12 ( .A1(u_1_0[2]), .A2(maj_246_n24), .ZN(maj_246_n20) );
  NAND2_X1 maj_246_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_246_n21) );
  NAND2_X1 maj_246_U10 ( .A1(maj_246_n21), .A2(maj_246_n20), .ZN(maj_246_n23)
         );
  XOR2_X1 maj_246_U9 ( .A(u_1_0[2]), .B(maj_246_n24), .Z(maj_246_n26) );
  XOR2_X1 maj_246_U8 ( .A(u_1_0[5]), .B(maj_246_n25), .Z(maj_246_n27) );
  XOR2_X1 maj_246_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_246_n24) );
  XOR2_X1 maj_246_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_246_n25) );
  OR2_X1 maj_246_U5 ( .A1(maj_246_n23), .A2(maj_246_n22), .ZN(maj_246_n32) );
  NAND2_X1 maj_246_U4 ( .A1(maj_246_n22), .A2(maj_246_n23), .ZN(maj_246_n34)
         );
  NAND2_X1 maj_246_U3 ( .A1(maj_246_n32), .A2(maj_246_n31), .ZN(maj_246_n33)
         );
  NAND2_X1 maj_246_U2 ( .A1(maj_246_n34), .A2(maj_246_n33), .ZN(maj_246_port_o) );
  OR2_X1 maj_247_U19 ( .A1(maj_247_n27), .A2(maj_247_n26), .ZN(maj_247_n28) );
  NAND2_X1 maj_247_U18 ( .A1(v_1_0[6]), .A2(maj_247_n28), .ZN(maj_247_n29) );
  NAND2_X1 maj_247_U17 ( .A1(maj_247_n26), .A2(maj_247_n27), .ZN(maj_247_n30)
         );
  NAND2_X1 maj_247_U16 ( .A1(maj_247_n30), .A2(maj_247_n29), .ZN(maj_247_n31)
         );
  NAND2_X1 maj_247_U15 ( .A1(v_1_0[5]), .A2(maj_247_n25), .ZN(maj_247_n18) );
  NAND2_X1 maj_247_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_247_n19) );
  NAND2_X1 maj_247_U13 ( .A1(maj_247_n19), .A2(maj_247_n18), .ZN(maj_247_n22)
         );
  NAND2_X1 maj_247_U12 ( .A1(v_1_0[2]), .A2(maj_247_n24), .ZN(maj_247_n20) );
  NAND2_X1 maj_247_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_247_n21) );
  NAND2_X1 maj_247_U10 ( .A1(maj_247_n21), .A2(maj_247_n20), .ZN(maj_247_n23)
         );
  XOR2_X1 maj_247_U9 ( .A(v_1_0[2]), .B(maj_247_n24), .Z(maj_247_n26) );
  XOR2_X1 maj_247_U8 ( .A(v_1_0[5]), .B(maj_247_n25), .Z(maj_247_n27) );
  XOR2_X1 maj_247_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_247_n24) );
  XOR2_X1 maj_247_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_247_n25) );
  OR2_X1 maj_247_U5 ( .A1(maj_247_n23), .A2(maj_247_n22), .ZN(maj_247_n32) );
  NAND2_X1 maj_247_U4 ( .A1(maj_247_n22), .A2(maj_247_n23), .ZN(maj_247_n34)
         );
  NAND2_X1 maj_247_U3 ( .A1(maj_247_n32), .A2(maj_247_n31), .ZN(maj_247_n33)
         );
  NAND2_X1 maj_247_U2 ( .A1(maj_247_n34), .A2(maj_247_n33), .ZN(maj_247_port_o) );
  OR2_X1 maj_248_U19 ( .A1(maj_248_n27), .A2(maj_248_n26), .ZN(maj_248_n28) );
  NAND2_X1 maj_248_U18 ( .A1(u_1_1[6]), .A2(maj_248_n28), .ZN(maj_248_n29) );
  NAND2_X1 maj_248_U17 ( .A1(maj_248_n26), .A2(maj_248_n27), .ZN(maj_248_n30)
         );
  NAND2_X1 maj_248_U16 ( .A1(maj_248_n30), .A2(maj_248_n29), .ZN(maj_248_n31)
         );
  NAND2_X1 maj_248_U15 ( .A1(u_1_1[5]), .A2(maj_248_n25), .ZN(maj_248_n18) );
  NAND2_X1 maj_248_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_248_n19) );
  NAND2_X1 maj_248_U13 ( .A1(maj_248_n19), .A2(maj_248_n18), .ZN(maj_248_n22)
         );
  NAND2_X1 maj_248_U12 ( .A1(u_1_1[2]), .A2(maj_248_n24), .ZN(maj_248_n20) );
  NAND2_X1 maj_248_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_248_n21) );
  NAND2_X1 maj_248_U10 ( .A1(maj_248_n21), .A2(maj_248_n20), .ZN(maj_248_n23)
         );
  XOR2_X1 maj_248_U9 ( .A(u_1_1[2]), .B(maj_248_n24), .Z(maj_248_n26) );
  XOR2_X1 maj_248_U8 ( .A(u_1_1[5]), .B(maj_248_n25), .Z(maj_248_n27) );
  XOR2_X1 maj_248_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_248_n24) );
  XOR2_X1 maj_248_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_248_n25) );
  OR2_X1 maj_248_U5 ( .A1(maj_248_n23), .A2(maj_248_n22), .ZN(maj_248_n32) );
  NAND2_X1 maj_248_U4 ( .A1(maj_248_n22), .A2(maj_248_n23), .ZN(maj_248_n34)
         );
  NAND2_X1 maj_248_U3 ( .A1(maj_248_n32), .A2(maj_248_n31), .ZN(maj_248_n33)
         );
  NAND2_X1 maj_248_U2 ( .A1(maj_248_n34), .A2(maj_248_n33), .ZN(maj_248_port_o) );
  OR2_X1 maj_249_U19 ( .A1(maj_249_n27), .A2(maj_249_n26), .ZN(maj_249_n28) );
  NAND2_X1 maj_249_U18 ( .A1(v_1_1[6]), .A2(maj_249_n28), .ZN(maj_249_n29) );
  NAND2_X1 maj_249_U17 ( .A1(maj_249_n26), .A2(maj_249_n27), .ZN(maj_249_n30)
         );
  NAND2_X1 maj_249_U16 ( .A1(maj_249_n30), .A2(maj_249_n29), .ZN(maj_249_n31)
         );
  NAND2_X1 maj_249_U15 ( .A1(v_1_1[5]), .A2(maj_249_n25), .ZN(maj_249_n18) );
  NAND2_X1 maj_249_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_249_n19) );
  NAND2_X1 maj_249_U13 ( .A1(maj_249_n19), .A2(maj_249_n18), .ZN(maj_249_n22)
         );
  NAND2_X1 maj_249_U12 ( .A1(v_1_1[2]), .A2(maj_249_n24), .ZN(maj_249_n20) );
  NAND2_X1 maj_249_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_249_n21) );
  NAND2_X1 maj_249_U10 ( .A1(maj_249_n21), .A2(maj_249_n20), .ZN(maj_249_n23)
         );
  XOR2_X1 maj_249_U9 ( .A(v_1_1[2]), .B(maj_249_n24), .Z(maj_249_n26) );
  XOR2_X1 maj_249_U8 ( .A(v_1_1[5]), .B(maj_249_n25), .Z(maj_249_n27) );
  XOR2_X1 maj_249_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_249_n24) );
  XOR2_X1 maj_249_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_249_n25) );
  OR2_X1 maj_249_U5 ( .A1(maj_249_n23), .A2(maj_249_n22), .ZN(maj_249_n32) );
  NAND2_X1 maj_249_U4 ( .A1(maj_249_n22), .A2(maj_249_n23), .ZN(maj_249_n34)
         );
  NAND2_X1 maj_249_U3 ( .A1(maj_249_n32), .A2(maj_249_n31), .ZN(maj_249_n33)
         );
  NAND2_X1 maj_249_U2 ( .A1(maj_249_n34), .A2(maj_249_n33), .ZN(maj_249_port_o) );
  OR2_X1 maj_250_U19 ( .A1(maj_250_n27), .A2(maj_250_n26), .ZN(maj_250_n28) );
  NAND2_X1 maj_250_U18 ( .A1(u_1_2[6]), .A2(maj_250_n28), .ZN(maj_250_n29) );
  NAND2_X1 maj_250_U17 ( .A1(maj_250_n26), .A2(maj_250_n27), .ZN(maj_250_n30)
         );
  NAND2_X1 maj_250_U16 ( .A1(maj_250_n30), .A2(maj_250_n29), .ZN(maj_250_n31)
         );
  NAND2_X1 maj_250_U15 ( .A1(u_1_2[5]), .A2(maj_250_n25), .ZN(maj_250_n18) );
  NAND2_X1 maj_250_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_250_n19) );
  NAND2_X1 maj_250_U13 ( .A1(maj_250_n19), .A2(maj_250_n18), .ZN(maj_250_n22)
         );
  NAND2_X1 maj_250_U12 ( .A1(u_1_2[2]), .A2(maj_250_n24), .ZN(maj_250_n20) );
  NAND2_X1 maj_250_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_250_n21) );
  NAND2_X1 maj_250_U10 ( .A1(maj_250_n21), .A2(maj_250_n20), .ZN(maj_250_n23)
         );
  XOR2_X1 maj_250_U9 ( .A(u_1_2[2]), .B(maj_250_n24), .Z(maj_250_n26) );
  XOR2_X1 maj_250_U8 ( .A(u_1_2[5]), .B(maj_250_n25), .Z(maj_250_n27) );
  XOR2_X1 maj_250_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_250_n24) );
  XOR2_X1 maj_250_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_250_n25) );
  OR2_X1 maj_250_U5 ( .A1(maj_250_n23), .A2(maj_250_n22), .ZN(maj_250_n32) );
  NAND2_X1 maj_250_U4 ( .A1(maj_250_n22), .A2(maj_250_n23), .ZN(maj_250_n34)
         );
  NAND2_X1 maj_250_U3 ( .A1(maj_250_n32), .A2(maj_250_n31), .ZN(maj_250_n33)
         );
  NAND2_X1 maj_250_U2 ( .A1(maj_250_n34), .A2(maj_250_n33), .ZN(maj_250_port_o) );
  OR2_X1 maj_251_U19 ( .A1(maj_251_n27), .A2(maj_251_n26), .ZN(maj_251_n28) );
  NAND2_X1 maj_251_U18 ( .A1(v_1_2[6]), .A2(maj_251_n28), .ZN(maj_251_n29) );
  NAND2_X1 maj_251_U17 ( .A1(maj_251_n26), .A2(maj_251_n27), .ZN(maj_251_n30)
         );
  NAND2_X1 maj_251_U16 ( .A1(maj_251_n30), .A2(maj_251_n29), .ZN(maj_251_n31)
         );
  NAND2_X1 maj_251_U15 ( .A1(v_1_2[5]), .A2(maj_251_n25), .ZN(maj_251_n18) );
  NAND2_X1 maj_251_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_251_n19) );
  NAND2_X1 maj_251_U13 ( .A1(maj_251_n19), .A2(maj_251_n18), .ZN(maj_251_n22)
         );
  NAND2_X1 maj_251_U12 ( .A1(v_1_2[2]), .A2(maj_251_n24), .ZN(maj_251_n20) );
  NAND2_X1 maj_251_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_251_n21) );
  NAND2_X1 maj_251_U10 ( .A1(maj_251_n21), .A2(maj_251_n20), .ZN(maj_251_n23)
         );
  XOR2_X1 maj_251_U9 ( .A(v_1_2[2]), .B(maj_251_n24), .Z(maj_251_n26) );
  XOR2_X1 maj_251_U8 ( .A(v_1_2[5]), .B(maj_251_n25), .Z(maj_251_n27) );
  XOR2_X1 maj_251_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_251_n24) );
  XOR2_X1 maj_251_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_251_n25) );
  OR2_X1 maj_251_U5 ( .A1(maj_251_n23), .A2(maj_251_n22), .ZN(maj_251_n32) );
  NAND2_X1 maj_251_U4 ( .A1(maj_251_n22), .A2(maj_251_n23), .ZN(maj_251_n34)
         );
  NAND2_X1 maj_251_U3 ( .A1(maj_251_n32), .A2(maj_251_n31), .ZN(maj_251_n33)
         );
  NAND2_X1 maj_251_U2 ( .A1(maj_251_n34), .A2(maj_251_n33), .ZN(maj_251_port_o) );
  OR2_X1 maj_252_U19 ( .A1(maj_252_n27), .A2(maj_252_n26), .ZN(maj_252_n28) );
  NAND2_X1 maj_252_U18 ( .A1(u_2_0[6]), .A2(maj_252_n28), .ZN(maj_252_n29) );
  NAND2_X1 maj_252_U17 ( .A1(maj_252_n26), .A2(maj_252_n27), .ZN(maj_252_n30)
         );
  NAND2_X1 maj_252_U16 ( .A1(maj_252_n30), .A2(maj_252_n29), .ZN(maj_252_n31)
         );
  NAND2_X1 maj_252_U15 ( .A1(u_2_0[5]), .A2(maj_252_n25), .ZN(maj_252_n18) );
  NAND2_X1 maj_252_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_252_n19) );
  NAND2_X1 maj_252_U13 ( .A1(maj_252_n19), .A2(maj_252_n18), .ZN(maj_252_n22)
         );
  NAND2_X1 maj_252_U12 ( .A1(u_2_0[2]), .A2(maj_252_n24), .ZN(maj_252_n20) );
  NAND2_X1 maj_252_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_252_n21) );
  NAND2_X1 maj_252_U10 ( .A1(maj_252_n21), .A2(maj_252_n20), .ZN(maj_252_n23)
         );
  XOR2_X1 maj_252_U9 ( .A(u_2_0[2]), .B(maj_252_n24), .Z(maj_252_n26) );
  XOR2_X1 maj_252_U8 ( .A(u_2_0[5]), .B(maj_252_n25), .Z(maj_252_n27) );
  XOR2_X1 maj_252_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_252_n24) );
  XOR2_X1 maj_252_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_252_n25) );
  OR2_X1 maj_252_U5 ( .A1(maj_252_n23), .A2(maj_252_n22), .ZN(maj_252_n32) );
  NAND2_X1 maj_252_U4 ( .A1(maj_252_n22), .A2(maj_252_n23), .ZN(maj_252_n34)
         );
  NAND2_X1 maj_252_U3 ( .A1(maj_252_n32), .A2(maj_252_n31), .ZN(maj_252_n33)
         );
  NAND2_X1 maj_252_U2 ( .A1(maj_252_n34), .A2(maj_252_n33), .ZN(maj_252_port_o) );
  OR2_X1 maj_253_U19 ( .A1(maj_253_n27), .A2(maj_253_n26), .ZN(maj_253_n28) );
  NAND2_X1 maj_253_U18 ( .A1(v_2_0[6]), .A2(maj_253_n28), .ZN(maj_253_n29) );
  NAND2_X1 maj_253_U17 ( .A1(maj_253_n26), .A2(maj_253_n27), .ZN(maj_253_n30)
         );
  NAND2_X1 maj_253_U16 ( .A1(maj_253_n30), .A2(maj_253_n29), .ZN(maj_253_n31)
         );
  NAND2_X1 maj_253_U15 ( .A1(v_2_0[5]), .A2(maj_253_n25), .ZN(maj_253_n18) );
  NAND2_X1 maj_253_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_253_n19) );
  NAND2_X1 maj_253_U13 ( .A1(maj_253_n19), .A2(maj_253_n18), .ZN(maj_253_n22)
         );
  NAND2_X1 maj_253_U12 ( .A1(v_2_0[2]), .A2(maj_253_n24), .ZN(maj_253_n20) );
  NAND2_X1 maj_253_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_253_n21) );
  NAND2_X1 maj_253_U10 ( .A1(maj_253_n21), .A2(maj_253_n20), .ZN(maj_253_n23)
         );
  XOR2_X1 maj_253_U9 ( .A(v_2_0[2]), .B(maj_253_n24), .Z(maj_253_n26) );
  XOR2_X1 maj_253_U8 ( .A(v_2_0[5]), .B(maj_253_n25), .Z(maj_253_n27) );
  XOR2_X1 maj_253_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_253_n24) );
  XOR2_X1 maj_253_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_253_n25) );
  OR2_X1 maj_253_U5 ( .A1(maj_253_n23), .A2(maj_253_n22), .ZN(maj_253_n32) );
  NAND2_X1 maj_253_U4 ( .A1(maj_253_n22), .A2(maj_253_n23), .ZN(maj_253_n34)
         );
  NAND2_X1 maj_253_U3 ( .A1(maj_253_n32), .A2(maj_253_n31), .ZN(maj_253_n33)
         );
  NAND2_X1 maj_253_U2 ( .A1(maj_253_n34), .A2(maj_253_n33), .ZN(maj_253_port_o) );
  OR2_X1 maj_254_U19 ( .A1(maj_254_n27), .A2(maj_254_n26), .ZN(maj_254_n28) );
  NAND2_X1 maj_254_U18 ( .A1(u_2_1[6]), .A2(maj_254_n28), .ZN(maj_254_n29) );
  NAND2_X1 maj_254_U17 ( .A1(maj_254_n26), .A2(maj_254_n27), .ZN(maj_254_n30)
         );
  NAND2_X1 maj_254_U16 ( .A1(maj_254_n30), .A2(maj_254_n29), .ZN(maj_254_n31)
         );
  NAND2_X1 maj_254_U15 ( .A1(u_2_1[5]), .A2(maj_254_n25), .ZN(maj_254_n18) );
  NAND2_X1 maj_254_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_254_n19) );
  NAND2_X1 maj_254_U13 ( .A1(maj_254_n19), .A2(maj_254_n18), .ZN(maj_254_n22)
         );
  NAND2_X1 maj_254_U12 ( .A1(u_2_1[2]), .A2(maj_254_n24), .ZN(maj_254_n20) );
  NAND2_X1 maj_254_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_254_n21) );
  NAND2_X1 maj_254_U10 ( .A1(maj_254_n21), .A2(maj_254_n20), .ZN(maj_254_n23)
         );
  XOR2_X1 maj_254_U9 ( .A(u_2_1[2]), .B(maj_254_n24), .Z(maj_254_n26) );
  XOR2_X1 maj_254_U8 ( .A(u_2_1[5]), .B(maj_254_n25), .Z(maj_254_n27) );
  XOR2_X1 maj_254_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_254_n24) );
  XOR2_X1 maj_254_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_254_n25) );
  OR2_X1 maj_254_U5 ( .A1(maj_254_n23), .A2(maj_254_n22), .ZN(maj_254_n32) );
  NAND2_X1 maj_254_U4 ( .A1(maj_254_n22), .A2(maj_254_n23), .ZN(maj_254_n34)
         );
  NAND2_X1 maj_254_U3 ( .A1(maj_254_n32), .A2(maj_254_n31), .ZN(maj_254_n33)
         );
  NAND2_X1 maj_254_U2 ( .A1(maj_254_n34), .A2(maj_254_n33), .ZN(maj_254_port_o) );
  OR2_X1 maj_255_U19 ( .A1(maj_255_n27), .A2(maj_255_n26), .ZN(maj_255_n28) );
  NAND2_X1 maj_255_U18 ( .A1(v_2_1[6]), .A2(maj_255_n28), .ZN(maj_255_n29) );
  NAND2_X1 maj_255_U17 ( .A1(maj_255_n26), .A2(maj_255_n27), .ZN(maj_255_n30)
         );
  NAND2_X1 maj_255_U16 ( .A1(maj_255_n30), .A2(maj_255_n29), .ZN(maj_255_n31)
         );
  NAND2_X1 maj_255_U15 ( .A1(v_2_1[5]), .A2(maj_255_n25), .ZN(maj_255_n18) );
  NAND2_X1 maj_255_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_255_n19) );
  NAND2_X1 maj_255_U13 ( .A1(maj_255_n19), .A2(maj_255_n18), .ZN(maj_255_n22)
         );
  NAND2_X1 maj_255_U12 ( .A1(v_2_1[2]), .A2(maj_255_n24), .ZN(maj_255_n20) );
  NAND2_X1 maj_255_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_255_n21) );
  NAND2_X1 maj_255_U10 ( .A1(maj_255_n21), .A2(maj_255_n20), .ZN(maj_255_n23)
         );
  XOR2_X1 maj_255_U9 ( .A(v_2_1[2]), .B(maj_255_n24), .Z(maj_255_n26) );
  XOR2_X1 maj_255_U8 ( .A(v_2_1[5]), .B(maj_255_n25), .Z(maj_255_n27) );
  XOR2_X1 maj_255_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_255_n24) );
  XOR2_X1 maj_255_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_255_n25) );
  OR2_X1 maj_255_U5 ( .A1(maj_255_n23), .A2(maj_255_n22), .ZN(maj_255_n32) );
  NAND2_X1 maj_255_U4 ( .A1(maj_255_n22), .A2(maj_255_n23), .ZN(maj_255_n34)
         );
  NAND2_X1 maj_255_U3 ( .A1(maj_255_n32), .A2(maj_255_n31), .ZN(maj_255_n33)
         );
  NAND2_X1 maj_255_U2 ( .A1(maj_255_n34), .A2(maj_255_n33), .ZN(maj_255_port_o) );
  OR2_X1 maj_256_U19 ( .A1(maj_256_n27), .A2(maj_256_n26), .ZN(maj_256_n28) );
  NAND2_X1 maj_256_U18 ( .A1(u_2_2[6]), .A2(maj_256_n28), .ZN(maj_256_n29) );
  NAND2_X1 maj_256_U17 ( .A1(maj_256_n26), .A2(maj_256_n27), .ZN(maj_256_n30)
         );
  NAND2_X1 maj_256_U16 ( .A1(maj_256_n30), .A2(maj_256_n29), .ZN(maj_256_n31)
         );
  NAND2_X1 maj_256_U15 ( .A1(u_2_2[5]), .A2(maj_256_n25), .ZN(maj_256_n18) );
  NAND2_X1 maj_256_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_256_n19) );
  NAND2_X1 maj_256_U13 ( .A1(maj_256_n19), .A2(maj_256_n18), .ZN(maj_256_n22)
         );
  NAND2_X1 maj_256_U12 ( .A1(u_2_2[2]), .A2(maj_256_n24), .ZN(maj_256_n20) );
  NAND2_X1 maj_256_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_256_n21) );
  NAND2_X1 maj_256_U10 ( .A1(maj_256_n21), .A2(maj_256_n20), .ZN(maj_256_n23)
         );
  XOR2_X1 maj_256_U9 ( .A(u_2_2[2]), .B(maj_256_n24), .Z(maj_256_n26) );
  XOR2_X1 maj_256_U8 ( .A(u_2_2[5]), .B(maj_256_n25), .Z(maj_256_n27) );
  XOR2_X1 maj_256_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_256_n24) );
  XOR2_X1 maj_256_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_256_n25) );
  OR2_X1 maj_256_U5 ( .A1(maj_256_n23), .A2(maj_256_n22), .ZN(maj_256_n32) );
  NAND2_X1 maj_256_U4 ( .A1(maj_256_n22), .A2(maj_256_n23), .ZN(maj_256_n34)
         );
  NAND2_X1 maj_256_U3 ( .A1(maj_256_n32), .A2(maj_256_n31), .ZN(maj_256_n33)
         );
  NAND2_X1 maj_256_U2 ( .A1(maj_256_n34), .A2(maj_256_n33), .ZN(maj_256_port_o) );
  OR2_X1 maj_257_U19 ( .A1(maj_257_n27), .A2(maj_257_n26), .ZN(maj_257_n28) );
  NAND2_X1 maj_257_U18 ( .A1(v_2_2[6]), .A2(maj_257_n28), .ZN(maj_257_n29) );
  NAND2_X1 maj_257_U17 ( .A1(maj_257_n26), .A2(maj_257_n27), .ZN(maj_257_n30)
         );
  NAND2_X1 maj_257_U16 ( .A1(maj_257_n30), .A2(maj_257_n29), .ZN(maj_257_n31)
         );
  NAND2_X1 maj_257_U15 ( .A1(v_2_2[5]), .A2(maj_257_n25), .ZN(maj_257_n18) );
  NAND2_X1 maj_257_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_257_n19) );
  NAND2_X1 maj_257_U13 ( .A1(maj_257_n19), .A2(maj_257_n18), .ZN(maj_257_n22)
         );
  NAND2_X1 maj_257_U12 ( .A1(v_2_2[2]), .A2(maj_257_n24), .ZN(maj_257_n20) );
  NAND2_X1 maj_257_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_257_n21) );
  NAND2_X1 maj_257_U10 ( .A1(maj_257_n21), .A2(maj_257_n20), .ZN(maj_257_n23)
         );
  XOR2_X1 maj_257_U9 ( .A(v_2_2[2]), .B(maj_257_n24), .Z(maj_257_n26) );
  XOR2_X1 maj_257_U8 ( .A(v_2_2[5]), .B(maj_257_n25), .Z(maj_257_n27) );
  XOR2_X1 maj_257_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_257_n24) );
  XOR2_X1 maj_257_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_257_n25) );
  OR2_X1 maj_257_U5 ( .A1(maj_257_n23), .A2(maj_257_n22), .ZN(maj_257_n32) );
  NAND2_X1 maj_257_U4 ( .A1(maj_257_n22), .A2(maj_257_n23), .ZN(maj_257_n34)
         );
  NAND2_X1 maj_257_U3 ( .A1(maj_257_n32), .A2(maj_257_n31), .ZN(maj_257_n33)
         );
  NAND2_X1 maj_257_U2 ( .A1(maj_257_n34), .A2(maj_257_n33), .ZN(maj_257_port_o) );
  OR2_X1 maj_258_U19 ( .A1(maj_258_n27), .A2(maj_258_n26), .ZN(maj_258_n28) );
  NAND2_X1 maj_258_U18 ( .A1(u_3_0[6]), .A2(maj_258_n28), .ZN(maj_258_n29) );
  NAND2_X1 maj_258_U17 ( .A1(maj_258_n26), .A2(maj_258_n27), .ZN(maj_258_n30)
         );
  NAND2_X1 maj_258_U16 ( .A1(maj_258_n30), .A2(maj_258_n29), .ZN(maj_258_n31)
         );
  NAND2_X1 maj_258_U15 ( .A1(u_3_0[5]), .A2(maj_258_n25), .ZN(maj_258_n18) );
  NAND2_X1 maj_258_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_258_n19) );
  NAND2_X1 maj_258_U13 ( .A1(maj_258_n19), .A2(maj_258_n18), .ZN(maj_258_n22)
         );
  NAND2_X1 maj_258_U12 ( .A1(u_3_0[2]), .A2(maj_258_n24), .ZN(maj_258_n20) );
  NAND2_X1 maj_258_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_258_n21) );
  NAND2_X1 maj_258_U10 ( .A1(maj_258_n21), .A2(maj_258_n20), .ZN(maj_258_n23)
         );
  XOR2_X1 maj_258_U9 ( .A(u_3_0[2]), .B(maj_258_n24), .Z(maj_258_n26) );
  XOR2_X1 maj_258_U8 ( .A(u_3_0[5]), .B(maj_258_n25), .Z(maj_258_n27) );
  XOR2_X1 maj_258_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_258_n24) );
  XOR2_X1 maj_258_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_258_n25) );
  OR2_X1 maj_258_U5 ( .A1(maj_258_n23), .A2(maj_258_n22), .ZN(maj_258_n32) );
  NAND2_X1 maj_258_U4 ( .A1(maj_258_n22), .A2(maj_258_n23), .ZN(maj_258_n34)
         );
  NAND2_X1 maj_258_U3 ( .A1(maj_258_n32), .A2(maj_258_n31), .ZN(maj_258_n33)
         );
  NAND2_X1 maj_258_U2 ( .A1(maj_258_n34), .A2(maj_258_n33), .ZN(maj_258_port_o) );
  OR2_X1 maj_259_U19 ( .A1(maj_259_n27), .A2(maj_259_n26), .ZN(maj_259_n28) );
  NAND2_X1 maj_259_U18 ( .A1(v_3_0[6]), .A2(maj_259_n28), .ZN(maj_259_n29) );
  NAND2_X1 maj_259_U17 ( .A1(maj_259_n26), .A2(maj_259_n27), .ZN(maj_259_n30)
         );
  NAND2_X1 maj_259_U16 ( .A1(maj_259_n30), .A2(maj_259_n29), .ZN(maj_259_n31)
         );
  NAND2_X1 maj_259_U15 ( .A1(v_3_0[5]), .A2(maj_259_n25), .ZN(maj_259_n18) );
  NAND2_X1 maj_259_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_259_n19) );
  NAND2_X1 maj_259_U13 ( .A1(maj_259_n19), .A2(maj_259_n18), .ZN(maj_259_n22)
         );
  NAND2_X1 maj_259_U12 ( .A1(v_3_0[2]), .A2(maj_259_n24), .ZN(maj_259_n20) );
  NAND2_X1 maj_259_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_259_n21) );
  NAND2_X1 maj_259_U10 ( .A1(maj_259_n21), .A2(maj_259_n20), .ZN(maj_259_n23)
         );
  XOR2_X1 maj_259_U9 ( .A(v_3_0[2]), .B(maj_259_n24), .Z(maj_259_n26) );
  XOR2_X1 maj_259_U8 ( .A(v_3_0[5]), .B(maj_259_n25), .Z(maj_259_n27) );
  XOR2_X1 maj_259_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_259_n24) );
  XOR2_X1 maj_259_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_259_n25) );
  OR2_X1 maj_259_U5 ( .A1(maj_259_n23), .A2(maj_259_n22), .ZN(maj_259_n32) );
  NAND2_X1 maj_259_U4 ( .A1(maj_259_n22), .A2(maj_259_n23), .ZN(maj_259_n34)
         );
  NAND2_X1 maj_259_U3 ( .A1(maj_259_n32), .A2(maj_259_n31), .ZN(maj_259_n33)
         );
  NAND2_X1 maj_259_U2 ( .A1(maj_259_n34), .A2(maj_259_n33), .ZN(maj_259_port_o) );
  OR2_X1 maj_260_U19 ( .A1(maj_260_n27), .A2(maj_260_n26), .ZN(maj_260_n28) );
  NAND2_X1 maj_260_U18 ( .A1(u_3_1[6]), .A2(maj_260_n28), .ZN(maj_260_n29) );
  NAND2_X1 maj_260_U17 ( .A1(maj_260_n26), .A2(maj_260_n27), .ZN(maj_260_n30)
         );
  NAND2_X1 maj_260_U16 ( .A1(maj_260_n30), .A2(maj_260_n29), .ZN(maj_260_n31)
         );
  NAND2_X1 maj_260_U15 ( .A1(u_3_1[5]), .A2(maj_260_n25), .ZN(maj_260_n18) );
  NAND2_X1 maj_260_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_260_n19) );
  NAND2_X1 maj_260_U13 ( .A1(maj_260_n19), .A2(maj_260_n18), .ZN(maj_260_n22)
         );
  NAND2_X1 maj_260_U12 ( .A1(u_3_1[2]), .A2(maj_260_n24), .ZN(maj_260_n20) );
  NAND2_X1 maj_260_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_260_n21) );
  NAND2_X1 maj_260_U10 ( .A1(maj_260_n21), .A2(maj_260_n20), .ZN(maj_260_n23)
         );
  XOR2_X1 maj_260_U9 ( .A(u_3_1[2]), .B(maj_260_n24), .Z(maj_260_n26) );
  XOR2_X1 maj_260_U8 ( .A(u_3_1[5]), .B(maj_260_n25), .Z(maj_260_n27) );
  XOR2_X1 maj_260_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_260_n24) );
  XOR2_X1 maj_260_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_260_n25) );
  OR2_X1 maj_260_U5 ( .A1(maj_260_n23), .A2(maj_260_n22), .ZN(maj_260_n32) );
  NAND2_X1 maj_260_U4 ( .A1(maj_260_n22), .A2(maj_260_n23), .ZN(maj_260_n34)
         );
  NAND2_X1 maj_260_U3 ( .A1(maj_260_n32), .A2(maj_260_n31), .ZN(maj_260_n33)
         );
  NAND2_X1 maj_260_U2 ( .A1(maj_260_n34), .A2(maj_260_n33), .ZN(maj_260_port_o) );
  OR2_X1 maj_261_U19 ( .A1(maj_261_n27), .A2(maj_261_n26), .ZN(maj_261_n28) );
  NAND2_X1 maj_261_U18 ( .A1(v_3_1[6]), .A2(maj_261_n28), .ZN(maj_261_n29) );
  NAND2_X1 maj_261_U17 ( .A1(maj_261_n26), .A2(maj_261_n27), .ZN(maj_261_n30)
         );
  NAND2_X1 maj_261_U16 ( .A1(maj_261_n30), .A2(maj_261_n29), .ZN(maj_261_n31)
         );
  NAND2_X1 maj_261_U15 ( .A1(v_3_1[5]), .A2(maj_261_n25), .ZN(maj_261_n18) );
  NAND2_X1 maj_261_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_261_n19) );
  NAND2_X1 maj_261_U13 ( .A1(maj_261_n19), .A2(maj_261_n18), .ZN(maj_261_n22)
         );
  NAND2_X1 maj_261_U12 ( .A1(v_3_1[2]), .A2(maj_261_n24), .ZN(maj_261_n20) );
  NAND2_X1 maj_261_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_261_n21) );
  NAND2_X1 maj_261_U10 ( .A1(maj_261_n21), .A2(maj_261_n20), .ZN(maj_261_n23)
         );
  XOR2_X1 maj_261_U9 ( .A(v_3_1[2]), .B(maj_261_n24), .Z(maj_261_n26) );
  XOR2_X1 maj_261_U8 ( .A(v_3_1[5]), .B(maj_261_n25), .Z(maj_261_n27) );
  XOR2_X1 maj_261_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_261_n24) );
  XOR2_X1 maj_261_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_261_n25) );
  OR2_X1 maj_261_U5 ( .A1(maj_261_n23), .A2(maj_261_n22), .ZN(maj_261_n32) );
  NAND2_X1 maj_261_U4 ( .A1(maj_261_n22), .A2(maj_261_n23), .ZN(maj_261_n34)
         );
  NAND2_X1 maj_261_U3 ( .A1(maj_261_n32), .A2(maj_261_n31), .ZN(maj_261_n33)
         );
  NAND2_X1 maj_261_U2 ( .A1(maj_261_n34), .A2(maj_261_n33), .ZN(maj_261_port_o) );
  OR2_X1 maj_262_U19 ( .A1(maj_262_n27), .A2(maj_262_n26), .ZN(maj_262_n28) );
  NAND2_X1 maj_262_U18 ( .A1(u_3_2[6]), .A2(maj_262_n28), .ZN(maj_262_n29) );
  NAND2_X1 maj_262_U17 ( .A1(maj_262_n26), .A2(maj_262_n27), .ZN(maj_262_n30)
         );
  NAND2_X1 maj_262_U16 ( .A1(maj_262_n30), .A2(maj_262_n29), .ZN(maj_262_n31)
         );
  NAND2_X1 maj_262_U15 ( .A1(u_3_2[5]), .A2(maj_262_n25), .ZN(maj_262_n18) );
  NAND2_X1 maj_262_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_262_n19) );
  NAND2_X1 maj_262_U13 ( .A1(maj_262_n19), .A2(maj_262_n18), .ZN(maj_262_n22)
         );
  NAND2_X1 maj_262_U12 ( .A1(u_3_2[2]), .A2(maj_262_n24), .ZN(maj_262_n20) );
  NAND2_X1 maj_262_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_262_n21) );
  NAND2_X1 maj_262_U10 ( .A1(maj_262_n21), .A2(maj_262_n20), .ZN(maj_262_n23)
         );
  XOR2_X1 maj_262_U9 ( .A(u_3_2[2]), .B(maj_262_n24), .Z(maj_262_n26) );
  XOR2_X1 maj_262_U8 ( .A(u_3_2[5]), .B(maj_262_n25), .Z(maj_262_n27) );
  XOR2_X1 maj_262_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_262_n24) );
  XOR2_X1 maj_262_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_262_n25) );
  OR2_X1 maj_262_U5 ( .A1(maj_262_n23), .A2(maj_262_n22), .ZN(maj_262_n32) );
  NAND2_X1 maj_262_U4 ( .A1(maj_262_n22), .A2(maj_262_n23), .ZN(maj_262_n34)
         );
  NAND2_X1 maj_262_U3 ( .A1(maj_262_n32), .A2(maj_262_n31), .ZN(maj_262_n33)
         );
  NAND2_X1 maj_262_U2 ( .A1(maj_262_n34), .A2(maj_262_n33), .ZN(maj_262_port_o) );
  OR2_X1 maj_263_U19 ( .A1(maj_263_n27), .A2(maj_263_n26), .ZN(maj_263_n28) );
  NAND2_X1 maj_263_U18 ( .A1(v_3_2[6]), .A2(maj_263_n28), .ZN(maj_263_n29) );
  NAND2_X1 maj_263_U17 ( .A1(maj_263_n26), .A2(maj_263_n27), .ZN(maj_263_n30)
         );
  NAND2_X1 maj_263_U16 ( .A1(maj_263_n30), .A2(maj_263_n29), .ZN(maj_263_n31)
         );
  NAND2_X1 maj_263_U15 ( .A1(v_3_2[5]), .A2(maj_263_n25), .ZN(maj_263_n18) );
  NAND2_X1 maj_263_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_263_n19) );
  NAND2_X1 maj_263_U13 ( .A1(maj_263_n19), .A2(maj_263_n18), .ZN(maj_263_n22)
         );
  NAND2_X1 maj_263_U12 ( .A1(v_3_2[2]), .A2(maj_263_n24), .ZN(maj_263_n20) );
  NAND2_X1 maj_263_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_263_n21) );
  NAND2_X1 maj_263_U10 ( .A1(maj_263_n21), .A2(maj_263_n20), .ZN(maj_263_n23)
         );
  XOR2_X1 maj_263_U9 ( .A(v_3_2[2]), .B(maj_263_n24), .Z(maj_263_n26) );
  XOR2_X1 maj_263_U8 ( .A(v_3_2[5]), .B(maj_263_n25), .Z(maj_263_n27) );
  XOR2_X1 maj_263_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_263_n24) );
  XOR2_X1 maj_263_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_263_n25) );
  OR2_X1 maj_263_U5 ( .A1(maj_263_n23), .A2(maj_263_n22), .ZN(maj_263_n32) );
  NAND2_X1 maj_263_U4 ( .A1(maj_263_n22), .A2(maj_263_n23), .ZN(maj_263_n34)
         );
  NAND2_X1 maj_263_U3 ( .A1(maj_263_n32), .A2(maj_263_n31), .ZN(maj_263_n33)
         );
  NAND2_X1 maj_263_U2 ( .A1(maj_263_n34), .A2(maj_263_n33), .ZN(maj_263_port_o) );
  OR2_X1 maj_264_U19 ( .A1(maj_264_n27), .A2(maj_264_n26), .ZN(maj_264_n28) );
  NAND2_X1 maj_264_U18 ( .A1(u_0_0[6]), .A2(maj_264_n28), .ZN(maj_264_n29) );
  NAND2_X1 maj_264_U17 ( .A1(maj_264_n26), .A2(maj_264_n27), .ZN(maj_264_n30)
         );
  NAND2_X1 maj_264_U16 ( .A1(maj_264_n30), .A2(maj_264_n29), .ZN(maj_264_n31)
         );
  NAND2_X1 maj_264_U15 ( .A1(u_0_0[5]), .A2(maj_264_n25), .ZN(maj_264_n18) );
  NAND2_X1 maj_264_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_264_n19) );
  NAND2_X1 maj_264_U13 ( .A1(maj_264_n19), .A2(maj_264_n18), .ZN(maj_264_n22)
         );
  NAND2_X1 maj_264_U12 ( .A1(u_0_0[2]), .A2(maj_264_n24), .ZN(maj_264_n20) );
  NAND2_X1 maj_264_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_264_n21) );
  NAND2_X1 maj_264_U10 ( .A1(maj_264_n21), .A2(maj_264_n20), .ZN(maj_264_n23)
         );
  XOR2_X1 maj_264_U9 ( .A(u_0_0[2]), .B(maj_264_n24), .Z(maj_264_n26) );
  XOR2_X1 maj_264_U8 ( .A(u_0_0[5]), .B(maj_264_n25), .Z(maj_264_n27) );
  XOR2_X1 maj_264_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_264_n24) );
  XOR2_X1 maj_264_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_264_n25) );
  OR2_X1 maj_264_U5 ( .A1(maj_264_n23), .A2(maj_264_n22), .ZN(maj_264_n32) );
  NAND2_X1 maj_264_U4 ( .A1(maj_264_n22), .A2(maj_264_n23), .ZN(maj_264_n34)
         );
  NAND2_X1 maj_264_U3 ( .A1(maj_264_n32), .A2(maj_264_n31), .ZN(maj_264_n33)
         );
  NAND2_X1 maj_264_U2 ( .A1(maj_264_n34), .A2(maj_264_n33), .ZN(maj_264_port_o) );
  OR2_X1 maj_265_U19 ( .A1(maj_265_n27), .A2(maj_265_n26), .ZN(maj_265_n28) );
  NAND2_X1 maj_265_U18 ( .A1(v_0_0[6]), .A2(maj_265_n28), .ZN(maj_265_n29) );
  NAND2_X1 maj_265_U17 ( .A1(maj_265_n26), .A2(maj_265_n27), .ZN(maj_265_n30)
         );
  NAND2_X1 maj_265_U16 ( .A1(maj_265_n30), .A2(maj_265_n29), .ZN(maj_265_n31)
         );
  NAND2_X1 maj_265_U15 ( .A1(v_0_0[5]), .A2(maj_265_n25), .ZN(maj_265_n18) );
  NAND2_X1 maj_265_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_265_n19) );
  NAND2_X1 maj_265_U13 ( .A1(maj_265_n19), .A2(maj_265_n18), .ZN(maj_265_n22)
         );
  NAND2_X1 maj_265_U12 ( .A1(v_0_0[2]), .A2(maj_265_n24), .ZN(maj_265_n20) );
  NAND2_X1 maj_265_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_265_n21) );
  NAND2_X1 maj_265_U10 ( .A1(maj_265_n21), .A2(maj_265_n20), .ZN(maj_265_n23)
         );
  XOR2_X1 maj_265_U9 ( .A(v_0_0[2]), .B(maj_265_n24), .Z(maj_265_n26) );
  XOR2_X1 maj_265_U8 ( .A(v_0_0[5]), .B(maj_265_n25), .Z(maj_265_n27) );
  XOR2_X1 maj_265_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_265_n24) );
  XOR2_X1 maj_265_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_265_n25) );
  OR2_X1 maj_265_U5 ( .A1(maj_265_n23), .A2(maj_265_n22), .ZN(maj_265_n32) );
  NAND2_X1 maj_265_U4 ( .A1(maj_265_n22), .A2(maj_265_n23), .ZN(maj_265_n34)
         );
  NAND2_X1 maj_265_U3 ( .A1(maj_265_n32), .A2(maj_265_n31), .ZN(maj_265_n33)
         );
  NAND2_X1 maj_265_U2 ( .A1(maj_265_n34), .A2(maj_265_n33), .ZN(maj_265_port_o) );
  OR2_X1 maj_266_U19 ( .A1(maj_266_n27), .A2(maj_266_n26), .ZN(maj_266_n28) );
  NAND2_X1 maj_266_U18 ( .A1(u_0_1[6]), .A2(maj_266_n28), .ZN(maj_266_n29) );
  NAND2_X1 maj_266_U17 ( .A1(maj_266_n26), .A2(maj_266_n27), .ZN(maj_266_n30)
         );
  NAND2_X1 maj_266_U16 ( .A1(maj_266_n30), .A2(maj_266_n29), .ZN(maj_266_n31)
         );
  NAND2_X1 maj_266_U15 ( .A1(u_0_1[5]), .A2(maj_266_n25), .ZN(maj_266_n18) );
  NAND2_X1 maj_266_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_266_n19) );
  NAND2_X1 maj_266_U13 ( .A1(maj_266_n19), .A2(maj_266_n18), .ZN(maj_266_n22)
         );
  NAND2_X1 maj_266_U12 ( .A1(u_0_1[2]), .A2(maj_266_n24), .ZN(maj_266_n20) );
  NAND2_X1 maj_266_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_266_n21) );
  NAND2_X1 maj_266_U10 ( .A1(maj_266_n21), .A2(maj_266_n20), .ZN(maj_266_n23)
         );
  XOR2_X1 maj_266_U9 ( .A(u_0_1[2]), .B(maj_266_n24), .Z(maj_266_n26) );
  XOR2_X1 maj_266_U8 ( .A(u_0_1[5]), .B(maj_266_n25), .Z(maj_266_n27) );
  XOR2_X1 maj_266_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_266_n24) );
  XOR2_X1 maj_266_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_266_n25) );
  OR2_X1 maj_266_U5 ( .A1(maj_266_n23), .A2(maj_266_n22), .ZN(maj_266_n32) );
  NAND2_X1 maj_266_U4 ( .A1(maj_266_n22), .A2(maj_266_n23), .ZN(maj_266_n34)
         );
  NAND2_X1 maj_266_U3 ( .A1(maj_266_n32), .A2(maj_266_n31), .ZN(maj_266_n33)
         );
  NAND2_X1 maj_266_U2 ( .A1(maj_266_n34), .A2(maj_266_n33), .ZN(maj_266_port_o) );
  OR2_X1 maj_267_U19 ( .A1(maj_267_n27), .A2(maj_267_n26), .ZN(maj_267_n28) );
  NAND2_X1 maj_267_U18 ( .A1(v_0_1[6]), .A2(maj_267_n28), .ZN(maj_267_n29) );
  NAND2_X1 maj_267_U17 ( .A1(maj_267_n26), .A2(maj_267_n27), .ZN(maj_267_n30)
         );
  NAND2_X1 maj_267_U16 ( .A1(maj_267_n30), .A2(maj_267_n29), .ZN(maj_267_n31)
         );
  NAND2_X1 maj_267_U15 ( .A1(v_0_1[5]), .A2(maj_267_n25), .ZN(maj_267_n18) );
  NAND2_X1 maj_267_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_267_n19) );
  NAND2_X1 maj_267_U13 ( .A1(maj_267_n19), .A2(maj_267_n18), .ZN(maj_267_n22)
         );
  NAND2_X1 maj_267_U12 ( .A1(v_0_1[2]), .A2(maj_267_n24), .ZN(maj_267_n20) );
  NAND2_X1 maj_267_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_267_n21) );
  NAND2_X1 maj_267_U10 ( .A1(maj_267_n21), .A2(maj_267_n20), .ZN(maj_267_n23)
         );
  XOR2_X1 maj_267_U9 ( .A(v_0_1[2]), .B(maj_267_n24), .Z(maj_267_n26) );
  XOR2_X1 maj_267_U8 ( .A(v_0_1[5]), .B(maj_267_n25), .Z(maj_267_n27) );
  XOR2_X1 maj_267_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_267_n24) );
  XOR2_X1 maj_267_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_267_n25) );
  OR2_X1 maj_267_U5 ( .A1(maj_267_n23), .A2(maj_267_n22), .ZN(maj_267_n32) );
  NAND2_X1 maj_267_U4 ( .A1(maj_267_n22), .A2(maj_267_n23), .ZN(maj_267_n34)
         );
  NAND2_X1 maj_267_U3 ( .A1(maj_267_n32), .A2(maj_267_n31), .ZN(maj_267_n33)
         );
  NAND2_X1 maj_267_U2 ( .A1(maj_267_n34), .A2(maj_267_n33), .ZN(maj_267_port_o) );
  OR2_X1 maj_268_U19 ( .A1(maj_268_n27), .A2(maj_268_n26), .ZN(maj_268_n28) );
  NAND2_X1 maj_268_U18 ( .A1(u_0_2[6]), .A2(maj_268_n28), .ZN(maj_268_n29) );
  NAND2_X1 maj_268_U17 ( .A1(maj_268_n26), .A2(maj_268_n27), .ZN(maj_268_n30)
         );
  NAND2_X1 maj_268_U16 ( .A1(maj_268_n30), .A2(maj_268_n29), .ZN(maj_268_n31)
         );
  NAND2_X1 maj_268_U15 ( .A1(u_0_2[5]), .A2(maj_268_n25), .ZN(maj_268_n18) );
  NAND2_X1 maj_268_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_268_n19) );
  NAND2_X1 maj_268_U13 ( .A1(maj_268_n19), .A2(maj_268_n18), .ZN(maj_268_n22)
         );
  NAND2_X1 maj_268_U12 ( .A1(u_0_2[2]), .A2(maj_268_n24), .ZN(maj_268_n20) );
  NAND2_X1 maj_268_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_268_n21) );
  NAND2_X1 maj_268_U10 ( .A1(maj_268_n21), .A2(maj_268_n20), .ZN(maj_268_n23)
         );
  XOR2_X1 maj_268_U9 ( .A(u_0_2[2]), .B(maj_268_n24), .Z(maj_268_n26) );
  XOR2_X1 maj_268_U8 ( .A(u_0_2[5]), .B(maj_268_n25), .Z(maj_268_n27) );
  XOR2_X1 maj_268_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_268_n24) );
  XOR2_X1 maj_268_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_268_n25) );
  OR2_X1 maj_268_U5 ( .A1(maj_268_n23), .A2(maj_268_n22), .ZN(maj_268_n32) );
  NAND2_X1 maj_268_U4 ( .A1(maj_268_n22), .A2(maj_268_n23), .ZN(maj_268_n34)
         );
  NAND2_X1 maj_268_U3 ( .A1(maj_268_n32), .A2(maj_268_n31), .ZN(maj_268_n33)
         );
  NAND2_X1 maj_268_U2 ( .A1(maj_268_n34), .A2(maj_268_n33), .ZN(maj_268_port_o) );
  OR2_X1 maj_269_U19 ( .A1(maj_269_n27), .A2(maj_269_n26), .ZN(maj_269_n28) );
  NAND2_X1 maj_269_U18 ( .A1(v_0_2[6]), .A2(maj_269_n28), .ZN(maj_269_n29) );
  NAND2_X1 maj_269_U17 ( .A1(maj_269_n26), .A2(maj_269_n27), .ZN(maj_269_n30)
         );
  NAND2_X1 maj_269_U16 ( .A1(maj_269_n30), .A2(maj_269_n29), .ZN(maj_269_n31)
         );
  NAND2_X1 maj_269_U15 ( .A1(v_0_2[5]), .A2(maj_269_n25), .ZN(maj_269_n18) );
  NAND2_X1 maj_269_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_269_n19) );
  NAND2_X1 maj_269_U13 ( .A1(maj_269_n19), .A2(maj_269_n18), .ZN(maj_269_n22)
         );
  NAND2_X1 maj_269_U12 ( .A1(v_0_2[2]), .A2(maj_269_n24), .ZN(maj_269_n20) );
  NAND2_X1 maj_269_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_269_n21) );
  NAND2_X1 maj_269_U10 ( .A1(maj_269_n21), .A2(maj_269_n20), .ZN(maj_269_n23)
         );
  XOR2_X1 maj_269_U9 ( .A(v_0_2[2]), .B(maj_269_n24), .Z(maj_269_n26) );
  XOR2_X1 maj_269_U8 ( .A(v_0_2[5]), .B(maj_269_n25), .Z(maj_269_n27) );
  XOR2_X1 maj_269_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_269_n24) );
  XOR2_X1 maj_269_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_269_n25) );
  OR2_X1 maj_269_U5 ( .A1(maj_269_n23), .A2(maj_269_n22), .ZN(maj_269_n32) );
  NAND2_X1 maj_269_U4 ( .A1(maj_269_n22), .A2(maj_269_n23), .ZN(maj_269_n34)
         );
  NAND2_X1 maj_269_U3 ( .A1(maj_269_n32), .A2(maj_269_n31), .ZN(maj_269_n33)
         );
  NAND2_X1 maj_269_U2 ( .A1(maj_269_n34), .A2(maj_269_n33), .ZN(maj_269_port_o) );
  OR2_X1 maj_270_U19 ( .A1(maj_270_n27), .A2(maj_270_n26), .ZN(maj_270_n28) );
  NAND2_X1 maj_270_U18 ( .A1(u_1_0[6]), .A2(maj_270_n28), .ZN(maj_270_n29) );
  NAND2_X1 maj_270_U17 ( .A1(maj_270_n26), .A2(maj_270_n27), .ZN(maj_270_n30)
         );
  NAND2_X1 maj_270_U16 ( .A1(maj_270_n30), .A2(maj_270_n29), .ZN(maj_270_n31)
         );
  NAND2_X1 maj_270_U15 ( .A1(u_1_0[5]), .A2(maj_270_n25), .ZN(maj_270_n18) );
  NAND2_X1 maj_270_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_270_n19) );
  NAND2_X1 maj_270_U13 ( .A1(maj_270_n19), .A2(maj_270_n18), .ZN(maj_270_n22)
         );
  NAND2_X1 maj_270_U12 ( .A1(u_1_0[2]), .A2(maj_270_n24), .ZN(maj_270_n20) );
  NAND2_X1 maj_270_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_270_n21) );
  NAND2_X1 maj_270_U10 ( .A1(maj_270_n21), .A2(maj_270_n20), .ZN(maj_270_n23)
         );
  XOR2_X1 maj_270_U9 ( .A(u_1_0[2]), .B(maj_270_n24), .Z(maj_270_n26) );
  XOR2_X1 maj_270_U8 ( .A(u_1_0[5]), .B(maj_270_n25), .Z(maj_270_n27) );
  XOR2_X1 maj_270_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_270_n24) );
  XOR2_X1 maj_270_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_270_n25) );
  OR2_X1 maj_270_U5 ( .A1(maj_270_n23), .A2(maj_270_n22), .ZN(maj_270_n32) );
  NAND2_X1 maj_270_U4 ( .A1(maj_270_n22), .A2(maj_270_n23), .ZN(maj_270_n34)
         );
  NAND2_X1 maj_270_U3 ( .A1(maj_270_n32), .A2(maj_270_n31), .ZN(maj_270_n33)
         );
  NAND2_X1 maj_270_U2 ( .A1(maj_270_n34), .A2(maj_270_n33), .ZN(maj_270_port_o) );
  OR2_X1 maj_271_U19 ( .A1(maj_271_n27), .A2(maj_271_n26), .ZN(maj_271_n28) );
  NAND2_X1 maj_271_U18 ( .A1(v_1_0[6]), .A2(maj_271_n28), .ZN(maj_271_n29) );
  NAND2_X1 maj_271_U17 ( .A1(maj_271_n26), .A2(maj_271_n27), .ZN(maj_271_n30)
         );
  NAND2_X1 maj_271_U16 ( .A1(maj_271_n30), .A2(maj_271_n29), .ZN(maj_271_n31)
         );
  NAND2_X1 maj_271_U15 ( .A1(v_1_0[5]), .A2(maj_271_n25), .ZN(maj_271_n18) );
  NAND2_X1 maj_271_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_271_n19) );
  NAND2_X1 maj_271_U13 ( .A1(maj_271_n19), .A2(maj_271_n18), .ZN(maj_271_n22)
         );
  NAND2_X1 maj_271_U12 ( .A1(v_1_0[2]), .A2(maj_271_n24), .ZN(maj_271_n20) );
  NAND2_X1 maj_271_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_271_n21) );
  NAND2_X1 maj_271_U10 ( .A1(maj_271_n21), .A2(maj_271_n20), .ZN(maj_271_n23)
         );
  XOR2_X1 maj_271_U9 ( .A(v_1_0[2]), .B(maj_271_n24), .Z(maj_271_n26) );
  XOR2_X1 maj_271_U8 ( .A(v_1_0[5]), .B(maj_271_n25), .Z(maj_271_n27) );
  XOR2_X1 maj_271_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_271_n24) );
  XOR2_X1 maj_271_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_271_n25) );
  OR2_X1 maj_271_U5 ( .A1(maj_271_n23), .A2(maj_271_n22), .ZN(maj_271_n32) );
  NAND2_X1 maj_271_U4 ( .A1(maj_271_n22), .A2(maj_271_n23), .ZN(maj_271_n34)
         );
  NAND2_X1 maj_271_U3 ( .A1(maj_271_n32), .A2(maj_271_n31), .ZN(maj_271_n33)
         );
  NAND2_X1 maj_271_U2 ( .A1(maj_271_n34), .A2(maj_271_n33), .ZN(maj_271_port_o) );
  OR2_X1 maj_272_U19 ( .A1(maj_272_n27), .A2(maj_272_n26), .ZN(maj_272_n28) );
  NAND2_X1 maj_272_U18 ( .A1(u_1_1[6]), .A2(maj_272_n28), .ZN(maj_272_n29) );
  NAND2_X1 maj_272_U17 ( .A1(maj_272_n26), .A2(maj_272_n27), .ZN(maj_272_n30)
         );
  NAND2_X1 maj_272_U16 ( .A1(maj_272_n30), .A2(maj_272_n29), .ZN(maj_272_n31)
         );
  NAND2_X1 maj_272_U15 ( .A1(u_1_1[5]), .A2(maj_272_n25), .ZN(maj_272_n18) );
  NAND2_X1 maj_272_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_272_n19) );
  NAND2_X1 maj_272_U13 ( .A1(maj_272_n19), .A2(maj_272_n18), .ZN(maj_272_n22)
         );
  NAND2_X1 maj_272_U12 ( .A1(u_1_1[2]), .A2(maj_272_n24), .ZN(maj_272_n20) );
  NAND2_X1 maj_272_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_272_n21) );
  NAND2_X1 maj_272_U10 ( .A1(maj_272_n21), .A2(maj_272_n20), .ZN(maj_272_n23)
         );
  XOR2_X1 maj_272_U9 ( .A(u_1_1[2]), .B(maj_272_n24), .Z(maj_272_n26) );
  XOR2_X1 maj_272_U8 ( .A(u_1_1[5]), .B(maj_272_n25), .Z(maj_272_n27) );
  XOR2_X1 maj_272_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_272_n24) );
  XOR2_X1 maj_272_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_272_n25) );
  OR2_X1 maj_272_U5 ( .A1(maj_272_n23), .A2(maj_272_n22), .ZN(maj_272_n32) );
  NAND2_X1 maj_272_U4 ( .A1(maj_272_n22), .A2(maj_272_n23), .ZN(maj_272_n34)
         );
  NAND2_X1 maj_272_U3 ( .A1(maj_272_n32), .A2(maj_272_n31), .ZN(maj_272_n33)
         );
  NAND2_X1 maj_272_U2 ( .A1(maj_272_n34), .A2(maj_272_n33), .ZN(maj_272_port_o) );
  OR2_X1 maj_273_U19 ( .A1(maj_273_n27), .A2(maj_273_n26), .ZN(maj_273_n28) );
  NAND2_X1 maj_273_U18 ( .A1(v_1_1[6]), .A2(maj_273_n28), .ZN(maj_273_n29) );
  NAND2_X1 maj_273_U17 ( .A1(maj_273_n26), .A2(maj_273_n27), .ZN(maj_273_n30)
         );
  NAND2_X1 maj_273_U16 ( .A1(maj_273_n30), .A2(maj_273_n29), .ZN(maj_273_n31)
         );
  NAND2_X1 maj_273_U15 ( .A1(v_1_1[5]), .A2(maj_273_n25), .ZN(maj_273_n18) );
  NAND2_X1 maj_273_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_273_n19) );
  NAND2_X1 maj_273_U13 ( .A1(maj_273_n19), .A2(maj_273_n18), .ZN(maj_273_n22)
         );
  NAND2_X1 maj_273_U12 ( .A1(v_1_1[2]), .A2(maj_273_n24), .ZN(maj_273_n20) );
  NAND2_X1 maj_273_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_273_n21) );
  NAND2_X1 maj_273_U10 ( .A1(maj_273_n21), .A2(maj_273_n20), .ZN(maj_273_n23)
         );
  XOR2_X1 maj_273_U9 ( .A(v_1_1[2]), .B(maj_273_n24), .Z(maj_273_n26) );
  XOR2_X1 maj_273_U8 ( .A(v_1_1[5]), .B(maj_273_n25), .Z(maj_273_n27) );
  XOR2_X1 maj_273_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_273_n24) );
  XOR2_X1 maj_273_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_273_n25) );
  OR2_X1 maj_273_U5 ( .A1(maj_273_n23), .A2(maj_273_n22), .ZN(maj_273_n32) );
  NAND2_X1 maj_273_U4 ( .A1(maj_273_n22), .A2(maj_273_n23), .ZN(maj_273_n34)
         );
  NAND2_X1 maj_273_U3 ( .A1(maj_273_n32), .A2(maj_273_n31), .ZN(maj_273_n33)
         );
  NAND2_X1 maj_273_U2 ( .A1(maj_273_n34), .A2(maj_273_n33), .ZN(maj_273_port_o) );
  OR2_X1 maj_274_U19 ( .A1(maj_274_n27), .A2(maj_274_n26), .ZN(maj_274_n28) );
  NAND2_X1 maj_274_U18 ( .A1(u_1_2[6]), .A2(maj_274_n28), .ZN(maj_274_n29) );
  NAND2_X1 maj_274_U17 ( .A1(maj_274_n26), .A2(maj_274_n27), .ZN(maj_274_n30)
         );
  NAND2_X1 maj_274_U16 ( .A1(maj_274_n30), .A2(maj_274_n29), .ZN(maj_274_n31)
         );
  NAND2_X1 maj_274_U15 ( .A1(u_1_2[5]), .A2(maj_274_n25), .ZN(maj_274_n18) );
  NAND2_X1 maj_274_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_274_n19) );
  NAND2_X1 maj_274_U13 ( .A1(maj_274_n19), .A2(maj_274_n18), .ZN(maj_274_n22)
         );
  NAND2_X1 maj_274_U12 ( .A1(u_1_2[2]), .A2(maj_274_n24), .ZN(maj_274_n20) );
  NAND2_X1 maj_274_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_274_n21) );
  NAND2_X1 maj_274_U10 ( .A1(maj_274_n21), .A2(maj_274_n20), .ZN(maj_274_n23)
         );
  XOR2_X1 maj_274_U9 ( .A(u_1_2[2]), .B(maj_274_n24), .Z(maj_274_n26) );
  XOR2_X1 maj_274_U8 ( .A(u_1_2[5]), .B(maj_274_n25), .Z(maj_274_n27) );
  XOR2_X1 maj_274_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_274_n24) );
  XOR2_X1 maj_274_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_274_n25) );
  OR2_X1 maj_274_U5 ( .A1(maj_274_n23), .A2(maj_274_n22), .ZN(maj_274_n32) );
  NAND2_X1 maj_274_U4 ( .A1(maj_274_n22), .A2(maj_274_n23), .ZN(maj_274_n34)
         );
  NAND2_X1 maj_274_U3 ( .A1(maj_274_n32), .A2(maj_274_n31), .ZN(maj_274_n33)
         );
  NAND2_X1 maj_274_U2 ( .A1(maj_274_n34), .A2(maj_274_n33), .ZN(maj_274_port_o) );
  OR2_X1 maj_275_U19 ( .A1(maj_275_n27), .A2(maj_275_n26), .ZN(maj_275_n28) );
  NAND2_X1 maj_275_U18 ( .A1(v_1_2[6]), .A2(maj_275_n28), .ZN(maj_275_n29) );
  NAND2_X1 maj_275_U17 ( .A1(maj_275_n26), .A2(maj_275_n27), .ZN(maj_275_n30)
         );
  NAND2_X1 maj_275_U16 ( .A1(maj_275_n30), .A2(maj_275_n29), .ZN(maj_275_n31)
         );
  NAND2_X1 maj_275_U15 ( .A1(v_1_2[5]), .A2(maj_275_n25), .ZN(maj_275_n18) );
  NAND2_X1 maj_275_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_275_n19) );
  NAND2_X1 maj_275_U13 ( .A1(maj_275_n19), .A2(maj_275_n18), .ZN(maj_275_n22)
         );
  NAND2_X1 maj_275_U12 ( .A1(v_1_2[2]), .A2(maj_275_n24), .ZN(maj_275_n20) );
  NAND2_X1 maj_275_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_275_n21) );
  NAND2_X1 maj_275_U10 ( .A1(maj_275_n21), .A2(maj_275_n20), .ZN(maj_275_n23)
         );
  XOR2_X1 maj_275_U9 ( .A(v_1_2[2]), .B(maj_275_n24), .Z(maj_275_n26) );
  XOR2_X1 maj_275_U8 ( .A(v_1_2[5]), .B(maj_275_n25), .Z(maj_275_n27) );
  XOR2_X1 maj_275_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_275_n24) );
  XOR2_X1 maj_275_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_275_n25) );
  OR2_X1 maj_275_U5 ( .A1(maj_275_n23), .A2(maj_275_n22), .ZN(maj_275_n32) );
  NAND2_X1 maj_275_U4 ( .A1(maj_275_n22), .A2(maj_275_n23), .ZN(maj_275_n34)
         );
  NAND2_X1 maj_275_U3 ( .A1(maj_275_n32), .A2(maj_275_n31), .ZN(maj_275_n33)
         );
  NAND2_X1 maj_275_U2 ( .A1(maj_275_n34), .A2(maj_275_n33), .ZN(maj_275_port_o) );
  OR2_X1 maj_276_U19 ( .A1(maj_276_n27), .A2(maj_276_n26), .ZN(maj_276_n28) );
  NAND2_X1 maj_276_U18 ( .A1(u_2_0[6]), .A2(maj_276_n28), .ZN(maj_276_n29) );
  NAND2_X1 maj_276_U17 ( .A1(maj_276_n26), .A2(maj_276_n27), .ZN(maj_276_n30)
         );
  NAND2_X1 maj_276_U16 ( .A1(maj_276_n30), .A2(maj_276_n29), .ZN(maj_276_n31)
         );
  NAND2_X1 maj_276_U15 ( .A1(u_2_0[5]), .A2(maj_276_n25), .ZN(maj_276_n18) );
  NAND2_X1 maj_276_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_276_n19) );
  NAND2_X1 maj_276_U13 ( .A1(maj_276_n19), .A2(maj_276_n18), .ZN(maj_276_n22)
         );
  NAND2_X1 maj_276_U12 ( .A1(u_2_0[2]), .A2(maj_276_n24), .ZN(maj_276_n20) );
  NAND2_X1 maj_276_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_276_n21) );
  NAND2_X1 maj_276_U10 ( .A1(maj_276_n21), .A2(maj_276_n20), .ZN(maj_276_n23)
         );
  XOR2_X1 maj_276_U9 ( .A(u_2_0[2]), .B(maj_276_n24), .Z(maj_276_n26) );
  XOR2_X1 maj_276_U8 ( .A(u_2_0[5]), .B(maj_276_n25), .Z(maj_276_n27) );
  XOR2_X1 maj_276_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_276_n24) );
  XOR2_X1 maj_276_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_276_n25) );
  OR2_X1 maj_276_U5 ( .A1(maj_276_n23), .A2(maj_276_n22), .ZN(maj_276_n32) );
  NAND2_X1 maj_276_U4 ( .A1(maj_276_n22), .A2(maj_276_n23), .ZN(maj_276_n34)
         );
  NAND2_X1 maj_276_U3 ( .A1(maj_276_n32), .A2(maj_276_n31), .ZN(maj_276_n33)
         );
  NAND2_X1 maj_276_U2 ( .A1(maj_276_n34), .A2(maj_276_n33), .ZN(maj_276_port_o) );
  OR2_X1 maj_277_U19 ( .A1(maj_277_n27), .A2(maj_277_n26), .ZN(maj_277_n28) );
  NAND2_X1 maj_277_U18 ( .A1(v_2_0[6]), .A2(maj_277_n28), .ZN(maj_277_n29) );
  NAND2_X1 maj_277_U17 ( .A1(maj_277_n26), .A2(maj_277_n27), .ZN(maj_277_n30)
         );
  NAND2_X1 maj_277_U16 ( .A1(maj_277_n30), .A2(maj_277_n29), .ZN(maj_277_n31)
         );
  NAND2_X1 maj_277_U15 ( .A1(v_2_0[5]), .A2(maj_277_n25), .ZN(maj_277_n18) );
  NAND2_X1 maj_277_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_277_n19) );
  NAND2_X1 maj_277_U13 ( .A1(maj_277_n19), .A2(maj_277_n18), .ZN(maj_277_n22)
         );
  NAND2_X1 maj_277_U12 ( .A1(v_2_0[2]), .A2(maj_277_n24), .ZN(maj_277_n20) );
  NAND2_X1 maj_277_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_277_n21) );
  NAND2_X1 maj_277_U10 ( .A1(maj_277_n21), .A2(maj_277_n20), .ZN(maj_277_n23)
         );
  XOR2_X1 maj_277_U9 ( .A(v_2_0[2]), .B(maj_277_n24), .Z(maj_277_n26) );
  XOR2_X1 maj_277_U8 ( .A(v_2_0[5]), .B(maj_277_n25), .Z(maj_277_n27) );
  XOR2_X1 maj_277_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_277_n24) );
  XOR2_X1 maj_277_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_277_n25) );
  OR2_X1 maj_277_U5 ( .A1(maj_277_n23), .A2(maj_277_n22), .ZN(maj_277_n32) );
  NAND2_X1 maj_277_U4 ( .A1(maj_277_n22), .A2(maj_277_n23), .ZN(maj_277_n34)
         );
  NAND2_X1 maj_277_U3 ( .A1(maj_277_n32), .A2(maj_277_n31), .ZN(maj_277_n33)
         );
  NAND2_X1 maj_277_U2 ( .A1(maj_277_n34), .A2(maj_277_n33), .ZN(maj_277_port_o) );
  OR2_X1 maj_278_U19 ( .A1(maj_278_n27), .A2(maj_278_n26), .ZN(maj_278_n28) );
  NAND2_X1 maj_278_U18 ( .A1(u_2_1[6]), .A2(maj_278_n28), .ZN(maj_278_n29) );
  NAND2_X1 maj_278_U17 ( .A1(maj_278_n26), .A2(maj_278_n27), .ZN(maj_278_n30)
         );
  NAND2_X1 maj_278_U16 ( .A1(maj_278_n30), .A2(maj_278_n29), .ZN(maj_278_n31)
         );
  NAND2_X1 maj_278_U15 ( .A1(u_2_1[5]), .A2(maj_278_n25), .ZN(maj_278_n18) );
  NAND2_X1 maj_278_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_278_n19) );
  NAND2_X1 maj_278_U13 ( .A1(maj_278_n19), .A2(maj_278_n18), .ZN(maj_278_n22)
         );
  NAND2_X1 maj_278_U12 ( .A1(u_2_1[2]), .A2(maj_278_n24), .ZN(maj_278_n20) );
  NAND2_X1 maj_278_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_278_n21) );
  NAND2_X1 maj_278_U10 ( .A1(maj_278_n21), .A2(maj_278_n20), .ZN(maj_278_n23)
         );
  XOR2_X1 maj_278_U9 ( .A(u_2_1[2]), .B(maj_278_n24), .Z(maj_278_n26) );
  XOR2_X1 maj_278_U8 ( .A(u_2_1[5]), .B(maj_278_n25), .Z(maj_278_n27) );
  XOR2_X1 maj_278_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_278_n24) );
  XOR2_X1 maj_278_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_278_n25) );
  OR2_X1 maj_278_U5 ( .A1(maj_278_n23), .A2(maj_278_n22), .ZN(maj_278_n32) );
  NAND2_X1 maj_278_U4 ( .A1(maj_278_n22), .A2(maj_278_n23), .ZN(maj_278_n34)
         );
  NAND2_X1 maj_278_U3 ( .A1(maj_278_n32), .A2(maj_278_n31), .ZN(maj_278_n33)
         );
  NAND2_X1 maj_278_U2 ( .A1(maj_278_n34), .A2(maj_278_n33), .ZN(maj_278_port_o) );
  OR2_X1 maj_279_U19 ( .A1(maj_279_n27), .A2(maj_279_n26), .ZN(maj_279_n28) );
  NAND2_X1 maj_279_U18 ( .A1(v_2_1[6]), .A2(maj_279_n28), .ZN(maj_279_n29) );
  NAND2_X1 maj_279_U17 ( .A1(maj_279_n26), .A2(maj_279_n27), .ZN(maj_279_n30)
         );
  NAND2_X1 maj_279_U16 ( .A1(maj_279_n30), .A2(maj_279_n29), .ZN(maj_279_n31)
         );
  NAND2_X1 maj_279_U15 ( .A1(v_2_1[5]), .A2(maj_279_n25), .ZN(maj_279_n18) );
  NAND2_X1 maj_279_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_279_n19) );
  NAND2_X1 maj_279_U13 ( .A1(maj_279_n19), .A2(maj_279_n18), .ZN(maj_279_n22)
         );
  NAND2_X1 maj_279_U12 ( .A1(v_2_1[2]), .A2(maj_279_n24), .ZN(maj_279_n20) );
  NAND2_X1 maj_279_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_279_n21) );
  NAND2_X1 maj_279_U10 ( .A1(maj_279_n21), .A2(maj_279_n20), .ZN(maj_279_n23)
         );
  XOR2_X1 maj_279_U9 ( .A(v_2_1[2]), .B(maj_279_n24), .Z(maj_279_n26) );
  XOR2_X1 maj_279_U8 ( .A(v_2_1[5]), .B(maj_279_n25), .Z(maj_279_n27) );
  XOR2_X1 maj_279_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_279_n24) );
  XOR2_X1 maj_279_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_279_n25) );
  OR2_X1 maj_279_U5 ( .A1(maj_279_n23), .A2(maj_279_n22), .ZN(maj_279_n32) );
  NAND2_X1 maj_279_U4 ( .A1(maj_279_n22), .A2(maj_279_n23), .ZN(maj_279_n34)
         );
  NAND2_X1 maj_279_U3 ( .A1(maj_279_n32), .A2(maj_279_n31), .ZN(maj_279_n33)
         );
  NAND2_X1 maj_279_U2 ( .A1(maj_279_n34), .A2(maj_279_n33), .ZN(maj_279_port_o) );
  OR2_X1 maj_280_U19 ( .A1(maj_280_n27), .A2(maj_280_n26), .ZN(maj_280_n28) );
  NAND2_X1 maj_280_U18 ( .A1(u_2_2[6]), .A2(maj_280_n28), .ZN(maj_280_n29) );
  NAND2_X1 maj_280_U17 ( .A1(maj_280_n26), .A2(maj_280_n27), .ZN(maj_280_n30)
         );
  NAND2_X1 maj_280_U16 ( .A1(maj_280_n30), .A2(maj_280_n29), .ZN(maj_280_n31)
         );
  NAND2_X1 maj_280_U15 ( .A1(u_2_2[5]), .A2(maj_280_n25), .ZN(maj_280_n18) );
  NAND2_X1 maj_280_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_280_n19) );
  NAND2_X1 maj_280_U13 ( .A1(maj_280_n19), .A2(maj_280_n18), .ZN(maj_280_n22)
         );
  NAND2_X1 maj_280_U12 ( .A1(u_2_2[2]), .A2(maj_280_n24), .ZN(maj_280_n20) );
  NAND2_X1 maj_280_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_280_n21) );
  NAND2_X1 maj_280_U10 ( .A1(maj_280_n21), .A2(maj_280_n20), .ZN(maj_280_n23)
         );
  XOR2_X1 maj_280_U9 ( .A(u_2_2[2]), .B(maj_280_n24), .Z(maj_280_n26) );
  XOR2_X1 maj_280_U8 ( .A(u_2_2[5]), .B(maj_280_n25), .Z(maj_280_n27) );
  XOR2_X1 maj_280_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_280_n24) );
  XOR2_X1 maj_280_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_280_n25) );
  OR2_X1 maj_280_U5 ( .A1(maj_280_n23), .A2(maj_280_n22), .ZN(maj_280_n32) );
  NAND2_X1 maj_280_U4 ( .A1(maj_280_n22), .A2(maj_280_n23), .ZN(maj_280_n34)
         );
  NAND2_X1 maj_280_U3 ( .A1(maj_280_n32), .A2(maj_280_n31), .ZN(maj_280_n33)
         );
  NAND2_X1 maj_280_U2 ( .A1(maj_280_n34), .A2(maj_280_n33), .ZN(maj_280_port_o) );
  OR2_X1 maj_281_U19 ( .A1(maj_281_n27), .A2(maj_281_n26), .ZN(maj_281_n28) );
  NAND2_X1 maj_281_U18 ( .A1(v_2_2[6]), .A2(maj_281_n28), .ZN(maj_281_n29) );
  NAND2_X1 maj_281_U17 ( .A1(maj_281_n26), .A2(maj_281_n27), .ZN(maj_281_n30)
         );
  NAND2_X1 maj_281_U16 ( .A1(maj_281_n30), .A2(maj_281_n29), .ZN(maj_281_n31)
         );
  NAND2_X1 maj_281_U15 ( .A1(v_2_2[5]), .A2(maj_281_n25), .ZN(maj_281_n18) );
  NAND2_X1 maj_281_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_281_n19) );
  NAND2_X1 maj_281_U13 ( .A1(maj_281_n19), .A2(maj_281_n18), .ZN(maj_281_n22)
         );
  NAND2_X1 maj_281_U12 ( .A1(v_2_2[2]), .A2(maj_281_n24), .ZN(maj_281_n20) );
  NAND2_X1 maj_281_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_281_n21) );
  NAND2_X1 maj_281_U10 ( .A1(maj_281_n21), .A2(maj_281_n20), .ZN(maj_281_n23)
         );
  XOR2_X1 maj_281_U9 ( .A(v_2_2[2]), .B(maj_281_n24), .Z(maj_281_n26) );
  XOR2_X1 maj_281_U8 ( .A(v_2_2[5]), .B(maj_281_n25), .Z(maj_281_n27) );
  XOR2_X1 maj_281_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_281_n24) );
  XOR2_X1 maj_281_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_281_n25) );
  OR2_X1 maj_281_U5 ( .A1(maj_281_n23), .A2(maj_281_n22), .ZN(maj_281_n32) );
  NAND2_X1 maj_281_U4 ( .A1(maj_281_n22), .A2(maj_281_n23), .ZN(maj_281_n34)
         );
  NAND2_X1 maj_281_U3 ( .A1(maj_281_n32), .A2(maj_281_n31), .ZN(maj_281_n33)
         );
  NAND2_X1 maj_281_U2 ( .A1(maj_281_n34), .A2(maj_281_n33), .ZN(maj_281_port_o) );
  OR2_X1 maj_282_U19 ( .A1(maj_282_n27), .A2(maj_282_n26), .ZN(maj_282_n28) );
  NAND2_X1 maj_282_U18 ( .A1(u_3_0[6]), .A2(maj_282_n28), .ZN(maj_282_n29) );
  NAND2_X1 maj_282_U17 ( .A1(maj_282_n26), .A2(maj_282_n27), .ZN(maj_282_n30)
         );
  NAND2_X1 maj_282_U16 ( .A1(maj_282_n30), .A2(maj_282_n29), .ZN(maj_282_n31)
         );
  NAND2_X1 maj_282_U15 ( .A1(u_3_0[5]), .A2(maj_282_n25), .ZN(maj_282_n18) );
  NAND2_X1 maj_282_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_282_n19) );
  NAND2_X1 maj_282_U13 ( .A1(maj_282_n19), .A2(maj_282_n18), .ZN(maj_282_n22)
         );
  NAND2_X1 maj_282_U12 ( .A1(u_3_0[2]), .A2(maj_282_n24), .ZN(maj_282_n20) );
  NAND2_X1 maj_282_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_282_n21) );
  NAND2_X1 maj_282_U10 ( .A1(maj_282_n21), .A2(maj_282_n20), .ZN(maj_282_n23)
         );
  XOR2_X1 maj_282_U9 ( .A(u_3_0[2]), .B(maj_282_n24), .Z(maj_282_n26) );
  XOR2_X1 maj_282_U8 ( .A(u_3_0[5]), .B(maj_282_n25), .Z(maj_282_n27) );
  XOR2_X1 maj_282_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_282_n24) );
  XOR2_X1 maj_282_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_282_n25) );
  OR2_X1 maj_282_U5 ( .A1(maj_282_n23), .A2(maj_282_n22), .ZN(maj_282_n32) );
  NAND2_X1 maj_282_U4 ( .A1(maj_282_n22), .A2(maj_282_n23), .ZN(maj_282_n34)
         );
  NAND2_X1 maj_282_U3 ( .A1(maj_282_n32), .A2(maj_282_n31), .ZN(maj_282_n33)
         );
  NAND2_X1 maj_282_U2 ( .A1(maj_282_n34), .A2(maj_282_n33), .ZN(maj_282_port_o) );
  OR2_X1 maj_283_U19 ( .A1(maj_283_n27), .A2(maj_283_n26), .ZN(maj_283_n28) );
  NAND2_X1 maj_283_U18 ( .A1(v_3_0[6]), .A2(maj_283_n28), .ZN(maj_283_n29) );
  NAND2_X1 maj_283_U17 ( .A1(maj_283_n26), .A2(maj_283_n27), .ZN(maj_283_n30)
         );
  NAND2_X1 maj_283_U16 ( .A1(maj_283_n30), .A2(maj_283_n29), .ZN(maj_283_n31)
         );
  NAND2_X1 maj_283_U15 ( .A1(v_3_0[5]), .A2(maj_283_n25), .ZN(maj_283_n18) );
  NAND2_X1 maj_283_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_283_n19) );
  NAND2_X1 maj_283_U13 ( .A1(maj_283_n19), .A2(maj_283_n18), .ZN(maj_283_n22)
         );
  NAND2_X1 maj_283_U12 ( .A1(v_3_0[2]), .A2(maj_283_n24), .ZN(maj_283_n20) );
  NAND2_X1 maj_283_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_283_n21) );
  NAND2_X1 maj_283_U10 ( .A1(maj_283_n21), .A2(maj_283_n20), .ZN(maj_283_n23)
         );
  XOR2_X1 maj_283_U9 ( .A(v_3_0[2]), .B(maj_283_n24), .Z(maj_283_n26) );
  XOR2_X1 maj_283_U8 ( .A(v_3_0[5]), .B(maj_283_n25), .Z(maj_283_n27) );
  XOR2_X1 maj_283_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_283_n24) );
  XOR2_X1 maj_283_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_283_n25) );
  OR2_X1 maj_283_U5 ( .A1(maj_283_n23), .A2(maj_283_n22), .ZN(maj_283_n32) );
  NAND2_X1 maj_283_U4 ( .A1(maj_283_n22), .A2(maj_283_n23), .ZN(maj_283_n34)
         );
  NAND2_X1 maj_283_U3 ( .A1(maj_283_n32), .A2(maj_283_n31), .ZN(maj_283_n33)
         );
  NAND2_X1 maj_283_U2 ( .A1(maj_283_n34), .A2(maj_283_n33), .ZN(maj_283_port_o) );
  OR2_X1 maj_284_U19 ( .A1(maj_284_n27), .A2(maj_284_n26), .ZN(maj_284_n28) );
  NAND2_X1 maj_284_U18 ( .A1(u_3_1[6]), .A2(maj_284_n28), .ZN(maj_284_n29) );
  NAND2_X1 maj_284_U17 ( .A1(maj_284_n26), .A2(maj_284_n27), .ZN(maj_284_n30)
         );
  NAND2_X1 maj_284_U16 ( .A1(maj_284_n30), .A2(maj_284_n29), .ZN(maj_284_n31)
         );
  NAND2_X1 maj_284_U15 ( .A1(u_3_1[5]), .A2(maj_284_n25), .ZN(maj_284_n18) );
  NAND2_X1 maj_284_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_284_n19) );
  NAND2_X1 maj_284_U13 ( .A1(maj_284_n19), .A2(maj_284_n18), .ZN(maj_284_n22)
         );
  NAND2_X1 maj_284_U12 ( .A1(u_3_1[2]), .A2(maj_284_n24), .ZN(maj_284_n20) );
  NAND2_X1 maj_284_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_284_n21) );
  NAND2_X1 maj_284_U10 ( .A1(maj_284_n21), .A2(maj_284_n20), .ZN(maj_284_n23)
         );
  XOR2_X1 maj_284_U9 ( .A(u_3_1[2]), .B(maj_284_n24), .Z(maj_284_n26) );
  XOR2_X1 maj_284_U8 ( .A(u_3_1[5]), .B(maj_284_n25), .Z(maj_284_n27) );
  XOR2_X1 maj_284_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_284_n24) );
  XOR2_X1 maj_284_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_284_n25) );
  OR2_X1 maj_284_U5 ( .A1(maj_284_n23), .A2(maj_284_n22), .ZN(maj_284_n32) );
  NAND2_X1 maj_284_U4 ( .A1(maj_284_n22), .A2(maj_284_n23), .ZN(maj_284_n34)
         );
  NAND2_X1 maj_284_U3 ( .A1(maj_284_n32), .A2(maj_284_n31), .ZN(maj_284_n33)
         );
  NAND2_X1 maj_284_U2 ( .A1(maj_284_n34), .A2(maj_284_n33), .ZN(maj_284_port_o) );
  OR2_X1 maj_285_U19 ( .A1(maj_285_n27), .A2(maj_285_n26), .ZN(maj_285_n28) );
  NAND2_X1 maj_285_U18 ( .A1(v_3_1[6]), .A2(maj_285_n28), .ZN(maj_285_n29) );
  NAND2_X1 maj_285_U17 ( .A1(maj_285_n26), .A2(maj_285_n27), .ZN(maj_285_n30)
         );
  NAND2_X1 maj_285_U16 ( .A1(maj_285_n30), .A2(maj_285_n29), .ZN(maj_285_n31)
         );
  NAND2_X1 maj_285_U15 ( .A1(v_3_1[5]), .A2(maj_285_n25), .ZN(maj_285_n18) );
  NAND2_X1 maj_285_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_285_n19) );
  NAND2_X1 maj_285_U13 ( .A1(maj_285_n19), .A2(maj_285_n18), .ZN(maj_285_n22)
         );
  NAND2_X1 maj_285_U12 ( .A1(v_3_1[2]), .A2(maj_285_n24), .ZN(maj_285_n20) );
  NAND2_X1 maj_285_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_285_n21) );
  NAND2_X1 maj_285_U10 ( .A1(maj_285_n21), .A2(maj_285_n20), .ZN(maj_285_n23)
         );
  XOR2_X1 maj_285_U9 ( .A(v_3_1[2]), .B(maj_285_n24), .Z(maj_285_n26) );
  XOR2_X1 maj_285_U8 ( .A(v_3_1[5]), .B(maj_285_n25), .Z(maj_285_n27) );
  XOR2_X1 maj_285_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_285_n24) );
  XOR2_X1 maj_285_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_285_n25) );
  OR2_X1 maj_285_U5 ( .A1(maj_285_n23), .A2(maj_285_n22), .ZN(maj_285_n32) );
  NAND2_X1 maj_285_U4 ( .A1(maj_285_n22), .A2(maj_285_n23), .ZN(maj_285_n34)
         );
  NAND2_X1 maj_285_U3 ( .A1(maj_285_n32), .A2(maj_285_n31), .ZN(maj_285_n33)
         );
  NAND2_X1 maj_285_U2 ( .A1(maj_285_n34), .A2(maj_285_n33), .ZN(maj_285_port_o) );
  OR2_X1 maj_286_U19 ( .A1(maj_286_n27), .A2(maj_286_n26), .ZN(maj_286_n28) );
  NAND2_X1 maj_286_U18 ( .A1(u_3_2[6]), .A2(maj_286_n28), .ZN(maj_286_n29) );
  NAND2_X1 maj_286_U17 ( .A1(maj_286_n26), .A2(maj_286_n27), .ZN(maj_286_n30)
         );
  NAND2_X1 maj_286_U16 ( .A1(maj_286_n30), .A2(maj_286_n29), .ZN(maj_286_n31)
         );
  NAND2_X1 maj_286_U15 ( .A1(u_3_2[5]), .A2(maj_286_n25), .ZN(maj_286_n18) );
  NAND2_X1 maj_286_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_286_n19) );
  NAND2_X1 maj_286_U13 ( .A1(maj_286_n19), .A2(maj_286_n18), .ZN(maj_286_n22)
         );
  NAND2_X1 maj_286_U12 ( .A1(u_3_2[2]), .A2(maj_286_n24), .ZN(maj_286_n20) );
  NAND2_X1 maj_286_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_286_n21) );
  NAND2_X1 maj_286_U10 ( .A1(maj_286_n21), .A2(maj_286_n20), .ZN(maj_286_n23)
         );
  XOR2_X1 maj_286_U9 ( .A(u_3_2[2]), .B(maj_286_n24), .Z(maj_286_n26) );
  XOR2_X1 maj_286_U8 ( .A(u_3_2[5]), .B(maj_286_n25), .Z(maj_286_n27) );
  XOR2_X1 maj_286_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_286_n24) );
  XOR2_X1 maj_286_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_286_n25) );
  OR2_X1 maj_286_U5 ( .A1(maj_286_n23), .A2(maj_286_n22), .ZN(maj_286_n32) );
  NAND2_X1 maj_286_U4 ( .A1(maj_286_n22), .A2(maj_286_n23), .ZN(maj_286_n34)
         );
  NAND2_X1 maj_286_U3 ( .A1(maj_286_n32), .A2(maj_286_n31), .ZN(maj_286_n33)
         );
  NAND2_X1 maj_286_U2 ( .A1(maj_286_n34), .A2(maj_286_n33), .ZN(maj_286_port_o) );
  OR2_X1 maj_287_U19 ( .A1(maj_287_n27), .A2(maj_287_n26), .ZN(maj_287_n28) );
  NAND2_X1 maj_287_U18 ( .A1(v_3_2[6]), .A2(maj_287_n28), .ZN(maj_287_n29) );
  NAND2_X1 maj_287_U17 ( .A1(maj_287_n26), .A2(maj_287_n27), .ZN(maj_287_n30)
         );
  NAND2_X1 maj_287_U16 ( .A1(maj_287_n30), .A2(maj_287_n29), .ZN(maj_287_n31)
         );
  NAND2_X1 maj_287_U15 ( .A1(v_3_2[5]), .A2(maj_287_n25), .ZN(maj_287_n18) );
  NAND2_X1 maj_287_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_287_n19) );
  NAND2_X1 maj_287_U13 ( .A1(maj_287_n19), .A2(maj_287_n18), .ZN(maj_287_n22)
         );
  NAND2_X1 maj_287_U12 ( .A1(v_3_2[2]), .A2(maj_287_n24), .ZN(maj_287_n20) );
  NAND2_X1 maj_287_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_287_n21) );
  NAND2_X1 maj_287_U10 ( .A1(maj_287_n21), .A2(maj_287_n20), .ZN(maj_287_n23)
         );
  XOR2_X1 maj_287_U9 ( .A(v_3_2[2]), .B(maj_287_n24), .Z(maj_287_n26) );
  XOR2_X1 maj_287_U8 ( .A(v_3_2[5]), .B(maj_287_n25), .Z(maj_287_n27) );
  XOR2_X1 maj_287_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_287_n24) );
  XOR2_X1 maj_287_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_287_n25) );
  OR2_X1 maj_287_U5 ( .A1(maj_287_n23), .A2(maj_287_n22), .ZN(maj_287_n32) );
  NAND2_X1 maj_287_U4 ( .A1(maj_287_n22), .A2(maj_287_n23), .ZN(maj_287_n34)
         );
  NAND2_X1 maj_287_U3 ( .A1(maj_287_n32), .A2(maj_287_n31), .ZN(maj_287_n33)
         );
  NAND2_X1 maj_287_U2 ( .A1(maj_287_n34), .A2(maj_287_n33), .ZN(maj_287_port_o) );
  OR2_X1 maj_288_U19 ( .A1(maj_288_n27), .A2(maj_288_n26), .ZN(maj_288_n28) );
  NAND2_X1 maj_288_U18 ( .A1(u_0_0[6]), .A2(maj_288_n28), .ZN(maj_288_n29) );
  NAND2_X1 maj_288_U17 ( .A1(maj_288_n26), .A2(maj_288_n27), .ZN(maj_288_n30)
         );
  NAND2_X1 maj_288_U16 ( .A1(maj_288_n30), .A2(maj_288_n29), .ZN(maj_288_n31)
         );
  NAND2_X1 maj_288_U15 ( .A1(u_0_0[5]), .A2(maj_288_n25), .ZN(maj_288_n18) );
  NAND2_X1 maj_288_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_288_n19) );
  NAND2_X1 maj_288_U13 ( .A1(maj_288_n19), .A2(maj_288_n18), .ZN(maj_288_n22)
         );
  NAND2_X1 maj_288_U12 ( .A1(u_0_0[2]), .A2(maj_288_n24), .ZN(maj_288_n20) );
  NAND2_X1 maj_288_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_288_n21) );
  NAND2_X1 maj_288_U10 ( .A1(maj_288_n21), .A2(maj_288_n20), .ZN(maj_288_n23)
         );
  XOR2_X1 maj_288_U9 ( .A(u_0_0[2]), .B(maj_288_n24), .Z(maj_288_n26) );
  XOR2_X1 maj_288_U8 ( .A(u_0_0[5]), .B(maj_288_n25), .Z(maj_288_n27) );
  XOR2_X1 maj_288_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_288_n24) );
  XOR2_X1 maj_288_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_288_n25) );
  OR2_X1 maj_288_U5 ( .A1(maj_288_n23), .A2(maj_288_n22), .ZN(maj_288_n32) );
  NAND2_X1 maj_288_U4 ( .A1(maj_288_n22), .A2(maj_288_n23), .ZN(maj_288_n34)
         );
  NAND2_X1 maj_288_U3 ( .A1(maj_288_n32), .A2(maj_288_n31), .ZN(maj_288_n33)
         );
  NAND2_X1 maj_288_U2 ( .A1(maj_288_n34), .A2(maj_288_n33), .ZN(maj_288_port_o) );
  OR2_X1 maj_289_U19 ( .A1(maj_289_n27), .A2(maj_289_n26), .ZN(maj_289_n28) );
  NAND2_X1 maj_289_U18 ( .A1(v_0_0[6]), .A2(maj_289_n28), .ZN(maj_289_n29) );
  NAND2_X1 maj_289_U17 ( .A1(maj_289_n26), .A2(maj_289_n27), .ZN(maj_289_n30)
         );
  NAND2_X1 maj_289_U16 ( .A1(maj_289_n30), .A2(maj_289_n29), .ZN(maj_289_n31)
         );
  NAND2_X1 maj_289_U15 ( .A1(v_0_0[5]), .A2(maj_289_n25), .ZN(maj_289_n18) );
  NAND2_X1 maj_289_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_289_n19) );
  NAND2_X1 maj_289_U13 ( .A1(maj_289_n19), .A2(maj_289_n18), .ZN(maj_289_n22)
         );
  NAND2_X1 maj_289_U12 ( .A1(v_0_0[2]), .A2(maj_289_n24), .ZN(maj_289_n20) );
  NAND2_X1 maj_289_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_289_n21) );
  NAND2_X1 maj_289_U10 ( .A1(maj_289_n21), .A2(maj_289_n20), .ZN(maj_289_n23)
         );
  XOR2_X1 maj_289_U9 ( .A(v_0_0[2]), .B(maj_289_n24), .Z(maj_289_n26) );
  XOR2_X1 maj_289_U8 ( .A(v_0_0[5]), .B(maj_289_n25), .Z(maj_289_n27) );
  XOR2_X1 maj_289_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_289_n24) );
  XOR2_X1 maj_289_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_289_n25) );
  OR2_X1 maj_289_U5 ( .A1(maj_289_n23), .A2(maj_289_n22), .ZN(maj_289_n32) );
  NAND2_X1 maj_289_U4 ( .A1(maj_289_n22), .A2(maj_289_n23), .ZN(maj_289_n34)
         );
  NAND2_X1 maj_289_U3 ( .A1(maj_289_n32), .A2(maj_289_n31), .ZN(maj_289_n33)
         );
  NAND2_X1 maj_289_U2 ( .A1(maj_289_n34), .A2(maj_289_n33), .ZN(maj_289_port_o) );
  OR2_X1 maj_290_U19 ( .A1(maj_290_n27), .A2(maj_290_n26), .ZN(maj_290_n28) );
  NAND2_X1 maj_290_U18 ( .A1(u_0_1[6]), .A2(maj_290_n28), .ZN(maj_290_n29) );
  NAND2_X1 maj_290_U17 ( .A1(maj_290_n26), .A2(maj_290_n27), .ZN(maj_290_n30)
         );
  NAND2_X1 maj_290_U16 ( .A1(maj_290_n30), .A2(maj_290_n29), .ZN(maj_290_n31)
         );
  NAND2_X1 maj_290_U15 ( .A1(u_0_1[5]), .A2(maj_290_n25), .ZN(maj_290_n18) );
  NAND2_X1 maj_290_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_290_n19) );
  NAND2_X1 maj_290_U13 ( .A1(maj_290_n19), .A2(maj_290_n18), .ZN(maj_290_n22)
         );
  NAND2_X1 maj_290_U12 ( .A1(u_0_1[2]), .A2(maj_290_n24), .ZN(maj_290_n20) );
  NAND2_X1 maj_290_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_290_n21) );
  NAND2_X1 maj_290_U10 ( .A1(maj_290_n21), .A2(maj_290_n20), .ZN(maj_290_n23)
         );
  XOR2_X1 maj_290_U9 ( .A(u_0_1[2]), .B(maj_290_n24), .Z(maj_290_n26) );
  XOR2_X1 maj_290_U8 ( .A(u_0_1[5]), .B(maj_290_n25), .Z(maj_290_n27) );
  XOR2_X1 maj_290_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_290_n24) );
  XOR2_X1 maj_290_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_290_n25) );
  OR2_X1 maj_290_U5 ( .A1(maj_290_n23), .A2(maj_290_n22), .ZN(maj_290_n32) );
  NAND2_X1 maj_290_U4 ( .A1(maj_290_n22), .A2(maj_290_n23), .ZN(maj_290_n34)
         );
  NAND2_X1 maj_290_U3 ( .A1(maj_290_n32), .A2(maj_290_n31), .ZN(maj_290_n33)
         );
  NAND2_X1 maj_290_U2 ( .A1(maj_290_n34), .A2(maj_290_n33), .ZN(maj_290_port_o) );
  OR2_X1 maj_291_U19 ( .A1(maj_291_n27), .A2(maj_291_n26), .ZN(maj_291_n28) );
  NAND2_X1 maj_291_U18 ( .A1(v_0_1[6]), .A2(maj_291_n28), .ZN(maj_291_n29) );
  NAND2_X1 maj_291_U17 ( .A1(maj_291_n26), .A2(maj_291_n27), .ZN(maj_291_n30)
         );
  NAND2_X1 maj_291_U16 ( .A1(maj_291_n30), .A2(maj_291_n29), .ZN(maj_291_n31)
         );
  NAND2_X1 maj_291_U15 ( .A1(v_0_1[5]), .A2(maj_291_n25), .ZN(maj_291_n18) );
  NAND2_X1 maj_291_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_291_n19) );
  NAND2_X1 maj_291_U13 ( .A1(maj_291_n19), .A2(maj_291_n18), .ZN(maj_291_n22)
         );
  NAND2_X1 maj_291_U12 ( .A1(v_0_1[2]), .A2(maj_291_n24), .ZN(maj_291_n20) );
  NAND2_X1 maj_291_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_291_n21) );
  NAND2_X1 maj_291_U10 ( .A1(maj_291_n21), .A2(maj_291_n20), .ZN(maj_291_n23)
         );
  XOR2_X1 maj_291_U9 ( .A(v_0_1[2]), .B(maj_291_n24), .Z(maj_291_n26) );
  XOR2_X1 maj_291_U8 ( .A(v_0_1[5]), .B(maj_291_n25), .Z(maj_291_n27) );
  XOR2_X1 maj_291_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_291_n24) );
  XOR2_X1 maj_291_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_291_n25) );
  OR2_X1 maj_291_U5 ( .A1(maj_291_n23), .A2(maj_291_n22), .ZN(maj_291_n32) );
  NAND2_X1 maj_291_U4 ( .A1(maj_291_n22), .A2(maj_291_n23), .ZN(maj_291_n34)
         );
  NAND2_X1 maj_291_U3 ( .A1(maj_291_n32), .A2(maj_291_n31), .ZN(maj_291_n33)
         );
  NAND2_X1 maj_291_U2 ( .A1(maj_291_n34), .A2(maj_291_n33), .ZN(maj_291_port_o) );
  OR2_X1 maj_292_U19 ( .A1(maj_292_n27), .A2(maj_292_n26), .ZN(maj_292_n28) );
  NAND2_X1 maj_292_U18 ( .A1(u_0_2[6]), .A2(maj_292_n28), .ZN(maj_292_n29) );
  NAND2_X1 maj_292_U17 ( .A1(maj_292_n26), .A2(maj_292_n27), .ZN(maj_292_n30)
         );
  NAND2_X1 maj_292_U16 ( .A1(maj_292_n30), .A2(maj_292_n29), .ZN(maj_292_n31)
         );
  NAND2_X1 maj_292_U15 ( .A1(u_0_2[5]), .A2(maj_292_n25), .ZN(maj_292_n18) );
  NAND2_X1 maj_292_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_292_n19) );
  NAND2_X1 maj_292_U13 ( .A1(maj_292_n19), .A2(maj_292_n18), .ZN(maj_292_n22)
         );
  NAND2_X1 maj_292_U12 ( .A1(u_0_2[2]), .A2(maj_292_n24), .ZN(maj_292_n20) );
  NAND2_X1 maj_292_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_292_n21) );
  NAND2_X1 maj_292_U10 ( .A1(maj_292_n21), .A2(maj_292_n20), .ZN(maj_292_n23)
         );
  XOR2_X1 maj_292_U9 ( .A(u_0_2[2]), .B(maj_292_n24), .Z(maj_292_n26) );
  XOR2_X1 maj_292_U8 ( .A(u_0_2[5]), .B(maj_292_n25), .Z(maj_292_n27) );
  XOR2_X1 maj_292_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_292_n24) );
  XOR2_X1 maj_292_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_292_n25) );
  OR2_X1 maj_292_U5 ( .A1(maj_292_n23), .A2(maj_292_n22), .ZN(maj_292_n32) );
  NAND2_X1 maj_292_U4 ( .A1(maj_292_n22), .A2(maj_292_n23), .ZN(maj_292_n34)
         );
  NAND2_X1 maj_292_U3 ( .A1(maj_292_n32), .A2(maj_292_n31), .ZN(maj_292_n33)
         );
  NAND2_X1 maj_292_U2 ( .A1(maj_292_n34), .A2(maj_292_n33), .ZN(maj_292_port_o) );
  OR2_X1 maj_293_U19 ( .A1(maj_293_n27), .A2(maj_293_n26), .ZN(maj_293_n28) );
  NAND2_X1 maj_293_U18 ( .A1(v_0_2[6]), .A2(maj_293_n28), .ZN(maj_293_n29) );
  NAND2_X1 maj_293_U17 ( .A1(maj_293_n26), .A2(maj_293_n27), .ZN(maj_293_n30)
         );
  NAND2_X1 maj_293_U16 ( .A1(maj_293_n30), .A2(maj_293_n29), .ZN(maj_293_n31)
         );
  NAND2_X1 maj_293_U15 ( .A1(v_0_2[5]), .A2(maj_293_n25), .ZN(maj_293_n18) );
  NAND2_X1 maj_293_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_293_n19) );
  NAND2_X1 maj_293_U13 ( .A1(maj_293_n19), .A2(maj_293_n18), .ZN(maj_293_n22)
         );
  NAND2_X1 maj_293_U12 ( .A1(v_0_2[2]), .A2(maj_293_n24), .ZN(maj_293_n20) );
  NAND2_X1 maj_293_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_293_n21) );
  NAND2_X1 maj_293_U10 ( .A1(maj_293_n21), .A2(maj_293_n20), .ZN(maj_293_n23)
         );
  XOR2_X1 maj_293_U9 ( .A(v_0_2[2]), .B(maj_293_n24), .Z(maj_293_n26) );
  XOR2_X1 maj_293_U8 ( .A(v_0_2[5]), .B(maj_293_n25), .Z(maj_293_n27) );
  XOR2_X1 maj_293_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_293_n24) );
  XOR2_X1 maj_293_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_293_n25) );
  OR2_X1 maj_293_U5 ( .A1(maj_293_n23), .A2(maj_293_n22), .ZN(maj_293_n32) );
  NAND2_X1 maj_293_U4 ( .A1(maj_293_n22), .A2(maj_293_n23), .ZN(maj_293_n34)
         );
  NAND2_X1 maj_293_U3 ( .A1(maj_293_n32), .A2(maj_293_n31), .ZN(maj_293_n33)
         );
  NAND2_X1 maj_293_U2 ( .A1(maj_293_n34), .A2(maj_293_n33), .ZN(maj_293_port_o) );
  OR2_X1 maj_294_U19 ( .A1(maj_294_n27), .A2(maj_294_n26), .ZN(maj_294_n28) );
  NAND2_X1 maj_294_U18 ( .A1(u_1_0[6]), .A2(maj_294_n28), .ZN(maj_294_n29) );
  NAND2_X1 maj_294_U17 ( .A1(maj_294_n26), .A2(maj_294_n27), .ZN(maj_294_n30)
         );
  NAND2_X1 maj_294_U16 ( .A1(maj_294_n30), .A2(maj_294_n29), .ZN(maj_294_n31)
         );
  NAND2_X1 maj_294_U15 ( .A1(u_1_0[5]), .A2(maj_294_n25), .ZN(maj_294_n18) );
  NAND2_X1 maj_294_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_294_n19) );
  NAND2_X1 maj_294_U13 ( .A1(maj_294_n19), .A2(maj_294_n18), .ZN(maj_294_n22)
         );
  NAND2_X1 maj_294_U12 ( .A1(u_1_0[2]), .A2(maj_294_n24), .ZN(maj_294_n20) );
  NAND2_X1 maj_294_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_294_n21) );
  NAND2_X1 maj_294_U10 ( .A1(maj_294_n21), .A2(maj_294_n20), .ZN(maj_294_n23)
         );
  XOR2_X1 maj_294_U9 ( .A(u_1_0[2]), .B(maj_294_n24), .Z(maj_294_n26) );
  XOR2_X1 maj_294_U8 ( .A(u_1_0[5]), .B(maj_294_n25), .Z(maj_294_n27) );
  XOR2_X1 maj_294_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_294_n24) );
  XOR2_X1 maj_294_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_294_n25) );
  OR2_X1 maj_294_U5 ( .A1(maj_294_n23), .A2(maj_294_n22), .ZN(maj_294_n32) );
  NAND2_X1 maj_294_U4 ( .A1(maj_294_n22), .A2(maj_294_n23), .ZN(maj_294_n34)
         );
  NAND2_X1 maj_294_U3 ( .A1(maj_294_n32), .A2(maj_294_n31), .ZN(maj_294_n33)
         );
  NAND2_X1 maj_294_U2 ( .A1(maj_294_n34), .A2(maj_294_n33), .ZN(maj_294_port_o) );
  OR2_X1 maj_295_U19 ( .A1(maj_295_n27), .A2(maj_295_n26), .ZN(maj_295_n28) );
  NAND2_X1 maj_295_U18 ( .A1(v_1_0[6]), .A2(maj_295_n28), .ZN(maj_295_n29) );
  NAND2_X1 maj_295_U17 ( .A1(maj_295_n26), .A2(maj_295_n27), .ZN(maj_295_n30)
         );
  NAND2_X1 maj_295_U16 ( .A1(maj_295_n30), .A2(maj_295_n29), .ZN(maj_295_n31)
         );
  NAND2_X1 maj_295_U15 ( .A1(v_1_0[5]), .A2(maj_295_n25), .ZN(maj_295_n18) );
  NAND2_X1 maj_295_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_295_n19) );
  NAND2_X1 maj_295_U13 ( .A1(maj_295_n19), .A2(maj_295_n18), .ZN(maj_295_n22)
         );
  NAND2_X1 maj_295_U12 ( .A1(v_1_0[2]), .A2(maj_295_n24), .ZN(maj_295_n20) );
  NAND2_X1 maj_295_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_295_n21) );
  NAND2_X1 maj_295_U10 ( .A1(maj_295_n21), .A2(maj_295_n20), .ZN(maj_295_n23)
         );
  XOR2_X1 maj_295_U9 ( .A(v_1_0[2]), .B(maj_295_n24), .Z(maj_295_n26) );
  XOR2_X1 maj_295_U8 ( .A(v_1_0[5]), .B(maj_295_n25), .Z(maj_295_n27) );
  XOR2_X1 maj_295_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_295_n24) );
  XOR2_X1 maj_295_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_295_n25) );
  OR2_X1 maj_295_U5 ( .A1(maj_295_n23), .A2(maj_295_n22), .ZN(maj_295_n32) );
  NAND2_X1 maj_295_U4 ( .A1(maj_295_n22), .A2(maj_295_n23), .ZN(maj_295_n34)
         );
  NAND2_X1 maj_295_U3 ( .A1(maj_295_n32), .A2(maj_295_n31), .ZN(maj_295_n33)
         );
  NAND2_X1 maj_295_U2 ( .A1(maj_295_n34), .A2(maj_295_n33), .ZN(maj_295_port_o) );
  OR2_X1 maj_296_U19 ( .A1(maj_296_n27), .A2(maj_296_n26), .ZN(maj_296_n28) );
  NAND2_X1 maj_296_U18 ( .A1(u_1_1[6]), .A2(maj_296_n28), .ZN(maj_296_n29) );
  NAND2_X1 maj_296_U17 ( .A1(maj_296_n26), .A2(maj_296_n27), .ZN(maj_296_n30)
         );
  NAND2_X1 maj_296_U16 ( .A1(maj_296_n30), .A2(maj_296_n29), .ZN(maj_296_n31)
         );
  NAND2_X1 maj_296_U15 ( .A1(u_1_1[5]), .A2(maj_296_n25), .ZN(maj_296_n18) );
  NAND2_X1 maj_296_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_296_n19) );
  NAND2_X1 maj_296_U13 ( .A1(maj_296_n19), .A2(maj_296_n18), .ZN(maj_296_n22)
         );
  NAND2_X1 maj_296_U12 ( .A1(u_1_1[2]), .A2(maj_296_n24), .ZN(maj_296_n20) );
  NAND2_X1 maj_296_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_296_n21) );
  NAND2_X1 maj_296_U10 ( .A1(maj_296_n21), .A2(maj_296_n20), .ZN(maj_296_n23)
         );
  XOR2_X1 maj_296_U9 ( .A(u_1_1[2]), .B(maj_296_n24), .Z(maj_296_n26) );
  XOR2_X1 maj_296_U8 ( .A(u_1_1[5]), .B(maj_296_n25), .Z(maj_296_n27) );
  XOR2_X1 maj_296_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_296_n24) );
  XOR2_X1 maj_296_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_296_n25) );
  OR2_X1 maj_296_U5 ( .A1(maj_296_n23), .A2(maj_296_n22), .ZN(maj_296_n32) );
  NAND2_X1 maj_296_U4 ( .A1(maj_296_n22), .A2(maj_296_n23), .ZN(maj_296_n34)
         );
  NAND2_X1 maj_296_U3 ( .A1(maj_296_n32), .A2(maj_296_n31), .ZN(maj_296_n33)
         );
  NAND2_X1 maj_296_U2 ( .A1(maj_296_n34), .A2(maj_296_n33), .ZN(maj_296_port_o) );
  OR2_X1 maj_297_U19 ( .A1(maj_297_n27), .A2(maj_297_n26), .ZN(maj_297_n28) );
  NAND2_X1 maj_297_U18 ( .A1(v_1_1[6]), .A2(maj_297_n28), .ZN(maj_297_n29) );
  NAND2_X1 maj_297_U17 ( .A1(maj_297_n26), .A2(maj_297_n27), .ZN(maj_297_n30)
         );
  NAND2_X1 maj_297_U16 ( .A1(maj_297_n30), .A2(maj_297_n29), .ZN(maj_297_n31)
         );
  NAND2_X1 maj_297_U15 ( .A1(v_1_1[5]), .A2(maj_297_n25), .ZN(maj_297_n18) );
  NAND2_X1 maj_297_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_297_n19) );
  NAND2_X1 maj_297_U13 ( .A1(maj_297_n19), .A2(maj_297_n18), .ZN(maj_297_n22)
         );
  NAND2_X1 maj_297_U12 ( .A1(v_1_1[2]), .A2(maj_297_n24), .ZN(maj_297_n20) );
  NAND2_X1 maj_297_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_297_n21) );
  NAND2_X1 maj_297_U10 ( .A1(maj_297_n21), .A2(maj_297_n20), .ZN(maj_297_n23)
         );
  XOR2_X1 maj_297_U9 ( .A(v_1_1[2]), .B(maj_297_n24), .Z(maj_297_n26) );
  XOR2_X1 maj_297_U8 ( .A(v_1_1[5]), .B(maj_297_n25), .Z(maj_297_n27) );
  XOR2_X1 maj_297_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_297_n24) );
  XOR2_X1 maj_297_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_297_n25) );
  OR2_X1 maj_297_U5 ( .A1(maj_297_n23), .A2(maj_297_n22), .ZN(maj_297_n32) );
  NAND2_X1 maj_297_U4 ( .A1(maj_297_n22), .A2(maj_297_n23), .ZN(maj_297_n34)
         );
  NAND2_X1 maj_297_U3 ( .A1(maj_297_n32), .A2(maj_297_n31), .ZN(maj_297_n33)
         );
  NAND2_X1 maj_297_U2 ( .A1(maj_297_n34), .A2(maj_297_n33), .ZN(maj_297_port_o) );
  OR2_X1 maj_298_U19 ( .A1(maj_298_n27), .A2(maj_298_n26), .ZN(maj_298_n28) );
  NAND2_X1 maj_298_U18 ( .A1(u_1_2[6]), .A2(maj_298_n28), .ZN(maj_298_n29) );
  NAND2_X1 maj_298_U17 ( .A1(maj_298_n26), .A2(maj_298_n27), .ZN(maj_298_n30)
         );
  NAND2_X1 maj_298_U16 ( .A1(maj_298_n30), .A2(maj_298_n29), .ZN(maj_298_n31)
         );
  NAND2_X1 maj_298_U15 ( .A1(u_1_2[5]), .A2(maj_298_n25), .ZN(maj_298_n18) );
  NAND2_X1 maj_298_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_298_n19) );
  NAND2_X1 maj_298_U13 ( .A1(maj_298_n19), .A2(maj_298_n18), .ZN(maj_298_n22)
         );
  NAND2_X1 maj_298_U12 ( .A1(u_1_2[2]), .A2(maj_298_n24), .ZN(maj_298_n20) );
  NAND2_X1 maj_298_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_298_n21) );
  NAND2_X1 maj_298_U10 ( .A1(maj_298_n21), .A2(maj_298_n20), .ZN(maj_298_n23)
         );
  XOR2_X1 maj_298_U9 ( .A(u_1_2[2]), .B(maj_298_n24), .Z(maj_298_n26) );
  XOR2_X1 maj_298_U8 ( .A(u_1_2[5]), .B(maj_298_n25), .Z(maj_298_n27) );
  XOR2_X1 maj_298_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_298_n24) );
  XOR2_X1 maj_298_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_298_n25) );
  OR2_X1 maj_298_U5 ( .A1(maj_298_n23), .A2(maj_298_n22), .ZN(maj_298_n32) );
  NAND2_X1 maj_298_U4 ( .A1(maj_298_n22), .A2(maj_298_n23), .ZN(maj_298_n34)
         );
  NAND2_X1 maj_298_U3 ( .A1(maj_298_n32), .A2(maj_298_n31), .ZN(maj_298_n33)
         );
  NAND2_X1 maj_298_U2 ( .A1(maj_298_n34), .A2(maj_298_n33), .ZN(maj_298_port_o) );
  OR2_X1 maj_299_U19 ( .A1(maj_299_n27), .A2(maj_299_n26), .ZN(maj_299_n28) );
  NAND2_X1 maj_299_U18 ( .A1(v_1_2[6]), .A2(maj_299_n28), .ZN(maj_299_n29) );
  NAND2_X1 maj_299_U17 ( .A1(maj_299_n26), .A2(maj_299_n27), .ZN(maj_299_n30)
         );
  NAND2_X1 maj_299_U16 ( .A1(maj_299_n30), .A2(maj_299_n29), .ZN(maj_299_n31)
         );
  NAND2_X1 maj_299_U15 ( .A1(v_1_2[5]), .A2(maj_299_n25), .ZN(maj_299_n18) );
  NAND2_X1 maj_299_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_299_n19) );
  NAND2_X1 maj_299_U13 ( .A1(maj_299_n19), .A2(maj_299_n18), .ZN(maj_299_n22)
         );
  NAND2_X1 maj_299_U12 ( .A1(v_1_2[2]), .A2(maj_299_n24), .ZN(maj_299_n20) );
  NAND2_X1 maj_299_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_299_n21) );
  NAND2_X1 maj_299_U10 ( .A1(maj_299_n21), .A2(maj_299_n20), .ZN(maj_299_n23)
         );
  XOR2_X1 maj_299_U9 ( .A(v_1_2[2]), .B(maj_299_n24), .Z(maj_299_n26) );
  XOR2_X1 maj_299_U8 ( .A(v_1_2[5]), .B(maj_299_n25), .Z(maj_299_n27) );
  XOR2_X1 maj_299_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_299_n24) );
  XOR2_X1 maj_299_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_299_n25) );
  OR2_X1 maj_299_U5 ( .A1(maj_299_n23), .A2(maj_299_n22), .ZN(maj_299_n32) );
  NAND2_X1 maj_299_U4 ( .A1(maj_299_n22), .A2(maj_299_n23), .ZN(maj_299_n34)
         );
  NAND2_X1 maj_299_U3 ( .A1(maj_299_n32), .A2(maj_299_n31), .ZN(maj_299_n33)
         );
  NAND2_X1 maj_299_U2 ( .A1(maj_299_n34), .A2(maj_299_n33), .ZN(maj_299_port_o) );
  OR2_X1 maj_300_U19 ( .A1(maj_300_n27), .A2(maj_300_n26), .ZN(maj_300_n28) );
  NAND2_X1 maj_300_U18 ( .A1(u_2_0[6]), .A2(maj_300_n28), .ZN(maj_300_n29) );
  NAND2_X1 maj_300_U17 ( .A1(maj_300_n26), .A2(maj_300_n27), .ZN(maj_300_n30)
         );
  NAND2_X1 maj_300_U16 ( .A1(maj_300_n30), .A2(maj_300_n29), .ZN(maj_300_n31)
         );
  NAND2_X1 maj_300_U15 ( .A1(u_2_0[5]), .A2(maj_300_n25), .ZN(maj_300_n18) );
  NAND2_X1 maj_300_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_300_n19) );
  NAND2_X1 maj_300_U13 ( .A1(maj_300_n19), .A2(maj_300_n18), .ZN(maj_300_n22)
         );
  NAND2_X1 maj_300_U12 ( .A1(u_2_0[2]), .A2(maj_300_n24), .ZN(maj_300_n20) );
  NAND2_X1 maj_300_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_300_n21) );
  NAND2_X1 maj_300_U10 ( .A1(maj_300_n21), .A2(maj_300_n20), .ZN(maj_300_n23)
         );
  XOR2_X1 maj_300_U9 ( .A(u_2_0[2]), .B(maj_300_n24), .Z(maj_300_n26) );
  XOR2_X1 maj_300_U8 ( .A(u_2_0[5]), .B(maj_300_n25), .Z(maj_300_n27) );
  XOR2_X1 maj_300_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_300_n24) );
  XOR2_X1 maj_300_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_300_n25) );
  OR2_X1 maj_300_U5 ( .A1(maj_300_n23), .A2(maj_300_n22), .ZN(maj_300_n32) );
  NAND2_X1 maj_300_U4 ( .A1(maj_300_n22), .A2(maj_300_n23), .ZN(maj_300_n34)
         );
  NAND2_X1 maj_300_U3 ( .A1(maj_300_n32), .A2(maj_300_n31), .ZN(maj_300_n33)
         );
  NAND2_X1 maj_300_U2 ( .A1(maj_300_n34), .A2(maj_300_n33), .ZN(maj_300_port_o) );
  OR2_X1 maj_301_U19 ( .A1(maj_301_n27), .A2(maj_301_n26), .ZN(maj_301_n28) );
  NAND2_X1 maj_301_U18 ( .A1(v_2_0[6]), .A2(maj_301_n28), .ZN(maj_301_n29) );
  NAND2_X1 maj_301_U17 ( .A1(maj_301_n26), .A2(maj_301_n27), .ZN(maj_301_n30)
         );
  NAND2_X1 maj_301_U16 ( .A1(maj_301_n30), .A2(maj_301_n29), .ZN(maj_301_n31)
         );
  NAND2_X1 maj_301_U15 ( .A1(v_2_0[5]), .A2(maj_301_n25), .ZN(maj_301_n18) );
  NAND2_X1 maj_301_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_301_n19) );
  NAND2_X1 maj_301_U13 ( .A1(maj_301_n19), .A2(maj_301_n18), .ZN(maj_301_n22)
         );
  NAND2_X1 maj_301_U12 ( .A1(v_2_0[2]), .A2(maj_301_n24), .ZN(maj_301_n20) );
  NAND2_X1 maj_301_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_301_n21) );
  NAND2_X1 maj_301_U10 ( .A1(maj_301_n21), .A2(maj_301_n20), .ZN(maj_301_n23)
         );
  XOR2_X1 maj_301_U9 ( .A(v_2_0[2]), .B(maj_301_n24), .Z(maj_301_n26) );
  XOR2_X1 maj_301_U8 ( .A(v_2_0[5]), .B(maj_301_n25), .Z(maj_301_n27) );
  XOR2_X1 maj_301_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_301_n24) );
  XOR2_X1 maj_301_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_301_n25) );
  OR2_X1 maj_301_U5 ( .A1(maj_301_n23), .A2(maj_301_n22), .ZN(maj_301_n32) );
  NAND2_X1 maj_301_U4 ( .A1(maj_301_n22), .A2(maj_301_n23), .ZN(maj_301_n34)
         );
  NAND2_X1 maj_301_U3 ( .A1(maj_301_n32), .A2(maj_301_n31), .ZN(maj_301_n33)
         );
  NAND2_X1 maj_301_U2 ( .A1(maj_301_n34), .A2(maj_301_n33), .ZN(maj_301_port_o) );
  OR2_X1 maj_302_U19 ( .A1(maj_302_n27), .A2(maj_302_n26), .ZN(maj_302_n28) );
  NAND2_X1 maj_302_U18 ( .A1(u_2_1[6]), .A2(maj_302_n28), .ZN(maj_302_n29) );
  NAND2_X1 maj_302_U17 ( .A1(maj_302_n26), .A2(maj_302_n27), .ZN(maj_302_n30)
         );
  NAND2_X1 maj_302_U16 ( .A1(maj_302_n30), .A2(maj_302_n29), .ZN(maj_302_n31)
         );
  NAND2_X1 maj_302_U15 ( .A1(u_2_1[5]), .A2(maj_302_n25), .ZN(maj_302_n18) );
  NAND2_X1 maj_302_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_302_n19) );
  NAND2_X1 maj_302_U13 ( .A1(maj_302_n19), .A2(maj_302_n18), .ZN(maj_302_n22)
         );
  NAND2_X1 maj_302_U12 ( .A1(u_2_1[2]), .A2(maj_302_n24), .ZN(maj_302_n20) );
  NAND2_X1 maj_302_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_302_n21) );
  NAND2_X1 maj_302_U10 ( .A1(maj_302_n21), .A2(maj_302_n20), .ZN(maj_302_n23)
         );
  XOR2_X1 maj_302_U9 ( .A(u_2_1[2]), .B(maj_302_n24), .Z(maj_302_n26) );
  XOR2_X1 maj_302_U8 ( .A(u_2_1[5]), .B(maj_302_n25), .Z(maj_302_n27) );
  XOR2_X1 maj_302_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_302_n24) );
  XOR2_X1 maj_302_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_302_n25) );
  OR2_X1 maj_302_U5 ( .A1(maj_302_n23), .A2(maj_302_n22), .ZN(maj_302_n32) );
  NAND2_X1 maj_302_U4 ( .A1(maj_302_n22), .A2(maj_302_n23), .ZN(maj_302_n34)
         );
  NAND2_X1 maj_302_U3 ( .A1(maj_302_n32), .A2(maj_302_n31), .ZN(maj_302_n33)
         );
  NAND2_X1 maj_302_U2 ( .A1(maj_302_n34), .A2(maj_302_n33), .ZN(maj_302_port_o) );
  OR2_X1 maj_303_U19 ( .A1(maj_303_n27), .A2(maj_303_n26), .ZN(maj_303_n28) );
  NAND2_X1 maj_303_U18 ( .A1(v_2_1[6]), .A2(maj_303_n28), .ZN(maj_303_n29) );
  NAND2_X1 maj_303_U17 ( .A1(maj_303_n26), .A2(maj_303_n27), .ZN(maj_303_n30)
         );
  NAND2_X1 maj_303_U16 ( .A1(maj_303_n30), .A2(maj_303_n29), .ZN(maj_303_n31)
         );
  NAND2_X1 maj_303_U15 ( .A1(v_2_1[5]), .A2(maj_303_n25), .ZN(maj_303_n18) );
  NAND2_X1 maj_303_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_303_n19) );
  NAND2_X1 maj_303_U13 ( .A1(maj_303_n19), .A2(maj_303_n18), .ZN(maj_303_n22)
         );
  NAND2_X1 maj_303_U12 ( .A1(v_2_1[2]), .A2(maj_303_n24), .ZN(maj_303_n20) );
  NAND2_X1 maj_303_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_303_n21) );
  NAND2_X1 maj_303_U10 ( .A1(maj_303_n21), .A2(maj_303_n20), .ZN(maj_303_n23)
         );
  XOR2_X1 maj_303_U9 ( .A(v_2_1[2]), .B(maj_303_n24), .Z(maj_303_n26) );
  XOR2_X1 maj_303_U8 ( .A(v_2_1[5]), .B(maj_303_n25), .Z(maj_303_n27) );
  XOR2_X1 maj_303_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_303_n24) );
  XOR2_X1 maj_303_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_303_n25) );
  OR2_X1 maj_303_U5 ( .A1(maj_303_n23), .A2(maj_303_n22), .ZN(maj_303_n32) );
  NAND2_X1 maj_303_U4 ( .A1(maj_303_n22), .A2(maj_303_n23), .ZN(maj_303_n34)
         );
  NAND2_X1 maj_303_U3 ( .A1(maj_303_n32), .A2(maj_303_n31), .ZN(maj_303_n33)
         );
  NAND2_X1 maj_303_U2 ( .A1(maj_303_n34), .A2(maj_303_n33), .ZN(maj_303_port_o) );
  OR2_X1 maj_304_U19 ( .A1(maj_304_n27), .A2(maj_304_n26), .ZN(maj_304_n28) );
  NAND2_X1 maj_304_U18 ( .A1(u_2_2[6]), .A2(maj_304_n28), .ZN(maj_304_n29) );
  NAND2_X1 maj_304_U17 ( .A1(maj_304_n26), .A2(maj_304_n27), .ZN(maj_304_n30)
         );
  NAND2_X1 maj_304_U16 ( .A1(maj_304_n30), .A2(maj_304_n29), .ZN(maj_304_n31)
         );
  NAND2_X1 maj_304_U15 ( .A1(u_2_2[5]), .A2(maj_304_n25), .ZN(maj_304_n18) );
  NAND2_X1 maj_304_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_304_n19) );
  NAND2_X1 maj_304_U13 ( .A1(maj_304_n19), .A2(maj_304_n18), .ZN(maj_304_n22)
         );
  NAND2_X1 maj_304_U12 ( .A1(u_2_2[2]), .A2(maj_304_n24), .ZN(maj_304_n20) );
  NAND2_X1 maj_304_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_304_n21) );
  NAND2_X1 maj_304_U10 ( .A1(maj_304_n21), .A2(maj_304_n20), .ZN(maj_304_n23)
         );
  XOR2_X1 maj_304_U9 ( .A(u_2_2[2]), .B(maj_304_n24), .Z(maj_304_n26) );
  XOR2_X1 maj_304_U8 ( .A(u_2_2[5]), .B(maj_304_n25), .Z(maj_304_n27) );
  XOR2_X1 maj_304_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_304_n24) );
  XOR2_X1 maj_304_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_304_n25) );
  OR2_X1 maj_304_U5 ( .A1(maj_304_n23), .A2(maj_304_n22), .ZN(maj_304_n32) );
  NAND2_X1 maj_304_U4 ( .A1(maj_304_n22), .A2(maj_304_n23), .ZN(maj_304_n34)
         );
  NAND2_X1 maj_304_U3 ( .A1(maj_304_n32), .A2(maj_304_n31), .ZN(maj_304_n33)
         );
  NAND2_X1 maj_304_U2 ( .A1(maj_304_n34), .A2(maj_304_n33), .ZN(maj_304_port_o) );
  OR2_X1 maj_305_U19 ( .A1(maj_305_n27), .A2(maj_305_n26), .ZN(maj_305_n28) );
  NAND2_X1 maj_305_U18 ( .A1(v_2_2[6]), .A2(maj_305_n28), .ZN(maj_305_n29) );
  NAND2_X1 maj_305_U17 ( .A1(maj_305_n26), .A2(maj_305_n27), .ZN(maj_305_n30)
         );
  NAND2_X1 maj_305_U16 ( .A1(maj_305_n30), .A2(maj_305_n29), .ZN(maj_305_n31)
         );
  NAND2_X1 maj_305_U15 ( .A1(v_2_2[5]), .A2(maj_305_n25), .ZN(maj_305_n18) );
  NAND2_X1 maj_305_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_305_n19) );
  NAND2_X1 maj_305_U13 ( .A1(maj_305_n19), .A2(maj_305_n18), .ZN(maj_305_n22)
         );
  NAND2_X1 maj_305_U12 ( .A1(v_2_2[2]), .A2(maj_305_n24), .ZN(maj_305_n20) );
  NAND2_X1 maj_305_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_305_n21) );
  NAND2_X1 maj_305_U10 ( .A1(maj_305_n21), .A2(maj_305_n20), .ZN(maj_305_n23)
         );
  XOR2_X1 maj_305_U9 ( .A(v_2_2[2]), .B(maj_305_n24), .Z(maj_305_n26) );
  XOR2_X1 maj_305_U8 ( .A(v_2_2[5]), .B(maj_305_n25), .Z(maj_305_n27) );
  XOR2_X1 maj_305_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_305_n24) );
  XOR2_X1 maj_305_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_305_n25) );
  OR2_X1 maj_305_U5 ( .A1(maj_305_n23), .A2(maj_305_n22), .ZN(maj_305_n32) );
  NAND2_X1 maj_305_U4 ( .A1(maj_305_n22), .A2(maj_305_n23), .ZN(maj_305_n34)
         );
  NAND2_X1 maj_305_U3 ( .A1(maj_305_n32), .A2(maj_305_n31), .ZN(maj_305_n33)
         );
  NAND2_X1 maj_305_U2 ( .A1(maj_305_n34), .A2(maj_305_n33), .ZN(maj_305_port_o) );
  OR2_X1 maj_306_U19 ( .A1(maj_306_n27), .A2(maj_306_n26), .ZN(maj_306_n28) );
  NAND2_X1 maj_306_U18 ( .A1(u_3_0[6]), .A2(maj_306_n28), .ZN(maj_306_n29) );
  NAND2_X1 maj_306_U17 ( .A1(maj_306_n26), .A2(maj_306_n27), .ZN(maj_306_n30)
         );
  NAND2_X1 maj_306_U16 ( .A1(maj_306_n30), .A2(maj_306_n29), .ZN(maj_306_n31)
         );
  NAND2_X1 maj_306_U15 ( .A1(u_3_0[5]), .A2(maj_306_n25), .ZN(maj_306_n18) );
  NAND2_X1 maj_306_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_306_n19) );
  NAND2_X1 maj_306_U13 ( .A1(maj_306_n19), .A2(maj_306_n18), .ZN(maj_306_n22)
         );
  NAND2_X1 maj_306_U12 ( .A1(u_3_0[2]), .A2(maj_306_n24), .ZN(maj_306_n20) );
  NAND2_X1 maj_306_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_306_n21) );
  NAND2_X1 maj_306_U10 ( .A1(maj_306_n21), .A2(maj_306_n20), .ZN(maj_306_n23)
         );
  XOR2_X1 maj_306_U9 ( .A(u_3_0[2]), .B(maj_306_n24), .Z(maj_306_n26) );
  XOR2_X1 maj_306_U8 ( .A(u_3_0[5]), .B(maj_306_n25), .Z(maj_306_n27) );
  XOR2_X1 maj_306_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_306_n24) );
  XOR2_X1 maj_306_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_306_n25) );
  OR2_X1 maj_306_U5 ( .A1(maj_306_n23), .A2(maj_306_n22), .ZN(maj_306_n32) );
  NAND2_X1 maj_306_U4 ( .A1(maj_306_n22), .A2(maj_306_n23), .ZN(maj_306_n34)
         );
  NAND2_X1 maj_306_U3 ( .A1(maj_306_n32), .A2(maj_306_n31), .ZN(maj_306_n33)
         );
  NAND2_X1 maj_306_U2 ( .A1(maj_306_n34), .A2(maj_306_n33), .ZN(maj_306_port_o) );
  OR2_X1 maj_307_U19 ( .A1(maj_307_n27), .A2(maj_307_n26), .ZN(maj_307_n28) );
  NAND2_X1 maj_307_U18 ( .A1(v_3_0[6]), .A2(maj_307_n28), .ZN(maj_307_n29) );
  NAND2_X1 maj_307_U17 ( .A1(maj_307_n26), .A2(maj_307_n27), .ZN(maj_307_n30)
         );
  NAND2_X1 maj_307_U16 ( .A1(maj_307_n30), .A2(maj_307_n29), .ZN(maj_307_n31)
         );
  NAND2_X1 maj_307_U15 ( .A1(v_3_0[5]), .A2(maj_307_n25), .ZN(maj_307_n18) );
  NAND2_X1 maj_307_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_307_n19) );
  NAND2_X1 maj_307_U13 ( .A1(maj_307_n19), .A2(maj_307_n18), .ZN(maj_307_n22)
         );
  NAND2_X1 maj_307_U12 ( .A1(v_3_0[2]), .A2(maj_307_n24), .ZN(maj_307_n20) );
  NAND2_X1 maj_307_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_307_n21) );
  NAND2_X1 maj_307_U10 ( .A1(maj_307_n21), .A2(maj_307_n20), .ZN(maj_307_n23)
         );
  XOR2_X1 maj_307_U9 ( .A(v_3_0[2]), .B(maj_307_n24), .Z(maj_307_n26) );
  XOR2_X1 maj_307_U8 ( .A(v_3_0[5]), .B(maj_307_n25), .Z(maj_307_n27) );
  XOR2_X1 maj_307_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_307_n24) );
  XOR2_X1 maj_307_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_307_n25) );
  OR2_X1 maj_307_U5 ( .A1(maj_307_n23), .A2(maj_307_n22), .ZN(maj_307_n32) );
  NAND2_X1 maj_307_U4 ( .A1(maj_307_n22), .A2(maj_307_n23), .ZN(maj_307_n34)
         );
  NAND2_X1 maj_307_U3 ( .A1(maj_307_n32), .A2(maj_307_n31), .ZN(maj_307_n33)
         );
  NAND2_X1 maj_307_U2 ( .A1(maj_307_n34), .A2(maj_307_n33), .ZN(maj_307_port_o) );
  OR2_X1 maj_308_U19 ( .A1(maj_308_n27), .A2(maj_308_n26), .ZN(maj_308_n28) );
  NAND2_X1 maj_308_U18 ( .A1(u_3_1[6]), .A2(maj_308_n28), .ZN(maj_308_n29) );
  NAND2_X1 maj_308_U17 ( .A1(maj_308_n26), .A2(maj_308_n27), .ZN(maj_308_n30)
         );
  NAND2_X1 maj_308_U16 ( .A1(maj_308_n30), .A2(maj_308_n29), .ZN(maj_308_n31)
         );
  NAND2_X1 maj_308_U15 ( .A1(u_3_1[5]), .A2(maj_308_n25), .ZN(maj_308_n18) );
  NAND2_X1 maj_308_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_308_n19) );
  NAND2_X1 maj_308_U13 ( .A1(maj_308_n19), .A2(maj_308_n18), .ZN(maj_308_n22)
         );
  NAND2_X1 maj_308_U12 ( .A1(u_3_1[2]), .A2(maj_308_n24), .ZN(maj_308_n20) );
  NAND2_X1 maj_308_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_308_n21) );
  NAND2_X1 maj_308_U10 ( .A1(maj_308_n21), .A2(maj_308_n20), .ZN(maj_308_n23)
         );
  XOR2_X1 maj_308_U9 ( .A(u_3_1[2]), .B(maj_308_n24), .Z(maj_308_n26) );
  XOR2_X1 maj_308_U8 ( .A(u_3_1[5]), .B(maj_308_n25), .Z(maj_308_n27) );
  XOR2_X1 maj_308_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_308_n24) );
  XOR2_X1 maj_308_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_308_n25) );
  OR2_X1 maj_308_U5 ( .A1(maj_308_n23), .A2(maj_308_n22), .ZN(maj_308_n32) );
  NAND2_X1 maj_308_U4 ( .A1(maj_308_n22), .A2(maj_308_n23), .ZN(maj_308_n34)
         );
  NAND2_X1 maj_308_U3 ( .A1(maj_308_n32), .A2(maj_308_n31), .ZN(maj_308_n33)
         );
  NAND2_X1 maj_308_U2 ( .A1(maj_308_n34), .A2(maj_308_n33), .ZN(maj_308_port_o) );
  OR2_X1 maj_309_U19 ( .A1(maj_309_n27), .A2(maj_309_n26), .ZN(maj_309_n28) );
  NAND2_X1 maj_309_U18 ( .A1(v_3_1[6]), .A2(maj_309_n28), .ZN(maj_309_n29) );
  NAND2_X1 maj_309_U17 ( .A1(maj_309_n26), .A2(maj_309_n27), .ZN(maj_309_n30)
         );
  NAND2_X1 maj_309_U16 ( .A1(maj_309_n30), .A2(maj_309_n29), .ZN(maj_309_n31)
         );
  NAND2_X1 maj_309_U15 ( .A1(v_3_1[5]), .A2(maj_309_n25), .ZN(maj_309_n18) );
  NAND2_X1 maj_309_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_309_n19) );
  NAND2_X1 maj_309_U13 ( .A1(maj_309_n19), .A2(maj_309_n18), .ZN(maj_309_n22)
         );
  NAND2_X1 maj_309_U12 ( .A1(v_3_1[2]), .A2(maj_309_n24), .ZN(maj_309_n20) );
  NAND2_X1 maj_309_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_309_n21) );
  NAND2_X1 maj_309_U10 ( .A1(maj_309_n21), .A2(maj_309_n20), .ZN(maj_309_n23)
         );
  XOR2_X1 maj_309_U9 ( .A(v_3_1[2]), .B(maj_309_n24), .Z(maj_309_n26) );
  XOR2_X1 maj_309_U8 ( .A(v_3_1[5]), .B(maj_309_n25), .Z(maj_309_n27) );
  XOR2_X1 maj_309_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_309_n24) );
  XOR2_X1 maj_309_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_309_n25) );
  OR2_X1 maj_309_U5 ( .A1(maj_309_n23), .A2(maj_309_n22), .ZN(maj_309_n32) );
  NAND2_X1 maj_309_U4 ( .A1(maj_309_n22), .A2(maj_309_n23), .ZN(maj_309_n34)
         );
  NAND2_X1 maj_309_U3 ( .A1(maj_309_n32), .A2(maj_309_n31), .ZN(maj_309_n33)
         );
  NAND2_X1 maj_309_U2 ( .A1(maj_309_n34), .A2(maj_309_n33), .ZN(maj_309_port_o) );
  OR2_X1 maj_310_U19 ( .A1(maj_310_n27), .A2(maj_310_n26), .ZN(maj_310_n28) );
  NAND2_X1 maj_310_U18 ( .A1(u_3_2[6]), .A2(maj_310_n28), .ZN(maj_310_n29) );
  NAND2_X1 maj_310_U17 ( .A1(maj_310_n26), .A2(maj_310_n27), .ZN(maj_310_n30)
         );
  NAND2_X1 maj_310_U16 ( .A1(maj_310_n30), .A2(maj_310_n29), .ZN(maj_310_n31)
         );
  NAND2_X1 maj_310_U15 ( .A1(u_3_2[5]), .A2(maj_310_n25), .ZN(maj_310_n18) );
  NAND2_X1 maj_310_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_310_n19) );
  NAND2_X1 maj_310_U13 ( .A1(maj_310_n19), .A2(maj_310_n18), .ZN(maj_310_n22)
         );
  NAND2_X1 maj_310_U12 ( .A1(u_3_2[2]), .A2(maj_310_n24), .ZN(maj_310_n20) );
  NAND2_X1 maj_310_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_310_n21) );
  NAND2_X1 maj_310_U10 ( .A1(maj_310_n21), .A2(maj_310_n20), .ZN(maj_310_n23)
         );
  XOR2_X1 maj_310_U9 ( .A(u_3_2[2]), .B(maj_310_n24), .Z(maj_310_n26) );
  XOR2_X1 maj_310_U8 ( .A(u_3_2[5]), .B(maj_310_n25), .Z(maj_310_n27) );
  XOR2_X1 maj_310_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_310_n24) );
  XOR2_X1 maj_310_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_310_n25) );
  OR2_X1 maj_310_U5 ( .A1(maj_310_n23), .A2(maj_310_n22), .ZN(maj_310_n32) );
  NAND2_X1 maj_310_U4 ( .A1(maj_310_n22), .A2(maj_310_n23), .ZN(maj_310_n34)
         );
  NAND2_X1 maj_310_U3 ( .A1(maj_310_n32), .A2(maj_310_n31), .ZN(maj_310_n33)
         );
  NAND2_X1 maj_310_U2 ( .A1(maj_310_n34), .A2(maj_310_n33), .ZN(maj_310_port_o) );
  OR2_X1 maj_311_U19 ( .A1(maj_311_n27), .A2(maj_311_n26), .ZN(maj_311_n28) );
  NAND2_X1 maj_311_U18 ( .A1(v_3_2[6]), .A2(maj_311_n28), .ZN(maj_311_n29) );
  NAND2_X1 maj_311_U17 ( .A1(maj_311_n26), .A2(maj_311_n27), .ZN(maj_311_n30)
         );
  NAND2_X1 maj_311_U16 ( .A1(maj_311_n30), .A2(maj_311_n29), .ZN(maj_311_n31)
         );
  NAND2_X1 maj_311_U15 ( .A1(v_3_2[5]), .A2(maj_311_n25), .ZN(maj_311_n18) );
  NAND2_X1 maj_311_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_311_n19) );
  NAND2_X1 maj_311_U13 ( .A1(maj_311_n19), .A2(maj_311_n18), .ZN(maj_311_n22)
         );
  NAND2_X1 maj_311_U12 ( .A1(v_3_2[2]), .A2(maj_311_n24), .ZN(maj_311_n20) );
  NAND2_X1 maj_311_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_311_n21) );
  NAND2_X1 maj_311_U10 ( .A1(maj_311_n21), .A2(maj_311_n20), .ZN(maj_311_n23)
         );
  XOR2_X1 maj_311_U9 ( .A(v_3_2[2]), .B(maj_311_n24), .Z(maj_311_n26) );
  XOR2_X1 maj_311_U8 ( .A(v_3_2[5]), .B(maj_311_n25), .Z(maj_311_n27) );
  XOR2_X1 maj_311_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_311_n24) );
  XOR2_X1 maj_311_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_311_n25) );
  OR2_X1 maj_311_U5 ( .A1(maj_311_n23), .A2(maj_311_n22), .ZN(maj_311_n32) );
  NAND2_X1 maj_311_U4 ( .A1(maj_311_n22), .A2(maj_311_n23), .ZN(maj_311_n34)
         );
  NAND2_X1 maj_311_U3 ( .A1(maj_311_n32), .A2(maj_311_n31), .ZN(maj_311_n33)
         );
  NAND2_X1 maj_311_U2 ( .A1(maj_311_n34), .A2(maj_311_n33), .ZN(maj_311_port_o) );
  OR2_X1 maj_312_U19 ( .A1(maj_312_n27), .A2(maj_312_n26), .ZN(maj_312_n28) );
  NAND2_X1 maj_312_U18 ( .A1(u_0_0[6]), .A2(maj_312_n28), .ZN(maj_312_n29) );
  NAND2_X1 maj_312_U17 ( .A1(maj_312_n26), .A2(maj_312_n27), .ZN(maj_312_n30)
         );
  NAND2_X1 maj_312_U16 ( .A1(maj_312_n30), .A2(maj_312_n29), .ZN(maj_312_n31)
         );
  NAND2_X1 maj_312_U15 ( .A1(u_0_0[5]), .A2(maj_312_n25), .ZN(maj_312_n18) );
  NAND2_X1 maj_312_U14 ( .A1(u_0_0[3]), .A2(u_0_0[4]), .ZN(maj_312_n19) );
  NAND2_X1 maj_312_U13 ( .A1(maj_312_n19), .A2(maj_312_n18), .ZN(maj_312_n22)
         );
  NAND2_X1 maj_312_U12 ( .A1(u_0_0[2]), .A2(maj_312_n24), .ZN(maj_312_n20) );
  NAND2_X1 maj_312_U11 ( .A1(u_0_0[0]), .A2(u_0_0[1]), .ZN(maj_312_n21) );
  NAND2_X1 maj_312_U10 ( .A1(maj_312_n21), .A2(maj_312_n20), .ZN(maj_312_n23)
         );
  XOR2_X1 maj_312_U9 ( .A(u_0_0[2]), .B(maj_312_n24), .Z(maj_312_n26) );
  XOR2_X1 maj_312_U8 ( .A(u_0_0[5]), .B(maj_312_n25), .Z(maj_312_n27) );
  XOR2_X1 maj_312_U7 ( .A(u_0_0[0]), .B(u_0_0[1]), .Z(maj_312_n24) );
  XOR2_X1 maj_312_U6 ( .A(u_0_0[3]), .B(u_0_0[4]), .Z(maj_312_n25) );
  OR2_X1 maj_312_U5 ( .A1(maj_312_n23), .A2(maj_312_n22), .ZN(maj_312_n32) );
  NAND2_X1 maj_312_U4 ( .A1(maj_312_n22), .A2(maj_312_n23), .ZN(maj_312_n34)
         );
  NAND2_X1 maj_312_U3 ( .A1(maj_312_n32), .A2(maj_312_n31), .ZN(maj_312_n33)
         );
  NAND2_X1 maj_312_U2 ( .A1(maj_312_n34), .A2(maj_312_n33), .ZN(maj_312_port_o) );
  OR2_X1 maj_313_U19 ( .A1(maj_313_n27), .A2(maj_313_n26), .ZN(maj_313_n28) );
  NAND2_X1 maj_313_U18 ( .A1(v_0_0[6]), .A2(maj_313_n28), .ZN(maj_313_n29) );
  NAND2_X1 maj_313_U17 ( .A1(maj_313_n26), .A2(maj_313_n27), .ZN(maj_313_n30)
         );
  NAND2_X1 maj_313_U16 ( .A1(maj_313_n30), .A2(maj_313_n29), .ZN(maj_313_n31)
         );
  NAND2_X1 maj_313_U15 ( .A1(v_0_0[5]), .A2(maj_313_n25), .ZN(maj_313_n18) );
  NAND2_X1 maj_313_U14 ( .A1(v_0_0[3]), .A2(v_0_0[4]), .ZN(maj_313_n19) );
  NAND2_X1 maj_313_U13 ( .A1(maj_313_n19), .A2(maj_313_n18), .ZN(maj_313_n22)
         );
  NAND2_X1 maj_313_U12 ( .A1(v_0_0[2]), .A2(maj_313_n24), .ZN(maj_313_n20) );
  NAND2_X1 maj_313_U11 ( .A1(v_0_0[0]), .A2(v_0_0[1]), .ZN(maj_313_n21) );
  NAND2_X1 maj_313_U10 ( .A1(maj_313_n21), .A2(maj_313_n20), .ZN(maj_313_n23)
         );
  XOR2_X1 maj_313_U9 ( .A(v_0_0[2]), .B(maj_313_n24), .Z(maj_313_n26) );
  XOR2_X1 maj_313_U8 ( .A(v_0_0[5]), .B(maj_313_n25), .Z(maj_313_n27) );
  XOR2_X1 maj_313_U7 ( .A(v_0_0[0]), .B(v_0_0[1]), .Z(maj_313_n24) );
  XOR2_X1 maj_313_U6 ( .A(v_0_0[3]), .B(v_0_0[4]), .Z(maj_313_n25) );
  OR2_X1 maj_313_U5 ( .A1(maj_313_n23), .A2(maj_313_n22), .ZN(maj_313_n32) );
  NAND2_X1 maj_313_U4 ( .A1(maj_313_n22), .A2(maj_313_n23), .ZN(maj_313_n34)
         );
  NAND2_X1 maj_313_U3 ( .A1(maj_313_n32), .A2(maj_313_n31), .ZN(maj_313_n33)
         );
  NAND2_X1 maj_313_U2 ( .A1(maj_313_n34), .A2(maj_313_n33), .ZN(maj_313_port_o) );
  OR2_X1 maj_314_U19 ( .A1(maj_314_n27), .A2(maj_314_n26), .ZN(maj_314_n28) );
  NAND2_X1 maj_314_U18 ( .A1(u_0_1[6]), .A2(maj_314_n28), .ZN(maj_314_n29) );
  NAND2_X1 maj_314_U17 ( .A1(maj_314_n26), .A2(maj_314_n27), .ZN(maj_314_n30)
         );
  NAND2_X1 maj_314_U16 ( .A1(maj_314_n30), .A2(maj_314_n29), .ZN(maj_314_n31)
         );
  NAND2_X1 maj_314_U15 ( .A1(u_0_1[5]), .A2(maj_314_n25), .ZN(maj_314_n18) );
  NAND2_X1 maj_314_U14 ( .A1(u_0_1[3]), .A2(u_0_1[4]), .ZN(maj_314_n19) );
  NAND2_X1 maj_314_U13 ( .A1(maj_314_n19), .A2(maj_314_n18), .ZN(maj_314_n22)
         );
  NAND2_X1 maj_314_U12 ( .A1(u_0_1[2]), .A2(maj_314_n24), .ZN(maj_314_n20) );
  NAND2_X1 maj_314_U11 ( .A1(u_0_1[0]), .A2(u_0_1[1]), .ZN(maj_314_n21) );
  NAND2_X1 maj_314_U10 ( .A1(maj_314_n21), .A2(maj_314_n20), .ZN(maj_314_n23)
         );
  XOR2_X1 maj_314_U9 ( .A(u_0_1[2]), .B(maj_314_n24), .Z(maj_314_n26) );
  XOR2_X1 maj_314_U8 ( .A(u_0_1[5]), .B(maj_314_n25), .Z(maj_314_n27) );
  XOR2_X1 maj_314_U7 ( .A(u_0_1[0]), .B(u_0_1[1]), .Z(maj_314_n24) );
  XOR2_X1 maj_314_U6 ( .A(u_0_1[3]), .B(u_0_1[4]), .Z(maj_314_n25) );
  OR2_X1 maj_314_U5 ( .A1(maj_314_n23), .A2(maj_314_n22), .ZN(maj_314_n32) );
  NAND2_X1 maj_314_U4 ( .A1(maj_314_n22), .A2(maj_314_n23), .ZN(maj_314_n34)
         );
  NAND2_X1 maj_314_U3 ( .A1(maj_314_n32), .A2(maj_314_n31), .ZN(maj_314_n33)
         );
  NAND2_X1 maj_314_U2 ( .A1(maj_314_n34), .A2(maj_314_n33), .ZN(maj_314_port_o) );
  OR2_X1 maj_315_U19 ( .A1(maj_315_n27), .A2(maj_315_n26), .ZN(maj_315_n28) );
  NAND2_X1 maj_315_U18 ( .A1(v_0_1[6]), .A2(maj_315_n28), .ZN(maj_315_n29) );
  NAND2_X1 maj_315_U17 ( .A1(maj_315_n26), .A2(maj_315_n27), .ZN(maj_315_n30)
         );
  NAND2_X1 maj_315_U16 ( .A1(maj_315_n30), .A2(maj_315_n29), .ZN(maj_315_n31)
         );
  NAND2_X1 maj_315_U15 ( .A1(v_0_1[5]), .A2(maj_315_n25), .ZN(maj_315_n18) );
  NAND2_X1 maj_315_U14 ( .A1(v_0_1[3]), .A2(v_0_1[4]), .ZN(maj_315_n19) );
  NAND2_X1 maj_315_U13 ( .A1(maj_315_n19), .A2(maj_315_n18), .ZN(maj_315_n22)
         );
  NAND2_X1 maj_315_U12 ( .A1(v_0_1[2]), .A2(maj_315_n24), .ZN(maj_315_n20) );
  NAND2_X1 maj_315_U11 ( .A1(v_0_1[0]), .A2(v_0_1[1]), .ZN(maj_315_n21) );
  NAND2_X1 maj_315_U10 ( .A1(maj_315_n21), .A2(maj_315_n20), .ZN(maj_315_n23)
         );
  XOR2_X1 maj_315_U9 ( .A(v_0_1[2]), .B(maj_315_n24), .Z(maj_315_n26) );
  XOR2_X1 maj_315_U8 ( .A(v_0_1[5]), .B(maj_315_n25), .Z(maj_315_n27) );
  XOR2_X1 maj_315_U7 ( .A(v_0_1[0]), .B(v_0_1[1]), .Z(maj_315_n24) );
  XOR2_X1 maj_315_U6 ( .A(v_0_1[3]), .B(v_0_1[4]), .Z(maj_315_n25) );
  OR2_X1 maj_315_U5 ( .A1(maj_315_n23), .A2(maj_315_n22), .ZN(maj_315_n32) );
  NAND2_X1 maj_315_U4 ( .A1(maj_315_n22), .A2(maj_315_n23), .ZN(maj_315_n34)
         );
  NAND2_X1 maj_315_U3 ( .A1(maj_315_n32), .A2(maj_315_n31), .ZN(maj_315_n33)
         );
  NAND2_X1 maj_315_U2 ( .A1(maj_315_n34), .A2(maj_315_n33), .ZN(maj_315_port_o) );
  OR2_X1 maj_316_U19 ( .A1(maj_316_n27), .A2(maj_316_n26), .ZN(maj_316_n28) );
  NAND2_X1 maj_316_U18 ( .A1(u_0_2[6]), .A2(maj_316_n28), .ZN(maj_316_n29) );
  NAND2_X1 maj_316_U17 ( .A1(maj_316_n26), .A2(maj_316_n27), .ZN(maj_316_n30)
         );
  NAND2_X1 maj_316_U16 ( .A1(maj_316_n30), .A2(maj_316_n29), .ZN(maj_316_n31)
         );
  NAND2_X1 maj_316_U15 ( .A1(u_0_2[5]), .A2(maj_316_n25), .ZN(maj_316_n18) );
  NAND2_X1 maj_316_U14 ( .A1(u_0_2[3]), .A2(u_0_2[4]), .ZN(maj_316_n19) );
  NAND2_X1 maj_316_U13 ( .A1(maj_316_n19), .A2(maj_316_n18), .ZN(maj_316_n22)
         );
  NAND2_X1 maj_316_U12 ( .A1(u_0_2[2]), .A2(maj_316_n24), .ZN(maj_316_n20) );
  NAND2_X1 maj_316_U11 ( .A1(u_0_2[0]), .A2(u_0_2[1]), .ZN(maj_316_n21) );
  NAND2_X1 maj_316_U10 ( .A1(maj_316_n21), .A2(maj_316_n20), .ZN(maj_316_n23)
         );
  XOR2_X1 maj_316_U9 ( .A(u_0_2[2]), .B(maj_316_n24), .Z(maj_316_n26) );
  XOR2_X1 maj_316_U8 ( .A(u_0_2[5]), .B(maj_316_n25), .Z(maj_316_n27) );
  XOR2_X1 maj_316_U7 ( .A(u_0_2[0]), .B(u_0_2[1]), .Z(maj_316_n24) );
  XOR2_X1 maj_316_U6 ( .A(u_0_2[3]), .B(u_0_2[4]), .Z(maj_316_n25) );
  OR2_X1 maj_316_U5 ( .A1(maj_316_n23), .A2(maj_316_n22), .ZN(maj_316_n32) );
  NAND2_X1 maj_316_U4 ( .A1(maj_316_n22), .A2(maj_316_n23), .ZN(maj_316_n34)
         );
  NAND2_X1 maj_316_U3 ( .A1(maj_316_n32), .A2(maj_316_n31), .ZN(maj_316_n33)
         );
  NAND2_X1 maj_316_U2 ( .A1(maj_316_n34), .A2(maj_316_n33), .ZN(maj_316_port_o) );
  OR2_X1 maj_317_U19 ( .A1(maj_317_n27), .A2(maj_317_n26), .ZN(maj_317_n28) );
  NAND2_X1 maj_317_U18 ( .A1(v_0_2[6]), .A2(maj_317_n28), .ZN(maj_317_n29) );
  NAND2_X1 maj_317_U17 ( .A1(maj_317_n26), .A2(maj_317_n27), .ZN(maj_317_n30)
         );
  NAND2_X1 maj_317_U16 ( .A1(maj_317_n30), .A2(maj_317_n29), .ZN(maj_317_n31)
         );
  NAND2_X1 maj_317_U15 ( .A1(v_0_2[5]), .A2(maj_317_n25), .ZN(maj_317_n18) );
  NAND2_X1 maj_317_U14 ( .A1(v_0_2[3]), .A2(v_0_2[4]), .ZN(maj_317_n19) );
  NAND2_X1 maj_317_U13 ( .A1(maj_317_n19), .A2(maj_317_n18), .ZN(maj_317_n22)
         );
  NAND2_X1 maj_317_U12 ( .A1(v_0_2[2]), .A2(maj_317_n24), .ZN(maj_317_n20) );
  NAND2_X1 maj_317_U11 ( .A1(v_0_2[0]), .A2(v_0_2[1]), .ZN(maj_317_n21) );
  NAND2_X1 maj_317_U10 ( .A1(maj_317_n21), .A2(maj_317_n20), .ZN(maj_317_n23)
         );
  XOR2_X1 maj_317_U9 ( .A(v_0_2[2]), .B(maj_317_n24), .Z(maj_317_n26) );
  XOR2_X1 maj_317_U8 ( .A(v_0_2[5]), .B(maj_317_n25), .Z(maj_317_n27) );
  XOR2_X1 maj_317_U7 ( .A(v_0_2[0]), .B(v_0_2[1]), .Z(maj_317_n24) );
  XOR2_X1 maj_317_U6 ( .A(v_0_2[3]), .B(v_0_2[4]), .Z(maj_317_n25) );
  OR2_X1 maj_317_U5 ( .A1(maj_317_n23), .A2(maj_317_n22), .ZN(maj_317_n32) );
  NAND2_X1 maj_317_U4 ( .A1(maj_317_n22), .A2(maj_317_n23), .ZN(maj_317_n34)
         );
  NAND2_X1 maj_317_U3 ( .A1(maj_317_n32), .A2(maj_317_n31), .ZN(maj_317_n33)
         );
  NAND2_X1 maj_317_U2 ( .A1(maj_317_n34), .A2(maj_317_n33), .ZN(maj_317_port_o) );
  OR2_X1 maj_318_U19 ( .A1(maj_318_n27), .A2(maj_318_n26), .ZN(maj_318_n28) );
  NAND2_X1 maj_318_U18 ( .A1(u_1_0[6]), .A2(maj_318_n28), .ZN(maj_318_n29) );
  NAND2_X1 maj_318_U17 ( .A1(maj_318_n26), .A2(maj_318_n27), .ZN(maj_318_n30)
         );
  NAND2_X1 maj_318_U16 ( .A1(maj_318_n30), .A2(maj_318_n29), .ZN(maj_318_n31)
         );
  NAND2_X1 maj_318_U15 ( .A1(u_1_0[5]), .A2(maj_318_n25), .ZN(maj_318_n18) );
  NAND2_X1 maj_318_U14 ( .A1(u_1_0[3]), .A2(u_1_0[4]), .ZN(maj_318_n19) );
  NAND2_X1 maj_318_U13 ( .A1(maj_318_n19), .A2(maj_318_n18), .ZN(maj_318_n22)
         );
  NAND2_X1 maj_318_U12 ( .A1(u_1_0[2]), .A2(maj_318_n24), .ZN(maj_318_n20) );
  NAND2_X1 maj_318_U11 ( .A1(u_1_0[0]), .A2(u_1_0[1]), .ZN(maj_318_n21) );
  NAND2_X1 maj_318_U10 ( .A1(maj_318_n21), .A2(maj_318_n20), .ZN(maj_318_n23)
         );
  XOR2_X1 maj_318_U9 ( .A(u_1_0[2]), .B(maj_318_n24), .Z(maj_318_n26) );
  XOR2_X1 maj_318_U8 ( .A(u_1_0[5]), .B(maj_318_n25), .Z(maj_318_n27) );
  XOR2_X1 maj_318_U7 ( .A(u_1_0[0]), .B(u_1_0[1]), .Z(maj_318_n24) );
  XOR2_X1 maj_318_U6 ( .A(u_1_0[3]), .B(u_1_0[4]), .Z(maj_318_n25) );
  OR2_X1 maj_318_U5 ( .A1(maj_318_n23), .A2(maj_318_n22), .ZN(maj_318_n32) );
  NAND2_X1 maj_318_U4 ( .A1(maj_318_n22), .A2(maj_318_n23), .ZN(maj_318_n34)
         );
  NAND2_X1 maj_318_U3 ( .A1(maj_318_n32), .A2(maj_318_n31), .ZN(maj_318_n33)
         );
  NAND2_X1 maj_318_U2 ( .A1(maj_318_n34), .A2(maj_318_n33), .ZN(maj_318_port_o) );
  OR2_X1 maj_319_U19 ( .A1(maj_319_n27), .A2(maj_319_n26), .ZN(maj_319_n28) );
  NAND2_X1 maj_319_U18 ( .A1(v_1_0[6]), .A2(maj_319_n28), .ZN(maj_319_n29) );
  NAND2_X1 maj_319_U17 ( .A1(maj_319_n26), .A2(maj_319_n27), .ZN(maj_319_n30)
         );
  NAND2_X1 maj_319_U16 ( .A1(maj_319_n30), .A2(maj_319_n29), .ZN(maj_319_n31)
         );
  NAND2_X1 maj_319_U15 ( .A1(v_1_0[5]), .A2(maj_319_n25), .ZN(maj_319_n18) );
  NAND2_X1 maj_319_U14 ( .A1(v_1_0[3]), .A2(v_1_0[4]), .ZN(maj_319_n19) );
  NAND2_X1 maj_319_U13 ( .A1(maj_319_n19), .A2(maj_319_n18), .ZN(maj_319_n22)
         );
  NAND2_X1 maj_319_U12 ( .A1(v_1_0[2]), .A2(maj_319_n24), .ZN(maj_319_n20) );
  NAND2_X1 maj_319_U11 ( .A1(v_1_0[0]), .A2(v_1_0[1]), .ZN(maj_319_n21) );
  NAND2_X1 maj_319_U10 ( .A1(maj_319_n21), .A2(maj_319_n20), .ZN(maj_319_n23)
         );
  XOR2_X1 maj_319_U9 ( .A(v_1_0[2]), .B(maj_319_n24), .Z(maj_319_n26) );
  XOR2_X1 maj_319_U8 ( .A(v_1_0[5]), .B(maj_319_n25), .Z(maj_319_n27) );
  XOR2_X1 maj_319_U7 ( .A(v_1_0[0]), .B(v_1_0[1]), .Z(maj_319_n24) );
  XOR2_X1 maj_319_U6 ( .A(v_1_0[3]), .B(v_1_0[4]), .Z(maj_319_n25) );
  OR2_X1 maj_319_U5 ( .A1(maj_319_n23), .A2(maj_319_n22), .ZN(maj_319_n32) );
  NAND2_X1 maj_319_U4 ( .A1(maj_319_n22), .A2(maj_319_n23), .ZN(maj_319_n34)
         );
  NAND2_X1 maj_319_U3 ( .A1(maj_319_n32), .A2(maj_319_n31), .ZN(maj_319_n33)
         );
  NAND2_X1 maj_319_U2 ( .A1(maj_319_n34), .A2(maj_319_n33), .ZN(maj_319_port_o) );
  OR2_X1 maj_320_U19 ( .A1(maj_320_n27), .A2(maj_320_n26), .ZN(maj_320_n28) );
  NAND2_X1 maj_320_U18 ( .A1(u_1_1[6]), .A2(maj_320_n28), .ZN(maj_320_n29) );
  NAND2_X1 maj_320_U17 ( .A1(maj_320_n26), .A2(maj_320_n27), .ZN(maj_320_n30)
         );
  NAND2_X1 maj_320_U16 ( .A1(maj_320_n30), .A2(maj_320_n29), .ZN(maj_320_n31)
         );
  NAND2_X1 maj_320_U15 ( .A1(u_1_1[5]), .A2(maj_320_n25), .ZN(maj_320_n18) );
  NAND2_X1 maj_320_U14 ( .A1(u_1_1[3]), .A2(u_1_1[4]), .ZN(maj_320_n19) );
  NAND2_X1 maj_320_U13 ( .A1(maj_320_n19), .A2(maj_320_n18), .ZN(maj_320_n22)
         );
  NAND2_X1 maj_320_U12 ( .A1(u_1_1[2]), .A2(maj_320_n24), .ZN(maj_320_n20) );
  NAND2_X1 maj_320_U11 ( .A1(u_1_1[0]), .A2(u_1_1[1]), .ZN(maj_320_n21) );
  NAND2_X1 maj_320_U10 ( .A1(maj_320_n21), .A2(maj_320_n20), .ZN(maj_320_n23)
         );
  XOR2_X1 maj_320_U9 ( .A(u_1_1[2]), .B(maj_320_n24), .Z(maj_320_n26) );
  XOR2_X1 maj_320_U8 ( .A(u_1_1[5]), .B(maj_320_n25), .Z(maj_320_n27) );
  XOR2_X1 maj_320_U7 ( .A(u_1_1[0]), .B(u_1_1[1]), .Z(maj_320_n24) );
  XOR2_X1 maj_320_U6 ( .A(u_1_1[3]), .B(u_1_1[4]), .Z(maj_320_n25) );
  OR2_X1 maj_320_U5 ( .A1(maj_320_n23), .A2(maj_320_n22), .ZN(maj_320_n32) );
  NAND2_X1 maj_320_U4 ( .A1(maj_320_n22), .A2(maj_320_n23), .ZN(maj_320_n34)
         );
  NAND2_X1 maj_320_U3 ( .A1(maj_320_n32), .A2(maj_320_n31), .ZN(maj_320_n33)
         );
  NAND2_X1 maj_320_U2 ( .A1(maj_320_n34), .A2(maj_320_n33), .ZN(maj_320_port_o) );
  OR2_X1 maj_321_U19 ( .A1(maj_321_n27), .A2(maj_321_n26), .ZN(maj_321_n28) );
  NAND2_X1 maj_321_U18 ( .A1(v_1_1[6]), .A2(maj_321_n28), .ZN(maj_321_n29) );
  NAND2_X1 maj_321_U17 ( .A1(maj_321_n26), .A2(maj_321_n27), .ZN(maj_321_n30)
         );
  NAND2_X1 maj_321_U16 ( .A1(maj_321_n30), .A2(maj_321_n29), .ZN(maj_321_n31)
         );
  NAND2_X1 maj_321_U15 ( .A1(v_1_1[5]), .A2(maj_321_n25), .ZN(maj_321_n18) );
  NAND2_X1 maj_321_U14 ( .A1(v_1_1[3]), .A2(v_1_1[4]), .ZN(maj_321_n19) );
  NAND2_X1 maj_321_U13 ( .A1(maj_321_n19), .A2(maj_321_n18), .ZN(maj_321_n22)
         );
  NAND2_X1 maj_321_U12 ( .A1(v_1_1[2]), .A2(maj_321_n24), .ZN(maj_321_n20) );
  NAND2_X1 maj_321_U11 ( .A1(v_1_1[0]), .A2(v_1_1[1]), .ZN(maj_321_n21) );
  NAND2_X1 maj_321_U10 ( .A1(maj_321_n21), .A2(maj_321_n20), .ZN(maj_321_n23)
         );
  XOR2_X1 maj_321_U9 ( .A(v_1_1[2]), .B(maj_321_n24), .Z(maj_321_n26) );
  XOR2_X1 maj_321_U8 ( .A(v_1_1[5]), .B(maj_321_n25), .Z(maj_321_n27) );
  XOR2_X1 maj_321_U7 ( .A(v_1_1[0]), .B(v_1_1[1]), .Z(maj_321_n24) );
  XOR2_X1 maj_321_U6 ( .A(v_1_1[3]), .B(v_1_1[4]), .Z(maj_321_n25) );
  OR2_X1 maj_321_U5 ( .A1(maj_321_n23), .A2(maj_321_n22), .ZN(maj_321_n32) );
  NAND2_X1 maj_321_U4 ( .A1(maj_321_n22), .A2(maj_321_n23), .ZN(maj_321_n34)
         );
  NAND2_X1 maj_321_U3 ( .A1(maj_321_n32), .A2(maj_321_n31), .ZN(maj_321_n33)
         );
  NAND2_X1 maj_321_U2 ( .A1(maj_321_n34), .A2(maj_321_n33), .ZN(maj_321_port_o) );
  OR2_X1 maj_322_U19 ( .A1(maj_322_n27), .A2(maj_322_n26), .ZN(maj_322_n28) );
  NAND2_X1 maj_322_U18 ( .A1(u_1_2[6]), .A2(maj_322_n28), .ZN(maj_322_n29) );
  NAND2_X1 maj_322_U17 ( .A1(maj_322_n26), .A2(maj_322_n27), .ZN(maj_322_n30)
         );
  NAND2_X1 maj_322_U16 ( .A1(maj_322_n30), .A2(maj_322_n29), .ZN(maj_322_n31)
         );
  NAND2_X1 maj_322_U15 ( .A1(u_1_2[5]), .A2(maj_322_n25), .ZN(maj_322_n18) );
  NAND2_X1 maj_322_U14 ( .A1(u_1_2[3]), .A2(u_1_2[4]), .ZN(maj_322_n19) );
  NAND2_X1 maj_322_U13 ( .A1(maj_322_n19), .A2(maj_322_n18), .ZN(maj_322_n22)
         );
  NAND2_X1 maj_322_U12 ( .A1(u_1_2[2]), .A2(maj_322_n24), .ZN(maj_322_n20) );
  NAND2_X1 maj_322_U11 ( .A1(u_1_2[0]), .A2(u_1_2[1]), .ZN(maj_322_n21) );
  NAND2_X1 maj_322_U10 ( .A1(maj_322_n21), .A2(maj_322_n20), .ZN(maj_322_n23)
         );
  XOR2_X1 maj_322_U9 ( .A(u_1_2[2]), .B(maj_322_n24), .Z(maj_322_n26) );
  XOR2_X1 maj_322_U8 ( .A(u_1_2[5]), .B(maj_322_n25), .Z(maj_322_n27) );
  XOR2_X1 maj_322_U7 ( .A(u_1_2[0]), .B(u_1_2[1]), .Z(maj_322_n24) );
  XOR2_X1 maj_322_U6 ( .A(u_1_2[3]), .B(u_1_2[4]), .Z(maj_322_n25) );
  OR2_X1 maj_322_U5 ( .A1(maj_322_n23), .A2(maj_322_n22), .ZN(maj_322_n32) );
  NAND2_X1 maj_322_U4 ( .A1(maj_322_n22), .A2(maj_322_n23), .ZN(maj_322_n34)
         );
  NAND2_X1 maj_322_U3 ( .A1(maj_322_n32), .A2(maj_322_n31), .ZN(maj_322_n33)
         );
  NAND2_X1 maj_322_U2 ( .A1(maj_322_n34), .A2(maj_322_n33), .ZN(maj_322_port_o) );
  OR2_X1 maj_323_U19 ( .A1(maj_323_n27), .A2(maj_323_n26), .ZN(maj_323_n28) );
  NAND2_X1 maj_323_U18 ( .A1(v_1_2[6]), .A2(maj_323_n28), .ZN(maj_323_n29) );
  NAND2_X1 maj_323_U17 ( .A1(maj_323_n26), .A2(maj_323_n27), .ZN(maj_323_n30)
         );
  NAND2_X1 maj_323_U16 ( .A1(maj_323_n30), .A2(maj_323_n29), .ZN(maj_323_n31)
         );
  NAND2_X1 maj_323_U15 ( .A1(v_1_2[5]), .A2(maj_323_n25), .ZN(maj_323_n18) );
  NAND2_X1 maj_323_U14 ( .A1(v_1_2[3]), .A2(v_1_2[4]), .ZN(maj_323_n19) );
  NAND2_X1 maj_323_U13 ( .A1(maj_323_n19), .A2(maj_323_n18), .ZN(maj_323_n22)
         );
  NAND2_X1 maj_323_U12 ( .A1(v_1_2[2]), .A2(maj_323_n24), .ZN(maj_323_n20) );
  NAND2_X1 maj_323_U11 ( .A1(v_1_2[0]), .A2(v_1_2[1]), .ZN(maj_323_n21) );
  NAND2_X1 maj_323_U10 ( .A1(maj_323_n21), .A2(maj_323_n20), .ZN(maj_323_n23)
         );
  XOR2_X1 maj_323_U9 ( .A(v_1_2[2]), .B(maj_323_n24), .Z(maj_323_n26) );
  XOR2_X1 maj_323_U8 ( .A(v_1_2[5]), .B(maj_323_n25), .Z(maj_323_n27) );
  XOR2_X1 maj_323_U7 ( .A(v_1_2[0]), .B(v_1_2[1]), .Z(maj_323_n24) );
  XOR2_X1 maj_323_U6 ( .A(v_1_2[3]), .B(v_1_2[4]), .Z(maj_323_n25) );
  OR2_X1 maj_323_U5 ( .A1(maj_323_n23), .A2(maj_323_n22), .ZN(maj_323_n32) );
  NAND2_X1 maj_323_U4 ( .A1(maj_323_n22), .A2(maj_323_n23), .ZN(maj_323_n34)
         );
  NAND2_X1 maj_323_U3 ( .A1(maj_323_n32), .A2(maj_323_n31), .ZN(maj_323_n33)
         );
  NAND2_X1 maj_323_U2 ( .A1(maj_323_n34), .A2(maj_323_n33), .ZN(maj_323_port_o) );
  OR2_X1 maj_324_U19 ( .A1(maj_324_n27), .A2(maj_324_n26), .ZN(maj_324_n28) );
  NAND2_X1 maj_324_U18 ( .A1(u_2_0[6]), .A2(maj_324_n28), .ZN(maj_324_n29) );
  NAND2_X1 maj_324_U17 ( .A1(maj_324_n26), .A2(maj_324_n27), .ZN(maj_324_n30)
         );
  NAND2_X1 maj_324_U16 ( .A1(maj_324_n30), .A2(maj_324_n29), .ZN(maj_324_n31)
         );
  NAND2_X1 maj_324_U15 ( .A1(u_2_0[5]), .A2(maj_324_n25), .ZN(maj_324_n18) );
  NAND2_X1 maj_324_U14 ( .A1(u_2_0[3]), .A2(u_2_0[4]), .ZN(maj_324_n19) );
  NAND2_X1 maj_324_U13 ( .A1(maj_324_n19), .A2(maj_324_n18), .ZN(maj_324_n22)
         );
  NAND2_X1 maj_324_U12 ( .A1(u_2_0[2]), .A2(maj_324_n24), .ZN(maj_324_n20) );
  NAND2_X1 maj_324_U11 ( .A1(u_2_0[0]), .A2(u_2_0[1]), .ZN(maj_324_n21) );
  NAND2_X1 maj_324_U10 ( .A1(maj_324_n21), .A2(maj_324_n20), .ZN(maj_324_n23)
         );
  XOR2_X1 maj_324_U9 ( .A(u_2_0[2]), .B(maj_324_n24), .Z(maj_324_n26) );
  XOR2_X1 maj_324_U8 ( .A(u_2_0[5]), .B(maj_324_n25), .Z(maj_324_n27) );
  XOR2_X1 maj_324_U7 ( .A(u_2_0[0]), .B(u_2_0[1]), .Z(maj_324_n24) );
  XOR2_X1 maj_324_U6 ( .A(u_2_0[3]), .B(u_2_0[4]), .Z(maj_324_n25) );
  OR2_X1 maj_324_U5 ( .A1(maj_324_n23), .A2(maj_324_n22), .ZN(maj_324_n32) );
  NAND2_X1 maj_324_U4 ( .A1(maj_324_n22), .A2(maj_324_n23), .ZN(maj_324_n34)
         );
  NAND2_X1 maj_324_U3 ( .A1(maj_324_n32), .A2(maj_324_n31), .ZN(maj_324_n33)
         );
  NAND2_X1 maj_324_U2 ( .A1(maj_324_n34), .A2(maj_324_n33), .ZN(maj_324_port_o) );
  OR2_X1 maj_325_U19 ( .A1(maj_325_n27), .A2(maj_325_n26), .ZN(maj_325_n28) );
  NAND2_X1 maj_325_U18 ( .A1(v_2_0[6]), .A2(maj_325_n28), .ZN(maj_325_n29) );
  NAND2_X1 maj_325_U17 ( .A1(maj_325_n26), .A2(maj_325_n27), .ZN(maj_325_n30)
         );
  NAND2_X1 maj_325_U16 ( .A1(maj_325_n30), .A2(maj_325_n29), .ZN(maj_325_n31)
         );
  NAND2_X1 maj_325_U15 ( .A1(v_2_0[5]), .A2(maj_325_n25), .ZN(maj_325_n18) );
  NAND2_X1 maj_325_U14 ( .A1(v_2_0[3]), .A2(v_2_0[4]), .ZN(maj_325_n19) );
  NAND2_X1 maj_325_U13 ( .A1(maj_325_n19), .A2(maj_325_n18), .ZN(maj_325_n22)
         );
  NAND2_X1 maj_325_U12 ( .A1(v_2_0[2]), .A2(maj_325_n24), .ZN(maj_325_n20) );
  NAND2_X1 maj_325_U11 ( .A1(v_2_0[0]), .A2(v_2_0[1]), .ZN(maj_325_n21) );
  NAND2_X1 maj_325_U10 ( .A1(maj_325_n21), .A2(maj_325_n20), .ZN(maj_325_n23)
         );
  XOR2_X1 maj_325_U9 ( .A(v_2_0[2]), .B(maj_325_n24), .Z(maj_325_n26) );
  XOR2_X1 maj_325_U8 ( .A(v_2_0[5]), .B(maj_325_n25), .Z(maj_325_n27) );
  XOR2_X1 maj_325_U7 ( .A(v_2_0[0]), .B(v_2_0[1]), .Z(maj_325_n24) );
  XOR2_X1 maj_325_U6 ( .A(v_2_0[3]), .B(v_2_0[4]), .Z(maj_325_n25) );
  OR2_X1 maj_325_U5 ( .A1(maj_325_n23), .A2(maj_325_n22), .ZN(maj_325_n32) );
  NAND2_X1 maj_325_U4 ( .A1(maj_325_n22), .A2(maj_325_n23), .ZN(maj_325_n34)
         );
  NAND2_X1 maj_325_U3 ( .A1(maj_325_n32), .A2(maj_325_n31), .ZN(maj_325_n33)
         );
  NAND2_X1 maj_325_U2 ( .A1(maj_325_n34), .A2(maj_325_n33), .ZN(maj_325_port_o) );
  OR2_X1 maj_326_U19 ( .A1(maj_326_n27), .A2(maj_326_n26), .ZN(maj_326_n28) );
  NAND2_X1 maj_326_U18 ( .A1(u_2_1[6]), .A2(maj_326_n28), .ZN(maj_326_n29) );
  NAND2_X1 maj_326_U17 ( .A1(maj_326_n26), .A2(maj_326_n27), .ZN(maj_326_n30)
         );
  NAND2_X1 maj_326_U16 ( .A1(maj_326_n30), .A2(maj_326_n29), .ZN(maj_326_n31)
         );
  NAND2_X1 maj_326_U15 ( .A1(u_2_1[5]), .A2(maj_326_n25), .ZN(maj_326_n18) );
  NAND2_X1 maj_326_U14 ( .A1(u_2_1[3]), .A2(u_2_1[4]), .ZN(maj_326_n19) );
  NAND2_X1 maj_326_U13 ( .A1(maj_326_n19), .A2(maj_326_n18), .ZN(maj_326_n22)
         );
  NAND2_X1 maj_326_U12 ( .A1(u_2_1[2]), .A2(maj_326_n24), .ZN(maj_326_n20) );
  NAND2_X1 maj_326_U11 ( .A1(u_2_1[0]), .A2(u_2_1[1]), .ZN(maj_326_n21) );
  NAND2_X1 maj_326_U10 ( .A1(maj_326_n21), .A2(maj_326_n20), .ZN(maj_326_n23)
         );
  XOR2_X1 maj_326_U9 ( .A(u_2_1[2]), .B(maj_326_n24), .Z(maj_326_n26) );
  XOR2_X1 maj_326_U8 ( .A(u_2_1[5]), .B(maj_326_n25), .Z(maj_326_n27) );
  XOR2_X1 maj_326_U7 ( .A(u_2_1[0]), .B(u_2_1[1]), .Z(maj_326_n24) );
  XOR2_X1 maj_326_U6 ( .A(u_2_1[3]), .B(u_2_1[4]), .Z(maj_326_n25) );
  OR2_X1 maj_326_U5 ( .A1(maj_326_n23), .A2(maj_326_n22), .ZN(maj_326_n32) );
  NAND2_X1 maj_326_U4 ( .A1(maj_326_n22), .A2(maj_326_n23), .ZN(maj_326_n34)
         );
  NAND2_X1 maj_326_U3 ( .A1(maj_326_n32), .A2(maj_326_n31), .ZN(maj_326_n33)
         );
  NAND2_X1 maj_326_U2 ( .A1(maj_326_n34), .A2(maj_326_n33), .ZN(maj_326_port_o) );
  OR2_X1 maj_327_U19 ( .A1(maj_327_n27), .A2(maj_327_n26), .ZN(maj_327_n28) );
  NAND2_X1 maj_327_U18 ( .A1(v_2_1[6]), .A2(maj_327_n28), .ZN(maj_327_n29) );
  NAND2_X1 maj_327_U17 ( .A1(maj_327_n26), .A2(maj_327_n27), .ZN(maj_327_n30)
         );
  NAND2_X1 maj_327_U16 ( .A1(maj_327_n30), .A2(maj_327_n29), .ZN(maj_327_n31)
         );
  NAND2_X1 maj_327_U15 ( .A1(v_2_1[5]), .A2(maj_327_n25), .ZN(maj_327_n18) );
  NAND2_X1 maj_327_U14 ( .A1(v_2_1[3]), .A2(v_2_1[4]), .ZN(maj_327_n19) );
  NAND2_X1 maj_327_U13 ( .A1(maj_327_n19), .A2(maj_327_n18), .ZN(maj_327_n22)
         );
  NAND2_X1 maj_327_U12 ( .A1(v_2_1[2]), .A2(maj_327_n24), .ZN(maj_327_n20) );
  NAND2_X1 maj_327_U11 ( .A1(v_2_1[0]), .A2(v_2_1[1]), .ZN(maj_327_n21) );
  NAND2_X1 maj_327_U10 ( .A1(maj_327_n21), .A2(maj_327_n20), .ZN(maj_327_n23)
         );
  XOR2_X1 maj_327_U9 ( .A(v_2_1[2]), .B(maj_327_n24), .Z(maj_327_n26) );
  XOR2_X1 maj_327_U8 ( .A(v_2_1[5]), .B(maj_327_n25), .Z(maj_327_n27) );
  XOR2_X1 maj_327_U7 ( .A(v_2_1[0]), .B(v_2_1[1]), .Z(maj_327_n24) );
  XOR2_X1 maj_327_U6 ( .A(v_2_1[3]), .B(v_2_1[4]), .Z(maj_327_n25) );
  OR2_X1 maj_327_U5 ( .A1(maj_327_n23), .A2(maj_327_n22), .ZN(maj_327_n32) );
  NAND2_X1 maj_327_U4 ( .A1(maj_327_n22), .A2(maj_327_n23), .ZN(maj_327_n34)
         );
  NAND2_X1 maj_327_U3 ( .A1(maj_327_n32), .A2(maj_327_n31), .ZN(maj_327_n33)
         );
  NAND2_X1 maj_327_U2 ( .A1(maj_327_n34), .A2(maj_327_n33), .ZN(maj_327_port_o) );
  OR2_X1 maj_328_U19 ( .A1(maj_328_n27), .A2(maj_328_n26), .ZN(maj_328_n28) );
  NAND2_X1 maj_328_U18 ( .A1(u_2_2[6]), .A2(maj_328_n28), .ZN(maj_328_n29) );
  NAND2_X1 maj_328_U17 ( .A1(maj_328_n26), .A2(maj_328_n27), .ZN(maj_328_n30)
         );
  NAND2_X1 maj_328_U16 ( .A1(maj_328_n30), .A2(maj_328_n29), .ZN(maj_328_n31)
         );
  NAND2_X1 maj_328_U15 ( .A1(u_2_2[5]), .A2(maj_328_n25), .ZN(maj_328_n18) );
  NAND2_X1 maj_328_U14 ( .A1(u_2_2[3]), .A2(u_2_2[4]), .ZN(maj_328_n19) );
  NAND2_X1 maj_328_U13 ( .A1(maj_328_n19), .A2(maj_328_n18), .ZN(maj_328_n22)
         );
  NAND2_X1 maj_328_U12 ( .A1(u_2_2[2]), .A2(maj_328_n24), .ZN(maj_328_n20) );
  NAND2_X1 maj_328_U11 ( .A1(u_2_2[0]), .A2(u_2_2[1]), .ZN(maj_328_n21) );
  NAND2_X1 maj_328_U10 ( .A1(maj_328_n21), .A2(maj_328_n20), .ZN(maj_328_n23)
         );
  XOR2_X1 maj_328_U9 ( .A(u_2_2[2]), .B(maj_328_n24), .Z(maj_328_n26) );
  XOR2_X1 maj_328_U8 ( .A(u_2_2[5]), .B(maj_328_n25), .Z(maj_328_n27) );
  XOR2_X1 maj_328_U7 ( .A(u_2_2[0]), .B(u_2_2[1]), .Z(maj_328_n24) );
  XOR2_X1 maj_328_U6 ( .A(u_2_2[3]), .B(u_2_2[4]), .Z(maj_328_n25) );
  OR2_X1 maj_328_U5 ( .A1(maj_328_n23), .A2(maj_328_n22), .ZN(maj_328_n32) );
  NAND2_X1 maj_328_U4 ( .A1(maj_328_n22), .A2(maj_328_n23), .ZN(maj_328_n34)
         );
  NAND2_X1 maj_328_U3 ( .A1(maj_328_n32), .A2(maj_328_n31), .ZN(maj_328_n33)
         );
  NAND2_X1 maj_328_U2 ( .A1(maj_328_n34), .A2(maj_328_n33), .ZN(maj_328_port_o) );
  OR2_X1 maj_329_U19 ( .A1(maj_329_n27), .A2(maj_329_n26), .ZN(maj_329_n28) );
  NAND2_X1 maj_329_U18 ( .A1(v_2_2[6]), .A2(maj_329_n28), .ZN(maj_329_n29) );
  NAND2_X1 maj_329_U17 ( .A1(maj_329_n26), .A2(maj_329_n27), .ZN(maj_329_n30)
         );
  NAND2_X1 maj_329_U16 ( .A1(maj_329_n30), .A2(maj_329_n29), .ZN(maj_329_n31)
         );
  NAND2_X1 maj_329_U15 ( .A1(v_2_2[5]), .A2(maj_329_n25), .ZN(maj_329_n18) );
  NAND2_X1 maj_329_U14 ( .A1(v_2_2[3]), .A2(v_2_2[4]), .ZN(maj_329_n19) );
  NAND2_X1 maj_329_U13 ( .A1(maj_329_n19), .A2(maj_329_n18), .ZN(maj_329_n22)
         );
  NAND2_X1 maj_329_U12 ( .A1(v_2_2[2]), .A2(maj_329_n24), .ZN(maj_329_n20) );
  NAND2_X1 maj_329_U11 ( .A1(v_2_2[0]), .A2(v_2_2[1]), .ZN(maj_329_n21) );
  NAND2_X1 maj_329_U10 ( .A1(maj_329_n21), .A2(maj_329_n20), .ZN(maj_329_n23)
         );
  XOR2_X1 maj_329_U9 ( .A(v_2_2[2]), .B(maj_329_n24), .Z(maj_329_n26) );
  XOR2_X1 maj_329_U8 ( .A(v_2_2[5]), .B(maj_329_n25), .Z(maj_329_n27) );
  XOR2_X1 maj_329_U7 ( .A(v_2_2[0]), .B(v_2_2[1]), .Z(maj_329_n24) );
  XOR2_X1 maj_329_U6 ( .A(v_2_2[3]), .B(v_2_2[4]), .Z(maj_329_n25) );
  OR2_X1 maj_329_U5 ( .A1(maj_329_n23), .A2(maj_329_n22), .ZN(maj_329_n32) );
  NAND2_X1 maj_329_U4 ( .A1(maj_329_n22), .A2(maj_329_n23), .ZN(maj_329_n34)
         );
  NAND2_X1 maj_329_U3 ( .A1(maj_329_n32), .A2(maj_329_n31), .ZN(maj_329_n33)
         );
  NAND2_X1 maj_329_U2 ( .A1(maj_329_n34), .A2(maj_329_n33), .ZN(maj_329_port_o) );
  OR2_X1 maj_330_U19 ( .A1(maj_330_n27), .A2(maj_330_n26), .ZN(maj_330_n28) );
  NAND2_X1 maj_330_U18 ( .A1(u_3_0[6]), .A2(maj_330_n28), .ZN(maj_330_n29) );
  NAND2_X1 maj_330_U17 ( .A1(maj_330_n26), .A2(maj_330_n27), .ZN(maj_330_n30)
         );
  NAND2_X1 maj_330_U16 ( .A1(maj_330_n30), .A2(maj_330_n29), .ZN(maj_330_n31)
         );
  NAND2_X1 maj_330_U15 ( .A1(u_3_0[5]), .A2(maj_330_n25), .ZN(maj_330_n18) );
  NAND2_X1 maj_330_U14 ( .A1(u_3_0[3]), .A2(u_3_0[4]), .ZN(maj_330_n19) );
  NAND2_X1 maj_330_U13 ( .A1(maj_330_n19), .A2(maj_330_n18), .ZN(maj_330_n22)
         );
  NAND2_X1 maj_330_U12 ( .A1(u_3_0[2]), .A2(maj_330_n24), .ZN(maj_330_n20) );
  NAND2_X1 maj_330_U11 ( .A1(u_3_0[0]), .A2(u_3_0[1]), .ZN(maj_330_n21) );
  NAND2_X1 maj_330_U10 ( .A1(maj_330_n21), .A2(maj_330_n20), .ZN(maj_330_n23)
         );
  XOR2_X1 maj_330_U9 ( .A(u_3_0[2]), .B(maj_330_n24), .Z(maj_330_n26) );
  XOR2_X1 maj_330_U8 ( .A(u_3_0[5]), .B(maj_330_n25), .Z(maj_330_n27) );
  XOR2_X1 maj_330_U7 ( .A(u_3_0[0]), .B(u_3_0[1]), .Z(maj_330_n24) );
  XOR2_X1 maj_330_U6 ( .A(u_3_0[3]), .B(u_3_0[4]), .Z(maj_330_n25) );
  OR2_X1 maj_330_U5 ( .A1(maj_330_n23), .A2(maj_330_n22), .ZN(maj_330_n32) );
  NAND2_X1 maj_330_U4 ( .A1(maj_330_n22), .A2(maj_330_n23), .ZN(maj_330_n34)
         );
  NAND2_X1 maj_330_U3 ( .A1(maj_330_n32), .A2(maj_330_n31), .ZN(maj_330_n33)
         );
  NAND2_X1 maj_330_U2 ( .A1(maj_330_n34), .A2(maj_330_n33), .ZN(maj_330_port_o) );
  OR2_X1 maj_331_U19 ( .A1(maj_331_n27), .A2(maj_331_n26), .ZN(maj_331_n28) );
  NAND2_X1 maj_331_U18 ( .A1(v_3_0[6]), .A2(maj_331_n28), .ZN(maj_331_n29) );
  NAND2_X1 maj_331_U17 ( .A1(maj_331_n26), .A2(maj_331_n27), .ZN(maj_331_n30)
         );
  NAND2_X1 maj_331_U16 ( .A1(maj_331_n30), .A2(maj_331_n29), .ZN(maj_331_n31)
         );
  NAND2_X1 maj_331_U15 ( .A1(v_3_0[5]), .A2(maj_331_n25), .ZN(maj_331_n18) );
  NAND2_X1 maj_331_U14 ( .A1(v_3_0[3]), .A2(v_3_0[4]), .ZN(maj_331_n19) );
  NAND2_X1 maj_331_U13 ( .A1(maj_331_n19), .A2(maj_331_n18), .ZN(maj_331_n22)
         );
  NAND2_X1 maj_331_U12 ( .A1(v_3_0[2]), .A2(maj_331_n24), .ZN(maj_331_n20) );
  NAND2_X1 maj_331_U11 ( .A1(v_3_0[0]), .A2(v_3_0[1]), .ZN(maj_331_n21) );
  NAND2_X1 maj_331_U10 ( .A1(maj_331_n21), .A2(maj_331_n20), .ZN(maj_331_n23)
         );
  XOR2_X1 maj_331_U9 ( .A(v_3_0[2]), .B(maj_331_n24), .Z(maj_331_n26) );
  XOR2_X1 maj_331_U8 ( .A(v_3_0[5]), .B(maj_331_n25), .Z(maj_331_n27) );
  XOR2_X1 maj_331_U7 ( .A(v_3_0[0]), .B(v_3_0[1]), .Z(maj_331_n24) );
  XOR2_X1 maj_331_U6 ( .A(v_3_0[3]), .B(v_3_0[4]), .Z(maj_331_n25) );
  OR2_X1 maj_331_U5 ( .A1(maj_331_n23), .A2(maj_331_n22), .ZN(maj_331_n32) );
  NAND2_X1 maj_331_U4 ( .A1(maj_331_n22), .A2(maj_331_n23), .ZN(maj_331_n34)
         );
  NAND2_X1 maj_331_U3 ( .A1(maj_331_n32), .A2(maj_331_n31), .ZN(maj_331_n33)
         );
  NAND2_X1 maj_331_U2 ( .A1(maj_331_n34), .A2(maj_331_n33), .ZN(maj_331_port_o) );
  OR2_X1 maj_332_U19 ( .A1(maj_332_n27), .A2(maj_332_n26), .ZN(maj_332_n28) );
  NAND2_X1 maj_332_U18 ( .A1(u_3_1[6]), .A2(maj_332_n28), .ZN(maj_332_n29) );
  NAND2_X1 maj_332_U17 ( .A1(maj_332_n26), .A2(maj_332_n27), .ZN(maj_332_n30)
         );
  NAND2_X1 maj_332_U16 ( .A1(maj_332_n30), .A2(maj_332_n29), .ZN(maj_332_n31)
         );
  NAND2_X1 maj_332_U15 ( .A1(u_3_1[5]), .A2(maj_332_n25), .ZN(maj_332_n18) );
  NAND2_X1 maj_332_U14 ( .A1(u_3_1[3]), .A2(u_3_1[4]), .ZN(maj_332_n19) );
  NAND2_X1 maj_332_U13 ( .A1(maj_332_n19), .A2(maj_332_n18), .ZN(maj_332_n22)
         );
  NAND2_X1 maj_332_U12 ( .A1(u_3_1[2]), .A2(maj_332_n24), .ZN(maj_332_n20) );
  NAND2_X1 maj_332_U11 ( .A1(u_3_1[0]), .A2(u_3_1[1]), .ZN(maj_332_n21) );
  NAND2_X1 maj_332_U10 ( .A1(maj_332_n21), .A2(maj_332_n20), .ZN(maj_332_n23)
         );
  XOR2_X1 maj_332_U9 ( .A(u_3_1[2]), .B(maj_332_n24), .Z(maj_332_n26) );
  XOR2_X1 maj_332_U8 ( .A(u_3_1[5]), .B(maj_332_n25), .Z(maj_332_n27) );
  XOR2_X1 maj_332_U7 ( .A(u_3_1[0]), .B(u_3_1[1]), .Z(maj_332_n24) );
  XOR2_X1 maj_332_U6 ( .A(u_3_1[3]), .B(u_3_1[4]), .Z(maj_332_n25) );
  OR2_X1 maj_332_U5 ( .A1(maj_332_n23), .A2(maj_332_n22), .ZN(maj_332_n32) );
  NAND2_X1 maj_332_U4 ( .A1(maj_332_n22), .A2(maj_332_n23), .ZN(maj_332_n34)
         );
  NAND2_X1 maj_332_U3 ( .A1(maj_332_n32), .A2(maj_332_n31), .ZN(maj_332_n33)
         );
  NAND2_X1 maj_332_U2 ( .A1(maj_332_n34), .A2(maj_332_n33), .ZN(maj_332_port_o) );
  OR2_X1 maj_333_U19 ( .A1(maj_333_n27), .A2(maj_333_n26), .ZN(maj_333_n28) );
  NAND2_X1 maj_333_U18 ( .A1(v_3_1[6]), .A2(maj_333_n28), .ZN(maj_333_n29) );
  NAND2_X1 maj_333_U17 ( .A1(maj_333_n26), .A2(maj_333_n27), .ZN(maj_333_n30)
         );
  NAND2_X1 maj_333_U16 ( .A1(maj_333_n30), .A2(maj_333_n29), .ZN(maj_333_n31)
         );
  NAND2_X1 maj_333_U15 ( .A1(v_3_1[5]), .A2(maj_333_n25), .ZN(maj_333_n18) );
  NAND2_X1 maj_333_U14 ( .A1(v_3_1[3]), .A2(v_3_1[4]), .ZN(maj_333_n19) );
  NAND2_X1 maj_333_U13 ( .A1(maj_333_n19), .A2(maj_333_n18), .ZN(maj_333_n22)
         );
  NAND2_X1 maj_333_U12 ( .A1(v_3_1[2]), .A2(maj_333_n24), .ZN(maj_333_n20) );
  NAND2_X1 maj_333_U11 ( .A1(v_3_1[0]), .A2(v_3_1[1]), .ZN(maj_333_n21) );
  NAND2_X1 maj_333_U10 ( .A1(maj_333_n21), .A2(maj_333_n20), .ZN(maj_333_n23)
         );
  XOR2_X1 maj_333_U9 ( .A(v_3_1[2]), .B(maj_333_n24), .Z(maj_333_n26) );
  XOR2_X1 maj_333_U8 ( .A(v_3_1[5]), .B(maj_333_n25), .Z(maj_333_n27) );
  XOR2_X1 maj_333_U7 ( .A(v_3_1[0]), .B(v_3_1[1]), .Z(maj_333_n24) );
  XOR2_X1 maj_333_U6 ( .A(v_3_1[3]), .B(v_3_1[4]), .Z(maj_333_n25) );
  OR2_X1 maj_333_U5 ( .A1(maj_333_n23), .A2(maj_333_n22), .ZN(maj_333_n32) );
  NAND2_X1 maj_333_U4 ( .A1(maj_333_n22), .A2(maj_333_n23), .ZN(maj_333_n34)
         );
  NAND2_X1 maj_333_U3 ( .A1(maj_333_n32), .A2(maj_333_n31), .ZN(maj_333_n33)
         );
  NAND2_X1 maj_333_U2 ( .A1(maj_333_n34), .A2(maj_333_n33), .ZN(maj_333_port_o) );
  OR2_X1 maj_334_U19 ( .A1(maj_334_n27), .A2(maj_334_n26), .ZN(maj_334_n28) );
  NAND2_X1 maj_334_U18 ( .A1(u_3_2[6]), .A2(maj_334_n28), .ZN(maj_334_n29) );
  NAND2_X1 maj_334_U17 ( .A1(maj_334_n26), .A2(maj_334_n27), .ZN(maj_334_n30)
         );
  NAND2_X1 maj_334_U16 ( .A1(maj_334_n30), .A2(maj_334_n29), .ZN(maj_334_n31)
         );
  NAND2_X1 maj_334_U15 ( .A1(u_3_2[5]), .A2(maj_334_n25), .ZN(maj_334_n18) );
  NAND2_X1 maj_334_U14 ( .A1(u_3_2[3]), .A2(u_3_2[4]), .ZN(maj_334_n19) );
  NAND2_X1 maj_334_U13 ( .A1(maj_334_n19), .A2(maj_334_n18), .ZN(maj_334_n22)
         );
  NAND2_X1 maj_334_U12 ( .A1(u_3_2[2]), .A2(maj_334_n24), .ZN(maj_334_n20) );
  NAND2_X1 maj_334_U11 ( .A1(u_3_2[0]), .A2(u_3_2[1]), .ZN(maj_334_n21) );
  NAND2_X1 maj_334_U10 ( .A1(maj_334_n21), .A2(maj_334_n20), .ZN(maj_334_n23)
         );
  XOR2_X1 maj_334_U9 ( .A(u_3_2[2]), .B(maj_334_n24), .Z(maj_334_n26) );
  XOR2_X1 maj_334_U8 ( .A(u_3_2[5]), .B(maj_334_n25), .Z(maj_334_n27) );
  XOR2_X1 maj_334_U7 ( .A(u_3_2[0]), .B(u_3_2[1]), .Z(maj_334_n24) );
  XOR2_X1 maj_334_U6 ( .A(u_3_2[3]), .B(u_3_2[4]), .Z(maj_334_n25) );
  OR2_X1 maj_334_U5 ( .A1(maj_334_n23), .A2(maj_334_n22), .ZN(maj_334_n32) );
  NAND2_X1 maj_334_U4 ( .A1(maj_334_n22), .A2(maj_334_n23), .ZN(maj_334_n34)
         );
  NAND2_X1 maj_334_U3 ( .A1(maj_334_n32), .A2(maj_334_n31), .ZN(maj_334_n33)
         );
  NAND2_X1 maj_334_U2 ( .A1(maj_334_n34), .A2(maj_334_n33), .ZN(maj_334_port_o) );
  OR2_X1 maj_335_U19 ( .A1(maj_335_n27), .A2(maj_335_n26), .ZN(maj_335_n28) );
  NAND2_X1 maj_335_U18 ( .A1(v_3_2[6]), .A2(maj_335_n28), .ZN(maj_335_n29) );
  NAND2_X1 maj_335_U17 ( .A1(maj_335_n26), .A2(maj_335_n27), .ZN(maj_335_n30)
         );
  NAND2_X1 maj_335_U16 ( .A1(maj_335_n30), .A2(maj_335_n29), .ZN(maj_335_n31)
         );
  NAND2_X1 maj_335_U15 ( .A1(v_3_2[5]), .A2(maj_335_n25), .ZN(maj_335_n18) );
  NAND2_X1 maj_335_U14 ( .A1(v_3_2[3]), .A2(v_3_2[4]), .ZN(maj_335_n19) );
  NAND2_X1 maj_335_U13 ( .A1(maj_335_n19), .A2(maj_335_n18), .ZN(maj_335_n22)
         );
  NAND2_X1 maj_335_U12 ( .A1(v_3_2[2]), .A2(maj_335_n24), .ZN(maj_335_n20) );
  NAND2_X1 maj_335_U11 ( .A1(v_3_2[0]), .A2(v_3_2[1]), .ZN(maj_335_n21) );
  NAND2_X1 maj_335_U10 ( .A1(maj_335_n21), .A2(maj_335_n20), .ZN(maj_335_n23)
         );
  XOR2_X1 maj_335_U9 ( .A(v_3_2[2]), .B(maj_335_n24), .Z(maj_335_n26) );
  XOR2_X1 maj_335_U8 ( .A(v_3_2[5]), .B(maj_335_n25), .Z(maj_335_n27) );
  XOR2_X1 maj_335_U7 ( .A(v_3_2[0]), .B(v_3_2[1]), .Z(maj_335_n24) );
  XOR2_X1 maj_335_U6 ( .A(v_3_2[3]), .B(v_3_2[4]), .Z(maj_335_n25) );
  OR2_X1 maj_335_U5 ( .A1(maj_335_n23), .A2(maj_335_n22), .ZN(maj_335_n32) );
  NAND2_X1 maj_335_U4 ( .A1(maj_335_n22), .A2(maj_335_n23), .ZN(maj_335_n34)
         );
  NAND2_X1 maj_335_U3 ( .A1(maj_335_n32), .A2(maj_335_n31), .ZN(maj_335_n33)
         );
  NAND2_X1 maj_335_U2 ( .A1(maj_335_n34), .A2(maj_335_n33), .ZN(maj_335_port_o) );
endmodule

