
module And_gate ( clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, 
        clock_6, reset_0, reset_1, reset_2, reset_3, reset_4, reset_5, reset_6, 
        io_i0_s0_d0, io_i0_s0_d1, io_i0_s0_d2, io_i0_s0_d3, io_i0_s0_d4, 
        io_i0_s0_d5, io_i0_s0_d6, io_i0_s1_d0, io_i0_s1_d1, io_i0_s1_d2, 
        io_i0_s1_d3, io_i0_s1_d4, io_i0_s1_d5, io_i0_s1_d6, io_i0_s2_d0, 
        io_i0_s2_d1, io_i0_s2_d2, io_i0_s2_d3, io_i0_s2_d4, io_i0_s2_d5, 
        io_i0_s2_d6, io_i1_s0_d0, io_i1_s0_d1, io_i1_s0_d2, io_i1_s0_d3, 
        io_i1_s0_d4, io_i1_s0_d5, io_i1_s0_d6, io_i1_s1_d0, io_i1_s1_d1, 
        io_i1_s1_d2, io_i1_s1_d3, io_i1_s1_d4, io_i1_s1_d5, io_i1_s1_d6, 
        io_i1_s2_d0, io_i1_s2_d1, io_i1_s2_d2, io_i1_s2_d3, io_i1_s2_d4, 
        io_i1_s2_d5, io_i1_s2_d6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, 
        p_rand_4, p_rand_5, io_o0_s0_d0, io_o0_s0_d1, io_o0_s0_d2, io_o0_s0_d3, 
        io_o0_s0_d4, io_o0_s0_d5, io_o0_s0_d6, io_o0_s1_d0, io_o0_s1_d1, 
        io_o0_s1_d2, io_o0_s1_d3, io_o0_s1_d4, io_o0_s1_d5, io_o0_s1_d6, 
        io_o0_s2_d0, io_o0_s2_d1, io_o0_s2_d2, io_o0_s2_d3, io_o0_s2_d4, 
        io_o0_s2_d5, io_o0_s2_d6 );
  input clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, clock_6, reset_0,
         reset_1, reset_2, reset_3, reset_4, reset_5, reset_6, io_i0_s0_d0,
         io_i0_s0_d1, io_i0_s0_d2, io_i0_s0_d3, io_i0_s0_d4, io_i0_s0_d5,
         io_i0_s0_d6, io_i0_s1_d0, io_i0_s1_d1, io_i0_s1_d2, io_i0_s1_d3,
         io_i0_s1_d4, io_i0_s1_d5, io_i0_s1_d6, io_i0_s2_d0, io_i0_s2_d1,
         io_i0_s2_d2, io_i0_s2_d3, io_i0_s2_d4, io_i0_s2_d5, io_i0_s2_d6,
         io_i1_s0_d0, io_i1_s0_d1, io_i1_s0_d2, io_i1_s0_d3, io_i1_s0_d4,
         io_i1_s0_d5, io_i1_s0_d6, io_i1_s1_d0, io_i1_s1_d1, io_i1_s1_d2,
         io_i1_s1_d3, io_i1_s1_d4, io_i1_s1_d5, io_i1_s1_d6, io_i1_s2_d0,
         io_i1_s2_d1, io_i1_s2_d2, io_i1_s2_d3, io_i1_s2_d4, io_i1_s2_d5,
         io_i1_s2_d6, p_rand_0, p_rand_1, p_rand_2, p_rand_3, p_rand_4,
         p_rand_5;
  output io_o0_s0_d0, io_o0_s0_d1, io_o0_s0_d2, io_o0_s0_d3, io_o0_s0_d4,
         io_o0_s0_d5, io_o0_s0_d6, io_o0_s1_d0, io_o0_s1_d1, io_o0_s1_d2,
         io_o0_s1_d3, io_o0_s1_d4, io_o0_s1_d5, io_o0_s1_d6, io_o0_s2_d0,
         io_o0_s2_d1, io_o0_s2_d2, io_o0_s2_d3, io_o0_s2_d4, io_o0_s2_d5,
         io_o0_s2_d6;
  wire   n_xor_module_1_res, n_xor_module_2_res, n_xor_module_3_res,
         n_xor_module_4_res, n_xor_module_5_res, n_xor_module_6_res,
         n_xor_module_7_res, n_xor_module_8_res, n_xor_module_9_res,
         n_xor_module_10_res, n_xor_module_11_res, n_xor_module_12_res,
         n_xor_module_13_res, n_xor_module_14_res, n_xor_module_15_res,
         n_xor_module_16_res, n_xor_module_17_res, n_xor_module_18_res,
         n_xor_module_19_res, n_xor_module_20_res, n_xor_module_21_res,
         n_xor_module_22_res, n_xor_module_23_res, n_xor_module_24_res,
         n_xor_module_25_res, n_xor_module_26_res, n_xor_module_27_res,
         n_xor_module_28_res, n_xor_module_29_res, n_xor_module_30_res,
         n_xor_module_31_res, n_xor_module_32_res, n_xor_module_33_res,
         n_xor_module_34_res, n_xor_module_35_res, n_xor_module_36_res,
         n_xor_module_37_res, n_xor_module_38_res, n_xor_module_39_res,
         n_xor_module_40_res, n_xor_module_41_res, n_xor_module_42_res,
         n_majority7_module_0_res, n_reg_module_1_res,
         n_majority7_module_1_res, n_reg_module_2_res,
         n_majority7_module_2_res, n_reg_module_3_res,
         n_majority7_module_3_res, n_reg_module_4_res,
         n_majority7_module_4_res, n_reg_module_5_res,
         n_majority7_module_5_res, n_reg_module_6_res,
         n_majority7_module_6_res, n_reg_module_7_res,
         n_majority7_module_7_res, n_reg_module_8_res,
         n_majority7_module_8_res, n_reg_module_9_res,
         n_majority7_module_9_res, n_reg_module_10_res,
         n_majority7_module_10_res, n_reg_module_11_res,
         n_majority7_module_11_res, n_reg_module_12_res,
         n_majority7_module_12_res, n_reg_module_13_res,
         n_majority7_module_13_res, n_reg_module_14_res,
         n_majority7_module_14_res, n_reg_module_15_res,
         n_majority7_module_15_res, n_reg_module_16_res,
         n_majority7_module_16_res, n_reg_module_17_res,
         n_majority7_module_17_res, n_reg_module_18_res,
         n_majority7_module_18_res, n_reg_module_19_res,
         n_majority7_module_19_res, n_reg_module_20_res,
         n_majority7_module_20_res, n_reg_module_21_res,
         n_majority7_module_21_res, n_reg_module_22_res,
         n_majority7_module_22_res, n_reg_module_23_res,
         n_majority7_module_23_res, n_reg_module_24_res,
         n_majority7_module_24_res, n_reg_module_25_res,
         n_majority7_module_25_res, n_reg_module_26_res,
         n_majority7_module_26_res, n_reg_module_27_res,
         n_majority7_module_27_res, n_reg_module_28_res,
         n_majority7_module_28_res, n_reg_module_29_res,
         n_majority7_module_29_res, n_reg_module_30_res,
         n_majority7_module_30_res, n_reg_module_31_res,
         n_majority7_module_31_res, n_reg_module_32_res,
         n_majority7_module_32_res, n_reg_module_33_res,
         n_majority7_module_33_res, n_reg_module_34_res,
         n_majority7_module_34_res, n_reg_module_35_res,
         n_majority7_module_35_res, n_reg_module_36_res,
         n_majority7_module_36_res, n_reg_module_37_res,
         n_majority7_module_37_res, n_reg_module_38_res,
         n_majority7_module_38_res, n_reg_module_39_res,
         n_majority7_module_39_res, n_reg_module_40_res,
         n_majority7_module_40_res, n_reg_module_41_res,
         n_majority7_module_41_res, n_reg_module_42_res,
         n_majority7_module_42_res, n_reg_module_43_res,
         n_majority7_module_43_res, n_reg_module_44_res,
         n_majority7_module_44_res, n_reg_module_45_res,
         n_majority7_module_45_res, n_reg_module_46_res,
         n_majority7_module_46_res, n_reg_module_47_res,
         n_majority7_module_47_res, n_reg_module_48_res,
         n_majority7_module_48_res, n_reg_module_49_res,
         n_majority7_module_49_res, n_reg_module_50_res,
         n_majority7_module_50_res, n_reg_module_51_res,
         n_majority7_module_51_res, n_reg_module_52_res,
         n_majority7_module_52_res, n_reg_module_53_res,
         n_majority7_module_53_res, n_reg_module_54_res,
         n_majority7_module_54_res, n_reg_module_55_res,
         n_majority7_module_55_res, n_reg_module_56_res,
         n_majority7_module_56_res, n_reg_module_57_res,
         n_majority7_module_57_res, n_reg_module_58_res,
         n_majority7_module_58_res, n_reg_module_59_res,
         n_majority7_module_59_res, n_reg_module_60_res,
         n_majority7_module_60_res, n_reg_module_61_res,
         n_majority7_module_61_res, n_reg_module_62_res,
         n_majority7_module_62_res, n_reg_module_63_res, n_and_module_1_res,
         n_reg_module_64_res, n_and_module_2_res, n_xor_module_43_res,
         n_reg_module_65_res, n_and_module_3_res, n_xor_module_44_res,
         n_reg_module_66_res, n_and_module_4_res, n_xor_module_45_res,
         n_reg_module_67_res, n_and_module_5_res, n_reg_module_68_res,
         n_and_module_6_res, n_xor_module_46_res, n_reg_module_69_res,
         n_and_module_7_res, n_xor_module_47_res, n_reg_module_70_res,
         n_and_module_8_res, n_xor_module_48_res, n_reg_module_71_res,
         n_and_module_9_res, n_reg_module_72_res, n_and_module_10_res,
         n_reg_module_73_res, n_and_module_11_res, n_xor_module_49_res,
         n_reg_module_74_res, n_and_module_12_res, n_xor_module_50_res,
         n_reg_module_75_res, n_and_module_13_res, n_xor_module_51_res,
         n_reg_module_76_res, n_and_module_14_res, n_reg_module_77_res,
         n_and_module_15_res, n_xor_module_52_res, n_reg_module_78_res,
         n_and_module_16_res, n_xor_module_53_res, n_reg_module_79_res,
         n_and_module_17_res, n_xor_module_54_res, n_reg_module_80_res,
         n_and_module_18_res, n_reg_module_81_res, n_and_module_19_res,
         n_reg_module_82_res, n_and_module_20_res, n_xor_module_55_res,
         n_reg_module_83_res, n_and_module_21_res, n_xor_module_56_res,
         n_reg_module_84_res, n_and_module_22_res, n_xor_module_57_res,
         n_reg_module_85_res, n_and_module_23_res, n_reg_module_86_res,
         n_and_module_24_res, n_xor_module_58_res, n_reg_module_87_res,
         n_and_module_25_res, n_xor_module_59_res, n_reg_module_88_res,
         n_and_module_26_res, n_xor_module_60_res, n_reg_module_89_res,
         n_and_module_27_res, n_reg_module_90_res, n_and_module_28_res,
         n_reg_module_91_res, n_and_module_29_res, n_xor_module_61_res,
         n_reg_module_92_res, n_and_module_30_res, n_xor_module_62_res,
         n_reg_module_93_res, n_and_module_31_res, n_xor_module_63_res,
         n_reg_module_94_res, n_and_module_32_res, n_reg_module_95_res,
         n_and_module_33_res, n_xor_module_64_res, n_reg_module_96_res,
         n_and_module_34_res, n_xor_module_65_res, n_reg_module_97_res,
         n_and_module_35_res, n_xor_module_66_res, n_reg_module_98_res,
         n_and_module_36_res, n_reg_module_99_res, n_and_module_37_res,
         n_reg_module_100_res, n_and_module_38_res, n_xor_module_67_res,
         n_reg_module_101_res, n_and_module_39_res, n_xor_module_68_res,
         n_reg_module_102_res, n_and_module_40_res, n_xor_module_69_res,
         n_reg_module_103_res, n_and_module_41_res, n_reg_module_104_res,
         n_and_module_42_res, n_xor_module_70_res, n_reg_module_105_res,
         n_and_module_43_res, n_xor_module_71_res, n_reg_module_106_res,
         n_and_module_44_res, n_xor_module_72_res, n_reg_module_107_res,
         n_and_module_45_res, n_reg_module_108_res, n_and_module_46_res,
         n_reg_module_109_res, n_and_module_47_res, n_xor_module_73_res,
         n_reg_module_110_res, n_and_module_48_res, n_xor_module_74_res,
         n_reg_module_111_res, n_and_module_49_res, n_xor_module_75_res,
         n_reg_module_112_res, n_and_module_50_res, n_reg_module_113_res,
         n_and_module_51_res, n_xor_module_76_res, n_reg_module_114_res,
         n_and_module_52_res, n_xor_module_77_res, n_reg_module_115_res,
         n_and_module_53_res, n_xor_module_78_res, n_reg_module_116_res,
         n_and_module_54_res, n_reg_module_117_res, n_and_module_55_res,
         n_reg_module_118_res, n_and_module_56_res, n_xor_module_79_res,
         n_reg_module_119_res, n_and_module_57_res, n_xor_module_80_res,
         n_reg_module_120_res, n_and_module_58_res, n_xor_module_81_res,
         n_reg_module_121_res, n_and_module_59_res, n_reg_module_122_res,
         n_and_module_60_res, n_xor_module_82_res, n_reg_module_123_res,
         n_and_module_61_res, n_xor_module_83_res, n_reg_module_124_res,
         n_and_module_62_res, n_xor_module_84_res, n_reg_module_125_res,
         n_and_module_63_res, n_reg_module_126_res, n_xor_module_85_res,
         n_xor_module_87_res, n_xor_module_89_res, n_xor_module_91_res,
         n_xor_module_93_res, n_xor_module_95_res, n_xor_module_97_res,
         n_xor_module_99_res, n_xor_module_101_res, n_xor_module_103_res,
         n_xor_module_105_res, n_xor_module_107_res, n_xor_module_109_res,
         n_xor_module_111_res, n_xor_module_113_res, n_xor_module_115_res,
         n_xor_module_117_res, n_xor_module_119_res, n_xor_module_121_res,
         n_xor_module_123_res, n_xor_module_125_res, n_majority7_module_0_n7,
         n_majority7_module_0_n6, n_majority7_module_0_n5,
         n_majority7_module_0_n4, n_majority7_module_0_n3,
         n_majority7_module_0_n2, n_majority7_module_0_n1,
         n_majority7_module_0__and_module_10_res,
         n_majority7_module_0__or_module_11_res,
         n_majority7_module_0__and_module_9_res,
         n_majority7_module_0__or_module_10_res,
         n_majority7_module_0__or_module_9_res,
         n_majority7_module_0__and_module_8_res,
         n_majority7_module_0__or_module_8_res,
         n_majority7_module_0__and_module_7_res,
         n_majority7_module_0__or_module_7_res,
         n_majority7_module_0__or_module_6_res,
         n_majority7_module_0__and_module_6_res,
         n_majority7_module_0__or_module_5_res,
         n_majority7_module_0__and_module_5_res,
         n_majority7_module_0__or_module_4_res,
         n_majority7_module_0__and_module_4_res,
         n_majority7_module_0__or_module_3_res,
         n_majority7_module_0__and_module_3_res,
         n_majority7_module_0__or_module_2_res,
         n_majority7_module_0__and_module_2_res,
         n_majority7_module_0__or_module_1_res,
         n_majority7_module_0__and_module_1_res, n_majority7_module_1_n7,
         n_majority7_module_1_n6, n_majority7_module_1_n5,
         n_majority7_module_1_n4, n_majority7_module_1_n3,
         n_majority7_module_1_n2, n_majority7_module_1_n1,
         n_majority7_module_1__and_module_10_res,
         n_majority7_module_1__or_module_11_res,
         n_majority7_module_1__and_module_9_res,
         n_majority7_module_1__or_module_10_res,
         n_majority7_module_1__or_module_9_res,
         n_majority7_module_1__and_module_8_res,
         n_majority7_module_1__or_module_8_res,
         n_majority7_module_1__and_module_7_res,
         n_majority7_module_1__or_module_7_res,
         n_majority7_module_1__or_module_6_res,
         n_majority7_module_1__and_module_6_res,
         n_majority7_module_1__or_module_5_res,
         n_majority7_module_1__and_module_5_res,
         n_majority7_module_1__or_module_4_res,
         n_majority7_module_1__and_module_4_res,
         n_majority7_module_1__or_module_3_res,
         n_majority7_module_1__and_module_3_res,
         n_majority7_module_1__or_module_2_res,
         n_majority7_module_1__and_module_2_res,
         n_majority7_module_1__or_module_1_res,
         n_majority7_module_1__and_module_1_res, n_majority7_module_2_n7,
         n_majority7_module_2_n6, n_majority7_module_2_n5,
         n_majority7_module_2_n4, n_majority7_module_2_n3,
         n_majority7_module_2_n2, n_majority7_module_2_n1,
         n_majority7_module_2__and_module_10_res,
         n_majority7_module_2__or_module_11_res,
         n_majority7_module_2__and_module_9_res,
         n_majority7_module_2__or_module_10_res,
         n_majority7_module_2__or_module_9_res,
         n_majority7_module_2__and_module_8_res,
         n_majority7_module_2__or_module_8_res,
         n_majority7_module_2__and_module_7_res,
         n_majority7_module_2__or_module_7_res,
         n_majority7_module_2__or_module_6_res,
         n_majority7_module_2__and_module_6_res,
         n_majority7_module_2__or_module_5_res,
         n_majority7_module_2__and_module_5_res,
         n_majority7_module_2__or_module_4_res,
         n_majority7_module_2__and_module_4_res,
         n_majority7_module_2__or_module_3_res,
         n_majority7_module_2__and_module_3_res,
         n_majority7_module_2__or_module_2_res,
         n_majority7_module_2__and_module_2_res,
         n_majority7_module_2__or_module_1_res,
         n_majority7_module_2__and_module_1_res, n_majority7_module_3_n7,
         n_majority7_module_3_n6, n_majority7_module_3_n5,
         n_majority7_module_3_n4, n_majority7_module_3_n3,
         n_majority7_module_3_n2, n_majority7_module_3_n1,
         n_majority7_module_3__and_module_10_res,
         n_majority7_module_3__or_module_11_res,
         n_majority7_module_3__and_module_9_res,
         n_majority7_module_3__or_module_10_res,
         n_majority7_module_3__or_module_9_res,
         n_majority7_module_3__and_module_8_res,
         n_majority7_module_3__or_module_8_res,
         n_majority7_module_3__and_module_7_res,
         n_majority7_module_3__or_module_7_res,
         n_majority7_module_3__or_module_6_res,
         n_majority7_module_3__and_module_6_res,
         n_majority7_module_3__or_module_5_res,
         n_majority7_module_3__and_module_5_res,
         n_majority7_module_3__or_module_4_res,
         n_majority7_module_3__and_module_4_res,
         n_majority7_module_3__or_module_3_res,
         n_majority7_module_3__and_module_3_res,
         n_majority7_module_3__or_module_2_res,
         n_majority7_module_3__and_module_2_res,
         n_majority7_module_3__or_module_1_res,
         n_majority7_module_3__and_module_1_res, n_majority7_module_4_n7,
         n_majority7_module_4_n6, n_majority7_module_4_n5,
         n_majority7_module_4_n4, n_majority7_module_4_n3,
         n_majority7_module_4_n2, n_majority7_module_4_n1,
         n_majority7_module_4__and_module_10_res,
         n_majority7_module_4__or_module_11_res,
         n_majority7_module_4__and_module_9_res,
         n_majority7_module_4__or_module_10_res,
         n_majority7_module_4__or_module_9_res,
         n_majority7_module_4__and_module_8_res,
         n_majority7_module_4__or_module_8_res,
         n_majority7_module_4__and_module_7_res,
         n_majority7_module_4__or_module_7_res,
         n_majority7_module_4__or_module_6_res,
         n_majority7_module_4__and_module_6_res,
         n_majority7_module_4__or_module_5_res,
         n_majority7_module_4__and_module_5_res,
         n_majority7_module_4__or_module_4_res,
         n_majority7_module_4__and_module_4_res,
         n_majority7_module_4__or_module_3_res,
         n_majority7_module_4__and_module_3_res,
         n_majority7_module_4__or_module_2_res,
         n_majority7_module_4__and_module_2_res,
         n_majority7_module_4__or_module_1_res,
         n_majority7_module_4__and_module_1_res, n_majority7_module_5_n7,
         n_majority7_module_5_n6, n_majority7_module_5_n5,
         n_majority7_module_5_n4, n_majority7_module_5_n3,
         n_majority7_module_5_n2, n_majority7_module_5_n1,
         n_majority7_module_5__and_module_10_res,
         n_majority7_module_5__or_module_11_res,
         n_majority7_module_5__and_module_9_res,
         n_majority7_module_5__or_module_10_res,
         n_majority7_module_5__or_module_9_res,
         n_majority7_module_5__and_module_8_res,
         n_majority7_module_5__or_module_8_res,
         n_majority7_module_5__and_module_7_res,
         n_majority7_module_5__or_module_7_res,
         n_majority7_module_5__or_module_6_res,
         n_majority7_module_5__and_module_6_res,
         n_majority7_module_5__or_module_5_res,
         n_majority7_module_5__and_module_5_res,
         n_majority7_module_5__or_module_4_res,
         n_majority7_module_5__and_module_4_res,
         n_majority7_module_5__or_module_3_res,
         n_majority7_module_5__and_module_3_res,
         n_majority7_module_5__or_module_2_res,
         n_majority7_module_5__and_module_2_res,
         n_majority7_module_5__or_module_1_res,
         n_majority7_module_5__and_module_1_res, n_majority7_module_6_n7,
         n_majority7_module_6_n6, n_majority7_module_6_n5,
         n_majority7_module_6_n4, n_majority7_module_6_n3,
         n_majority7_module_6_n2, n_majority7_module_6_n1,
         n_majority7_module_6__and_module_10_res,
         n_majority7_module_6__or_module_11_res,
         n_majority7_module_6__and_module_9_res,
         n_majority7_module_6__or_module_10_res,
         n_majority7_module_6__or_module_9_res,
         n_majority7_module_6__and_module_8_res,
         n_majority7_module_6__or_module_8_res,
         n_majority7_module_6__and_module_7_res,
         n_majority7_module_6__or_module_7_res,
         n_majority7_module_6__or_module_6_res,
         n_majority7_module_6__and_module_6_res,
         n_majority7_module_6__or_module_5_res,
         n_majority7_module_6__and_module_5_res,
         n_majority7_module_6__or_module_4_res,
         n_majority7_module_6__and_module_4_res,
         n_majority7_module_6__or_module_3_res,
         n_majority7_module_6__and_module_3_res,
         n_majority7_module_6__or_module_2_res,
         n_majority7_module_6__and_module_2_res,
         n_majority7_module_6__or_module_1_res,
         n_majority7_module_6__and_module_1_res, n_majority7_module_7_n7,
         n_majority7_module_7_n6, n_majority7_module_7_n5,
         n_majority7_module_7_n4, n_majority7_module_7_n3,
         n_majority7_module_7_n2, n_majority7_module_7_n1,
         n_majority7_module_7__and_module_10_res,
         n_majority7_module_7__or_module_11_res,
         n_majority7_module_7__and_module_9_res,
         n_majority7_module_7__or_module_10_res,
         n_majority7_module_7__or_module_9_res,
         n_majority7_module_7__and_module_8_res,
         n_majority7_module_7__or_module_8_res,
         n_majority7_module_7__and_module_7_res,
         n_majority7_module_7__or_module_7_res,
         n_majority7_module_7__or_module_6_res,
         n_majority7_module_7__and_module_6_res,
         n_majority7_module_7__or_module_5_res,
         n_majority7_module_7__and_module_5_res,
         n_majority7_module_7__or_module_4_res,
         n_majority7_module_7__and_module_4_res,
         n_majority7_module_7__or_module_3_res,
         n_majority7_module_7__and_module_3_res,
         n_majority7_module_7__or_module_2_res,
         n_majority7_module_7__and_module_2_res,
         n_majority7_module_7__or_module_1_res,
         n_majority7_module_7__and_module_1_res, n_majority7_module_8_n7,
         n_majority7_module_8_n6, n_majority7_module_8_n5,
         n_majority7_module_8_n4, n_majority7_module_8_n3,
         n_majority7_module_8_n2, n_majority7_module_8_n1,
         n_majority7_module_8__and_module_10_res,
         n_majority7_module_8__or_module_11_res,
         n_majority7_module_8__and_module_9_res,
         n_majority7_module_8__or_module_10_res,
         n_majority7_module_8__or_module_9_res,
         n_majority7_module_8__and_module_8_res,
         n_majority7_module_8__or_module_8_res,
         n_majority7_module_8__and_module_7_res,
         n_majority7_module_8__or_module_7_res,
         n_majority7_module_8__or_module_6_res,
         n_majority7_module_8__and_module_6_res,
         n_majority7_module_8__or_module_5_res,
         n_majority7_module_8__and_module_5_res,
         n_majority7_module_8__or_module_4_res,
         n_majority7_module_8__and_module_4_res,
         n_majority7_module_8__or_module_3_res,
         n_majority7_module_8__and_module_3_res,
         n_majority7_module_8__or_module_2_res,
         n_majority7_module_8__and_module_2_res,
         n_majority7_module_8__or_module_1_res,
         n_majority7_module_8__and_module_1_res, n_majority7_module_9_n7,
         n_majority7_module_9_n6, n_majority7_module_9_n5,
         n_majority7_module_9_n4, n_majority7_module_9_n3,
         n_majority7_module_9_n2, n_majority7_module_9_n1,
         n_majority7_module_9__and_module_10_res,
         n_majority7_module_9__or_module_11_res,
         n_majority7_module_9__and_module_9_res,
         n_majority7_module_9__or_module_10_res,
         n_majority7_module_9__or_module_9_res,
         n_majority7_module_9__and_module_8_res,
         n_majority7_module_9__or_module_8_res,
         n_majority7_module_9__and_module_7_res,
         n_majority7_module_9__or_module_7_res,
         n_majority7_module_9__or_module_6_res,
         n_majority7_module_9__and_module_6_res,
         n_majority7_module_9__or_module_5_res,
         n_majority7_module_9__and_module_5_res,
         n_majority7_module_9__or_module_4_res,
         n_majority7_module_9__and_module_4_res,
         n_majority7_module_9__or_module_3_res,
         n_majority7_module_9__and_module_3_res,
         n_majority7_module_9__or_module_2_res,
         n_majority7_module_9__and_module_2_res,
         n_majority7_module_9__or_module_1_res,
         n_majority7_module_9__and_module_1_res, n_majority7_module_10_n7,
         n_majority7_module_10_n6, n_majority7_module_10_n5,
         n_majority7_module_10_n4, n_majority7_module_10_n3,
         n_majority7_module_10_n2, n_majority7_module_10_n1,
         n_majority7_module_10__and_module_10_res,
         n_majority7_module_10__or_module_11_res,
         n_majority7_module_10__and_module_9_res,
         n_majority7_module_10__or_module_10_res,
         n_majority7_module_10__or_module_9_res,
         n_majority7_module_10__and_module_8_res,
         n_majority7_module_10__or_module_8_res,
         n_majority7_module_10__and_module_7_res,
         n_majority7_module_10__or_module_7_res,
         n_majority7_module_10__or_module_6_res,
         n_majority7_module_10__and_module_6_res,
         n_majority7_module_10__or_module_5_res,
         n_majority7_module_10__and_module_5_res,
         n_majority7_module_10__or_module_4_res,
         n_majority7_module_10__and_module_4_res,
         n_majority7_module_10__or_module_3_res,
         n_majority7_module_10__and_module_3_res,
         n_majority7_module_10__or_module_2_res,
         n_majority7_module_10__and_module_2_res,
         n_majority7_module_10__or_module_1_res,
         n_majority7_module_10__and_module_1_res, n_majority7_module_11_n7,
         n_majority7_module_11_n6, n_majority7_module_11_n5,
         n_majority7_module_11_n4, n_majority7_module_11_n3,
         n_majority7_module_11_n2, n_majority7_module_11_n1,
         n_majority7_module_11__and_module_10_res,
         n_majority7_module_11__or_module_11_res,
         n_majority7_module_11__and_module_9_res,
         n_majority7_module_11__or_module_10_res,
         n_majority7_module_11__or_module_9_res,
         n_majority7_module_11__and_module_8_res,
         n_majority7_module_11__or_module_8_res,
         n_majority7_module_11__and_module_7_res,
         n_majority7_module_11__or_module_7_res,
         n_majority7_module_11__or_module_6_res,
         n_majority7_module_11__and_module_6_res,
         n_majority7_module_11__or_module_5_res,
         n_majority7_module_11__and_module_5_res,
         n_majority7_module_11__or_module_4_res,
         n_majority7_module_11__and_module_4_res,
         n_majority7_module_11__or_module_3_res,
         n_majority7_module_11__and_module_3_res,
         n_majority7_module_11__or_module_2_res,
         n_majority7_module_11__and_module_2_res,
         n_majority7_module_11__or_module_1_res,
         n_majority7_module_11__and_module_1_res, n_majority7_module_12_n7,
         n_majority7_module_12_n6, n_majority7_module_12_n5,
         n_majority7_module_12_n4, n_majority7_module_12_n3,
         n_majority7_module_12_n2, n_majority7_module_12_n1,
         n_majority7_module_12__and_module_10_res,
         n_majority7_module_12__or_module_11_res,
         n_majority7_module_12__and_module_9_res,
         n_majority7_module_12__or_module_10_res,
         n_majority7_module_12__or_module_9_res,
         n_majority7_module_12__and_module_8_res,
         n_majority7_module_12__or_module_8_res,
         n_majority7_module_12__and_module_7_res,
         n_majority7_module_12__or_module_7_res,
         n_majority7_module_12__or_module_6_res,
         n_majority7_module_12__and_module_6_res,
         n_majority7_module_12__or_module_5_res,
         n_majority7_module_12__and_module_5_res,
         n_majority7_module_12__or_module_4_res,
         n_majority7_module_12__and_module_4_res,
         n_majority7_module_12__or_module_3_res,
         n_majority7_module_12__and_module_3_res,
         n_majority7_module_12__or_module_2_res,
         n_majority7_module_12__and_module_2_res,
         n_majority7_module_12__or_module_1_res,
         n_majority7_module_12__and_module_1_res, n_majority7_module_13_n7,
         n_majority7_module_13_n6, n_majority7_module_13_n5,
         n_majority7_module_13_n4, n_majority7_module_13_n3,
         n_majority7_module_13_n2, n_majority7_module_13_n1,
         n_majority7_module_13__and_module_10_res,
         n_majority7_module_13__or_module_11_res,
         n_majority7_module_13__and_module_9_res,
         n_majority7_module_13__or_module_10_res,
         n_majority7_module_13__or_module_9_res,
         n_majority7_module_13__and_module_8_res,
         n_majority7_module_13__or_module_8_res,
         n_majority7_module_13__and_module_7_res,
         n_majority7_module_13__or_module_7_res,
         n_majority7_module_13__or_module_6_res,
         n_majority7_module_13__and_module_6_res,
         n_majority7_module_13__or_module_5_res,
         n_majority7_module_13__and_module_5_res,
         n_majority7_module_13__or_module_4_res,
         n_majority7_module_13__and_module_4_res,
         n_majority7_module_13__or_module_3_res,
         n_majority7_module_13__and_module_3_res,
         n_majority7_module_13__or_module_2_res,
         n_majority7_module_13__and_module_2_res,
         n_majority7_module_13__or_module_1_res,
         n_majority7_module_13__and_module_1_res, n_majority7_module_14_n7,
         n_majority7_module_14_n6, n_majority7_module_14_n5,
         n_majority7_module_14_n4, n_majority7_module_14_n3,
         n_majority7_module_14_n2, n_majority7_module_14_n1,
         n_majority7_module_14__and_module_10_res,
         n_majority7_module_14__or_module_11_res,
         n_majority7_module_14__and_module_9_res,
         n_majority7_module_14__or_module_10_res,
         n_majority7_module_14__or_module_9_res,
         n_majority7_module_14__and_module_8_res,
         n_majority7_module_14__or_module_8_res,
         n_majority7_module_14__and_module_7_res,
         n_majority7_module_14__or_module_7_res,
         n_majority7_module_14__or_module_6_res,
         n_majority7_module_14__and_module_6_res,
         n_majority7_module_14__or_module_5_res,
         n_majority7_module_14__and_module_5_res,
         n_majority7_module_14__or_module_4_res,
         n_majority7_module_14__and_module_4_res,
         n_majority7_module_14__or_module_3_res,
         n_majority7_module_14__and_module_3_res,
         n_majority7_module_14__or_module_2_res,
         n_majority7_module_14__and_module_2_res,
         n_majority7_module_14__or_module_1_res,
         n_majority7_module_14__and_module_1_res, n_majority7_module_15_n7,
         n_majority7_module_15_n6, n_majority7_module_15_n5,
         n_majority7_module_15_n4, n_majority7_module_15_n3,
         n_majority7_module_15_n2, n_majority7_module_15_n1,
         n_majority7_module_15__and_module_10_res,
         n_majority7_module_15__or_module_11_res,
         n_majority7_module_15__and_module_9_res,
         n_majority7_module_15__or_module_10_res,
         n_majority7_module_15__or_module_9_res,
         n_majority7_module_15__and_module_8_res,
         n_majority7_module_15__or_module_8_res,
         n_majority7_module_15__and_module_7_res,
         n_majority7_module_15__or_module_7_res,
         n_majority7_module_15__or_module_6_res,
         n_majority7_module_15__and_module_6_res,
         n_majority7_module_15__or_module_5_res,
         n_majority7_module_15__and_module_5_res,
         n_majority7_module_15__or_module_4_res,
         n_majority7_module_15__and_module_4_res,
         n_majority7_module_15__or_module_3_res,
         n_majority7_module_15__and_module_3_res,
         n_majority7_module_15__or_module_2_res,
         n_majority7_module_15__and_module_2_res,
         n_majority7_module_15__or_module_1_res,
         n_majority7_module_15__and_module_1_res, n_majority7_module_16_n7,
         n_majority7_module_16_n6, n_majority7_module_16_n5,
         n_majority7_module_16_n4, n_majority7_module_16_n3,
         n_majority7_module_16_n2, n_majority7_module_16_n1,
         n_majority7_module_16__and_module_10_res,
         n_majority7_module_16__or_module_11_res,
         n_majority7_module_16__and_module_9_res,
         n_majority7_module_16__or_module_10_res,
         n_majority7_module_16__or_module_9_res,
         n_majority7_module_16__and_module_8_res,
         n_majority7_module_16__or_module_8_res,
         n_majority7_module_16__and_module_7_res,
         n_majority7_module_16__or_module_7_res,
         n_majority7_module_16__or_module_6_res,
         n_majority7_module_16__and_module_6_res,
         n_majority7_module_16__or_module_5_res,
         n_majority7_module_16__and_module_5_res,
         n_majority7_module_16__or_module_4_res,
         n_majority7_module_16__and_module_4_res,
         n_majority7_module_16__or_module_3_res,
         n_majority7_module_16__and_module_3_res,
         n_majority7_module_16__or_module_2_res,
         n_majority7_module_16__and_module_2_res,
         n_majority7_module_16__or_module_1_res,
         n_majority7_module_16__and_module_1_res, n_majority7_module_17_n7,
         n_majority7_module_17_n6, n_majority7_module_17_n5,
         n_majority7_module_17_n4, n_majority7_module_17_n3,
         n_majority7_module_17_n2, n_majority7_module_17_n1,
         n_majority7_module_17__and_module_10_res,
         n_majority7_module_17__or_module_11_res,
         n_majority7_module_17__and_module_9_res,
         n_majority7_module_17__or_module_10_res,
         n_majority7_module_17__or_module_9_res,
         n_majority7_module_17__and_module_8_res,
         n_majority7_module_17__or_module_8_res,
         n_majority7_module_17__and_module_7_res,
         n_majority7_module_17__or_module_7_res,
         n_majority7_module_17__or_module_6_res,
         n_majority7_module_17__and_module_6_res,
         n_majority7_module_17__or_module_5_res,
         n_majority7_module_17__and_module_5_res,
         n_majority7_module_17__or_module_4_res,
         n_majority7_module_17__and_module_4_res,
         n_majority7_module_17__or_module_3_res,
         n_majority7_module_17__and_module_3_res,
         n_majority7_module_17__or_module_2_res,
         n_majority7_module_17__and_module_2_res,
         n_majority7_module_17__or_module_1_res,
         n_majority7_module_17__and_module_1_res, n_majority7_module_18_n7,
         n_majority7_module_18_n6, n_majority7_module_18_n5,
         n_majority7_module_18_n4, n_majority7_module_18_n3,
         n_majority7_module_18_n2, n_majority7_module_18_n1,
         n_majority7_module_18__and_module_10_res,
         n_majority7_module_18__or_module_11_res,
         n_majority7_module_18__and_module_9_res,
         n_majority7_module_18__or_module_10_res,
         n_majority7_module_18__or_module_9_res,
         n_majority7_module_18__and_module_8_res,
         n_majority7_module_18__or_module_8_res,
         n_majority7_module_18__and_module_7_res,
         n_majority7_module_18__or_module_7_res,
         n_majority7_module_18__or_module_6_res,
         n_majority7_module_18__and_module_6_res,
         n_majority7_module_18__or_module_5_res,
         n_majority7_module_18__and_module_5_res,
         n_majority7_module_18__or_module_4_res,
         n_majority7_module_18__and_module_4_res,
         n_majority7_module_18__or_module_3_res,
         n_majority7_module_18__and_module_3_res,
         n_majority7_module_18__or_module_2_res,
         n_majority7_module_18__and_module_2_res,
         n_majority7_module_18__or_module_1_res,
         n_majority7_module_18__and_module_1_res, n_majority7_module_19_n7,
         n_majority7_module_19_n6, n_majority7_module_19_n5,
         n_majority7_module_19_n4, n_majority7_module_19_n3,
         n_majority7_module_19_n2, n_majority7_module_19_n1,
         n_majority7_module_19__and_module_10_res,
         n_majority7_module_19__or_module_11_res,
         n_majority7_module_19__and_module_9_res,
         n_majority7_module_19__or_module_10_res,
         n_majority7_module_19__or_module_9_res,
         n_majority7_module_19__and_module_8_res,
         n_majority7_module_19__or_module_8_res,
         n_majority7_module_19__and_module_7_res,
         n_majority7_module_19__or_module_7_res,
         n_majority7_module_19__or_module_6_res,
         n_majority7_module_19__and_module_6_res,
         n_majority7_module_19__or_module_5_res,
         n_majority7_module_19__and_module_5_res,
         n_majority7_module_19__or_module_4_res,
         n_majority7_module_19__and_module_4_res,
         n_majority7_module_19__or_module_3_res,
         n_majority7_module_19__and_module_3_res,
         n_majority7_module_19__or_module_2_res,
         n_majority7_module_19__and_module_2_res,
         n_majority7_module_19__or_module_1_res,
         n_majority7_module_19__and_module_1_res, n_majority7_module_20_n7,
         n_majority7_module_20_n6, n_majority7_module_20_n5,
         n_majority7_module_20_n4, n_majority7_module_20_n3,
         n_majority7_module_20_n2, n_majority7_module_20_n1,
         n_majority7_module_20__and_module_10_res,
         n_majority7_module_20__or_module_11_res,
         n_majority7_module_20__and_module_9_res,
         n_majority7_module_20__or_module_10_res,
         n_majority7_module_20__or_module_9_res,
         n_majority7_module_20__and_module_8_res,
         n_majority7_module_20__or_module_8_res,
         n_majority7_module_20__and_module_7_res,
         n_majority7_module_20__or_module_7_res,
         n_majority7_module_20__or_module_6_res,
         n_majority7_module_20__and_module_6_res,
         n_majority7_module_20__or_module_5_res,
         n_majority7_module_20__and_module_5_res,
         n_majority7_module_20__or_module_4_res,
         n_majority7_module_20__and_module_4_res,
         n_majority7_module_20__or_module_3_res,
         n_majority7_module_20__and_module_3_res,
         n_majority7_module_20__or_module_2_res,
         n_majority7_module_20__and_module_2_res,
         n_majority7_module_20__or_module_1_res,
         n_majority7_module_20__and_module_1_res, n_majority7_module_21_n7,
         n_majority7_module_21_n6, n_majority7_module_21_n5,
         n_majority7_module_21_n4, n_majority7_module_21_n3,
         n_majority7_module_21_n2, n_majority7_module_21_n1,
         n_majority7_module_21__and_module_10_res,
         n_majority7_module_21__or_module_11_res,
         n_majority7_module_21__and_module_9_res,
         n_majority7_module_21__or_module_10_res,
         n_majority7_module_21__or_module_9_res,
         n_majority7_module_21__and_module_8_res,
         n_majority7_module_21__or_module_8_res,
         n_majority7_module_21__and_module_7_res,
         n_majority7_module_21__or_module_7_res,
         n_majority7_module_21__or_module_6_res,
         n_majority7_module_21__and_module_6_res,
         n_majority7_module_21__or_module_5_res,
         n_majority7_module_21__and_module_5_res,
         n_majority7_module_21__or_module_4_res,
         n_majority7_module_21__and_module_4_res,
         n_majority7_module_21__or_module_3_res,
         n_majority7_module_21__and_module_3_res,
         n_majority7_module_21__or_module_2_res,
         n_majority7_module_21__and_module_2_res,
         n_majority7_module_21__or_module_1_res,
         n_majority7_module_21__and_module_1_res, n_majority7_module_22_n7,
         n_majority7_module_22_n6, n_majority7_module_22_n5,
         n_majority7_module_22_n4, n_majority7_module_22_n3,
         n_majority7_module_22_n2, n_majority7_module_22_n1,
         n_majority7_module_22__and_module_10_res,
         n_majority7_module_22__or_module_11_res,
         n_majority7_module_22__and_module_9_res,
         n_majority7_module_22__or_module_10_res,
         n_majority7_module_22__or_module_9_res,
         n_majority7_module_22__and_module_8_res,
         n_majority7_module_22__or_module_8_res,
         n_majority7_module_22__and_module_7_res,
         n_majority7_module_22__or_module_7_res,
         n_majority7_module_22__or_module_6_res,
         n_majority7_module_22__and_module_6_res,
         n_majority7_module_22__or_module_5_res,
         n_majority7_module_22__and_module_5_res,
         n_majority7_module_22__or_module_4_res,
         n_majority7_module_22__and_module_4_res,
         n_majority7_module_22__or_module_3_res,
         n_majority7_module_22__and_module_3_res,
         n_majority7_module_22__or_module_2_res,
         n_majority7_module_22__and_module_2_res,
         n_majority7_module_22__or_module_1_res,
         n_majority7_module_22__and_module_1_res, n_majority7_module_23_n7,
         n_majority7_module_23_n6, n_majority7_module_23_n5,
         n_majority7_module_23_n4, n_majority7_module_23_n3,
         n_majority7_module_23_n2, n_majority7_module_23_n1,
         n_majority7_module_23__and_module_10_res,
         n_majority7_module_23__or_module_11_res,
         n_majority7_module_23__and_module_9_res,
         n_majority7_module_23__or_module_10_res,
         n_majority7_module_23__or_module_9_res,
         n_majority7_module_23__and_module_8_res,
         n_majority7_module_23__or_module_8_res,
         n_majority7_module_23__and_module_7_res,
         n_majority7_module_23__or_module_7_res,
         n_majority7_module_23__or_module_6_res,
         n_majority7_module_23__and_module_6_res,
         n_majority7_module_23__or_module_5_res,
         n_majority7_module_23__and_module_5_res,
         n_majority7_module_23__or_module_4_res,
         n_majority7_module_23__and_module_4_res,
         n_majority7_module_23__or_module_3_res,
         n_majority7_module_23__and_module_3_res,
         n_majority7_module_23__or_module_2_res,
         n_majority7_module_23__and_module_2_res,
         n_majority7_module_23__or_module_1_res,
         n_majority7_module_23__and_module_1_res, n_majority7_module_24_n7,
         n_majority7_module_24_n6, n_majority7_module_24_n5,
         n_majority7_module_24_n4, n_majority7_module_24_n3,
         n_majority7_module_24_n2, n_majority7_module_24_n1,
         n_majority7_module_24__and_module_10_res,
         n_majority7_module_24__or_module_11_res,
         n_majority7_module_24__and_module_9_res,
         n_majority7_module_24__or_module_10_res,
         n_majority7_module_24__or_module_9_res,
         n_majority7_module_24__and_module_8_res,
         n_majority7_module_24__or_module_8_res,
         n_majority7_module_24__and_module_7_res,
         n_majority7_module_24__or_module_7_res,
         n_majority7_module_24__or_module_6_res,
         n_majority7_module_24__and_module_6_res,
         n_majority7_module_24__or_module_5_res,
         n_majority7_module_24__and_module_5_res,
         n_majority7_module_24__or_module_4_res,
         n_majority7_module_24__and_module_4_res,
         n_majority7_module_24__or_module_3_res,
         n_majority7_module_24__and_module_3_res,
         n_majority7_module_24__or_module_2_res,
         n_majority7_module_24__and_module_2_res,
         n_majority7_module_24__or_module_1_res,
         n_majority7_module_24__and_module_1_res, n_majority7_module_25_n7,
         n_majority7_module_25_n6, n_majority7_module_25_n5,
         n_majority7_module_25_n4, n_majority7_module_25_n3,
         n_majority7_module_25_n2, n_majority7_module_25_n1,
         n_majority7_module_25__and_module_10_res,
         n_majority7_module_25__or_module_11_res,
         n_majority7_module_25__and_module_9_res,
         n_majority7_module_25__or_module_10_res,
         n_majority7_module_25__or_module_9_res,
         n_majority7_module_25__and_module_8_res,
         n_majority7_module_25__or_module_8_res,
         n_majority7_module_25__and_module_7_res,
         n_majority7_module_25__or_module_7_res,
         n_majority7_module_25__or_module_6_res,
         n_majority7_module_25__and_module_6_res,
         n_majority7_module_25__or_module_5_res,
         n_majority7_module_25__and_module_5_res,
         n_majority7_module_25__or_module_4_res,
         n_majority7_module_25__and_module_4_res,
         n_majority7_module_25__or_module_3_res,
         n_majority7_module_25__and_module_3_res,
         n_majority7_module_25__or_module_2_res,
         n_majority7_module_25__and_module_2_res,
         n_majority7_module_25__or_module_1_res,
         n_majority7_module_25__and_module_1_res, n_majority7_module_26_n7,
         n_majority7_module_26_n6, n_majority7_module_26_n5,
         n_majority7_module_26_n4, n_majority7_module_26_n3,
         n_majority7_module_26_n2, n_majority7_module_26_n1,
         n_majority7_module_26__and_module_10_res,
         n_majority7_module_26__or_module_11_res,
         n_majority7_module_26__and_module_9_res,
         n_majority7_module_26__or_module_10_res,
         n_majority7_module_26__or_module_9_res,
         n_majority7_module_26__and_module_8_res,
         n_majority7_module_26__or_module_8_res,
         n_majority7_module_26__and_module_7_res,
         n_majority7_module_26__or_module_7_res,
         n_majority7_module_26__or_module_6_res,
         n_majority7_module_26__and_module_6_res,
         n_majority7_module_26__or_module_5_res,
         n_majority7_module_26__and_module_5_res,
         n_majority7_module_26__or_module_4_res,
         n_majority7_module_26__and_module_4_res,
         n_majority7_module_26__or_module_3_res,
         n_majority7_module_26__and_module_3_res,
         n_majority7_module_26__or_module_2_res,
         n_majority7_module_26__and_module_2_res,
         n_majority7_module_26__or_module_1_res,
         n_majority7_module_26__and_module_1_res, n_majority7_module_27_n7,
         n_majority7_module_27_n6, n_majority7_module_27_n5,
         n_majority7_module_27_n4, n_majority7_module_27_n3,
         n_majority7_module_27_n2, n_majority7_module_27_n1,
         n_majority7_module_27__and_module_10_res,
         n_majority7_module_27__or_module_11_res,
         n_majority7_module_27__and_module_9_res,
         n_majority7_module_27__or_module_10_res,
         n_majority7_module_27__or_module_9_res,
         n_majority7_module_27__and_module_8_res,
         n_majority7_module_27__or_module_8_res,
         n_majority7_module_27__and_module_7_res,
         n_majority7_module_27__or_module_7_res,
         n_majority7_module_27__or_module_6_res,
         n_majority7_module_27__and_module_6_res,
         n_majority7_module_27__or_module_5_res,
         n_majority7_module_27__and_module_5_res,
         n_majority7_module_27__or_module_4_res,
         n_majority7_module_27__and_module_4_res,
         n_majority7_module_27__or_module_3_res,
         n_majority7_module_27__and_module_3_res,
         n_majority7_module_27__or_module_2_res,
         n_majority7_module_27__and_module_2_res,
         n_majority7_module_27__or_module_1_res,
         n_majority7_module_27__and_module_1_res, n_majority7_module_28_n7,
         n_majority7_module_28_n6, n_majority7_module_28_n5,
         n_majority7_module_28_n4, n_majority7_module_28_n3,
         n_majority7_module_28_n2, n_majority7_module_28_n1,
         n_majority7_module_28__and_module_10_res,
         n_majority7_module_28__or_module_11_res,
         n_majority7_module_28__and_module_9_res,
         n_majority7_module_28__or_module_10_res,
         n_majority7_module_28__or_module_9_res,
         n_majority7_module_28__and_module_8_res,
         n_majority7_module_28__or_module_8_res,
         n_majority7_module_28__and_module_7_res,
         n_majority7_module_28__or_module_7_res,
         n_majority7_module_28__or_module_6_res,
         n_majority7_module_28__and_module_6_res,
         n_majority7_module_28__or_module_5_res,
         n_majority7_module_28__and_module_5_res,
         n_majority7_module_28__or_module_4_res,
         n_majority7_module_28__and_module_4_res,
         n_majority7_module_28__or_module_3_res,
         n_majority7_module_28__and_module_3_res,
         n_majority7_module_28__or_module_2_res,
         n_majority7_module_28__and_module_2_res,
         n_majority7_module_28__or_module_1_res,
         n_majority7_module_28__and_module_1_res, n_majority7_module_29_n7,
         n_majority7_module_29_n6, n_majority7_module_29_n5,
         n_majority7_module_29_n4, n_majority7_module_29_n3,
         n_majority7_module_29_n2, n_majority7_module_29_n1,
         n_majority7_module_29__and_module_10_res,
         n_majority7_module_29__or_module_11_res,
         n_majority7_module_29__and_module_9_res,
         n_majority7_module_29__or_module_10_res,
         n_majority7_module_29__or_module_9_res,
         n_majority7_module_29__and_module_8_res,
         n_majority7_module_29__or_module_8_res,
         n_majority7_module_29__and_module_7_res,
         n_majority7_module_29__or_module_7_res,
         n_majority7_module_29__or_module_6_res,
         n_majority7_module_29__and_module_6_res,
         n_majority7_module_29__or_module_5_res,
         n_majority7_module_29__and_module_5_res,
         n_majority7_module_29__or_module_4_res,
         n_majority7_module_29__and_module_4_res,
         n_majority7_module_29__or_module_3_res,
         n_majority7_module_29__and_module_3_res,
         n_majority7_module_29__or_module_2_res,
         n_majority7_module_29__and_module_2_res,
         n_majority7_module_29__or_module_1_res,
         n_majority7_module_29__and_module_1_res, n_majority7_module_30_n7,
         n_majority7_module_30_n6, n_majority7_module_30_n5,
         n_majority7_module_30_n4, n_majority7_module_30_n3,
         n_majority7_module_30_n2, n_majority7_module_30_n1,
         n_majority7_module_30__and_module_10_res,
         n_majority7_module_30__or_module_11_res,
         n_majority7_module_30__and_module_9_res,
         n_majority7_module_30__or_module_10_res,
         n_majority7_module_30__or_module_9_res,
         n_majority7_module_30__and_module_8_res,
         n_majority7_module_30__or_module_8_res,
         n_majority7_module_30__and_module_7_res,
         n_majority7_module_30__or_module_7_res,
         n_majority7_module_30__or_module_6_res,
         n_majority7_module_30__and_module_6_res,
         n_majority7_module_30__or_module_5_res,
         n_majority7_module_30__and_module_5_res,
         n_majority7_module_30__or_module_4_res,
         n_majority7_module_30__and_module_4_res,
         n_majority7_module_30__or_module_3_res,
         n_majority7_module_30__and_module_3_res,
         n_majority7_module_30__or_module_2_res,
         n_majority7_module_30__and_module_2_res,
         n_majority7_module_30__or_module_1_res,
         n_majority7_module_30__and_module_1_res, n_majority7_module_31_n7,
         n_majority7_module_31_n6, n_majority7_module_31_n5,
         n_majority7_module_31_n4, n_majority7_module_31_n3,
         n_majority7_module_31_n2, n_majority7_module_31_n1,
         n_majority7_module_31__and_module_10_res,
         n_majority7_module_31__or_module_11_res,
         n_majority7_module_31__and_module_9_res,
         n_majority7_module_31__or_module_10_res,
         n_majority7_module_31__or_module_9_res,
         n_majority7_module_31__and_module_8_res,
         n_majority7_module_31__or_module_8_res,
         n_majority7_module_31__and_module_7_res,
         n_majority7_module_31__or_module_7_res,
         n_majority7_module_31__or_module_6_res,
         n_majority7_module_31__and_module_6_res,
         n_majority7_module_31__or_module_5_res,
         n_majority7_module_31__and_module_5_res,
         n_majority7_module_31__or_module_4_res,
         n_majority7_module_31__and_module_4_res,
         n_majority7_module_31__or_module_3_res,
         n_majority7_module_31__and_module_3_res,
         n_majority7_module_31__or_module_2_res,
         n_majority7_module_31__and_module_2_res,
         n_majority7_module_31__or_module_1_res,
         n_majority7_module_31__and_module_1_res, n_majority7_module_32_n7,
         n_majority7_module_32_n6, n_majority7_module_32_n5,
         n_majority7_module_32_n4, n_majority7_module_32_n3,
         n_majority7_module_32_n2, n_majority7_module_32_n1,
         n_majority7_module_32__and_module_10_res,
         n_majority7_module_32__or_module_11_res,
         n_majority7_module_32__and_module_9_res,
         n_majority7_module_32__or_module_10_res,
         n_majority7_module_32__or_module_9_res,
         n_majority7_module_32__and_module_8_res,
         n_majority7_module_32__or_module_8_res,
         n_majority7_module_32__and_module_7_res,
         n_majority7_module_32__or_module_7_res,
         n_majority7_module_32__or_module_6_res,
         n_majority7_module_32__and_module_6_res,
         n_majority7_module_32__or_module_5_res,
         n_majority7_module_32__and_module_5_res,
         n_majority7_module_32__or_module_4_res,
         n_majority7_module_32__and_module_4_res,
         n_majority7_module_32__or_module_3_res,
         n_majority7_module_32__and_module_3_res,
         n_majority7_module_32__or_module_2_res,
         n_majority7_module_32__and_module_2_res,
         n_majority7_module_32__or_module_1_res,
         n_majority7_module_32__and_module_1_res, n_majority7_module_33_n7,
         n_majority7_module_33_n6, n_majority7_module_33_n5,
         n_majority7_module_33_n4, n_majority7_module_33_n3,
         n_majority7_module_33_n2, n_majority7_module_33_n1,
         n_majority7_module_33__and_module_10_res,
         n_majority7_module_33__or_module_11_res,
         n_majority7_module_33__and_module_9_res,
         n_majority7_module_33__or_module_10_res,
         n_majority7_module_33__or_module_9_res,
         n_majority7_module_33__and_module_8_res,
         n_majority7_module_33__or_module_8_res,
         n_majority7_module_33__and_module_7_res,
         n_majority7_module_33__or_module_7_res,
         n_majority7_module_33__or_module_6_res,
         n_majority7_module_33__and_module_6_res,
         n_majority7_module_33__or_module_5_res,
         n_majority7_module_33__and_module_5_res,
         n_majority7_module_33__or_module_4_res,
         n_majority7_module_33__and_module_4_res,
         n_majority7_module_33__or_module_3_res,
         n_majority7_module_33__and_module_3_res,
         n_majority7_module_33__or_module_2_res,
         n_majority7_module_33__and_module_2_res,
         n_majority7_module_33__or_module_1_res,
         n_majority7_module_33__and_module_1_res, n_majority7_module_34_n7,
         n_majority7_module_34_n6, n_majority7_module_34_n5,
         n_majority7_module_34_n4, n_majority7_module_34_n3,
         n_majority7_module_34_n2, n_majority7_module_34_n1,
         n_majority7_module_34__and_module_10_res,
         n_majority7_module_34__or_module_11_res,
         n_majority7_module_34__and_module_9_res,
         n_majority7_module_34__or_module_10_res,
         n_majority7_module_34__or_module_9_res,
         n_majority7_module_34__and_module_8_res,
         n_majority7_module_34__or_module_8_res,
         n_majority7_module_34__and_module_7_res,
         n_majority7_module_34__or_module_7_res,
         n_majority7_module_34__or_module_6_res,
         n_majority7_module_34__and_module_6_res,
         n_majority7_module_34__or_module_5_res,
         n_majority7_module_34__and_module_5_res,
         n_majority7_module_34__or_module_4_res,
         n_majority7_module_34__and_module_4_res,
         n_majority7_module_34__or_module_3_res,
         n_majority7_module_34__and_module_3_res,
         n_majority7_module_34__or_module_2_res,
         n_majority7_module_34__and_module_2_res,
         n_majority7_module_34__or_module_1_res,
         n_majority7_module_34__and_module_1_res, n_majority7_module_35_n7,
         n_majority7_module_35_n6, n_majority7_module_35_n5,
         n_majority7_module_35_n4, n_majority7_module_35_n3,
         n_majority7_module_35_n2, n_majority7_module_35_n1,
         n_majority7_module_35__and_module_10_res,
         n_majority7_module_35__or_module_11_res,
         n_majority7_module_35__and_module_9_res,
         n_majority7_module_35__or_module_10_res,
         n_majority7_module_35__or_module_9_res,
         n_majority7_module_35__and_module_8_res,
         n_majority7_module_35__or_module_8_res,
         n_majority7_module_35__and_module_7_res,
         n_majority7_module_35__or_module_7_res,
         n_majority7_module_35__or_module_6_res,
         n_majority7_module_35__and_module_6_res,
         n_majority7_module_35__or_module_5_res,
         n_majority7_module_35__and_module_5_res,
         n_majority7_module_35__or_module_4_res,
         n_majority7_module_35__and_module_4_res,
         n_majority7_module_35__or_module_3_res,
         n_majority7_module_35__and_module_3_res,
         n_majority7_module_35__or_module_2_res,
         n_majority7_module_35__and_module_2_res,
         n_majority7_module_35__or_module_1_res,
         n_majority7_module_35__and_module_1_res, n_majority7_module_36_n7,
         n_majority7_module_36_n6, n_majority7_module_36_n5,
         n_majority7_module_36_n4, n_majority7_module_36_n3,
         n_majority7_module_36_n2, n_majority7_module_36_n1,
         n_majority7_module_36__and_module_10_res,
         n_majority7_module_36__or_module_11_res,
         n_majority7_module_36__and_module_9_res,
         n_majority7_module_36__or_module_10_res,
         n_majority7_module_36__or_module_9_res,
         n_majority7_module_36__and_module_8_res,
         n_majority7_module_36__or_module_8_res,
         n_majority7_module_36__and_module_7_res,
         n_majority7_module_36__or_module_7_res,
         n_majority7_module_36__or_module_6_res,
         n_majority7_module_36__and_module_6_res,
         n_majority7_module_36__or_module_5_res,
         n_majority7_module_36__and_module_5_res,
         n_majority7_module_36__or_module_4_res,
         n_majority7_module_36__and_module_4_res,
         n_majority7_module_36__or_module_3_res,
         n_majority7_module_36__and_module_3_res,
         n_majority7_module_36__or_module_2_res,
         n_majority7_module_36__and_module_2_res,
         n_majority7_module_36__or_module_1_res,
         n_majority7_module_36__and_module_1_res, n_majority7_module_37_n7,
         n_majority7_module_37_n6, n_majority7_module_37_n5,
         n_majority7_module_37_n4, n_majority7_module_37_n3,
         n_majority7_module_37_n2, n_majority7_module_37_n1,
         n_majority7_module_37__and_module_10_res,
         n_majority7_module_37__or_module_11_res,
         n_majority7_module_37__and_module_9_res,
         n_majority7_module_37__or_module_10_res,
         n_majority7_module_37__or_module_9_res,
         n_majority7_module_37__and_module_8_res,
         n_majority7_module_37__or_module_8_res,
         n_majority7_module_37__and_module_7_res,
         n_majority7_module_37__or_module_7_res,
         n_majority7_module_37__or_module_6_res,
         n_majority7_module_37__and_module_6_res,
         n_majority7_module_37__or_module_5_res,
         n_majority7_module_37__and_module_5_res,
         n_majority7_module_37__or_module_4_res,
         n_majority7_module_37__and_module_4_res,
         n_majority7_module_37__or_module_3_res,
         n_majority7_module_37__and_module_3_res,
         n_majority7_module_37__or_module_2_res,
         n_majority7_module_37__and_module_2_res,
         n_majority7_module_37__or_module_1_res,
         n_majority7_module_37__and_module_1_res, n_majority7_module_38_n7,
         n_majority7_module_38_n6, n_majority7_module_38_n5,
         n_majority7_module_38_n4, n_majority7_module_38_n3,
         n_majority7_module_38_n2, n_majority7_module_38_n1,
         n_majority7_module_38__and_module_10_res,
         n_majority7_module_38__or_module_11_res,
         n_majority7_module_38__and_module_9_res,
         n_majority7_module_38__or_module_10_res,
         n_majority7_module_38__or_module_9_res,
         n_majority7_module_38__and_module_8_res,
         n_majority7_module_38__or_module_8_res,
         n_majority7_module_38__and_module_7_res,
         n_majority7_module_38__or_module_7_res,
         n_majority7_module_38__or_module_6_res,
         n_majority7_module_38__and_module_6_res,
         n_majority7_module_38__or_module_5_res,
         n_majority7_module_38__and_module_5_res,
         n_majority7_module_38__or_module_4_res,
         n_majority7_module_38__and_module_4_res,
         n_majority7_module_38__or_module_3_res,
         n_majority7_module_38__and_module_3_res,
         n_majority7_module_38__or_module_2_res,
         n_majority7_module_38__and_module_2_res,
         n_majority7_module_38__or_module_1_res,
         n_majority7_module_38__and_module_1_res, n_majority7_module_39_n7,
         n_majority7_module_39_n6, n_majority7_module_39_n5,
         n_majority7_module_39_n4, n_majority7_module_39_n3,
         n_majority7_module_39_n2, n_majority7_module_39_n1,
         n_majority7_module_39__and_module_10_res,
         n_majority7_module_39__or_module_11_res,
         n_majority7_module_39__and_module_9_res,
         n_majority7_module_39__or_module_10_res,
         n_majority7_module_39__or_module_9_res,
         n_majority7_module_39__and_module_8_res,
         n_majority7_module_39__or_module_8_res,
         n_majority7_module_39__and_module_7_res,
         n_majority7_module_39__or_module_7_res,
         n_majority7_module_39__or_module_6_res,
         n_majority7_module_39__and_module_6_res,
         n_majority7_module_39__or_module_5_res,
         n_majority7_module_39__and_module_5_res,
         n_majority7_module_39__or_module_4_res,
         n_majority7_module_39__and_module_4_res,
         n_majority7_module_39__or_module_3_res,
         n_majority7_module_39__and_module_3_res,
         n_majority7_module_39__or_module_2_res,
         n_majority7_module_39__and_module_2_res,
         n_majority7_module_39__or_module_1_res,
         n_majority7_module_39__and_module_1_res, n_majority7_module_40_n7,
         n_majority7_module_40_n6, n_majority7_module_40_n5,
         n_majority7_module_40_n4, n_majority7_module_40_n3,
         n_majority7_module_40_n2, n_majority7_module_40_n1,
         n_majority7_module_40__and_module_10_res,
         n_majority7_module_40__or_module_11_res,
         n_majority7_module_40__and_module_9_res,
         n_majority7_module_40__or_module_10_res,
         n_majority7_module_40__or_module_9_res,
         n_majority7_module_40__and_module_8_res,
         n_majority7_module_40__or_module_8_res,
         n_majority7_module_40__and_module_7_res,
         n_majority7_module_40__or_module_7_res,
         n_majority7_module_40__or_module_6_res,
         n_majority7_module_40__and_module_6_res,
         n_majority7_module_40__or_module_5_res,
         n_majority7_module_40__and_module_5_res,
         n_majority7_module_40__or_module_4_res,
         n_majority7_module_40__and_module_4_res,
         n_majority7_module_40__or_module_3_res,
         n_majority7_module_40__and_module_3_res,
         n_majority7_module_40__or_module_2_res,
         n_majority7_module_40__and_module_2_res,
         n_majority7_module_40__or_module_1_res,
         n_majority7_module_40__and_module_1_res, n_majority7_module_41_n7,
         n_majority7_module_41_n6, n_majority7_module_41_n5,
         n_majority7_module_41_n4, n_majority7_module_41_n3,
         n_majority7_module_41_n2, n_majority7_module_41_n1,
         n_majority7_module_41__and_module_10_res,
         n_majority7_module_41__or_module_11_res,
         n_majority7_module_41__and_module_9_res,
         n_majority7_module_41__or_module_10_res,
         n_majority7_module_41__or_module_9_res,
         n_majority7_module_41__and_module_8_res,
         n_majority7_module_41__or_module_8_res,
         n_majority7_module_41__and_module_7_res,
         n_majority7_module_41__or_module_7_res,
         n_majority7_module_41__or_module_6_res,
         n_majority7_module_41__and_module_6_res,
         n_majority7_module_41__or_module_5_res,
         n_majority7_module_41__and_module_5_res,
         n_majority7_module_41__or_module_4_res,
         n_majority7_module_41__and_module_4_res,
         n_majority7_module_41__or_module_3_res,
         n_majority7_module_41__and_module_3_res,
         n_majority7_module_41__or_module_2_res,
         n_majority7_module_41__and_module_2_res,
         n_majority7_module_41__or_module_1_res,
         n_majority7_module_41__and_module_1_res, n_majority7_module_42_n7,
         n_majority7_module_42_n6, n_majority7_module_42_n5,
         n_majority7_module_42_n4, n_majority7_module_42_n3,
         n_majority7_module_42_n2, n_majority7_module_42_n1,
         n_majority7_module_42__and_module_10_res,
         n_majority7_module_42__or_module_11_res,
         n_majority7_module_42__and_module_9_res,
         n_majority7_module_42__or_module_10_res,
         n_majority7_module_42__or_module_9_res,
         n_majority7_module_42__and_module_8_res,
         n_majority7_module_42__or_module_8_res,
         n_majority7_module_42__and_module_7_res,
         n_majority7_module_42__or_module_7_res,
         n_majority7_module_42__or_module_6_res,
         n_majority7_module_42__and_module_6_res,
         n_majority7_module_42__or_module_5_res,
         n_majority7_module_42__and_module_5_res,
         n_majority7_module_42__or_module_4_res,
         n_majority7_module_42__and_module_4_res,
         n_majority7_module_42__or_module_3_res,
         n_majority7_module_42__and_module_3_res,
         n_majority7_module_42__or_module_2_res,
         n_majority7_module_42__and_module_2_res,
         n_majority7_module_42__or_module_1_res,
         n_majority7_module_42__and_module_1_res, n_majority7_module_43_n7,
         n_majority7_module_43_n6, n_majority7_module_43_n5,
         n_majority7_module_43_n4, n_majority7_module_43_n3,
         n_majority7_module_43_n2, n_majority7_module_43_n1,
         n_majority7_module_43__and_module_10_res,
         n_majority7_module_43__or_module_11_res,
         n_majority7_module_43__and_module_9_res,
         n_majority7_module_43__or_module_10_res,
         n_majority7_module_43__or_module_9_res,
         n_majority7_module_43__and_module_8_res,
         n_majority7_module_43__or_module_8_res,
         n_majority7_module_43__and_module_7_res,
         n_majority7_module_43__or_module_7_res,
         n_majority7_module_43__or_module_6_res,
         n_majority7_module_43__and_module_6_res,
         n_majority7_module_43__or_module_5_res,
         n_majority7_module_43__and_module_5_res,
         n_majority7_module_43__or_module_4_res,
         n_majority7_module_43__and_module_4_res,
         n_majority7_module_43__or_module_3_res,
         n_majority7_module_43__and_module_3_res,
         n_majority7_module_43__or_module_2_res,
         n_majority7_module_43__and_module_2_res,
         n_majority7_module_43__or_module_1_res,
         n_majority7_module_43__and_module_1_res, n_majority7_module_44_n7,
         n_majority7_module_44_n6, n_majority7_module_44_n5,
         n_majority7_module_44_n4, n_majority7_module_44_n3,
         n_majority7_module_44_n2, n_majority7_module_44_n1,
         n_majority7_module_44__and_module_10_res,
         n_majority7_module_44__or_module_11_res,
         n_majority7_module_44__and_module_9_res,
         n_majority7_module_44__or_module_10_res,
         n_majority7_module_44__or_module_9_res,
         n_majority7_module_44__and_module_8_res,
         n_majority7_module_44__or_module_8_res,
         n_majority7_module_44__and_module_7_res,
         n_majority7_module_44__or_module_7_res,
         n_majority7_module_44__or_module_6_res,
         n_majority7_module_44__and_module_6_res,
         n_majority7_module_44__or_module_5_res,
         n_majority7_module_44__and_module_5_res,
         n_majority7_module_44__or_module_4_res,
         n_majority7_module_44__and_module_4_res,
         n_majority7_module_44__or_module_3_res,
         n_majority7_module_44__and_module_3_res,
         n_majority7_module_44__or_module_2_res,
         n_majority7_module_44__and_module_2_res,
         n_majority7_module_44__or_module_1_res,
         n_majority7_module_44__and_module_1_res,
         n_majority7_module_45__and_module_10_res,
         n_majority7_module_45__or_module_11_res,
         n_majority7_module_45__and_module_9_res,
         n_majority7_module_45__or_module_10_res,
         n_majority7_module_45__or_module_9_res,
         n_majority7_module_45__and_module_8_res,
         n_majority7_module_45__or_module_8_res,
         n_majority7_module_45__and_module_7_res,
         n_majority7_module_45__or_module_7_res,
         n_majority7_module_45__or_module_6_res,
         n_majority7_module_45__and_module_6_res,
         n_majority7_module_45__or_module_5_res,
         n_majority7_module_45__and_module_5_res,
         n_majority7_module_45__or_module_4_res,
         n_majority7_module_45__and_module_4_res,
         n_majority7_module_45__or_module_3_res,
         n_majority7_module_45__and_module_3_res,
         n_majority7_module_45__or_module_2_res,
         n_majority7_module_45__and_module_2_res,
         n_majority7_module_45__or_module_1_res,
         n_majority7_module_45__and_module_1_res,
         n_majority7_module_46__and_module_10_res,
         n_majority7_module_46__or_module_11_res,
         n_majority7_module_46__and_module_9_res,
         n_majority7_module_46__or_module_10_res,
         n_majority7_module_46__or_module_9_res,
         n_majority7_module_46__and_module_8_res,
         n_majority7_module_46__or_module_8_res,
         n_majority7_module_46__and_module_7_res,
         n_majority7_module_46__or_module_7_res,
         n_majority7_module_46__or_module_6_res,
         n_majority7_module_46__and_module_6_res,
         n_majority7_module_46__or_module_5_res,
         n_majority7_module_46__and_module_5_res,
         n_majority7_module_46__or_module_4_res,
         n_majority7_module_46__and_module_4_res,
         n_majority7_module_46__or_module_3_res,
         n_majority7_module_46__and_module_3_res,
         n_majority7_module_46__or_module_2_res,
         n_majority7_module_46__and_module_2_res,
         n_majority7_module_46__or_module_1_res,
         n_majority7_module_46__and_module_1_res,
         n_majority7_module_47__and_module_10_res,
         n_majority7_module_47__or_module_11_res,
         n_majority7_module_47__and_module_9_res,
         n_majority7_module_47__or_module_10_res,
         n_majority7_module_47__or_module_9_res,
         n_majority7_module_47__and_module_8_res,
         n_majority7_module_47__or_module_8_res,
         n_majority7_module_47__and_module_7_res,
         n_majority7_module_47__or_module_7_res,
         n_majority7_module_47__or_module_6_res,
         n_majority7_module_47__and_module_6_res,
         n_majority7_module_47__or_module_5_res,
         n_majority7_module_47__and_module_5_res,
         n_majority7_module_47__or_module_4_res,
         n_majority7_module_47__and_module_4_res,
         n_majority7_module_47__or_module_3_res,
         n_majority7_module_47__and_module_3_res,
         n_majority7_module_47__or_module_2_res,
         n_majority7_module_47__and_module_2_res,
         n_majority7_module_47__or_module_1_res,
         n_majority7_module_47__and_module_1_res,
         n_majority7_module_48__and_module_10_res,
         n_majority7_module_48__or_module_11_res,
         n_majority7_module_48__and_module_9_res,
         n_majority7_module_48__or_module_10_res,
         n_majority7_module_48__or_module_9_res,
         n_majority7_module_48__and_module_8_res,
         n_majority7_module_48__or_module_8_res,
         n_majority7_module_48__and_module_7_res,
         n_majority7_module_48__or_module_7_res,
         n_majority7_module_48__or_module_6_res,
         n_majority7_module_48__and_module_6_res,
         n_majority7_module_48__or_module_5_res,
         n_majority7_module_48__and_module_5_res,
         n_majority7_module_48__or_module_4_res,
         n_majority7_module_48__and_module_4_res,
         n_majority7_module_48__or_module_3_res,
         n_majority7_module_48__and_module_3_res,
         n_majority7_module_48__or_module_2_res,
         n_majority7_module_48__and_module_2_res,
         n_majority7_module_48__or_module_1_res,
         n_majority7_module_48__and_module_1_res,
         n_majority7_module_49__and_module_10_res,
         n_majority7_module_49__or_module_11_res,
         n_majority7_module_49__and_module_9_res,
         n_majority7_module_49__or_module_10_res,
         n_majority7_module_49__or_module_9_res,
         n_majority7_module_49__and_module_8_res,
         n_majority7_module_49__or_module_8_res,
         n_majority7_module_49__and_module_7_res,
         n_majority7_module_49__or_module_7_res,
         n_majority7_module_49__or_module_6_res,
         n_majority7_module_49__and_module_6_res,
         n_majority7_module_49__or_module_5_res,
         n_majority7_module_49__and_module_5_res,
         n_majority7_module_49__or_module_4_res,
         n_majority7_module_49__and_module_4_res,
         n_majority7_module_49__or_module_3_res,
         n_majority7_module_49__and_module_3_res,
         n_majority7_module_49__or_module_2_res,
         n_majority7_module_49__and_module_2_res,
         n_majority7_module_49__or_module_1_res,
         n_majority7_module_49__and_module_1_res,
         n_majority7_module_50__and_module_10_res,
         n_majority7_module_50__or_module_11_res,
         n_majority7_module_50__and_module_9_res,
         n_majority7_module_50__or_module_10_res,
         n_majority7_module_50__or_module_9_res,
         n_majority7_module_50__and_module_8_res,
         n_majority7_module_50__or_module_8_res,
         n_majority7_module_50__and_module_7_res,
         n_majority7_module_50__or_module_7_res,
         n_majority7_module_50__or_module_6_res,
         n_majority7_module_50__and_module_6_res,
         n_majority7_module_50__or_module_5_res,
         n_majority7_module_50__and_module_5_res,
         n_majority7_module_50__or_module_4_res,
         n_majority7_module_50__and_module_4_res,
         n_majority7_module_50__or_module_3_res,
         n_majority7_module_50__and_module_3_res,
         n_majority7_module_50__or_module_2_res,
         n_majority7_module_50__and_module_2_res,
         n_majority7_module_50__or_module_1_res,
         n_majority7_module_50__and_module_1_res,
         n_majority7_module_51__and_module_10_res,
         n_majority7_module_51__or_module_11_res,
         n_majority7_module_51__and_module_9_res,
         n_majority7_module_51__or_module_10_res,
         n_majority7_module_51__or_module_9_res,
         n_majority7_module_51__and_module_8_res,
         n_majority7_module_51__or_module_8_res,
         n_majority7_module_51__and_module_7_res,
         n_majority7_module_51__or_module_7_res,
         n_majority7_module_51__or_module_6_res,
         n_majority7_module_51__and_module_6_res,
         n_majority7_module_51__or_module_5_res,
         n_majority7_module_51__and_module_5_res,
         n_majority7_module_51__or_module_4_res,
         n_majority7_module_51__and_module_4_res,
         n_majority7_module_51__or_module_3_res,
         n_majority7_module_51__and_module_3_res,
         n_majority7_module_51__or_module_2_res,
         n_majority7_module_51__and_module_2_res,
         n_majority7_module_51__or_module_1_res,
         n_majority7_module_51__and_module_1_res,
         n_majority7_module_52__and_module_10_res,
         n_majority7_module_52__or_module_11_res,
         n_majority7_module_52__and_module_9_res,
         n_majority7_module_52__or_module_10_res,
         n_majority7_module_52__or_module_9_res,
         n_majority7_module_52__and_module_8_res,
         n_majority7_module_52__or_module_8_res,
         n_majority7_module_52__and_module_7_res,
         n_majority7_module_52__or_module_7_res,
         n_majority7_module_52__or_module_6_res,
         n_majority7_module_52__and_module_6_res,
         n_majority7_module_52__or_module_5_res,
         n_majority7_module_52__and_module_5_res,
         n_majority7_module_52__or_module_4_res,
         n_majority7_module_52__and_module_4_res,
         n_majority7_module_52__or_module_3_res,
         n_majority7_module_52__and_module_3_res,
         n_majority7_module_52__or_module_2_res,
         n_majority7_module_52__and_module_2_res,
         n_majority7_module_52__or_module_1_res,
         n_majority7_module_52__and_module_1_res,
         n_majority7_module_53__and_module_10_res,
         n_majority7_module_53__or_module_11_res,
         n_majority7_module_53__and_module_9_res,
         n_majority7_module_53__or_module_10_res,
         n_majority7_module_53__or_module_9_res,
         n_majority7_module_53__and_module_8_res,
         n_majority7_module_53__or_module_8_res,
         n_majority7_module_53__and_module_7_res,
         n_majority7_module_53__or_module_7_res,
         n_majority7_module_53__or_module_6_res,
         n_majority7_module_53__and_module_6_res,
         n_majority7_module_53__or_module_5_res,
         n_majority7_module_53__and_module_5_res,
         n_majority7_module_53__or_module_4_res,
         n_majority7_module_53__and_module_4_res,
         n_majority7_module_53__or_module_3_res,
         n_majority7_module_53__and_module_3_res,
         n_majority7_module_53__or_module_2_res,
         n_majority7_module_53__and_module_2_res,
         n_majority7_module_53__or_module_1_res,
         n_majority7_module_53__and_module_1_res,
         n_majority7_module_54__and_module_10_res,
         n_majority7_module_54__or_module_11_res,
         n_majority7_module_54__and_module_9_res,
         n_majority7_module_54__or_module_10_res,
         n_majority7_module_54__or_module_9_res,
         n_majority7_module_54__and_module_8_res,
         n_majority7_module_54__or_module_8_res,
         n_majority7_module_54__and_module_7_res,
         n_majority7_module_54__or_module_7_res,
         n_majority7_module_54__or_module_6_res,
         n_majority7_module_54__and_module_6_res,
         n_majority7_module_54__or_module_5_res,
         n_majority7_module_54__and_module_5_res,
         n_majority7_module_54__or_module_4_res,
         n_majority7_module_54__and_module_4_res,
         n_majority7_module_54__or_module_3_res,
         n_majority7_module_54__and_module_3_res,
         n_majority7_module_54__or_module_2_res,
         n_majority7_module_54__and_module_2_res,
         n_majority7_module_54__or_module_1_res,
         n_majority7_module_54__and_module_1_res,
         n_majority7_module_55__and_module_10_res,
         n_majority7_module_55__or_module_11_res,
         n_majority7_module_55__and_module_9_res,
         n_majority7_module_55__or_module_10_res,
         n_majority7_module_55__or_module_9_res,
         n_majority7_module_55__and_module_8_res,
         n_majority7_module_55__or_module_8_res,
         n_majority7_module_55__and_module_7_res,
         n_majority7_module_55__or_module_7_res,
         n_majority7_module_55__or_module_6_res,
         n_majority7_module_55__and_module_6_res,
         n_majority7_module_55__or_module_5_res,
         n_majority7_module_55__and_module_5_res,
         n_majority7_module_55__or_module_4_res,
         n_majority7_module_55__and_module_4_res,
         n_majority7_module_55__or_module_3_res,
         n_majority7_module_55__and_module_3_res,
         n_majority7_module_55__or_module_2_res,
         n_majority7_module_55__and_module_2_res,
         n_majority7_module_55__or_module_1_res,
         n_majority7_module_55__and_module_1_res,
         n_majority7_module_56__and_module_10_res,
         n_majority7_module_56__or_module_11_res,
         n_majority7_module_56__and_module_9_res,
         n_majority7_module_56__or_module_10_res,
         n_majority7_module_56__or_module_9_res,
         n_majority7_module_56__and_module_8_res,
         n_majority7_module_56__or_module_8_res,
         n_majority7_module_56__and_module_7_res,
         n_majority7_module_56__or_module_7_res,
         n_majority7_module_56__or_module_6_res,
         n_majority7_module_56__and_module_6_res,
         n_majority7_module_56__or_module_5_res,
         n_majority7_module_56__and_module_5_res,
         n_majority7_module_56__or_module_4_res,
         n_majority7_module_56__and_module_4_res,
         n_majority7_module_56__or_module_3_res,
         n_majority7_module_56__and_module_3_res,
         n_majority7_module_56__or_module_2_res,
         n_majority7_module_56__and_module_2_res,
         n_majority7_module_56__or_module_1_res,
         n_majority7_module_56__and_module_1_res,
         n_majority7_module_57__and_module_10_res,
         n_majority7_module_57__or_module_11_res,
         n_majority7_module_57__and_module_9_res,
         n_majority7_module_57__or_module_10_res,
         n_majority7_module_57__or_module_9_res,
         n_majority7_module_57__and_module_8_res,
         n_majority7_module_57__or_module_8_res,
         n_majority7_module_57__and_module_7_res,
         n_majority7_module_57__or_module_7_res,
         n_majority7_module_57__or_module_6_res,
         n_majority7_module_57__and_module_6_res,
         n_majority7_module_57__or_module_5_res,
         n_majority7_module_57__and_module_5_res,
         n_majority7_module_57__or_module_4_res,
         n_majority7_module_57__and_module_4_res,
         n_majority7_module_57__or_module_3_res,
         n_majority7_module_57__and_module_3_res,
         n_majority7_module_57__or_module_2_res,
         n_majority7_module_57__and_module_2_res,
         n_majority7_module_57__or_module_1_res,
         n_majority7_module_57__and_module_1_res,
         n_majority7_module_58__and_module_10_res,
         n_majority7_module_58__or_module_11_res,
         n_majority7_module_58__and_module_9_res,
         n_majority7_module_58__or_module_10_res,
         n_majority7_module_58__or_module_9_res,
         n_majority7_module_58__and_module_8_res,
         n_majority7_module_58__or_module_8_res,
         n_majority7_module_58__and_module_7_res,
         n_majority7_module_58__or_module_7_res,
         n_majority7_module_58__or_module_6_res,
         n_majority7_module_58__and_module_6_res,
         n_majority7_module_58__or_module_5_res,
         n_majority7_module_58__and_module_5_res,
         n_majority7_module_58__or_module_4_res,
         n_majority7_module_58__and_module_4_res,
         n_majority7_module_58__or_module_3_res,
         n_majority7_module_58__and_module_3_res,
         n_majority7_module_58__or_module_2_res,
         n_majority7_module_58__and_module_2_res,
         n_majority7_module_58__or_module_1_res,
         n_majority7_module_58__and_module_1_res,
         n_majority7_module_59__and_module_10_res,
         n_majority7_module_59__or_module_11_res,
         n_majority7_module_59__and_module_9_res,
         n_majority7_module_59__or_module_10_res,
         n_majority7_module_59__or_module_9_res,
         n_majority7_module_59__and_module_8_res,
         n_majority7_module_59__or_module_8_res,
         n_majority7_module_59__and_module_7_res,
         n_majority7_module_59__or_module_7_res,
         n_majority7_module_59__or_module_6_res,
         n_majority7_module_59__and_module_6_res,
         n_majority7_module_59__or_module_5_res,
         n_majority7_module_59__and_module_5_res,
         n_majority7_module_59__or_module_4_res,
         n_majority7_module_59__and_module_4_res,
         n_majority7_module_59__or_module_3_res,
         n_majority7_module_59__and_module_3_res,
         n_majority7_module_59__or_module_2_res,
         n_majority7_module_59__and_module_2_res,
         n_majority7_module_59__or_module_1_res,
         n_majority7_module_59__and_module_1_res,
         n_majority7_module_60__and_module_10_res,
         n_majority7_module_60__or_module_11_res,
         n_majority7_module_60__and_module_9_res,
         n_majority7_module_60__or_module_10_res,
         n_majority7_module_60__or_module_9_res,
         n_majority7_module_60__and_module_8_res,
         n_majority7_module_60__or_module_8_res,
         n_majority7_module_60__and_module_7_res,
         n_majority7_module_60__or_module_7_res,
         n_majority7_module_60__or_module_6_res,
         n_majority7_module_60__and_module_6_res,
         n_majority7_module_60__or_module_5_res,
         n_majority7_module_60__and_module_5_res,
         n_majority7_module_60__or_module_4_res,
         n_majority7_module_60__and_module_4_res,
         n_majority7_module_60__or_module_3_res,
         n_majority7_module_60__and_module_3_res,
         n_majority7_module_60__or_module_2_res,
         n_majority7_module_60__and_module_2_res,
         n_majority7_module_60__or_module_1_res,
         n_majority7_module_60__and_module_1_res,
         n_majority7_module_61__and_module_10_res,
         n_majority7_module_61__or_module_11_res,
         n_majority7_module_61__and_module_9_res,
         n_majority7_module_61__or_module_10_res,
         n_majority7_module_61__or_module_9_res,
         n_majority7_module_61__and_module_8_res,
         n_majority7_module_61__or_module_8_res,
         n_majority7_module_61__and_module_7_res,
         n_majority7_module_61__or_module_7_res,
         n_majority7_module_61__or_module_6_res,
         n_majority7_module_61__and_module_6_res,
         n_majority7_module_61__or_module_5_res,
         n_majority7_module_61__and_module_5_res,
         n_majority7_module_61__or_module_4_res,
         n_majority7_module_61__and_module_4_res,
         n_majority7_module_61__or_module_3_res,
         n_majority7_module_61__and_module_3_res,
         n_majority7_module_61__or_module_2_res,
         n_majority7_module_61__and_module_2_res,
         n_majority7_module_61__or_module_1_res,
         n_majority7_module_61__and_module_1_res,
         n_majority7_module_62__and_module_10_res,
         n_majority7_module_62__or_module_11_res,
         n_majority7_module_62__and_module_9_res,
         n_majority7_module_62__or_module_10_res,
         n_majority7_module_62__or_module_9_res,
         n_majority7_module_62__and_module_8_res,
         n_majority7_module_62__or_module_8_res,
         n_majority7_module_62__and_module_7_res,
         n_majority7_module_62__or_module_7_res,
         n_majority7_module_62__or_module_6_res,
         n_majority7_module_62__and_module_6_res,
         n_majority7_module_62__or_module_5_res,
         n_majority7_module_62__and_module_5_res,
         n_majority7_module_62__or_module_4_res,
         n_majority7_module_62__and_module_4_res,
         n_majority7_module_62__or_module_3_res,
         n_majority7_module_62__and_module_3_res,
         n_majority7_module_62__or_module_2_res,
         n_majority7_module_62__and_module_2_res,
         n_majority7_module_62__or_module_1_res,
         n_majority7_module_62__and_module_1_res;

  XOR2_X1 u_xor_module_1_U1 ( .A(p_rand_0), .B(io_i1_s0_d0), .Z(
        n_xor_module_1_res) );
  XOR2_X2 u_xor_module_2_U1 ( .A(p_rand_1), .B(n_xor_module_1_res), .Z(
        n_xor_module_2_res) );
  XOR2_X1 u_xor_module_3_U1 ( .A(p_rand_0), .B(io_i1_s1_d0), .Z(
        n_xor_module_3_res) );
  XOR2_X2 u_xor_module_4_U1 ( .A(p_rand_2), .B(n_xor_module_3_res), .Z(
        n_xor_module_4_res) );
  XOR2_X1 u_xor_module_5_U1 ( .A(p_rand_1), .B(io_i1_s2_d0), .Z(
        n_xor_module_5_res) );
  XOR2_X2 u_xor_module_6_U1 ( .A(p_rand_2), .B(n_xor_module_5_res), .Z(
        n_xor_module_6_res) );
  XOR2_X1 u_xor_module_7_U1 ( .A(p_rand_0), .B(io_i1_s0_d1), .Z(
        n_xor_module_7_res) );
  XOR2_X2 u_xor_module_8_U1 ( .A(p_rand_1), .B(n_xor_module_7_res), .Z(
        n_xor_module_8_res) );
  XOR2_X1 u_xor_module_9_U1 ( .A(p_rand_0), .B(io_i1_s1_d1), .Z(
        n_xor_module_9_res) );
  XOR2_X2 u_xor_module_10_U1 ( .A(p_rand_2), .B(n_xor_module_9_res), .Z(
        n_xor_module_10_res) );
  XOR2_X1 u_xor_module_11_U1 ( .A(p_rand_1), .B(io_i1_s2_d1), .Z(
        n_xor_module_11_res) );
  XOR2_X2 u_xor_module_12_U1 ( .A(p_rand_2), .B(n_xor_module_11_res), .Z(
        n_xor_module_12_res) );
  XOR2_X1 u_xor_module_13_U1 ( .A(p_rand_0), .B(io_i1_s0_d2), .Z(
        n_xor_module_13_res) );
  XOR2_X2 u_xor_module_14_U1 ( .A(p_rand_1), .B(n_xor_module_13_res), .Z(
        n_xor_module_14_res) );
  XOR2_X1 u_xor_module_15_U1 ( .A(p_rand_0), .B(io_i1_s1_d2), .Z(
        n_xor_module_15_res) );
  XOR2_X2 u_xor_module_16_U1 ( .A(p_rand_2), .B(n_xor_module_15_res), .Z(
        n_xor_module_16_res) );
  XOR2_X1 u_xor_module_17_U1 ( .A(p_rand_1), .B(io_i1_s2_d2), .Z(
        n_xor_module_17_res) );
  XOR2_X2 u_xor_module_18_U1 ( .A(p_rand_2), .B(n_xor_module_17_res), .Z(
        n_xor_module_18_res) );
  XOR2_X1 u_xor_module_19_U1 ( .A(p_rand_0), .B(io_i1_s0_d3), .Z(
        n_xor_module_19_res) );
  XOR2_X2 u_xor_module_20_U1 ( .A(p_rand_1), .B(n_xor_module_19_res), .Z(
        n_xor_module_20_res) );
  XOR2_X1 u_xor_module_21_U1 ( .A(p_rand_0), .B(io_i1_s1_d3), .Z(
        n_xor_module_21_res) );
  XOR2_X2 u_xor_module_22_U1 ( .A(p_rand_2), .B(n_xor_module_21_res), .Z(
        n_xor_module_22_res) );
  XOR2_X1 u_xor_module_23_U1 ( .A(p_rand_1), .B(io_i1_s2_d3), .Z(
        n_xor_module_23_res) );
  XOR2_X2 u_xor_module_24_U1 ( .A(p_rand_2), .B(n_xor_module_23_res), .Z(
        n_xor_module_24_res) );
  XOR2_X1 u_xor_module_25_U1 ( .A(p_rand_0), .B(io_i1_s0_d4), .Z(
        n_xor_module_25_res) );
  XOR2_X2 u_xor_module_26_U1 ( .A(p_rand_1), .B(n_xor_module_25_res), .Z(
        n_xor_module_26_res) );
  XOR2_X1 u_xor_module_27_U1 ( .A(p_rand_0), .B(io_i1_s1_d4), .Z(
        n_xor_module_27_res) );
  XOR2_X2 u_xor_module_28_U1 ( .A(p_rand_2), .B(n_xor_module_27_res), .Z(
        n_xor_module_28_res) );
  XOR2_X1 u_xor_module_29_U1 ( .A(p_rand_1), .B(io_i1_s2_d4), .Z(
        n_xor_module_29_res) );
  XOR2_X2 u_xor_module_30_U1 ( .A(p_rand_2), .B(n_xor_module_29_res), .Z(
        n_xor_module_30_res) );
  XOR2_X1 u_xor_module_31_U1 ( .A(p_rand_0), .B(io_i1_s0_d5), .Z(
        n_xor_module_31_res) );
  XOR2_X2 u_xor_module_32_U1 ( .A(p_rand_1), .B(n_xor_module_31_res), .Z(
        n_xor_module_32_res) );
  XOR2_X1 u_xor_module_33_U1 ( .A(p_rand_0), .B(io_i1_s1_d5), .Z(
        n_xor_module_33_res) );
  XOR2_X2 u_xor_module_34_U1 ( .A(p_rand_2), .B(n_xor_module_33_res), .Z(
        n_xor_module_34_res) );
  XOR2_X1 u_xor_module_35_U1 ( .A(p_rand_1), .B(io_i1_s2_d5), .Z(
        n_xor_module_35_res) );
  XOR2_X2 u_xor_module_36_U1 ( .A(p_rand_2), .B(n_xor_module_35_res), .Z(
        n_xor_module_36_res) );
  XOR2_X1 u_xor_module_37_U1 ( .A(p_rand_0), .B(io_i1_s0_d6), .Z(
        n_xor_module_37_res) );
  XOR2_X2 u_xor_module_38_U1 ( .A(p_rand_1), .B(n_xor_module_37_res), .Z(
        n_xor_module_38_res) );
  XOR2_X1 u_xor_module_39_U1 ( .A(p_rand_0), .B(io_i1_s1_d6), .Z(
        n_xor_module_39_res) );
  XOR2_X2 u_xor_module_40_U1 ( .A(p_rand_2), .B(n_xor_module_39_res), .Z(
        n_xor_module_40_res) );
  XOR2_X1 u_xor_module_41_U1 ( .A(p_rand_1), .B(io_i1_s2_d6), .Z(
        n_xor_module_41_res) );
  XOR2_X2 u_xor_module_42_U1 ( .A(p_rand_2), .B(n_xor_module_41_res), .Z(
        n_xor_module_42_res) );
  BUF_X1 u_majority7_module_0_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_0_n7) );
  BUF_X1 u_majority7_module_0_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_0_n6) );
  BUF_X1 u_majority7_module_0_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_0_n5) );
  BUF_X1 u_majority7_module_0_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_0_n4) );
  BUF_X1 u_majority7_module_0_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_0_n3) );
  BUF_X1 u_majority7_module_0_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_0_n2) );
  BUF_X1 u_majority7_module_0_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_0_n1) );
  AND2_X1 u_majority7_module_0__and_module_1_U1 ( .A1(n_majority7_module_0_n5), 
        .A2(n_majority7_module_0_n4), .ZN(
        n_majority7_module_0__and_module_1_res) );
  OR2_X1 u_majority7_module_0__or_module_1_U1 ( .A1(n_majority7_module_0_n4), 
        .A2(n_majority7_module_0_n5), .ZN(
        n_majority7_module_0__or_module_1_res) );
  AND2_X1 u_majority7_module_0__and_module_2_U1 ( .A1(n_majority7_module_0_n7), 
        .A2(n_majority7_module_0_n2), .ZN(
        n_majority7_module_0__and_module_2_res) );
  OR2_X1 u_majority7_module_0__or_module_2_U1 ( .A1(n_majority7_module_0_n2), 
        .A2(n_majority7_module_0_n7), .ZN(
        n_majority7_module_0__or_module_2_res) );
  AND2_X1 u_majority7_module_0__and_module_3_U1 ( .A1(n_majority7_module_0_n6), 
        .A2(n_majority7_module_0_n1), .ZN(
        n_majority7_module_0__and_module_3_res) );
  OR2_X1 u_majority7_module_0__or_module_3_U1 ( .A1(n_majority7_module_0_n1), 
        .A2(n_majority7_module_0_n6), .ZN(
        n_majority7_module_0__or_module_3_res) );
  AND2_X1 u_majority7_module_0__and_module_4_U1 ( .A1(
        n_majority7_module_0__and_module_2_res), .A2(
        n_majority7_module_0__and_module_1_res), .ZN(
        n_majority7_module_0__and_module_4_res) );
  OR2_X1 u_majority7_module_0__or_module_4_U1 ( .A1(
        n_majority7_module_0__and_module_1_res), .A2(
        n_majority7_module_0__and_module_2_res), .ZN(
        n_majority7_module_0__or_module_4_res) );
  AND2_X1 u_majority7_module_0__and_module_5_U1 ( .A1(
        n_majority7_module_0__and_module_3_res), .A2(n_majority7_module_0_n3), 
        .ZN(n_majority7_module_0__and_module_5_res) );
  OR2_X1 u_majority7_module_0__or_module_5_U1 ( .A1(n_majority7_module_0_n3), 
        .A2(n_majority7_module_0__and_module_3_res), .ZN(
        n_majority7_module_0__or_module_5_res) );
  AND2_X1 u_majority7_module_0__and_module_6_U1 ( .A1(
        n_majority7_module_0__or_module_1_res), .A2(
        n_majority7_module_0__or_module_2_res), .ZN(
        n_majority7_module_0__and_module_6_res) );
  OR2_X1 u_majority7_module_0__or_module_6_U1 ( .A1(
        n_majority7_module_0__or_module_2_res), .A2(
        n_majority7_module_0__or_module_1_res), .ZN(
        n_majority7_module_0__or_module_6_res) );
  OR2_X1 u_majority7_module_0__or_module_7_U1 ( .A1(
        n_majority7_module_0__and_module_4_res), .A2(
        n_majority7_module_0__and_module_5_res), .ZN(
        n_majority7_module_0__or_module_7_res) );
  AND2_X1 u_majority7_module_0__and_module_7_U1 ( .A1(
        n_majority7_module_0__or_module_3_res), .A2(
        n_majority7_module_0__or_module_4_res), .ZN(
        n_majority7_module_0__and_module_7_res) );
  OR2_X1 u_majority7_module_0__or_module_8_U1 ( .A1(
        n_majority7_module_0__or_module_4_res), .A2(
        n_majority7_module_0__or_module_3_res), .ZN(
        n_majority7_module_0__or_module_8_res) );
  AND2_X1 u_majority7_module_0__and_module_8_U1 ( .A1(
        n_majority7_module_0__or_module_5_res), .A2(
        n_majority7_module_0__and_module_6_res), .ZN(
        n_majority7_module_0__and_module_8_res) );
  OR2_X1 u_majority7_module_0__or_module_9_U1 ( .A1(
        n_majority7_module_0__and_module_6_res), .A2(
        n_majority7_module_0__or_module_5_res), .ZN(
        n_majority7_module_0__or_module_9_res) );
  OR2_X1 u_majority7_module_0__or_module_10_U1 ( .A1(
        n_majority7_module_0__or_module_7_res), .A2(
        n_majority7_module_0__and_module_7_res), .ZN(
        n_majority7_module_0__or_module_10_res) );
  AND2_X1 u_majority7_module_0__and_module_9_U1 ( .A1(
        n_majority7_module_0__or_module_6_res), .A2(
        n_majority7_module_0__or_module_9_res), .ZN(
        n_majority7_module_0__and_module_9_res) );
  OR2_X1 u_majority7_module_0__or_module_11_U1 ( .A1(
        n_majority7_module_0__or_module_10_res), .A2(
        n_majority7_module_0__and_module_8_res), .ZN(
        n_majority7_module_0__or_module_11_res) );
  AND2_X1 u_majority7_module_0__and_module_10_U1 ( .A1(
        n_majority7_module_0__or_module_8_res), .A2(
        n_majority7_module_0__and_module_9_res), .ZN(
        n_majority7_module_0__and_module_10_res) );
  AND2_X1 u_majority7_module_0__and_module_11_U1 ( .A1(
        n_majority7_module_0__and_module_10_res), .A2(
        n_majority7_module_0__or_module_11_res), .ZN(n_majority7_module_0_res)
         );
  DFF_X1 u_reg_module_1__cini_mul_v000_reg ( .D(n_majority7_module_0_res), 
        .CK(clock_0), .Q(n_reg_module_1_res), .QN() );
  BUF_X1 u_majority7_module_1_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_1_n7) );
  BUF_X1 u_majority7_module_1_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_1_n6) );
  BUF_X1 u_majority7_module_1_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_1_n5) );
  BUF_X1 u_majority7_module_1_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_1_n4) );
  BUF_X1 u_majority7_module_1_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_1_n3) );
  BUF_X1 u_majority7_module_1_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_1_n2) );
  BUF_X1 u_majority7_module_1_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_1_n1) );
  AND2_X1 u_majority7_module_1__and_module_1_U1 ( .A1(n_majority7_module_1_n5), 
        .A2(n_majority7_module_1_n4), .ZN(
        n_majority7_module_1__and_module_1_res) );
  OR2_X1 u_majority7_module_1__or_module_1_U1 ( .A1(n_majority7_module_1_n4), 
        .A2(n_majority7_module_1_n5), .ZN(
        n_majority7_module_1__or_module_1_res) );
  AND2_X1 u_majority7_module_1__and_module_2_U1 ( .A1(n_majority7_module_1_n7), 
        .A2(n_majority7_module_1_n2), .ZN(
        n_majority7_module_1__and_module_2_res) );
  OR2_X1 u_majority7_module_1__or_module_2_U1 ( .A1(n_majority7_module_1_n2), 
        .A2(n_majority7_module_1_n7), .ZN(
        n_majority7_module_1__or_module_2_res) );
  AND2_X1 u_majority7_module_1__and_module_3_U1 ( .A1(n_majority7_module_1_n6), 
        .A2(n_majority7_module_1_n1), .ZN(
        n_majority7_module_1__and_module_3_res) );
  OR2_X1 u_majority7_module_1__or_module_3_U1 ( .A1(n_majority7_module_1_n1), 
        .A2(n_majority7_module_1_n6), .ZN(
        n_majority7_module_1__or_module_3_res) );
  AND2_X1 u_majority7_module_1__and_module_4_U1 ( .A1(
        n_majority7_module_1__and_module_2_res), .A2(
        n_majority7_module_1__and_module_1_res), .ZN(
        n_majority7_module_1__and_module_4_res) );
  OR2_X1 u_majority7_module_1__or_module_4_U1 ( .A1(
        n_majority7_module_1__and_module_1_res), .A2(
        n_majority7_module_1__and_module_2_res), .ZN(
        n_majority7_module_1__or_module_4_res) );
  AND2_X1 u_majority7_module_1__and_module_5_U1 ( .A1(
        n_majority7_module_1__and_module_3_res), .A2(n_majority7_module_1_n3), 
        .ZN(n_majority7_module_1__and_module_5_res) );
  OR2_X1 u_majority7_module_1__or_module_5_U1 ( .A1(n_majority7_module_1_n3), 
        .A2(n_majority7_module_1__and_module_3_res), .ZN(
        n_majority7_module_1__or_module_5_res) );
  AND2_X1 u_majority7_module_1__and_module_6_U1 ( .A1(
        n_majority7_module_1__or_module_1_res), .A2(
        n_majority7_module_1__or_module_2_res), .ZN(
        n_majority7_module_1__and_module_6_res) );
  OR2_X1 u_majority7_module_1__or_module_6_U1 ( .A1(
        n_majority7_module_1__or_module_2_res), .A2(
        n_majority7_module_1__or_module_1_res), .ZN(
        n_majority7_module_1__or_module_6_res) );
  OR2_X1 u_majority7_module_1__or_module_7_U1 ( .A1(
        n_majority7_module_1__and_module_4_res), .A2(
        n_majority7_module_1__and_module_5_res), .ZN(
        n_majority7_module_1__or_module_7_res) );
  AND2_X1 u_majority7_module_1__and_module_7_U1 ( .A1(
        n_majority7_module_1__or_module_3_res), .A2(
        n_majority7_module_1__or_module_4_res), .ZN(
        n_majority7_module_1__and_module_7_res) );
  OR2_X1 u_majority7_module_1__or_module_8_U1 ( .A1(
        n_majority7_module_1__or_module_4_res), .A2(
        n_majority7_module_1__or_module_3_res), .ZN(
        n_majority7_module_1__or_module_8_res) );
  AND2_X1 u_majority7_module_1__and_module_8_U1 ( .A1(
        n_majority7_module_1__or_module_5_res), .A2(
        n_majority7_module_1__and_module_6_res), .ZN(
        n_majority7_module_1__and_module_8_res) );
  OR2_X1 u_majority7_module_1__or_module_9_U1 ( .A1(
        n_majority7_module_1__and_module_6_res), .A2(
        n_majority7_module_1__or_module_5_res), .ZN(
        n_majority7_module_1__or_module_9_res) );
  OR2_X1 u_majority7_module_1__or_module_10_U1 ( .A1(
        n_majority7_module_1__or_module_7_res), .A2(
        n_majority7_module_1__and_module_7_res), .ZN(
        n_majority7_module_1__or_module_10_res) );
  AND2_X1 u_majority7_module_1__and_module_9_U1 ( .A1(
        n_majority7_module_1__or_module_6_res), .A2(
        n_majority7_module_1__or_module_9_res), .ZN(
        n_majority7_module_1__and_module_9_res) );
  OR2_X1 u_majority7_module_1__or_module_11_U1 ( .A1(
        n_majority7_module_1__or_module_10_res), .A2(
        n_majority7_module_1__and_module_8_res), .ZN(
        n_majority7_module_1__or_module_11_res) );
  AND2_X1 u_majority7_module_1__and_module_10_U1 ( .A1(
        n_majority7_module_1__or_module_8_res), .A2(
        n_majority7_module_1__and_module_9_res), .ZN(
        n_majority7_module_1__and_module_10_res) );
  AND2_X1 u_majority7_module_1__and_module_11_U1 ( .A1(
        n_majority7_module_1__and_module_10_res), .A2(
        n_majority7_module_1__or_module_11_res), .ZN(n_majority7_module_1_res)
         );
  DFF_X1 u_reg_module_2__cini_mul_v000_reg ( .D(n_majority7_module_1_res), 
        .CK(clock_0), .Q(n_reg_module_2_res), .QN() );
  BUF_X1 u_majority7_module_2_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_2_n7) );
  BUF_X1 u_majority7_module_2_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_2_n6) );
  BUF_X1 u_majority7_module_2_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_2_n5) );
  BUF_X1 u_majority7_module_2_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_2_n4) );
  BUF_X1 u_majority7_module_2_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_2_n3) );
  BUF_X1 u_majority7_module_2_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_2_n2) );
  BUF_X1 u_majority7_module_2_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_2_n1) );
  AND2_X1 u_majority7_module_2__and_module_1_U1 ( .A1(n_majority7_module_2_n5), 
        .A2(n_majority7_module_2_n4), .ZN(
        n_majority7_module_2__and_module_1_res) );
  OR2_X1 u_majority7_module_2__or_module_1_U1 ( .A1(n_majority7_module_2_n4), 
        .A2(n_majority7_module_2_n5), .ZN(
        n_majority7_module_2__or_module_1_res) );
  AND2_X1 u_majority7_module_2__and_module_2_U1 ( .A1(n_majority7_module_2_n7), 
        .A2(n_majority7_module_2_n2), .ZN(
        n_majority7_module_2__and_module_2_res) );
  OR2_X1 u_majority7_module_2__or_module_2_U1 ( .A1(n_majority7_module_2_n2), 
        .A2(n_majority7_module_2_n7), .ZN(
        n_majority7_module_2__or_module_2_res) );
  AND2_X1 u_majority7_module_2__and_module_3_U1 ( .A1(n_majority7_module_2_n6), 
        .A2(n_majority7_module_2_n1), .ZN(
        n_majority7_module_2__and_module_3_res) );
  OR2_X1 u_majority7_module_2__or_module_3_U1 ( .A1(n_majority7_module_2_n1), 
        .A2(n_majority7_module_2_n6), .ZN(
        n_majority7_module_2__or_module_3_res) );
  AND2_X1 u_majority7_module_2__and_module_4_U1 ( .A1(
        n_majority7_module_2__and_module_2_res), .A2(
        n_majority7_module_2__and_module_1_res), .ZN(
        n_majority7_module_2__and_module_4_res) );
  OR2_X1 u_majority7_module_2__or_module_4_U1 ( .A1(
        n_majority7_module_2__and_module_1_res), .A2(
        n_majority7_module_2__and_module_2_res), .ZN(
        n_majority7_module_2__or_module_4_res) );
  AND2_X1 u_majority7_module_2__and_module_5_U1 ( .A1(
        n_majority7_module_2__and_module_3_res), .A2(n_majority7_module_2_n3), 
        .ZN(n_majority7_module_2__and_module_5_res) );
  OR2_X1 u_majority7_module_2__or_module_5_U1 ( .A1(n_majority7_module_2_n3), 
        .A2(n_majority7_module_2__and_module_3_res), .ZN(
        n_majority7_module_2__or_module_5_res) );
  AND2_X1 u_majority7_module_2__and_module_6_U1 ( .A1(
        n_majority7_module_2__or_module_1_res), .A2(
        n_majority7_module_2__or_module_2_res), .ZN(
        n_majority7_module_2__and_module_6_res) );
  OR2_X1 u_majority7_module_2__or_module_6_U1 ( .A1(
        n_majority7_module_2__or_module_2_res), .A2(
        n_majority7_module_2__or_module_1_res), .ZN(
        n_majority7_module_2__or_module_6_res) );
  OR2_X1 u_majority7_module_2__or_module_7_U1 ( .A1(
        n_majority7_module_2__and_module_4_res), .A2(
        n_majority7_module_2__and_module_5_res), .ZN(
        n_majority7_module_2__or_module_7_res) );
  AND2_X1 u_majority7_module_2__and_module_7_U1 ( .A1(
        n_majority7_module_2__or_module_3_res), .A2(
        n_majority7_module_2__or_module_4_res), .ZN(
        n_majority7_module_2__and_module_7_res) );
  OR2_X1 u_majority7_module_2__or_module_8_U1 ( .A1(
        n_majority7_module_2__or_module_4_res), .A2(
        n_majority7_module_2__or_module_3_res), .ZN(
        n_majority7_module_2__or_module_8_res) );
  AND2_X1 u_majority7_module_2__and_module_8_U1 ( .A1(
        n_majority7_module_2__or_module_5_res), .A2(
        n_majority7_module_2__and_module_6_res), .ZN(
        n_majority7_module_2__and_module_8_res) );
  OR2_X1 u_majority7_module_2__or_module_9_U1 ( .A1(
        n_majority7_module_2__and_module_6_res), .A2(
        n_majority7_module_2__or_module_5_res), .ZN(
        n_majority7_module_2__or_module_9_res) );
  OR2_X1 u_majority7_module_2__or_module_10_U1 ( .A1(
        n_majority7_module_2__or_module_7_res), .A2(
        n_majority7_module_2__and_module_7_res), .ZN(
        n_majority7_module_2__or_module_10_res) );
  AND2_X1 u_majority7_module_2__and_module_9_U1 ( .A1(
        n_majority7_module_2__or_module_6_res), .A2(
        n_majority7_module_2__or_module_9_res), .ZN(
        n_majority7_module_2__and_module_9_res) );
  OR2_X1 u_majority7_module_2__or_module_11_U1 ( .A1(
        n_majority7_module_2__or_module_10_res), .A2(
        n_majority7_module_2__and_module_8_res), .ZN(
        n_majority7_module_2__or_module_11_res) );
  AND2_X1 u_majority7_module_2__and_module_10_U1 ( .A1(
        n_majority7_module_2__or_module_8_res), .A2(
        n_majority7_module_2__and_module_9_res), .ZN(
        n_majority7_module_2__and_module_10_res) );
  AND2_X1 u_majority7_module_2__and_module_11_U1 ( .A1(
        n_majority7_module_2__and_module_10_res), .A2(
        n_majority7_module_2__or_module_11_res), .ZN(n_majority7_module_2_res)
         );
  DFF_X1 u_reg_module_3__cini_mul_v000_reg ( .D(n_majority7_module_2_res), 
        .CK(clock_0), .Q(n_reg_module_3_res), .QN() );
  BUF_X1 u_majority7_module_3_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_3_n7) );
  BUF_X1 u_majority7_module_3_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_3_n6) );
  BUF_X1 u_majority7_module_3_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_3_n5) );
  BUF_X1 u_majority7_module_3_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_3_n4) );
  BUF_X1 u_majority7_module_3_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_3_n3) );
  BUF_X1 u_majority7_module_3_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_3_n2) );
  BUF_X1 u_majority7_module_3_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_3_n1) );
  AND2_X1 u_majority7_module_3__and_module_1_U1 ( .A1(n_majority7_module_3_n5), 
        .A2(n_majority7_module_3_n4), .ZN(
        n_majority7_module_3__and_module_1_res) );
  OR2_X1 u_majority7_module_3__or_module_1_U1 ( .A1(n_majority7_module_3_n4), 
        .A2(n_majority7_module_3_n5), .ZN(
        n_majority7_module_3__or_module_1_res) );
  AND2_X1 u_majority7_module_3__and_module_2_U1 ( .A1(n_majority7_module_3_n7), 
        .A2(n_majority7_module_3_n2), .ZN(
        n_majority7_module_3__and_module_2_res) );
  OR2_X1 u_majority7_module_3__or_module_2_U1 ( .A1(n_majority7_module_3_n2), 
        .A2(n_majority7_module_3_n7), .ZN(
        n_majority7_module_3__or_module_2_res) );
  AND2_X1 u_majority7_module_3__and_module_3_U1 ( .A1(n_majority7_module_3_n6), 
        .A2(n_majority7_module_3_n1), .ZN(
        n_majority7_module_3__and_module_3_res) );
  OR2_X1 u_majority7_module_3__or_module_3_U1 ( .A1(n_majority7_module_3_n1), 
        .A2(n_majority7_module_3_n6), .ZN(
        n_majority7_module_3__or_module_3_res) );
  AND2_X1 u_majority7_module_3__and_module_4_U1 ( .A1(
        n_majority7_module_3__and_module_2_res), .A2(
        n_majority7_module_3__and_module_1_res), .ZN(
        n_majority7_module_3__and_module_4_res) );
  OR2_X1 u_majority7_module_3__or_module_4_U1 ( .A1(
        n_majority7_module_3__and_module_1_res), .A2(
        n_majority7_module_3__and_module_2_res), .ZN(
        n_majority7_module_3__or_module_4_res) );
  AND2_X1 u_majority7_module_3__and_module_5_U1 ( .A1(
        n_majority7_module_3__and_module_3_res), .A2(n_majority7_module_3_n3), 
        .ZN(n_majority7_module_3__and_module_5_res) );
  OR2_X1 u_majority7_module_3__or_module_5_U1 ( .A1(n_majority7_module_3_n3), 
        .A2(n_majority7_module_3__and_module_3_res), .ZN(
        n_majority7_module_3__or_module_5_res) );
  AND2_X1 u_majority7_module_3__and_module_6_U1 ( .A1(
        n_majority7_module_3__or_module_1_res), .A2(
        n_majority7_module_3__or_module_2_res), .ZN(
        n_majority7_module_3__and_module_6_res) );
  OR2_X1 u_majority7_module_3__or_module_6_U1 ( .A1(
        n_majority7_module_3__or_module_2_res), .A2(
        n_majority7_module_3__or_module_1_res), .ZN(
        n_majority7_module_3__or_module_6_res) );
  OR2_X1 u_majority7_module_3__or_module_7_U1 ( .A1(
        n_majority7_module_3__and_module_4_res), .A2(
        n_majority7_module_3__and_module_5_res), .ZN(
        n_majority7_module_3__or_module_7_res) );
  AND2_X1 u_majority7_module_3__and_module_7_U1 ( .A1(
        n_majority7_module_3__or_module_3_res), .A2(
        n_majority7_module_3__or_module_4_res), .ZN(
        n_majority7_module_3__and_module_7_res) );
  OR2_X1 u_majority7_module_3__or_module_8_U1 ( .A1(
        n_majority7_module_3__or_module_4_res), .A2(
        n_majority7_module_3__or_module_3_res), .ZN(
        n_majority7_module_3__or_module_8_res) );
  AND2_X1 u_majority7_module_3__and_module_8_U1 ( .A1(
        n_majority7_module_3__or_module_5_res), .A2(
        n_majority7_module_3__and_module_6_res), .ZN(
        n_majority7_module_3__and_module_8_res) );
  OR2_X1 u_majority7_module_3__or_module_9_U1 ( .A1(
        n_majority7_module_3__and_module_6_res), .A2(
        n_majority7_module_3__or_module_5_res), .ZN(
        n_majority7_module_3__or_module_9_res) );
  OR2_X1 u_majority7_module_3__or_module_10_U1 ( .A1(
        n_majority7_module_3__or_module_7_res), .A2(
        n_majority7_module_3__and_module_7_res), .ZN(
        n_majority7_module_3__or_module_10_res) );
  AND2_X1 u_majority7_module_3__and_module_9_U1 ( .A1(
        n_majority7_module_3__or_module_6_res), .A2(
        n_majority7_module_3__or_module_9_res), .ZN(
        n_majority7_module_3__and_module_9_res) );
  OR2_X1 u_majority7_module_3__or_module_11_U1 ( .A1(
        n_majority7_module_3__or_module_10_res), .A2(
        n_majority7_module_3__and_module_8_res), .ZN(
        n_majority7_module_3__or_module_11_res) );
  AND2_X1 u_majority7_module_3__and_module_10_U1 ( .A1(
        n_majority7_module_3__or_module_8_res), .A2(
        n_majority7_module_3__and_module_9_res), .ZN(
        n_majority7_module_3__and_module_10_res) );
  AND2_X1 u_majority7_module_3__and_module_11_U1 ( .A1(
        n_majority7_module_3__and_module_10_res), .A2(
        n_majority7_module_3__or_module_11_res), .ZN(n_majority7_module_3_res)
         );
  DFF_X1 u_reg_module_4__cini_mul_v000_reg ( .D(n_majority7_module_3_res), 
        .CK(clock_0), .Q(n_reg_module_4_res), .QN() );
  BUF_X1 u_majority7_module_4_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_4_n7) );
  BUF_X1 u_majority7_module_4_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_4_n6) );
  BUF_X1 u_majority7_module_4_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_4_n5) );
  BUF_X1 u_majority7_module_4_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_4_n4) );
  BUF_X1 u_majority7_module_4_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_4_n3) );
  BUF_X1 u_majority7_module_4_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_4_n2) );
  BUF_X1 u_majority7_module_4_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_4_n1) );
  AND2_X1 u_majority7_module_4__and_module_1_U1 ( .A1(n_majority7_module_4_n5), 
        .A2(n_majority7_module_4_n4), .ZN(
        n_majority7_module_4__and_module_1_res) );
  OR2_X1 u_majority7_module_4__or_module_1_U1 ( .A1(n_majority7_module_4_n4), 
        .A2(n_majority7_module_4_n5), .ZN(
        n_majority7_module_4__or_module_1_res) );
  AND2_X1 u_majority7_module_4__and_module_2_U1 ( .A1(n_majority7_module_4_n7), 
        .A2(n_majority7_module_4_n2), .ZN(
        n_majority7_module_4__and_module_2_res) );
  OR2_X1 u_majority7_module_4__or_module_2_U1 ( .A1(n_majority7_module_4_n2), 
        .A2(n_majority7_module_4_n7), .ZN(
        n_majority7_module_4__or_module_2_res) );
  AND2_X1 u_majority7_module_4__and_module_3_U1 ( .A1(n_majority7_module_4_n6), 
        .A2(n_majority7_module_4_n1), .ZN(
        n_majority7_module_4__and_module_3_res) );
  OR2_X1 u_majority7_module_4__or_module_3_U1 ( .A1(n_majority7_module_4_n1), 
        .A2(n_majority7_module_4_n6), .ZN(
        n_majority7_module_4__or_module_3_res) );
  AND2_X1 u_majority7_module_4__and_module_4_U1 ( .A1(
        n_majority7_module_4__and_module_2_res), .A2(
        n_majority7_module_4__and_module_1_res), .ZN(
        n_majority7_module_4__and_module_4_res) );
  OR2_X1 u_majority7_module_4__or_module_4_U1 ( .A1(
        n_majority7_module_4__and_module_1_res), .A2(
        n_majority7_module_4__and_module_2_res), .ZN(
        n_majority7_module_4__or_module_4_res) );
  AND2_X1 u_majority7_module_4__and_module_5_U1 ( .A1(
        n_majority7_module_4__and_module_3_res), .A2(n_majority7_module_4_n3), 
        .ZN(n_majority7_module_4__and_module_5_res) );
  OR2_X1 u_majority7_module_4__or_module_5_U1 ( .A1(n_majority7_module_4_n3), 
        .A2(n_majority7_module_4__and_module_3_res), .ZN(
        n_majority7_module_4__or_module_5_res) );
  AND2_X1 u_majority7_module_4__and_module_6_U1 ( .A1(
        n_majority7_module_4__or_module_1_res), .A2(
        n_majority7_module_4__or_module_2_res), .ZN(
        n_majority7_module_4__and_module_6_res) );
  OR2_X1 u_majority7_module_4__or_module_6_U1 ( .A1(
        n_majority7_module_4__or_module_2_res), .A2(
        n_majority7_module_4__or_module_1_res), .ZN(
        n_majority7_module_4__or_module_6_res) );
  OR2_X1 u_majority7_module_4__or_module_7_U1 ( .A1(
        n_majority7_module_4__and_module_4_res), .A2(
        n_majority7_module_4__and_module_5_res), .ZN(
        n_majority7_module_4__or_module_7_res) );
  AND2_X1 u_majority7_module_4__and_module_7_U1 ( .A1(
        n_majority7_module_4__or_module_3_res), .A2(
        n_majority7_module_4__or_module_4_res), .ZN(
        n_majority7_module_4__and_module_7_res) );
  OR2_X1 u_majority7_module_4__or_module_8_U1 ( .A1(
        n_majority7_module_4__or_module_4_res), .A2(
        n_majority7_module_4__or_module_3_res), .ZN(
        n_majority7_module_4__or_module_8_res) );
  AND2_X1 u_majority7_module_4__and_module_8_U1 ( .A1(
        n_majority7_module_4__or_module_5_res), .A2(
        n_majority7_module_4__and_module_6_res), .ZN(
        n_majority7_module_4__and_module_8_res) );
  OR2_X1 u_majority7_module_4__or_module_9_U1 ( .A1(
        n_majority7_module_4__and_module_6_res), .A2(
        n_majority7_module_4__or_module_5_res), .ZN(
        n_majority7_module_4__or_module_9_res) );
  OR2_X1 u_majority7_module_4__or_module_10_U1 ( .A1(
        n_majority7_module_4__or_module_7_res), .A2(
        n_majority7_module_4__and_module_7_res), .ZN(
        n_majority7_module_4__or_module_10_res) );
  AND2_X1 u_majority7_module_4__and_module_9_U1 ( .A1(
        n_majority7_module_4__or_module_6_res), .A2(
        n_majority7_module_4__or_module_9_res), .ZN(
        n_majority7_module_4__and_module_9_res) );
  OR2_X1 u_majority7_module_4__or_module_11_U1 ( .A1(
        n_majority7_module_4__or_module_10_res), .A2(
        n_majority7_module_4__and_module_8_res), .ZN(
        n_majority7_module_4__or_module_11_res) );
  AND2_X1 u_majority7_module_4__and_module_10_U1 ( .A1(
        n_majority7_module_4__or_module_8_res), .A2(
        n_majority7_module_4__and_module_9_res), .ZN(
        n_majority7_module_4__and_module_10_res) );
  AND2_X1 u_majority7_module_4__and_module_11_U1 ( .A1(
        n_majority7_module_4__and_module_10_res), .A2(
        n_majority7_module_4__or_module_11_res), .ZN(n_majority7_module_4_res)
         );
  DFF_X1 u_reg_module_5__cini_mul_v000_reg ( .D(n_majority7_module_4_res), 
        .CK(clock_0), .Q(n_reg_module_5_res), .QN() );
  BUF_X1 u_majority7_module_5_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_5_n7) );
  BUF_X1 u_majority7_module_5_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_5_n6) );
  BUF_X1 u_majority7_module_5_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_5_n5) );
  BUF_X1 u_majority7_module_5_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_5_n4) );
  BUF_X1 u_majority7_module_5_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_5_n3) );
  BUF_X1 u_majority7_module_5_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_5_n2) );
  BUF_X1 u_majority7_module_5_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_5_n1) );
  AND2_X1 u_majority7_module_5__and_module_1_U1 ( .A1(n_majority7_module_5_n5), 
        .A2(n_majority7_module_5_n4), .ZN(
        n_majority7_module_5__and_module_1_res) );
  OR2_X1 u_majority7_module_5__or_module_1_U1 ( .A1(n_majority7_module_5_n4), 
        .A2(n_majority7_module_5_n5), .ZN(
        n_majority7_module_5__or_module_1_res) );
  AND2_X1 u_majority7_module_5__and_module_2_U1 ( .A1(n_majority7_module_5_n7), 
        .A2(n_majority7_module_5_n2), .ZN(
        n_majority7_module_5__and_module_2_res) );
  OR2_X1 u_majority7_module_5__or_module_2_U1 ( .A1(n_majority7_module_5_n2), 
        .A2(n_majority7_module_5_n7), .ZN(
        n_majority7_module_5__or_module_2_res) );
  AND2_X1 u_majority7_module_5__and_module_3_U1 ( .A1(n_majority7_module_5_n6), 
        .A2(n_majority7_module_5_n1), .ZN(
        n_majority7_module_5__and_module_3_res) );
  OR2_X1 u_majority7_module_5__or_module_3_U1 ( .A1(n_majority7_module_5_n1), 
        .A2(n_majority7_module_5_n6), .ZN(
        n_majority7_module_5__or_module_3_res) );
  AND2_X1 u_majority7_module_5__and_module_4_U1 ( .A1(
        n_majority7_module_5__and_module_2_res), .A2(
        n_majority7_module_5__and_module_1_res), .ZN(
        n_majority7_module_5__and_module_4_res) );
  OR2_X1 u_majority7_module_5__or_module_4_U1 ( .A1(
        n_majority7_module_5__and_module_1_res), .A2(
        n_majority7_module_5__and_module_2_res), .ZN(
        n_majority7_module_5__or_module_4_res) );
  AND2_X1 u_majority7_module_5__and_module_5_U1 ( .A1(
        n_majority7_module_5__and_module_3_res), .A2(n_majority7_module_5_n3), 
        .ZN(n_majority7_module_5__and_module_5_res) );
  OR2_X1 u_majority7_module_5__or_module_5_U1 ( .A1(n_majority7_module_5_n3), 
        .A2(n_majority7_module_5__and_module_3_res), .ZN(
        n_majority7_module_5__or_module_5_res) );
  AND2_X1 u_majority7_module_5__and_module_6_U1 ( .A1(
        n_majority7_module_5__or_module_1_res), .A2(
        n_majority7_module_5__or_module_2_res), .ZN(
        n_majority7_module_5__and_module_6_res) );
  OR2_X1 u_majority7_module_5__or_module_6_U1 ( .A1(
        n_majority7_module_5__or_module_2_res), .A2(
        n_majority7_module_5__or_module_1_res), .ZN(
        n_majority7_module_5__or_module_6_res) );
  OR2_X1 u_majority7_module_5__or_module_7_U1 ( .A1(
        n_majority7_module_5__and_module_4_res), .A2(
        n_majority7_module_5__and_module_5_res), .ZN(
        n_majority7_module_5__or_module_7_res) );
  AND2_X1 u_majority7_module_5__and_module_7_U1 ( .A1(
        n_majority7_module_5__or_module_3_res), .A2(
        n_majority7_module_5__or_module_4_res), .ZN(
        n_majority7_module_5__and_module_7_res) );
  OR2_X1 u_majority7_module_5__or_module_8_U1 ( .A1(
        n_majority7_module_5__or_module_4_res), .A2(
        n_majority7_module_5__or_module_3_res), .ZN(
        n_majority7_module_5__or_module_8_res) );
  AND2_X1 u_majority7_module_5__and_module_8_U1 ( .A1(
        n_majority7_module_5__or_module_5_res), .A2(
        n_majority7_module_5__and_module_6_res), .ZN(
        n_majority7_module_5__and_module_8_res) );
  OR2_X1 u_majority7_module_5__or_module_9_U1 ( .A1(
        n_majority7_module_5__and_module_6_res), .A2(
        n_majority7_module_5__or_module_5_res), .ZN(
        n_majority7_module_5__or_module_9_res) );
  OR2_X1 u_majority7_module_5__or_module_10_U1 ( .A1(
        n_majority7_module_5__or_module_7_res), .A2(
        n_majority7_module_5__and_module_7_res), .ZN(
        n_majority7_module_5__or_module_10_res) );
  AND2_X1 u_majority7_module_5__and_module_9_U1 ( .A1(
        n_majority7_module_5__or_module_6_res), .A2(
        n_majority7_module_5__or_module_9_res), .ZN(
        n_majority7_module_5__and_module_9_res) );
  OR2_X1 u_majority7_module_5__or_module_11_U1 ( .A1(
        n_majority7_module_5__or_module_10_res), .A2(
        n_majority7_module_5__and_module_8_res), .ZN(
        n_majority7_module_5__or_module_11_res) );
  AND2_X1 u_majority7_module_5__and_module_10_U1 ( .A1(
        n_majority7_module_5__or_module_8_res), .A2(
        n_majority7_module_5__and_module_9_res), .ZN(
        n_majority7_module_5__and_module_10_res) );
  AND2_X1 u_majority7_module_5__and_module_11_U1 ( .A1(
        n_majority7_module_5__and_module_10_res), .A2(
        n_majority7_module_5__or_module_11_res), .ZN(n_majority7_module_5_res)
         );
  DFF_X1 u_reg_module_6__cini_mul_v000_reg ( .D(n_majority7_module_5_res), 
        .CK(clock_0), .Q(n_reg_module_6_res), .QN() );
  BUF_X1 u_majority7_module_6_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_6_n7) );
  BUF_X1 u_majority7_module_6_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_6_n6) );
  BUF_X1 u_majority7_module_6_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_6_n5) );
  BUF_X1 u_majority7_module_6_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_6_n4) );
  BUF_X1 u_majority7_module_6_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_6_n3) );
  BUF_X1 u_majority7_module_6_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_6_n2) );
  BUF_X1 u_majority7_module_6_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_6_n1) );
  AND2_X1 u_majority7_module_6__and_module_1_U1 ( .A1(n_majority7_module_6_n5), 
        .A2(n_majority7_module_6_n4), .ZN(
        n_majority7_module_6__and_module_1_res) );
  OR2_X1 u_majority7_module_6__or_module_1_U1 ( .A1(n_majority7_module_6_n4), 
        .A2(n_majority7_module_6_n5), .ZN(
        n_majority7_module_6__or_module_1_res) );
  AND2_X1 u_majority7_module_6__and_module_2_U1 ( .A1(n_majority7_module_6_n7), 
        .A2(n_majority7_module_6_n2), .ZN(
        n_majority7_module_6__and_module_2_res) );
  OR2_X1 u_majority7_module_6__or_module_2_U1 ( .A1(n_majority7_module_6_n2), 
        .A2(n_majority7_module_6_n7), .ZN(
        n_majority7_module_6__or_module_2_res) );
  AND2_X1 u_majority7_module_6__and_module_3_U1 ( .A1(n_majority7_module_6_n6), 
        .A2(n_majority7_module_6_n1), .ZN(
        n_majority7_module_6__and_module_3_res) );
  OR2_X1 u_majority7_module_6__or_module_3_U1 ( .A1(n_majority7_module_6_n1), 
        .A2(n_majority7_module_6_n6), .ZN(
        n_majority7_module_6__or_module_3_res) );
  AND2_X1 u_majority7_module_6__and_module_4_U1 ( .A1(
        n_majority7_module_6__and_module_2_res), .A2(
        n_majority7_module_6__and_module_1_res), .ZN(
        n_majority7_module_6__and_module_4_res) );
  OR2_X1 u_majority7_module_6__or_module_4_U1 ( .A1(
        n_majority7_module_6__and_module_1_res), .A2(
        n_majority7_module_6__and_module_2_res), .ZN(
        n_majority7_module_6__or_module_4_res) );
  AND2_X1 u_majority7_module_6__and_module_5_U1 ( .A1(
        n_majority7_module_6__and_module_3_res), .A2(n_majority7_module_6_n3), 
        .ZN(n_majority7_module_6__and_module_5_res) );
  OR2_X1 u_majority7_module_6__or_module_5_U1 ( .A1(n_majority7_module_6_n3), 
        .A2(n_majority7_module_6__and_module_3_res), .ZN(
        n_majority7_module_6__or_module_5_res) );
  AND2_X1 u_majority7_module_6__and_module_6_U1 ( .A1(
        n_majority7_module_6__or_module_1_res), .A2(
        n_majority7_module_6__or_module_2_res), .ZN(
        n_majority7_module_6__and_module_6_res) );
  OR2_X1 u_majority7_module_6__or_module_6_U1 ( .A1(
        n_majority7_module_6__or_module_2_res), .A2(
        n_majority7_module_6__or_module_1_res), .ZN(
        n_majority7_module_6__or_module_6_res) );
  OR2_X1 u_majority7_module_6__or_module_7_U1 ( .A1(
        n_majority7_module_6__and_module_4_res), .A2(
        n_majority7_module_6__and_module_5_res), .ZN(
        n_majority7_module_6__or_module_7_res) );
  AND2_X1 u_majority7_module_6__and_module_7_U1 ( .A1(
        n_majority7_module_6__or_module_3_res), .A2(
        n_majority7_module_6__or_module_4_res), .ZN(
        n_majority7_module_6__and_module_7_res) );
  OR2_X1 u_majority7_module_6__or_module_8_U1 ( .A1(
        n_majority7_module_6__or_module_4_res), .A2(
        n_majority7_module_6__or_module_3_res), .ZN(
        n_majority7_module_6__or_module_8_res) );
  AND2_X1 u_majority7_module_6__and_module_8_U1 ( .A1(
        n_majority7_module_6__or_module_5_res), .A2(
        n_majority7_module_6__and_module_6_res), .ZN(
        n_majority7_module_6__and_module_8_res) );
  OR2_X1 u_majority7_module_6__or_module_9_U1 ( .A1(
        n_majority7_module_6__and_module_6_res), .A2(
        n_majority7_module_6__or_module_5_res), .ZN(
        n_majority7_module_6__or_module_9_res) );
  OR2_X1 u_majority7_module_6__or_module_10_U1 ( .A1(
        n_majority7_module_6__or_module_7_res), .A2(
        n_majority7_module_6__and_module_7_res), .ZN(
        n_majority7_module_6__or_module_10_res) );
  AND2_X1 u_majority7_module_6__and_module_9_U1 ( .A1(
        n_majority7_module_6__or_module_6_res), .A2(
        n_majority7_module_6__or_module_9_res), .ZN(
        n_majority7_module_6__and_module_9_res) );
  OR2_X1 u_majority7_module_6__or_module_11_U1 ( .A1(
        n_majority7_module_6__or_module_10_res), .A2(
        n_majority7_module_6__and_module_8_res), .ZN(
        n_majority7_module_6__or_module_11_res) );
  AND2_X1 u_majority7_module_6__and_module_10_U1 ( .A1(
        n_majority7_module_6__or_module_8_res), .A2(
        n_majority7_module_6__and_module_9_res), .ZN(
        n_majority7_module_6__and_module_10_res) );
  AND2_X1 u_majority7_module_6__and_module_11_U1 ( .A1(
        n_majority7_module_6__and_module_10_res), .A2(
        n_majority7_module_6__or_module_11_res), .ZN(n_majority7_module_6_res)
         );
  DFF_X1 u_reg_module_7__cini_mul_v000_reg ( .D(n_majority7_module_6_res), 
        .CK(clock_0), .Q(n_reg_module_7_res), .QN() );
  BUF_X1 u_majority7_module_7_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_7_n7) );
  BUF_X1 u_majority7_module_7_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_7_n6) );
  BUF_X1 u_majority7_module_7_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_7_n5) );
  BUF_X1 u_majority7_module_7_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_7_n4) );
  BUF_X1 u_majority7_module_7_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_7_n3) );
  BUF_X1 u_majority7_module_7_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_7_n2) );
  BUF_X1 u_majority7_module_7_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_7_n1) );
  AND2_X1 u_majority7_module_7__and_module_1_U1 ( .A1(n_majority7_module_7_n5), 
        .A2(n_majority7_module_7_n4), .ZN(
        n_majority7_module_7__and_module_1_res) );
  OR2_X1 u_majority7_module_7__or_module_1_U1 ( .A1(n_majority7_module_7_n4), 
        .A2(n_majority7_module_7_n5), .ZN(
        n_majority7_module_7__or_module_1_res) );
  AND2_X1 u_majority7_module_7__and_module_2_U1 ( .A1(n_majority7_module_7_n7), 
        .A2(n_majority7_module_7_n2), .ZN(
        n_majority7_module_7__and_module_2_res) );
  OR2_X1 u_majority7_module_7__or_module_2_U1 ( .A1(n_majority7_module_7_n2), 
        .A2(n_majority7_module_7_n7), .ZN(
        n_majority7_module_7__or_module_2_res) );
  AND2_X1 u_majority7_module_7__and_module_3_U1 ( .A1(n_majority7_module_7_n6), 
        .A2(n_majority7_module_7_n1), .ZN(
        n_majority7_module_7__and_module_3_res) );
  OR2_X1 u_majority7_module_7__or_module_3_U1 ( .A1(n_majority7_module_7_n1), 
        .A2(n_majority7_module_7_n6), .ZN(
        n_majority7_module_7__or_module_3_res) );
  AND2_X1 u_majority7_module_7__and_module_4_U1 ( .A1(
        n_majority7_module_7__and_module_2_res), .A2(
        n_majority7_module_7__and_module_1_res), .ZN(
        n_majority7_module_7__and_module_4_res) );
  OR2_X1 u_majority7_module_7__or_module_4_U1 ( .A1(
        n_majority7_module_7__and_module_1_res), .A2(
        n_majority7_module_7__and_module_2_res), .ZN(
        n_majority7_module_7__or_module_4_res) );
  AND2_X1 u_majority7_module_7__and_module_5_U1 ( .A1(
        n_majority7_module_7__and_module_3_res), .A2(n_majority7_module_7_n3), 
        .ZN(n_majority7_module_7__and_module_5_res) );
  OR2_X1 u_majority7_module_7__or_module_5_U1 ( .A1(n_majority7_module_7_n3), 
        .A2(n_majority7_module_7__and_module_3_res), .ZN(
        n_majority7_module_7__or_module_5_res) );
  AND2_X1 u_majority7_module_7__and_module_6_U1 ( .A1(
        n_majority7_module_7__or_module_1_res), .A2(
        n_majority7_module_7__or_module_2_res), .ZN(
        n_majority7_module_7__and_module_6_res) );
  OR2_X1 u_majority7_module_7__or_module_6_U1 ( .A1(
        n_majority7_module_7__or_module_2_res), .A2(
        n_majority7_module_7__or_module_1_res), .ZN(
        n_majority7_module_7__or_module_6_res) );
  OR2_X1 u_majority7_module_7__or_module_7_U1 ( .A1(
        n_majority7_module_7__and_module_4_res), .A2(
        n_majority7_module_7__and_module_5_res), .ZN(
        n_majority7_module_7__or_module_7_res) );
  AND2_X1 u_majority7_module_7__and_module_7_U1 ( .A1(
        n_majority7_module_7__or_module_3_res), .A2(
        n_majority7_module_7__or_module_4_res), .ZN(
        n_majority7_module_7__and_module_7_res) );
  OR2_X1 u_majority7_module_7__or_module_8_U1 ( .A1(
        n_majority7_module_7__or_module_4_res), .A2(
        n_majority7_module_7__or_module_3_res), .ZN(
        n_majority7_module_7__or_module_8_res) );
  AND2_X1 u_majority7_module_7__and_module_8_U1 ( .A1(
        n_majority7_module_7__or_module_5_res), .A2(
        n_majority7_module_7__and_module_6_res), .ZN(
        n_majority7_module_7__and_module_8_res) );
  OR2_X1 u_majority7_module_7__or_module_9_U1 ( .A1(
        n_majority7_module_7__and_module_6_res), .A2(
        n_majority7_module_7__or_module_5_res), .ZN(
        n_majority7_module_7__or_module_9_res) );
  OR2_X1 u_majority7_module_7__or_module_10_U1 ( .A1(
        n_majority7_module_7__or_module_7_res), .A2(
        n_majority7_module_7__and_module_7_res), .ZN(
        n_majority7_module_7__or_module_10_res) );
  AND2_X1 u_majority7_module_7__and_module_9_U1 ( .A1(
        n_majority7_module_7__or_module_6_res), .A2(
        n_majority7_module_7__or_module_9_res), .ZN(
        n_majority7_module_7__and_module_9_res) );
  OR2_X1 u_majority7_module_7__or_module_11_U1 ( .A1(
        n_majority7_module_7__or_module_10_res), .A2(
        n_majority7_module_7__and_module_8_res), .ZN(
        n_majority7_module_7__or_module_11_res) );
  AND2_X1 u_majority7_module_7__and_module_10_U1 ( .A1(
        n_majority7_module_7__or_module_8_res), .A2(
        n_majority7_module_7__and_module_9_res), .ZN(
        n_majority7_module_7__and_module_10_res) );
  AND2_X1 u_majority7_module_7__and_module_11_U1 ( .A1(
        n_majority7_module_7__and_module_10_res), .A2(
        n_majority7_module_7__or_module_11_res), .ZN(n_majority7_module_7_res)
         );
  DFF_X1 u_reg_module_8__cini_mul_v000_reg ( .D(n_majority7_module_7_res), 
        .CK(clock_0), .Q(n_reg_module_8_res), .QN() );
  BUF_X1 u_majority7_module_8_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_8_n7) );
  BUF_X1 u_majority7_module_8_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_8_n6) );
  BUF_X1 u_majority7_module_8_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_8_n5) );
  BUF_X1 u_majority7_module_8_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_8_n4) );
  BUF_X1 u_majority7_module_8_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_8_n3) );
  BUF_X1 u_majority7_module_8_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_8_n2) );
  BUF_X1 u_majority7_module_8_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_8_n1) );
  AND2_X1 u_majority7_module_8__and_module_1_U1 ( .A1(n_majority7_module_8_n5), 
        .A2(n_majority7_module_8_n4), .ZN(
        n_majority7_module_8__and_module_1_res) );
  OR2_X1 u_majority7_module_8__or_module_1_U1 ( .A1(n_majority7_module_8_n4), 
        .A2(n_majority7_module_8_n5), .ZN(
        n_majority7_module_8__or_module_1_res) );
  AND2_X1 u_majority7_module_8__and_module_2_U1 ( .A1(n_majority7_module_8_n7), 
        .A2(n_majority7_module_8_n2), .ZN(
        n_majority7_module_8__and_module_2_res) );
  OR2_X1 u_majority7_module_8__or_module_2_U1 ( .A1(n_majority7_module_8_n2), 
        .A2(n_majority7_module_8_n7), .ZN(
        n_majority7_module_8__or_module_2_res) );
  AND2_X1 u_majority7_module_8__and_module_3_U1 ( .A1(n_majority7_module_8_n6), 
        .A2(n_majority7_module_8_n1), .ZN(
        n_majority7_module_8__and_module_3_res) );
  OR2_X1 u_majority7_module_8__or_module_3_U1 ( .A1(n_majority7_module_8_n1), 
        .A2(n_majority7_module_8_n6), .ZN(
        n_majority7_module_8__or_module_3_res) );
  AND2_X1 u_majority7_module_8__and_module_4_U1 ( .A1(
        n_majority7_module_8__and_module_2_res), .A2(
        n_majority7_module_8__and_module_1_res), .ZN(
        n_majority7_module_8__and_module_4_res) );
  OR2_X1 u_majority7_module_8__or_module_4_U1 ( .A1(
        n_majority7_module_8__and_module_1_res), .A2(
        n_majority7_module_8__and_module_2_res), .ZN(
        n_majority7_module_8__or_module_4_res) );
  AND2_X1 u_majority7_module_8__and_module_5_U1 ( .A1(
        n_majority7_module_8__and_module_3_res), .A2(n_majority7_module_8_n3), 
        .ZN(n_majority7_module_8__and_module_5_res) );
  OR2_X1 u_majority7_module_8__or_module_5_U1 ( .A1(n_majority7_module_8_n3), 
        .A2(n_majority7_module_8__and_module_3_res), .ZN(
        n_majority7_module_8__or_module_5_res) );
  AND2_X1 u_majority7_module_8__and_module_6_U1 ( .A1(
        n_majority7_module_8__or_module_1_res), .A2(
        n_majority7_module_8__or_module_2_res), .ZN(
        n_majority7_module_8__and_module_6_res) );
  OR2_X1 u_majority7_module_8__or_module_6_U1 ( .A1(
        n_majority7_module_8__or_module_2_res), .A2(
        n_majority7_module_8__or_module_1_res), .ZN(
        n_majority7_module_8__or_module_6_res) );
  OR2_X1 u_majority7_module_8__or_module_7_U1 ( .A1(
        n_majority7_module_8__and_module_4_res), .A2(
        n_majority7_module_8__and_module_5_res), .ZN(
        n_majority7_module_8__or_module_7_res) );
  AND2_X1 u_majority7_module_8__and_module_7_U1 ( .A1(
        n_majority7_module_8__or_module_3_res), .A2(
        n_majority7_module_8__or_module_4_res), .ZN(
        n_majority7_module_8__and_module_7_res) );
  OR2_X1 u_majority7_module_8__or_module_8_U1 ( .A1(
        n_majority7_module_8__or_module_4_res), .A2(
        n_majority7_module_8__or_module_3_res), .ZN(
        n_majority7_module_8__or_module_8_res) );
  AND2_X1 u_majority7_module_8__and_module_8_U1 ( .A1(
        n_majority7_module_8__or_module_5_res), .A2(
        n_majority7_module_8__and_module_6_res), .ZN(
        n_majority7_module_8__and_module_8_res) );
  OR2_X1 u_majority7_module_8__or_module_9_U1 ( .A1(
        n_majority7_module_8__and_module_6_res), .A2(
        n_majority7_module_8__or_module_5_res), .ZN(
        n_majority7_module_8__or_module_9_res) );
  OR2_X1 u_majority7_module_8__or_module_10_U1 ( .A1(
        n_majority7_module_8__or_module_7_res), .A2(
        n_majority7_module_8__and_module_7_res), .ZN(
        n_majority7_module_8__or_module_10_res) );
  AND2_X1 u_majority7_module_8__and_module_9_U1 ( .A1(
        n_majority7_module_8__or_module_6_res), .A2(
        n_majority7_module_8__or_module_9_res), .ZN(
        n_majority7_module_8__and_module_9_res) );
  OR2_X1 u_majority7_module_8__or_module_11_U1 ( .A1(
        n_majority7_module_8__or_module_10_res), .A2(
        n_majority7_module_8__and_module_8_res), .ZN(
        n_majority7_module_8__or_module_11_res) );
  AND2_X1 u_majority7_module_8__and_module_10_U1 ( .A1(
        n_majority7_module_8__or_module_8_res), .A2(
        n_majority7_module_8__and_module_9_res), .ZN(
        n_majority7_module_8__and_module_10_res) );
  AND2_X1 u_majority7_module_8__and_module_11_U1 ( .A1(
        n_majority7_module_8__and_module_10_res), .A2(
        n_majority7_module_8__or_module_11_res), .ZN(n_majority7_module_8_res)
         );
  DFF_X1 u_reg_module_9__cini_mul_v000_reg ( .D(n_majority7_module_8_res), 
        .CK(clock_0), .Q(n_reg_module_9_res), .QN() );
  BUF_X1 u_majority7_module_9_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_9_n7) );
  BUF_X1 u_majority7_module_9_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_9_n6) );
  BUF_X1 u_majority7_module_9_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_9_n5) );
  BUF_X1 u_majority7_module_9_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_9_n4) );
  BUF_X1 u_majority7_module_9_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_9_n3) );
  BUF_X1 u_majority7_module_9_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_9_n2) );
  BUF_X1 u_majority7_module_9_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_9_n1) );
  AND2_X1 u_majority7_module_9__and_module_1_U1 ( .A1(n_majority7_module_9_n5), 
        .A2(n_majority7_module_9_n4), .ZN(
        n_majority7_module_9__and_module_1_res) );
  OR2_X1 u_majority7_module_9__or_module_1_U1 ( .A1(n_majority7_module_9_n4), 
        .A2(n_majority7_module_9_n5), .ZN(
        n_majority7_module_9__or_module_1_res) );
  AND2_X1 u_majority7_module_9__and_module_2_U1 ( .A1(n_majority7_module_9_n7), 
        .A2(n_majority7_module_9_n2), .ZN(
        n_majority7_module_9__and_module_2_res) );
  OR2_X1 u_majority7_module_9__or_module_2_U1 ( .A1(n_majority7_module_9_n2), 
        .A2(n_majority7_module_9_n7), .ZN(
        n_majority7_module_9__or_module_2_res) );
  AND2_X1 u_majority7_module_9__and_module_3_U1 ( .A1(n_majority7_module_9_n6), 
        .A2(n_majority7_module_9_n1), .ZN(
        n_majority7_module_9__and_module_3_res) );
  OR2_X1 u_majority7_module_9__or_module_3_U1 ( .A1(n_majority7_module_9_n1), 
        .A2(n_majority7_module_9_n6), .ZN(
        n_majority7_module_9__or_module_3_res) );
  AND2_X1 u_majority7_module_9__and_module_4_U1 ( .A1(
        n_majority7_module_9__and_module_2_res), .A2(
        n_majority7_module_9__and_module_1_res), .ZN(
        n_majority7_module_9__and_module_4_res) );
  OR2_X1 u_majority7_module_9__or_module_4_U1 ( .A1(
        n_majority7_module_9__and_module_1_res), .A2(
        n_majority7_module_9__and_module_2_res), .ZN(
        n_majority7_module_9__or_module_4_res) );
  AND2_X1 u_majority7_module_9__and_module_5_U1 ( .A1(
        n_majority7_module_9__and_module_3_res), .A2(n_majority7_module_9_n3), 
        .ZN(n_majority7_module_9__and_module_5_res) );
  OR2_X1 u_majority7_module_9__or_module_5_U1 ( .A1(n_majority7_module_9_n3), 
        .A2(n_majority7_module_9__and_module_3_res), .ZN(
        n_majority7_module_9__or_module_5_res) );
  AND2_X1 u_majority7_module_9__and_module_6_U1 ( .A1(
        n_majority7_module_9__or_module_1_res), .A2(
        n_majority7_module_9__or_module_2_res), .ZN(
        n_majority7_module_9__and_module_6_res) );
  OR2_X1 u_majority7_module_9__or_module_6_U1 ( .A1(
        n_majority7_module_9__or_module_2_res), .A2(
        n_majority7_module_9__or_module_1_res), .ZN(
        n_majority7_module_9__or_module_6_res) );
  OR2_X1 u_majority7_module_9__or_module_7_U1 ( .A1(
        n_majority7_module_9__and_module_4_res), .A2(
        n_majority7_module_9__and_module_5_res), .ZN(
        n_majority7_module_9__or_module_7_res) );
  AND2_X1 u_majority7_module_9__and_module_7_U1 ( .A1(
        n_majority7_module_9__or_module_3_res), .A2(
        n_majority7_module_9__or_module_4_res), .ZN(
        n_majority7_module_9__and_module_7_res) );
  OR2_X1 u_majority7_module_9__or_module_8_U1 ( .A1(
        n_majority7_module_9__or_module_4_res), .A2(
        n_majority7_module_9__or_module_3_res), .ZN(
        n_majority7_module_9__or_module_8_res) );
  AND2_X1 u_majority7_module_9__and_module_8_U1 ( .A1(
        n_majority7_module_9__or_module_5_res), .A2(
        n_majority7_module_9__and_module_6_res), .ZN(
        n_majority7_module_9__and_module_8_res) );
  OR2_X1 u_majority7_module_9__or_module_9_U1 ( .A1(
        n_majority7_module_9__and_module_6_res), .A2(
        n_majority7_module_9__or_module_5_res), .ZN(
        n_majority7_module_9__or_module_9_res) );
  OR2_X1 u_majority7_module_9__or_module_10_U1 ( .A1(
        n_majority7_module_9__or_module_7_res), .A2(
        n_majority7_module_9__and_module_7_res), .ZN(
        n_majority7_module_9__or_module_10_res) );
  AND2_X1 u_majority7_module_9__and_module_9_U1 ( .A1(
        n_majority7_module_9__or_module_6_res), .A2(
        n_majority7_module_9__or_module_9_res), .ZN(
        n_majority7_module_9__and_module_9_res) );
  OR2_X1 u_majority7_module_9__or_module_11_U1 ( .A1(
        n_majority7_module_9__or_module_10_res), .A2(
        n_majority7_module_9__and_module_8_res), .ZN(
        n_majority7_module_9__or_module_11_res) );
  AND2_X1 u_majority7_module_9__and_module_10_U1 ( .A1(
        n_majority7_module_9__or_module_8_res), .A2(
        n_majority7_module_9__and_module_9_res), .ZN(
        n_majority7_module_9__and_module_10_res) );
  AND2_X1 u_majority7_module_9__and_module_11_U1 ( .A1(
        n_majority7_module_9__and_module_10_res), .A2(
        n_majority7_module_9__or_module_11_res), .ZN(n_majority7_module_9_res)
         );
  DFF_X1 u_reg_module_10__cini_mul_v000_reg ( .D(n_majority7_module_9_res), 
        .CK(clock_1), .Q(n_reg_module_10_res), .QN() );
  BUF_X1 u_majority7_module_10_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_10_n7) );
  BUF_X1 u_majority7_module_10_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_10_n6) );
  BUF_X1 u_majority7_module_10_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_10_n5) );
  BUF_X1 u_majority7_module_10_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_10_n4) );
  BUF_X1 u_majority7_module_10_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_10_n3) );
  BUF_X1 u_majority7_module_10_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_10_n2) );
  BUF_X1 u_majority7_module_10_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_10_n1) );
  AND2_X1 u_majority7_module_10__and_module_1_U1 ( .A1(
        n_majority7_module_10_n5), .A2(n_majority7_module_10_n4), .ZN(
        n_majority7_module_10__and_module_1_res) );
  OR2_X1 u_majority7_module_10__or_module_1_U1 ( .A1(n_majority7_module_10_n4), 
        .A2(n_majority7_module_10_n5), .ZN(
        n_majority7_module_10__or_module_1_res) );
  AND2_X1 u_majority7_module_10__and_module_2_U1 ( .A1(
        n_majority7_module_10_n7), .A2(n_majority7_module_10_n2), .ZN(
        n_majority7_module_10__and_module_2_res) );
  OR2_X1 u_majority7_module_10__or_module_2_U1 ( .A1(n_majority7_module_10_n2), 
        .A2(n_majority7_module_10_n7), .ZN(
        n_majority7_module_10__or_module_2_res) );
  AND2_X1 u_majority7_module_10__and_module_3_U1 ( .A1(
        n_majority7_module_10_n6), .A2(n_majority7_module_10_n1), .ZN(
        n_majority7_module_10__and_module_3_res) );
  OR2_X1 u_majority7_module_10__or_module_3_U1 ( .A1(n_majority7_module_10_n1), 
        .A2(n_majority7_module_10_n6), .ZN(
        n_majority7_module_10__or_module_3_res) );
  AND2_X1 u_majority7_module_10__and_module_4_U1 ( .A1(
        n_majority7_module_10__and_module_2_res), .A2(
        n_majority7_module_10__and_module_1_res), .ZN(
        n_majority7_module_10__and_module_4_res) );
  OR2_X1 u_majority7_module_10__or_module_4_U1 ( .A1(
        n_majority7_module_10__and_module_1_res), .A2(
        n_majority7_module_10__and_module_2_res), .ZN(
        n_majority7_module_10__or_module_4_res) );
  AND2_X1 u_majority7_module_10__and_module_5_U1 ( .A1(
        n_majority7_module_10__and_module_3_res), .A2(n_majority7_module_10_n3), .ZN(n_majority7_module_10__and_module_5_res) );
  OR2_X1 u_majority7_module_10__or_module_5_U1 ( .A1(n_majority7_module_10_n3), 
        .A2(n_majority7_module_10__and_module_3_res), .ZN(
        n_majority7_module_10__or_module_5_res) );
  AND2_X1 u_majority7_module_10__and_module_6_U1 ( .A1(
        n_majority7_module_10__or_module_1_res), .A2(
        n_majority7_module_10__or_module_2_res), .ZN(
        n_majority7_module_10__and_module_6_res) );
  OR2_X1 u_majority7_module_10__or_module_6_U1 ( .A1(
        n_majority7_module_10__or_module_2_res), .A2(
        n_majority7_module_10__or_module_1_res), .ZN(
        n_majority7_module_10__or_module_6_res) );
  OR2_X1 u_majority7_module_10__or_module_7_U1 ( .A1(
        n_majority7_module_10__and_module_4_res), .A2(
        n_majority7_module_10__and_module_5_res), .ZN(
        n_majority7_module_10__or_module_7_res) );
  AND2_X1 u_majority7_module_10__and_module_7_U1 ( .A1(
        n_majority7_module_10__or_module_3_res), .A2(
        n_majority7_module_10__or_module_4_res), .ZN(
        n_majority7_module_10__and_module_7_res) );
  OR2_X1 u_majority7_module_10__or_module_8_U1 ( .A1(
        n_majority7_module_10__or_module_4_res), .A2(
        n_majority7_module_10__or_module_3_res), .ZN(
        n_majority7_module_10__or_module_8_res) );
  AND2_X1 u_majority7_module_10__and_module_8_U1 ( .A1(
        n_majority7_module_10__or_module_5_res), .A2(
        n_majority7_module_10__and_module_6_res), .ZN(
        n_majority7_module_10__and_module_8_res) );
  OR2_X1 u_majority7_module_10__or_module_9_U1 ( .A1(
        n_majority7_module_10__and_module_6_res), .A2(
        n_majority7_module_10__or_module_5_res), .ZN(
        n_majority7_module_10__or_module_9_res) );
  OR2_X1 u_majority7_module_10__or_module_10_U1 ( .A1(
        n_majority7_module_10__or_module_7_res), .A2(
        n_majority7_module_10__and_module_7_res), .ZN(
        n_majority7_module_10__or_module_10_res) );
  AND2_X1 u_majority7_module_10__and_module_9_U1 ( .A1(
        n_majority7_module_10__or_module_6_res), .A2(
        n_majority7_module_10__or_module_9_res), .ZN(
        n_majority7_module_10__and_module_9_res) );
  OR2_X1 u_majority7_module_10__or_module_11_U1 ( .A1(
        n_majority7_module_10__or_module_10_res), .A2(
        n_majority7_module_10__and_module_8_res), .ZN(
        n_majority7_module_10__or_module_11_res) );
  AND2_X1 u_majority7_module_10__and_module_10_U1 ( .A1(
        n_majority7_module_10__or_module_8_res), .A2(
        n_majority7_module_10__and_module_9_res), .ZN(
        n_majority7_module_10__and_module_10_res) );
  AND2_X1 u_majority7_module_10__and_module_11_U1 ( .A1(
        n_majority7_module_10__and_module_10_res), .A2(
        n_majority7_module_10__or_module_11_res), .ZN(
        n_majority7_module_10_res) );
  DFF_X1 u_reg_module_11__cini_mul_v000_reg ( .D(n_majority7_module_10_res), 
        .CK(clock_1), .Q(n_reg_module_11_res), .QN() );
  BUF_X1 u_majority7_module_11_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_11_n7) );
  BUF_X1 u_majority7_module_11_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_11_n6) );
  BUF_X1 u_majority7_module_11_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_11_n5) );
  BUF_X1 u_majority7_module_11_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_11_n4) );
  BUF_X1 u_majority7_module_11_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_11_n3) );
  BUF_X1 u_majority7_module_11_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_11_n2) );
  BUF_X1 u_majority7_module_11_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_11_n1) );
  AND2_X1 u_majority7_module_11__and_module_1_U1 ( .A1(
        n_majority7_module_11_n5), .A2(n_majority7_module_11_n4), .ZN(
        n_majority7_module_11__and_module_1_res) );
  OR2_X1 u_majority7_module_11__or_module_1_U1 ( .A1(n_majority7_module_11_n4), 
        .A2(n_majority7_module_11_n5), .ZN(
        n_majority7_module_11__or_module_1_res) );
  AND2_X1 u_majority7_module_11__and_module_2_U1 ( .A1(
        n_majority7_module_11_n7), .A2(n_majority7_module_11_n2), .ZN(
        n_majority7_module_11__and_module_2_res) );
  OR2_X1 u_majority7_module_11__or_module_2_U1 ( .A1(n_majority7_module_11_n2), 
        .A2(n_majority7_module_11_n7), .ZN(
        n_majority7_module_11__or_module_2_res) );
  AND2_X1 u_majority7_module_11__and_module_3_U1 ( .A1(
        n_majority7_module_11_n6), .A2(n_majority7_module_11_n1), .ZN(
        n_majority7_module_11__and_module_3_res) );
  OR2_X1 u_majority7_module_11__or_module_3_U1 ( .A1(n_majority7_module_11_n1), 
        .A2(n_majority7_module_11_n6), .ZN(
        n_majority7_module_11__or_module_3_res) );
  AND2_X1 u_majority7_module_11__and_module_4_U1 ( .A1(
        n_majority7_module_11__and_module_2_res), .A2(
        n_majority7_module_11__and_module_1_res), .ZN(
        n_majority7_module_11__and_module_4_res) );
  OR2_X1 u_majority7_module_11__or_module_4_U1 ( .A1(
        n_majority7_module_11__and_module_1_res), .A2(
        n_majority7_module_11__and_module_2_res), .ZN(
        n_majority7_module_11__or_module_4_res) );
  AND2_X1 u_majority7_module_11__and_module_5_U1 ( .A1(
        n_majority7_module_11__and_module_3_res), .A2(n_majority7_module_11_n3), .ZN(n_majority7_module_11__and_module_5_res) );
  OR2_X1 u_majority7_module_11__or_module_5_U1 ( .A1(n_majority7_module_11_n3), 
        .A2(n_majority7_module_11__and_module_3_res), .ZN(
        n_majority7_module_11__or_module_5_res) );
  AND2_X1 u_majority7_module_11__and_module_6_U1 ( .A1(
        n_majority7_module_11__or_module_1_res), .A2(
        n_majority7_module_11__or_module_2_res), .ZN(
        n_majority7_module_11__and_module_6_res) );
  OR2_X1 u_majority7_module_11__or_module_6_U1 ( .A1(
        n_majority7_module_11__or_module_2_res), .A2(
        n_majority7_module_11__or_module_1_res), .ZN(
        n_majority7_module_11__or_module_6_res) );
  OR2_X1 u_majority7_module_11__or_module_7_U1 ( .A1(
        n_majority7_module_11__and_module_4_res), .A2(
        n_majority7_module_11__and_module_5_res), .ZN(
        n_majority7_module_11__or_module_7_res) );
  AND2_X1 u_majority7_module_11__and_module_7_U1 ( .A1(
        n_majority7_module_11__or_module_3_res), .A2(
        n_majority7_module_11__or_module_4_res), .ZN(
        n_majority7_module_11__and_module_7_res) );
  OR2_X1 u_majority7_module_11__or_module_8_U1 ( .A1(
        n_majority7_module_11__or_module_4_res), .A2(
        n_majority7_module_11__or_module_3_res), .ZN(
        n_majority7_module_11__or_module_8_res) );
  AND2_X1 u_majority7_module_11__and_module_8_U1 ( .A1(
        n_majority7_module_11__or_module_5_res), .A2(
        n_majority7_module_11__and_module_6_res), .ZN(
        n_majority7_module_11__and_module_8_res) );
  OR2_X1 u_majority7_module_11__or_module_9_U1 ( .A1(
        n_majority7_module_11__and_module_6_res), .A2(
        n_majority7_module_11__or_module_5_res), .ZN(
        n_majority7_module_11__or_module_9_res) );
  OR2_X1 u_majority7_module_11__or_module_10_U1 ( .A1(
        n_majority7_module_11__or_module_7_res), .A2(
        n_majority7_module_11__and_module_7_res), .ZN(
        n_majority7_module_11__or_module_10_res) );
  AND2_X1 u_majority7_module_11__and_module_9_U1 ( .A1(
        n_majority7_module_11__or_module_6_res), .A2(
        n_majority7_module_11__or_module_9_res), .ZN(
        n_majority7_module_11__and_module_9_res) );
  OR2_X1 u_majority7_module_11__or_module_11_U1 ( .A1(
        n_majority7_module_11__or_module_10_res), .A2(
        n_majority7_module_11__and_module_8_res), .ZN(
        n_majority7_module_11__or_module_11_res) );
  AND2_X1 u_majority7_module_11__and_module_10_U1 ( .A1(
        n_majority7_module_11__or_module_8_res), .A2(
        n_majority7_module_11__and_module_9_res), .ZN(
        n_majority7_module_11__and_module_10_res) );
  AND2_X1 u_majority7_module_11__and_module_11_U1 ( .A1(
        n_majority7_module_11__and_module_10_res), .A2(
        n_majority7_module_11__or_module_11_res), .ZN(
        n_majority7_module_11_res) );
  DFF_X1 u_reg_module_12__cini_mul_v000_reg ( .D(n_majority7_module_11_res), 
        .CK(clock_1), .Q(n_reg_module_12_res), .QN() );
  BUF_X1 u_majority7_module_12_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_12_n7) );
  BUF_X1 u_majority7_module_12_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_12_n6) );
  BUF_X1 u_majority7_module_12_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_12_n5) );
  BUF_X1 u_majority7_module_12_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_12_n4) );
  BUF_X1 u_majority7_module_12_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_12_n3) );
  BUF_X1 u_majority7_module_12_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_12_n2) );
  BUF_X1 u_majority7_module_12_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_12_n1) );
  AND2_X1 u_majority7_module_12__and_module_1_U1 ( .A1(
        n_majority7_module_12_n5), .A2(n_majority7_module_12_n4), .ZN(
        n_majority7_module_12__and_module_1_res) );
  OR2_X1 u_majority7_module_12__or_module_1_U1 ( .A1(n_majority7_module_12_n4), 
        .A2(n_majority7_module_12_n5), .ZN(
        n_majority7_module_12__or_module_1_res) );
  AND2_X1 u_majority7_module_12__and_module_2_U1 ( .A1(
        n_majority7_module_12_n7), .A2(n_majority7_module_12_n2), .ZN(
        n_majority7_module_12__and_module_2_res) );
  OR2_X1 u_majority7_module_12__or_module_2_U1 ( .A1(n_majority7_module_12_n2), 
        .A2(n_majority7_module_12_n7), .ZN(
        n_majority7_module_12__or_module_2_res) );
  AND2_X1 u_majority7_module_12__and_module_3_U1 ( .A1(
        n_majority7_module_12_n6), .A2(n_majority7_module_12_n1), .ZN(
        n_majority7_module_12__and_module_3_res) );
  OR2_X1 u_majority7_module_12__or_module_3_U1 ( .A1(n_majority7_module_12_n1), 
        .A2(n_majority7_module_12_n6), .ZN(
        n_majority7_module_12__or_module_3_res) );
  AND2_X1 u_majority7_module_12__and_module_4_U1 ( .A1(
        n_majority7_module_12__and_module_2_res), .A2(
        n_majority7_module_12__and_module_1_res), .ZN(
        n_majority7_module_12__and_module_4_res) );
  OR2_X1 u_majority7_module_12__or_module_4_U1 ( .A1(
        n_majority7_module_12__and_module_1_res), .A2(
        n_majority7_module_12__and_module_2_res), .ZN(
        n_majority7_module_12__or_module_4_res) );
  AND2_X1 u_majority7_module_12__and_module_5_U1 ( .A1(
        n_majority7_module_12__and_module_3_res), .A2(n_majority7_module_12_n3), .ZN(n_majority7_module_12__and_module_5_res) );
  OR2_X1 u_majority7_module_12__or_module_5_U1 ( .A1(n_majority7_module_12_n3), 
        .A2(n_majority7_module_12__and_module_3_res), .ZN(
        n_majority7_module_12__or_module_5_res) );
  AND2_X1 u_majority7_module_12__and_module_6_U1 ( .A1(
        n_majority7_module_12__or_module_1_res), .A2(
        n_majority7_module_12__or_module_2_res), .ZN(
        n_majority7_module_12__and_module_6_res) );
  OR2_X1 u_majority7_module_12__or_module_6_U1 ( .A1(
        n_majority7_module_12__or_module_2_res), .A2(
        n_majority7_module_12__or_module_1_res), .ZN(
        n_majority7_module_12__or_module_6_res) );
  OR2_X1 u_majority7_module_12__or_module_7_U1 ( .A1(
        n_majority7_module_12__and_module_4_res), .A2(
        n_majority7_module_12__and_module_5_res), .ZN(
        n_majority7_module_12__or_module_7_res) );
  AND2_X1 u_majority7_module_12__and_module_7_U1 ( .A1(
        n_majority7_module_12__or_module_3_res), .A2(
        n_majority7_module_12__or_module_4_res), .ZN(
        n_majority7_module_12__and_module_7_res) );
  OR2_X1 u_majority7_module_12__or_module_8_U1 ( .A1(
        n_majority7_module_12__or_module_4_res), .A2(
        n_majority7_module_12__or_module_3_res), .ZN(
        n_majority7_module_12__or_module_8_res) );
  AND2_X1 u_majority7_module_12__and_module_8_U1 ( .A1(
        n_majority7_module_12__or_module_5_res), .A2(
        n_majority7_module_12__and_module_6_res), .ZN(
        n_majority7_module_12__and_module_8_res) );
  OR2_X1 u_majority7_module_12__or_module_9_U1 ( .A1(
        n_majority7_module_12__and_module_6_res), .A2(
        n_majority7_module_12__or_module_5_res), .ZN(
        n_majority7_module_12__or_module_9_res) );
  OR2_X1 u_majority7_module_12__or_module_10_U1 ( .A1(
        n_majority7_module_12__or_module_7_res), .A2(
        n_majority7_module_12__and_module_7_res), .ZN(
        n_majority7_module_12__or_module_10_res) );
  AND2_X1 u_majority7_module_12__and_module_9_U1 ( .A1(
        n_majority7_module_12__or_module_6_res), .A2(
        n_majority7_module_12__or_module_9_res), .ZN(
        n_majority7_module_12__and_module_9_res) );
  OR2_X1 u_majority7_module_12__or_module_11_U1 ( .A1(
        n_majority7_module_12__or_module_10_res), .A2(
        n_majority7_module_12__and_module_8_res), .ZN(
        n_majority7_module_12__or_module_11_res) );
  AND2_X1 u_majority7_module_12__and_module_10_U1 ( .A1(
        n_majority7_module_12__or_module_8_res), .A2(
        n_majority7_module_12__and_module_9_res), .ZN(
        n_majority7_module_12__and_module_10_res) );
  AND2_X1 u_majority7_module_12__and_module_11_U1 ( .A1(
        n_majority7_module_12__and_module_10_res), .A2(
        n_majority7_module_12__or_module_11_res), .ZN(
        n_majority7_module_12_res) );
  DFF_X1 u_reg_module_13__cini_mul_v000_reg ( .D(n_majority7_module_12_res), 
        .CK(clock_1), .Q(n_reg_module_13_res), .QN() );
  BUF_X1 u_majority7_module_13_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_13_n7) );
  BUF_X1 u_majority7_module_13_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_13_n6) );
  BUF_X1 u_majority7_module_13_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_13_n5) );
  BUF_X1 u_majority7_module_13_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_13_n4) );
  BUF_X1 u_majority7_module_13_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_13_n3) );
  BUF_X1 u_majority7_module_13_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_13_n2) );
  BUF_X1 u_majority7_module_13_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_13_n1) );
  AND2_X1 u_majority7_module_13__and_module_1_U1 ( .A1(
        n_majority7_module_13_n5), .A2(n_majority7_module_13_n4), .ZN(
        n_majority7_module_13__and_module_1_res) );
  OR2_X1 u_majority7_module_13__or_module_1_U1 ( .A1(n_majority7_module_13_n4), 
        .A2(n_majority7_module_13_n5), .ZN(
        n_majority7_module_13__or_module_1_res) );
  AND2_X1 u_majority7_module_13__and_module_2_U1 ( .A1(
        n_majority7_module_13_n7), .A2(n_majority7_module_13_n2), .ZN(
        n_majority7_module_13__and_module_2_res) );
  OR2_X1 u_majority7_module_13__or_module_2_U1 ( .A1(n_majority7_module_13_n2), 
        .A2(n_majority7_module_13_n7), .ZN(
        n_majority7_module_13__or_module_2_res) );
  AND2_X1 u_majority7_module_13__and_module_3_U1 ( .A1(
        n_majority7_module_13_n6), .A2(n_majority7_module_13_n1), .ZN(
        n_majority7_module_13__and_module_3_res) );
  OR2_X1 u_majority7_module_13__or_module_3_U1 ( .A1(n_majority7_module_13_n1), 
        .A2(n_majority7_module_13_n6), .ZN(
        n_majority7_module_13__or_module_3_res) );
  AND2_X1 u_majority7_module_13__and_module_4_U1 ( .A1(
        n_majority7_module_13__and_module_2_res), .A2(
        n_majority7_module_13__and_module_1_res), .ZN(
        n_majority7_module_13__and_module_4_res) );
  OR2_X1 u_majority7_module_13__or_module_4_U1 ( .A1(
        n_majority7_module_13__and_module_1_res), .A2(
        n_majority7_module_13__and_module_2_res), .ZN(
        n_majority7_module_13__or_module_4_res) );
  AND2_X1 u_majority7_module_13__and_module_5_U1 ( .A1(
        n_majority7_module_13__and_module_3_res), .A2(n_majority7_module_13_n3), .ZN(n_majority7_module_13__and_module_5_res) );
  OR2_X1 u_majority7_module_13__or_module_5_U1 ( .A1(n_majority7_module_13_n3), 
        .A2(n_majority7_module_13__and_module_3_res), .ZN(
        n_majority7_module_13__or_module_5_res) );
  AND2_X1 u_majority7_module_13__and_module_6_U1 ( .A1(
        n_majority7_module_13__or_module_1_res), .A2(
        n_majority7_module_13__or_module_2_res), .ZN(
        n_majority7_module_13__and_module_6_res) );
  OR2_X1 u_majority7_module_13__or_module_6_U1 ( .A1(
        n_majority7_module_13__or_module_2_res), .A2(
        n_majority7_module_13__or_module_1_res), .ZN(
        n_majority7_module_13__or_module_6_res) );
  OR2_X1 u_majority7_module_13__or_module_7_U1 ( .A1(
        n_majority7_module_13__and_module_4_res), .A2(
        n_majority7_module_13__and_module_5_res), .ZN(
        n_majority7_module_13__or_module_7_res) );
  AND2_X1 u_majority7_module_13__and_module_7_U1 ( .A1(
        n_majority7_module_13__or_module_3_res), .A2(
        n_majority7_module_13__or_module_4_res), .ZN(
        n_majority7_module_13__and_module_7_res) );
  OR2_X1 u_majority7_module_13__or_module_8_U1 ( .A1(
        n_majority7_module_13__or_module_4_res), .A2(
        n_majority7_module_13__or_module_3_res), .ZN(
        n_majority7_module_13__or_module_8_res) );
  AND2_X1 u_majority7_module_13__and_module_8_U1 ( .A1(
        n_majority7_module_13__or_module_5_res), .A2(
        n_majority7_module_13__and_module_6_res), .ZN(
        n_majority7_module_13__and_module_8_res) );
  OR2_X1 u_majority7_module_13__or_module_9_U1 ( .A1(
        n_majority7_module_13__and_module_6_res), .A2(
        n_majority7_module_13__or_module_5_res), .ZN(
        n_majority7_module_13__or_module_9_res) );
  OR2_X1 u_majority7_module_13__or_module_10_U1 ( .A1(
        n_majority7_module_13__or_module_7_res), .A2(
        n_majority7_module_13__and_module_7_res), .ZN(
        n_majority7_module_13__or_module_10_res) );
  AND2_X1 u_majority7_module_13__and_module_9_U1 ( .A1(
        n_majority7_module_13__or_module_6_res), .A2(
        n_majority7_module_13__or_module_9_res), .ZN(
        n_majority7_module_13__and_module_9_res) );
  OR2_X1 u_majority7_module_13__or_module_11_U1 ( .A1(
        n_majority7_module_13__or_module_10_res), .A2(
        n_majority7_module_13__and_module_8_res), .ZN(
        n_majority7_module_13__or_module_11_res) );
  AND2_X1 u_majority7_module_13__and_module_10_U1 ( .A1(
        n_majority7_module_13__or_module_8_res), .A2(
        n_majority7_module_13__and_module_9_res), .ZN(
        n_majority7_module_13__and_module_10_res) );
  AND2_X1 u_majority7_module_13__and_module_11_U1 ( .A1(
        n_majority7_module_13__and_module_10_res), .A2(
        n_majority7_module_13__or_module_11_res), .ZN(
        n_majority7_module_13_res) );
  DFF_X1 u_reg_module_14__cini_mul_v000_reg ( .D(n_majority7_module_13_res), 
        .CK(clock_1), .Q(n_reg_module_14_res), .QN() );
  BUF_X1 u_majority7_module_14_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_14_n7) );
  BUF_X1 u_majority7_module_14_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_14_n6) );
  BUF_X1 u_majority7_module_14_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_14_n5) );
  BUF_X1 u_majority7_module_14_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_14_n4) );
  BUF_X1 u_majority7_module_14_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_14_n3) );
  BUF_X1 u_majority7_module_14_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_14_n2) );
  BUF_X1 u_majority7_module_14_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_14_n1) );
  AND2_X1 u_majority7_module_14__and_module_1_U1 ( .A1(
        n_majority7_module_14_n5), .A2(n_majority7_module_14_n4), .ZN(
        n_majority7_module_14__and_module_1_res) );
  OR2_X1 u_majority7_module_14__or_module_1_U1 ( .A1(n_majority7_module_14_n4), 
        .A2(n_majority7_module_14_n5), .ZN(
        n_majority7_module_14__or_module_1_res) );
  AND2_X1 u_majority7_module_14__and_module_2_U1 ( .A1(
        n_majority7_module_14_n7), .A2(n_majority7_module_14_n2), .ZN(
        n_majority7_module_14__and_module_2_res) );
  OR2_X1 u_majority7_module_14__or_module_2_U1 ( .A1(n_majority7_module_14_n2), 
        .A2(n_majority7_module_14_n7), .ZN(
        n_majority7_module_14__or_module_2_res) );
  AND2_X1 u_majority7_module_14__and_module_3_U1 ( .A1(
        n_majority7_module_14_n6), .A2(n_majority7_module_14_n1), .ZN(
        n_majority7_module_14__and_module_3_res) );
  OR2_X1 u_majority7_module_14__or_module_3_U1 ( .A1(n_majority7_module_14_n1), 
        .A2(n_majority7_module_14_n6), .ZN(
        n_majority7_module_14__or_module_3_res) );
  AND2_X1 u_majority7_module_14__and_module_4_U1 ( .A1(
        n_majority7_module_14__and_module_2_res), .A2(
        n_majority7_module_14__and_module_1_res), .ZN(
        n_majority7_module_14__and_module_4_res) );
  OR2_X1 u_majority7_module_14__or_module_4_U1 ( .A1(
        n_majority7_module_14__and_module_1_res), .A2(
        n_majority7_module_14__and_module_2_res), .ZN(
        n_majority7_module_14__or_module_4_res) );
  AND2_X1 u_majority7_module_14__and_module_5_U1 ( .A1(
        n_majority7_module_14__and_module_3_res), .A2(n_majority7_module_14_n3), .ZN(n_majority7_module_14__and_module_5_res) );
  OR2_X1 u_majority7_module_14__or_module_5_U1 ( .A1(n_majority7_module_14_n3), 
        .A2(n_majority7_module_14__and_module_3_res), .ZN(
        n_majority7_module_14__or_module_5_res) );
  AND2_X1 u_majority7_module_14__and_module_6_U1 ( .A1(
        n_majority7_module_14__or_module_1_res), .A2(
        n_majority7_module_14__or_module_2_res), .ZN(
        n_majority7_module_14__and_module_6_res) );
  OR2_X1 u_majority7_module_14__or_module_6_U1 ( .A1(
        n_majority7_module_14__or_module_2_res), .A2(
        n_majority7_module_14__or_module_1_res), .ZN(
        n_majority7_module_14__or_module_6_res) );
  OR2_X1 u_majority7_module_14__or_module_7_U1 ( .A1(
        n_majority7_module_14__and_module_4_res), .A2(
        n_majority7_module_14__and_module_5_res), .ZN(
        n_majority7_module_14__or_module_7_res) );
  AND2_X1 u_majority7_module_14__and_module_7_U1 ( .A1(
        n_majority7_module_14__or_module_3_res), .A2(
        n_majority7_module_14__or_module_4_res), .ZN(
        n_majority7_module_14__and_module_7_res) );
  OR2_X1 u_majority7_module_14__or_module_8_U1 ( .A1(
        n_majority7_module_14__or_module_4_res), .A2(
        n_majority7_module_14__or_module_3_res), .ZN(
        n_majority7_module_14__or_module_8_res) );
  AND2_X1 u_majority7_module_14__and_module_8_U1 ( .A1(
        n_majority7_module_14__or_module_5_res), .A2(
        n_majority7_module_14__and_module_6_res), .ZN(
        n_majority7_module_14__and_module_8_res) );
  OR2_X1 u_majority7_module_14__or_module_9_U1 ( .A1(
        n_majority7_module_14__and_module_6_res), .A2(
        n_majority7_module_14__or_module_5_res), .ZN(
        n_majority7_module_14__or_module_9_res) );
  OR2_X1 u_majority7_module_14__or_module_10_U1 ( .A1(
        n_majority7_module_14__or_module_7_res), .A2(
        n_majority7_module_14__and_module_7_res), .ZN(
        n_majority7_module_14__or_module_10_res) );
  AND2_X1 u_majority7_module_14__and_module_9_U1 ( .A1(
        n_majority7_module_14__or_module_6_res), .A2(
        n_majority7_module_14__or_module_9_res), .ZN(
        n_majority7_module_14__and_module_9_res) );
  OR2_X1 u_majority7_module_14__or_module_11_U1 ( .A1(
        n_majority7_module_14__or_module_10_res), .A2(
        n_majority7_module_14__and_module_8_res), .ZN(
        n_majority7_module_14__or_module_11_res) );
  AND2_X1 u_majority7_module_14__and_module_10_U1 ( .A1(
        n_majority7_module_14__or_module_8_res), .A2(
        n_majority7_module_14__and_module_9_res), .ZN(
        n_majority7_module_14__and_module_10_res) );
  AND2_X1 u_majority7_module_14__and_module_11_U1 ( .A1(
        n_majority7_module_14__and_module_10_res), .A2(
        n_majority7_module_14__or_module_11_res), .ZN(
        n_majority7_module_14_res) );
  DFF_X1 u_reg_module_15__cini_mul_v000_reg ( .D(n_majority7_module_14_res), 
        .CK(clock_1), .Q(n_reg_module_15_res), .QN() );
  BUF_X1 u_majority7_module_15_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_15_n7) );
  BUF_X1 u_majority7_module_15_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_15_n6) );
  BUF_X1 u_majority7_module_15_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_15_n5) );
  BUF_X1 u_majority7_module_15_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_15_n4) );
  BUF_X1 u_majority7_module_15_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_15_n3) );
  BUF_X1 u_majority7_module_15_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_15_n2) );
  BUF_X1 u_majority7_module_15_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_15_n1) );
  AND2_X1 u_majority7_module_15__and_module_1_U1 ( .A1(
        n_majority7_module_15_n5), .A2(n_majority7_module_15_n4), .ZN(
        n_majority7_module_15__and_module_1_res) );
  OR2_X1 u_majority7_module_15__or_module_1_U1 ( .A1(n_majority7_module_15_n4), 
        .A2(n_majority7_module_15_n5), .ZN(
        n_majority7_module_15__or_module_1_res) );
  AND2_X1 u_majority7_module_15__and_module_2_U1 ( .A1(
        n_majority7_module_15_n7), .A2(n_majority7_module_15_n2), .ZN(
        n_majority7_module_15__and_module_2_res) );
  OR2_X1 u_majority7_module_15__or_module_2_U1 ( .A1(n_majority7_module_15_n2), 
        .A2(n_majority7_module_15_n7), .ZN(
        n_majority7_module_15__or_module_2_res) );
  AND2_X1 u_majority7_module_15__and_module_3_U1 ( .A1(
        n_majority7_module_15_n6), .A2(n_majority7_module_15_n1), .ZN(
        n_majority7_module_15__and_module_3_res) );
  OR2_X1 u_majority7_module_15__or_module_3_U1 ( .A1(n_majority7_module_15_n1), 
        .A2(n_majority7_module_15_n6), .ZN(
        n_majority7_module_15__or_module_3_res) );
  AND2_X1 u_majority7_module_15__and_module_4_U1 ( .A1(
        n_majority7_module_15__and_module_2_res), .A2(
        n_majority7_module_15__and_module_1_res), .ZN(
        n_majority7_module_15__and_module_4_res) );
  OR2_X1 u_majority7_module_15__or_module_4_U1 ( .A1(
        n_majority7_module_15__and_module_1_res), .A2(
        n_majority7_module_15__and_module_2_res), .ZN(
        n_majority7_module_15__or_module_4_res) );
  AND2_X1 u_majority7_module_15__and_module_5_U1 ( .A1(
        n_majority7_module_15__and_module_3_res), .A2(n_majority7_module_15_n3), .ZN(n_majority7_module_15__and_module_5_res) );
  OR2_X1 u_majority7_module_15__or_module_5_U1 ( .A1(n_majority7_module_15_n3), 
        .A2(n_majority7_module_15__and_module_3_res), .ZN(
        n_majority7_module_15__or_module_5_res) );
  AND2_X1 u_majority7_module_15__and_module_6_U1 ( .A1(
        n_majority7_module_15__or_module_1_res), .A2(
        n_majority7_module_15__or_module_2_res), .ZN(
        n_majority7_module_15__and_module_6_res) );
  OR2_X1 u_majority7_module_15__or_module_6_U1 ( .A1(
        n_majority7_module_15__or_module_2_res), .A2(
        n_majority7_module_15__or_module_1_res), .ZN(
        n_majority7_module_15__or_module_6_res) );
  OR2_X1 u_majority7_module_15__or_module_7_U1 ( .A1(
        n_majority7_module_15__and_module_4_res), .A2(
        n_majority7_module_15__and_module_5_res), .ZN(
        n_majority7_module_15__or_module_7_res) );
  AND2_X1 u_majority7_module_15__and_module_7_U1 ( .A1(
        n_majority7_module_15__or_module_3_res), .A2(
        n_majority7_module_15__or_module_4_res), .ZN(
        n_majority7_module_15__and_module_7_res) );
  OR2_X1 u_majority7_module_15__or_module_8_U1 ( .A1(
        n_majority7_module_15__or_module_4_res), .A2(
        n_majority7_module_15__or_module_3_res), .ZN(
        n_majority7_module_15__or_module_8_res) );
  AND2_X1 u_majority7_module_15__and_module_8_U1 ( .A1(
        n_majority7_module_15__or_module_5_res), .A2(
        n_majority7_module_15__and_module_6_res), .ZN(
        n_majority7_module_15__and_module_8_res) );
  OR2_X1 u_majority7_module_15__or_module_9_U1 ( .A1(
        n_majority7_module_15__and_module_6_res), .A2(
        n_majority7_module_15__or_module_5_res), .ZN(
        n_majority7_module_15__or_module_9_res) );
  OR2_X1 u_majority7_module_15__or_module_10_U1 ( .A1(
        n_majority7_module_15__or_module_7_res), .A2(
        n_majority7_module_15__and_module_7_res), .ZN(
        n_majority7_module_15__or_module_10_res) );
  AND2_X1 u_majority7_module_15__and_module_9_U1 ( .A1(
        n_majority7_module_15__or_module_6_res), .A2(
        n_majority7_module_15__or_module_9_res), .ZN(
        n_majority7_module_15__and_module_9_res) );
  OR2_X1 u_majority7_module_15__or_module_11_U1 ( .A1(
        n_majority7_module_15__or_module_10_res), .A2(
        n_majority7_module_15__and_module_8_res), .ZN(
        n_majority7_module_15__or_module_11_res) );
  AND2_X1 u_majority7_module_15__and_module_10_U1 ( .A1(
        n_majority7_module_15__or_module_8_res), .A2(
        n_majority7_module_15__and_module_9_res), .ZN(
        n_majority7_module_15__and_module_10_res) );
  AND2_X1 u_majority7_module_15__and_module_11_U1 ( .A1(
        n_majority7_module_15__and_module_10_res), .A2(
        n_majority7_module_15__or_module_11_res), .ZN(
        n_majority7_module_15_res) );
  DFF_X1 u_reg_module_16__cini_mul_v000_reg ( .D(n_majority7_module_15_res), 
        .CK(clock_1), .Q(n_reg_module_16_res), .QN() );
  BUF_X1 u_majority7_module_16_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_16_n7) );
  BUF_X1 u_majority7_module_16_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_16_n6) );
  BUF_X1 u_majority7_module_16_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_16_n5) );
  BUF_X1 u_majority7_module_16_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_16_n4) );
  BUF_X1 u_majority7_module_16_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_16_n3) );
  BUF_X1 u_majority7_module_16_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_16_n2) );
  BUF_X1 u_majority7_module_16_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_16_n1) );
  AND2_X1 u_majority7_module_16__and_module_1_U1 ( .A1(
        n_majority7_module_16_n5), .A2(n_majority7_module_16_n4), .ZN(
        n_majority7_module_16__and_module_1_res) );
  OR2_X1 u_majority7_module_16__or_module_1_U1 ( .A1(n_majority7_module_16_n4), 
        .A2(n_majority7_module_16_n5), .ZN(
        n_majority7_module_16__or_module_1_res) );
  AND2_X1 u_majority7_module_16__and_module_2_U1 ( .A1(
        n_majority7_module_16_n7), .A2(n_majority7_module_16_n2), .ZN(
        n_majority7_module_16__and_module_2_res) );
  OR2_X1 u_majority7_module_16__or_module_2_U1 ( .A1(n_majority7_module_16_n2), 
        .A2(n_majority7_module_16_n7), .ZN(
        n_majority7_module_16__or_module_2_res) );
  AND2_X1 u_majority7_module_16__and_module_3_U1 ( .A1(
        n_majority7_module_16_n6), .A2(n_majority7_module_16_n1), .ZN(
        n_majority7_module_16__and_module_3_res) );
  OR2_X1 u_majority7_module_16__or_module_3_U1 ( .A1(n_majority7_module_16_n1), 
        .A2(n_majority7_module_16_n6), .ZN(
        n_majority7_module_16__or_module_3_res) );
  AND2_X1 u_majority7_module_16__and_module_4_U1 ( .A1(
        n_majority7_module_16__and_module_2_res), .A2(
        n_majority7_module_16__and_module_1_res), .ZN(
        n_majority7_module_16__and_module_4_res) );
  OR2_X1 u_majority7_module_16__or_module_4_U1 ( .A1(
        n_majority7_module_16__and_module_1_res), .A2(
        n_majority7_module_16__and_module_2_res), .ZN(
        n_majority7_module_16__or_module_4_res) );
  AND2_X1 u_majority7_module_16__and_module_5_U1 ( .A1(
        n_majority7_module_16__and_module_3_res), .A2(n_majority7_module_16_n3), .ZN(n_majority7_module_16__and_module_5_res) );
  OR2_X1 u_majority7_module_16__or_module_5_U1 ( .A1(n_majority7_module_16_n3), 
        .A2(n_majority7_module_16__and_module_3_res), .ZN(
        n_majority7_module_16__or_module_5_res) );
  AND2_X1 u_majority7_module_16__and_module_6_U1 ( .A1(
        n_majority7_module_16__or_module_1_res), .A2(
        n_majority7_module_16__or_module_2_res), .ZN(
        n_majority7_module_16__and_module_6_res) );
  OR2_X1 u_majority7_module_16__or_module_6_U1 ( .A1(
        n_majority7_module_16__or_module_2_res), .A2(
        n_majority7_module_16__or_module_1_res), .ZN(
        n_majority7_module_16__or_module_6_res) );
  OR2_X1 u_majority7_module_16__or_module_7_U1 ( .A1(
        n_majority7_module_16__and_module_4_res), .A2(
        n_majority7_module_16__and_module_5_res), .ZN(
        n_majority7_module_16__or_module_7_res) );
  AND2_X1 u_majority7_module_16__and_module_7_U1 ( .A1(
        n_majority7_module_16__or_module_3_res), .A2(
        n_majority7_module_16__or_module_4_res), .ZN(
        n_majority7_module_16__and_module_7_res) );
  OR2_X1 u_majority7_module_16__or_module_8_U1 ( .A1(
        n_majority7_module_16__or_module_4_res), .A2(
        n_majority7_module_16__or_module_3_res), .ZN(
        n_majority7_module_16__or_module_8_res) );
  AND2_X1 u_majority7_module_16__and_module_8_U1 ( .A1(
        n_majority7_module_16__or_module_5_res), .A2(
        n_majority7_module_16__and_module_6_res), .ZN(
        n_majority7_module_16__and_module_8_res) );
  OR2_X1 u_majority7_module_16__or_module_9_U1 ( .A1(
        n_majority7_module_16__and_module_6_res), .A2(
        n_majority7_module_16__or_module_5_res), .ZN(
        n_majority7_module_16__or_module_9_res) );
  OR2_X1 u_majority7_module_16__or_module_10_U1 ( .A1(
        n_majority7_module_16__or_module_7_res), .A2(
        n_majority7_module_16__and_module_7_res), .ZN(
        n_majority7_module_16__or_module_10_res) );
  AND2_X1 u_majority7_module_16__and_module_9_U1 ( .A1(
        n_majority7_module_16__or_module_6_res), .A2(
        n_majority7_module_16__or_module_9_res), .ZN(
        n_majority7_module_16__and_module_9_res) );
  OR2_X1 u_majority7_module_16__or_module_11_U1 ( .A1(
        n_majority7_module_16__or_module_10_res), .A2(
        n_majority7_module_16__and_module_8_res), .ZN(
        n_majority7_module_16__or_module_11_res) );
  AND2_X1 u_majority7_module_16__and_module_10_U1 ( .A1(
        n_majority7_module_16__or_module_8_res), .A2(
        n_majority7_module_16__and_module_9_res), .ZN(
        n_majority7_module_16__and_module_10_res) );
  AND2_X1 u_majority7_module_16__and_module_11_U1 ( .A1(
        n_majority7_module_16__and_module_10_res), .A2(
        n_majority7_module_16__or_module_11_res), .ZN(
        n_majority7_module_16_res) );
  DFF_X1 u_reg_module_17__cini_mul_v000_reg ( .D(n_majority7_module_16_res), 
        .CK(clock_1), .Q(n_reg_module_17_res), .QN() );
  BUF_X1 u_majority7_module_17_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_17_n7) );
  BUF_X1 u_majority7_module_17_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_17_n6) );
  BUF_X1 u_majority7_module_17_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_17_n5) );
  BUF_X1 u_majority7_module_17_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_17_n4) );
  BUF_X1 u_majority7_module_17_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_17_n3) );
  BUF_X1 u_majority7_module_17_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_17_n2) );
  BUF_X1 u_majority7_module_17_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_17_n1) );
  AND2_X1 u_majority7_module_17__and_module_1_U1 ( .A1(
        n_majority7_module_17_n5), .A2(n_majority7_module_17_n4), .ZN(
        n_majority7_module_17__and_module_1_res) );
  OR2_X1 u_majority7_module_17__or_module_1_U1 ( .A1(n_majority7_module_17_n4), 
        .A2(n_majority7_module_17_n5), .ZN(
        n_majority7_module_17__or_module_1_res) );
  AND2_X1 u_majority7_module_17__and_module_2_U1 ( .A1(
        n_majority7_module_17_n7), .A2(n_majority7_module_17_n2), .ZN(
        n_majority7_module_17__and_module_2_res) );
  OR2_X1 u_majority7_module_17__or_module_2_U1 ( .A1(n_majority7_module_17_n2), 
        .A2(n_majority7_module_17_n7), .ZN(
        n_majority7_module_17__or_module_2_res) );
  AND2_X1 u_majority7_module_17__and_module_3_U1 ( .A1(
        n_majority7_module_17_n6), .A2(n_majority7_module_17_n1), .ZN(
        n_majority7_module_17__and_module_3_res) );
  OR2_X1 u_majority7_module_17__or_module_3_U1 ( .A1(n_majority7_module_17_n1), 
        .A2(n_majority7_module_17_n6), .ZN(
        n_majority7_module_17__or_module_3_res) );
  AND2_X1 u_majority7_module_17__and_module_4_U1 ( .A1(
        n_majority7_module_17__and_module_2_res), .A2(
        n_majority7_module_17__and_module_1_res), .ZN(
        n_majority7_module_17__and_module_4_res) );
  OR2_X1 u_majority7_module_17__or_module_4_U1 ( .A1(
        n_majority7_module_17__and_module_1_res), .A2(
        n_majority7_module_17__and_module_2_res), .ZN(
        n_majority7_module_17__or_module_4_res) );
  AND2_X1 u_majority7_module_17__and_module_5_U1 ( .A1(
        n_majority7_module_17__and_module_3_res), .A2(n_majority7_module_17_n3), .ZN(n_majority7_module_17__and_module_5_res) );
  OR2_X1 u_majority7_module_17__or_module_5_U1 ( .A1(n_majority7_module_17_n3), 
        .A2(n_majority7_module_17__and_module_3_res), .ZN(
        n_majority7_module_17__or_module_5_res) );
  AND2_X1 u_majority7_module_17__and_module_6_U1 ( .A1(
        n_majority7_module_17__or_module_1_res), .A2(
        n_majority7_module_17__or_module_2_res), .ZN(
        n_majority7_module_17__and_module_6_res) );
  OR2_X1 u_majority7_module_17__or_module_6_U1 ( .A1(
        n_majority7_module_17__or_module_2_res), .A2(
        n_majority7_module_17__or_module_1_res), .ZN(
        n_majority7_module_17__or_module_6_res) );
  OR2_X1 u_majority7_module_17__or_module_7_U1 ( .A1(
        n_majority7_module_17__and_module_4_res), .A2(
        n_majority7_module_17__and_module_5_res), .ZN(
        n_majority7_module_17__or_module_7_res) );
  AND2_X1 u_majority7_module_17__and_module_7_U1 ( .A1(
        n_majority7_module_17__or_module_3_res), .A2(
        n_majority7_module_17__or_module_4_res), .ZN(
        n_majority7_module_17__and_module_7_res) );
  OR2_X1 u_majority7_module_17__or_module_8_U1 ( .A1(
        n_majority7_module_17__or_module_4_res), .A2(
        n_majority7_module_17__or_module_3_res), .ZN(
        n_majority7_module_17__or_module_8_res) );
  AND2_X1 u_majority7_module_17__and_module_8_U1 ( .A1(
        n_majority7_module_17__or_module_5_res), .A2(
        n_majority7_module_17__and_module_6_res), .ZN(
        n_majority7_module_17__and_module_8_res) );
  OR2_X1 u_majority7_module_17__or_module_9_U1 ( .A1(
        n_majority7_module_17__and_module_6_res), .A2(
        n_majority7_module_17__or_module_5_res), .ZN(
        n_majority7_module_17__or_module_9_res) );
  OR2_X1 u_majority7_module_17__or_module_10_U1 ( .A1(
        n_majority7_module_17__or_module_7_res), .A2(
        n_majority7_module_17__and_module_7_res), .ZN(
        n_majority7_module_17__or_module_10_res) );
  AND2_X1 u_majority7_module_17__and_module_9_U1 ( .A1(
        n_majority7_module_17__or_module_6_res), .A2(
        n_majority7_module_17__or_module_9_res), .ZN(
        n_majority7_module_17__and_module_9_res) );
  OR2_X1 u_majority7_module_17__or_module_11_U1 ( .A1(
        n_majority7_module_17__or_module_10_res), .A2(
        n_majority7_module_17__and_module_8_res), .ZN(
        n_majority7_module_17__or_module_11_res) );
  AND2_X1 u_majority7_module_17__and_module_10_U1 ( .A1(
        n_majority7_module_17__or_module_8_res), .A2(
        n_majority7_module_17__and_module_9_res), .ZN(
        n_majority7_module_17__and_module_10_res) );
  AND2_X1 u_majority7_module_17__and_module_11_U1 ( .A1(
        n_majority7_module_17__and_module_10_res), .A2(
        n_majority7_module_17__or_module_11_res), .ZN(
        n_majority7_module_17_res) );
  DFF_X1 u_reg_module_18__cini_mul_v000_reg ( .D(n_majority7_module_17_res), 
        .CK(clock_1), .Q(n_reg_module_18_res), .QN() );
  BUF_X1 u_majority7_module_18_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_18_n7) );
  BUF_X1 u_majority7_module_18_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_18_n6) );
  BUF_X1 u_majority7_module_18_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_18_n5) );
  BUF_X1 u_majority7_module_18_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_18_n4) );
  BUF_X1 u_majority7_module_18_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_18_n3) );
  BUF_X1 u_majority7_module_18_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_18_n2) );
  BUF_X1 u_majority7_module_18_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_18_n1) );
  AND2_X1 u_majority7_module_18__and_module_1_U1 ( .A1(
        n_majority7_module_18_n5), .A2(n_majority7_module_18_n4), .ZN(
        n_majority7_module_18__and_module_1_res) );
  OR2_X1 u_majority7_module_18__or_module_1_U1 ( .A1(n_majority7_module_18_n4), 
        .A2(n_majority7_module_18_n5), .ZN(
        n_majority7_module_18__or_module_1_res) );
  AND2_X1 u_majority7_module_18__and_module_2_U1 ( .A1(
        n_majority7_module_18_n7), .A2(n_majority7_module_18_n2), .ZN(
        n_majority7_module_18__and_module_2_res) );
  OR2_X1 u_majority7_module_18__or_module_2_U1 ( .A1(n_majority7_module_18_n2), 
        .A2(n_majority7_module_18_n7), .ZN(
        n_majority7_module_18__or_module_2_res) );
  AND2_X1 u_majority7_module_18__and_module_3_U1 ( .A1(
        n_majority7_module_18_n6), .A2(n_majority7_module_18_n1), .ZN(
        n_majority7_module_18__and_module_3_res) );
  OR2_X1 u_majority7_module_18__or_module_3_U1 ( .A1(n_majority7_module_18_n1), 
        .A2(n_majority7_module_18_n6), .ZN(
        n_majority7_module_18__or_module_3_res) );
  AND2_X1 u_majority7_module_18__and_module_4_U1 ( .A1(
        n_majority7_module_18__and_module_2_res), .A2(
        n_majority7_module_18__and_module_1_res), .ZN(
        n_majority7_module_18__and_module_4_res) );
  OR2_X1 u_majority7_module_18__or_module_4_U1 ( .A1(
        n_majority7_module_18__and_module_1_res), .A2(
        n_majority7_module_18__and_module_2_res), .ZN(
        n_majority7_module_18__or_module_4_res) );
  AND2_X1 u_majority7_module_18__and_module_5_U1 ( .A1(
        n_majority7_module_18__and_module_3_res), .A2(n_majority7_module_18_n3), .ZN(n_majority7_module_18__and_module_5_res) );
  OR2_X1 u_majority7_module_18__or_module_5_U1 ( .A1(n_majority7_module_18_n3), 
        .A2(n_majority7_module_18__and_module_3_res), .ZN(
        n_majority7_module_18__or_module_5_res) );
  AND2_X1 u_majority7_module_18__and_module_6_U1 ( .A1(
        n_majority7_module_18__or_module_1_res), .A2(
        n_majority7_module_18__or_module_2_res), .ZN(
        n_majority7_module_18__and_module_6_res) );
  OR2_X1 u_majority7_module_18__or_module_6_U1 ( .A1(
        n_majority7_module_18__or_module_2_res), .A2(
        n_majority7_module_18__or_module_1_res), .ZN(
        n_majority7_module_18__or_module_6_res) );
  OR2_X1 u_majority7_module_18__or_module_7_U1 ( .A1(
        n_majority7_module_18__and_module_4_res), .A2(
        n_majority7_module_18__and_module_5_res), .ZN(
        n_majority7_module_18__or_module_7_res) );
  AND2_X1 u_majority7_module_18__and_module_7_U1 ( .A1(
        n_majority7_module_18__or_module_3_res), .A2(
        n_majority7_module_18__or_module_4_res), .ZN(
        n_majority7_module_18__and_module_7_res) );
  OR2_X1 u_majority7_module_18__or_module_8_U1 ( .A1(
        n_majority7_module_18__or_module_4_res), .A2(
        n_majority7_module_18__or_module_3_res), .ZN(
        n_majority7_module_18__or_module_8_res) );
  AND2_X1 u_majority7_module_18__and_module_8_U1 ( .A1(
        n_majority7_module_18__or_module_5_res), .A2(
        n_majority7_module_18__and_module_6_res), .ZN(
        n_majority7_module_18__and_module_8_res) );
  OR2_X1 u_majority7_module_18__or_module_9_U1 ( .A1(
        n_majority7_module_18__and_module_6_res), .A2(
        n_majority7_module_18__or_module_5_res), .ZN(
        n_majority7_module_18__or_module_9_res) );
  OR2_X1 u_majority7_module_18__or_module_10_U1 ( .A1(
        n_majority7_module_18__or_module_7_res), .A2(
        n_majority7_module_18__and_module_7_res), .ZN(
        n_majority7_module_18__or_module_10_res) );
  AND2_X1 u_majority7_module_18__and_module_9_U1 ( .A1(
        n_majority7_module_18__or_module_6_res), .A2(
        n_majority7_module_18__or_module_9_res), .ZN(
        n_majority7_module_18__and_module_9_res) );
  OR2_X1 u_majority7_module_18__or_module_11_U1 ( .A1(
        n_majority7_module_18__or_module_10_res), .A2(
        n_majority7_module_18__and_module_8_res), .ZN(
        n_majority7_module_18__or_module_11_res) );
  AND2_X1 u_majority7_module_18__and_module_10_U1 ( .A1(
        n_majority7_module_18__or_module_8_res), .A2(
        n_majority7_module_18__and_module_9_res), .ZN(
        n_majority7_module_18__and_module_10_res) );
  AND2_X1 u_majority7_module_18__and_module_11_U1 ( .A1(
        n_majority7_module_18__and_module_10_res), .A2(
        n_majority7_module_18__or_module_11_res), .ZN(
        n_majority7_module_18_res) );
  DFF_X1 u_reg_module_19__cini_mul_v000_reg ( .D(n_majority7_module_18_res), 
        .CK(clock_2), .Q(n_reg_module_19_res), .QN() );
  BUF_X1 u_majority7_module_19_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_19_n7) );
  BUF_X1 u_majority7_module_19_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_19_n6) );
  BUF_X1 u_majority7_module_19_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_19_n5) );
  BUF_X1 u_majority7_module_19_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_19_n4) );
  BUF_X1 u_majority7_module_19_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_19_n3) );
  BUF_X1 u_majority7_module_19_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_19_n2) );
  BUF_X1 u_majority7_module_19_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_19_n1) );
  AND2_X1 u_majority7_module_19__and_module_1_U1 ( .A1(
        n_majority7_module_19_n5), .A2(n_majority7_module_19_n4), .ZN(
        n_majority7_module_19__and_module_1_res) );
  OR2_X1 u_majority7_module_19__or_module_1_U1 ( .A1(n_majority7_module_19_n4), 
        .A2(n_majority7_module_19_n5), .ZN(
        n_majority7_module_19__or_module_1_res) );
  AND2_X1 u_majority7_module_19__and_module_2_U1 ( .A1(
        n_majority7_module_19_n7), .A2(n_majority7_module_19_n2), .ZN(
        n_majority7_module_19__and_module_2_res) );
  OR2_X1 u_majority7_module_19__or_module_2_U1 ( .A1(n_majority7_module_19_n2), 
        .A2(n_majority7_module_19_n7), .ZN(
        n_majority7_module_19__or_module_2_res) );
  AND2_X1 u_majority7_module_19__and_module_3_U1 ( .A1(
        n_majority7_module_19_n6), .A2(n_majority7_module_19_n1), .ZN(
        n_majority7_module_19__and_module_3_res) );
  OR2_X1 u_majority7_module_19__or_module_3_U1 ( .A1(n_majority7_module_19_n1), 
        .A2(n_majority7_module_19_n6), .ZN(
        n_majority7_module_19__or_module_3_res) );
  AND2_X1 u_majority7_module_19__and_module_4_U1 ( .A1(
        n_majority7_module_19__and_module_2_res), .A2(
        n_majority7_module_19__and_module_1_res), .ZN(
        n_majority7_module_19__and_module_4_res) );
  OR2_X1 u_majority7_module_19__or_module_4_U1 ( .A1(
        n_majority7_module_19__and_module_1_res), .A2(
        n_majority7_module_19__and_module_2_res), .ZN(
        n_majority7_module_19__or_module_4_res) );
  AND2_X1 u_majority7_module_19__and_module_5_U1 ( .A1(
        n_majority7_module_19__and_module_3_res), .A2(n_majority7_module_19_n3), .ZN(n_majority7_module_19__and_module_5_res) );
  OR2_X1 u_majority7_module_19__or_module_5_U1 ( .A1(n_majority7_module_19_n3), 
        .A2(n_majority7_module_19__and_module_3_res), .ZN(
        n_majority7_module_19__or_module_5_res) );
  AND2_X1 u_majority7_module_19__and_module_6_U1 ( .A1(
        n_majority7_module_19__or_module_1_res), .A2(
        n_majority7_module_19__or_module_2_res), .ZN(
        n_majority7_module_19__and_module_6_res) );
  OR2_X1 u_majority7_module_19__or_module_6_U1 ( .A1(
        n_majority7_module_19__or_module_2_res), .A2(
        n_majority7_module_19__or_module_1_res), .ZN(
        n_majority7_module_19__or_module_6_res) );
  OR2_X1 u_majority7_module_19__or_module_7_U1 ( .A1(
        n_majority7_module_19__and_module_4_res), .A2(
        n_majority7_module_19__and_module_5_res), .ZN(
        n_majority7_module_19__or_module_7_res) );
  AND2_X1 u_majority7_module_19__and_module_7_U1 ( .A1(
        n_majority7_module_19__or_module_3_res), .A2(
        n_majority7_module_19__or_module_4_res), .ZN(
        n_majority7_module_19__and_module_7_res) );
  OR2_X1 u_majority7_module_19__or_module_8_U1 ( .A1(
        n_majority7_module_19__or_module_4_res), .A2(
        n_majority7_module_19__or_module_3_res), .ZN(
        n_majority7_module_19__or_module_8_res) );
  AND2_X1 u_majority7_module_19__and_module_8_U1 ( .A1(
        n_majority7_module_19__or_module_5_res), .A2(
        n_majority7_module_19__and_module_6_res), .ZN(
        n_majority7_module_19__and_module_8_res) );
  OR2_X1 u_majority7_module_19__or_module_9_U1 ( .A1(
        n_majority7_module_19__and_module_6_res), .A2(
        n_majority7_module_19__or_module_5_res), .ZN(
        n_majority7_module_19__or_module_9_res) );
  OR2_X1 u_majority7_module_19__or_module_10_U1 ( .A1(
        n_majority7_module_19__or_module_7_res), .A2(
        n_majority7_module_19__and_module_7_res), .ZN(
        n_majority7_module_19__or_module_10_res) );
  AND2_X1 u_majority7_module_19__and_module_9_U1 ( .A1(
        n_majority7_module_19__or_module_6_res), .A2(
        n_majority7_module_19__or_module_9_res), .ZN(
        n_majority7_module_19__and_module_9_res) );
  OR2_X1 u_majority7_module_19__or_module_11_U1 ( .A1(
        n_majority7_module_19__or_module_10_res), .A2(
        n_majority7_module_19__and_module_8_res), .ZN(
        n_majority7_module_19__or_module_11_res) );
  AND2_X1 u_majority7_module_19__and_module_10_U1 ( .A1(
        n_majority7_module_19__or_module_8_res), .A2(
        n_majority7_module_19__and_module_9_res), .ZN(
        n_majority7_module_19__and_module_10_res) );
  AND2_X1 u_majority7_module_19__and_module_11_U1 ( .A1(
        n_majority7_module_19__and_module_10_res), .A2(
        n_majority7_module_19__or_module_11_res), .ZN(
        n_majority7_module_19_res) );
  DFF_X1 u_reg_module_20__cini_mul_v000_reg ( .D(n_majority7_module_19_res), 
        .CK(clock_2), .Q(n_reg_module_20_res), .QN() );
  BUF_X1 u_majority7_module_20_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_20_n7) );
  BUF_X1 u_majority7_module_20_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_20_n6) );
  BUF_X1 u_majority7_module_20_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_20_n5) );
  BUF_X1 u_majority7_module_20_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_20_n4) );
  BUF_X1 u_majority7_module_20_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_20_n3) );
  BUF_X1 u_majority7_module_20_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_20_n2) );
  BUF_X1 u_majority7_module_20_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_20_n1) );
  AND2_X1 u_majority7_module_20__and_module_1_U1 ( .A1(
        n_majority7_module_20_n5), .A2(n_majority7_module_20_n4), .ZN(
        n_majority7_module_20__and_module_1_res) );
  OR2_X1 u_majority7_module_20__or_module_1_U1 ( .A1(n_majority7_module_20_n4), 
        .A2(n_majority7_module_20_n5), .ZN(
        n_majority7_module_20__or_module_1_res) );
  AND2_X1 u_majority7_module_20__and_module_2_U1 ( .A1(
        n_majority7_module_20_n7), .A2(n_majority7_module_20_n2), .ZN(
        n_majority7_module_20__and_module_2_res) );
  OR2_X1 u_majority7_module_20__or_module_2_U1 ( .A1(n_majority7_module_20_n2), 
        .A2(n_majority7_module_20_n7), .ZN(
        n_majority7_module_20__or_module_2_res) );
  AND2_X1 u_majority7_module_20__and_module_3_U1 ( .A1(
        n_majority7_module_20_n6), .A2(n_majority7_module_20_n1), .ZN(
        n_majority7_module_20__and_module_3_res) );
  OR2_X1 u_majority7_module_20__or_module_3_U1 ( .A1(n_majority7_module_20_n1), 
        .A2(n_majority7_module_20_n6), .ZN(
        n_majority7_module_20__or_module_3_res) );
  AND2_X1 u_majority7_module_20__and_module_4_U1 ( .A1(
        n_majority7_module_20__and_module_2_res), .A2(
        n_majority7_module_20__and_module_1_res), .ZN(
        n_majority7_module_20__and_module_4_res) );
  OR2_X1 u_majority7_module_20__or_module_4_U1 ( .A1(
        n_majority7_module_20__and_module_1_res), .A2(
        n_majority7_module_20__and_module_2_res), .ZN(
        n_majority7_module_20__or_module_4_res) );
  AND2_X1 u_majority7_module_20__and_module_5_U1 ( .A1(
        n_majority7_module_20__and_module_3_res), .A2(n_majority7_module_20_n3), .ZN(n_majority7_module_20__and_module_5_res) );
  OR2_X1 u_majority7_module_20__or_module_5_U1 ( .A1(n_majority7_module_20_n3), 
        .A2(n_majority7_module_20__and_module_3_res), .ZN(
        n_majority7_module_20__or_module_5_res) );
  AND2_X1 u_majority7_module_20__and_module_6_U1 ( .A1(
        n_majority7_module_20__or_module_1_res), .A2(
        n_majority7_module_20__or_module_2_res), .ZN(
        n_majority7_module_20__and_module_6_res) );
  OR2_X1 u_majority7_module_20__or_module_6_U1 ( .A1(
        n_majority7_module_20__or_module_2_res), .A2(
        n_majority7_module_20__or_module_1_res), .ZN(
        n_majority7_module_20__or_module_6_res) );
  OR2_X1 u_majority7_module_20__or_module_7_U1 ( .A1(
        n_majority7_module_20__and_module_4_res), .A2(
        n_majority7_module_20__and_module_5_res), .ZN(
        n_majority7_module_20__or_module_7_res) );
  AND2_X1 u_majority7_module_20__and_module_7_U1 ( .A1(
        n_majority7_module_20__or_module_3_res), .A2(
        n_majority7_module_20__or_module_4_res), .ZN(
        n_majority7_module_20__and_module_7_res) );
  OR2_X1 u_majority7_module_20__or_module_8_U1 ( .A1(
        n_majority7_module_20__or_module_4_res), .A2(
        n_majority7_module_20__or_module_3_res), .ZN(
        n_majority7_module_20__or_module_8_res) );
  AND2_X1 u_majority7_module_20__and_module_8_U1 ( .A1(
        n_majority7_module_20__or_module_5_res), .A2(
        n_majority7_module_20__and_module_6_res), .ZN(
        n_majority7_module_20__and_module_8_res) );
  OR2_X1 u_majority7_module_20__or_module_9_U1 ( .A1(
        n_majority7_module_20__and_module_6_res), .A2(
        n_majority7_module_20__or_module_5_res), .ZN(
        n_majority7_module_20__or_module_9_res) );
  OR2_X1 u_majority7_module_20__or_module_10_U1 ( .A1(
        n_majority7_module_20__or_module_7_res), .A2(
        n_majority7_module_20__and_module_7_res), .ZN(
        n_majority7_module_20__or_module_10_res) );
  AND2_X1 u_majority7_module_20__and_module_9_U1 ( .A1(
        n_majority7_module_20__or_module_6_res), .A2(
        n_majority7_module_20__or_module_9_res), .ZN(
        n_majority7_module_20__and_module_9_res) );
  OR2_X1 u_majority7_module_20__or_module_11_U1 ( .A1(
        n_majority7_module_20__or_module_10_res), .A2(
        n_majority7_module_20__and_module_8_res), .ZN(
        n_majority7_module_20__or_module_11_res) );
  AND2_X1 u_majority7_module_20__and_module_10_U1 ( .A1(
        n_majority7_module_20__or_module_8_res), .A2(
        n_majority7_module_20__and_module_9_res), .ZN(
        n_majority7_module_20__and_module_10_res) );
  AND2_X1 u_majority7_module_20__and_module_11_U1 ( .A1(
        n_majority7_module_20__and_module_10_res), .A2(
        n_majority7_module_20__or_module_11_res), .ZN(
        n_majority7_module_20_res) );
  DFF_X1 u_reg_module_21__cini_mul_v000_reg ( .D(n_majority7_module_20_res), 
        .CK(clock_2), .Q(n_reg_module_21_res), .QN() );
  BUF_X1 u_majority7_module_21_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_21_n7) );
  BUF_X1 u_majority7_module_21_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_21_n6) );
  BUF_X1 u_majority7_module_21_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_21_n5) );
  BUF_X1 u_majority7_module_21_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_21_n4) );
  BUF_X1 u_majority7_module_21_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_21_n3) );
  BUF_X1 u_majority7_module_21_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_21_n2) );
  BUF_X1 u_majority7_module_21_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_21_n1) );
  AND2_X1 u_majority7_module_21__and_module_1_U1 ( .A1(
        n_majority7_module_21_n5), .A2(n_majority7_module_21_n4), .ZN(
        n_majority7_module_21__and_module_1_res) );
  OR2_X1 u_majority7_module_21__or_module_1_U1 ( .A1(n_majority7_module_21_n4), 
        .A2(n_majority7_module_21_n5), .ZN(
        n_majority7_module_21__or_module_1_res) );
  AND2_X1 u_majority7_module_21__and_module_2_U1 ( .A1(
        n_majority7_module_21_n7), .A2(n_majority7_module_21_n2), .ZN(
        n_majority7_module_21__and_module_2_res) );
  OR2_X1 u_majority7_module_21__or_module_2_U1 ( .A1(n_majority7_module_21_n2), 
        .A2(n_majority7_module_21_n7), .ZN(
        n_majority7_module_21__or_module_2_res) );
  AND2_X1 u_majority7_module_21__and_module_3_U1 ( .A1(
        n_majority7_module_21_n6), .A2(n_majority7_module_21_n1), .ZN(
        n_majority7_module_21__and_module_3_res) );
  OR2_X1 u_majority7_module_21__or_module_3_U1 ( .A1(n_majority7_module_21_n1), 
        .A2(n_majority7_module_21_n6), .ZN(
        n_majority7_module_21__or_module_3_res) );
  AND2_X1 u_majority7_module_21__and_module_4_U1 ( .A1(
        n_majority7_module_21__and_module_2_res), .A2(
        n_majority7_module_21__and_module_1_res), .ZN(
        n_majority7_module_21__and_module_4_res) );
  OR2_X1 u_majority7_module_21__or_module_4_U1 ( .A1(
        n_majority7_module_21__and_module_1_res), .A2(
        n_majority7_module_21__and_module_2_res), .ZN(
        n_majority7_module_21__or_module_4_res) );
  AND2_X1 u_majority7_module_21__and_module_5_U1 ( .A1(
        n_majority7_module_21__and_module_3_res), .A2(n_majority7_module_21_n3), .ZN(n_majority7_module_21__and_module_5_res) );
  OR2_X1 u_majority7_module_21__or_module_5_U1 ( .A1(n_majority7_module_21_n3), 
        .A2(n_majority7_module_21__and_module_3_res), .ZN(
        n_majority7_module_21__or_module_5_res) );
  AND2_X1 u_majority7_module_21__and_module_6_U1 ( .A1(
        n_majority7_module_21__or_module_1_res), .A2(
        n_majority7_module_21__or_module_2_res), .ZN(
        n_majority7_module_21__and_module_6_res) );
  OR2_X1 u_majority7_module_21__or_module_6_U1 ( .A1(
        n_majority7_module_21__or_module_2_res), .A2(
        n_majority7_module_21__or_module_1_res), .ZN(
        n_majority7_module_21__or_module_6_res) );
  OR2_X1 u_majority7_module_21__or_module_7_U1 ( .A1(
        n_majority7_module_21__and_module_4_res), .A2(
        n_majority7_module_21__and_module_5_res), .ZN(
        n_majority7_module_21__or_module_7_res) );
  AND2_X1 u_majority7_module_21__and_module_7_U1 ( .A1(
        n_majority7_module_21__or_module_3_res), .A2(
        n_majority7_module_21__or_module_4_res), .ZN(
        n_majority7_module_21__and_module_7_res) );
  OR2_X1 u_majority7_module_21__or_module_8_U1 ( .A1(
        n_majority7_module_21__or_module_4_res), .A2(
        n_majority7_module_21__or_module_3_res), .ZN(
        n_majority7_module_21__or_module_8_res) );
  AND2_X1 u_majority7_module_21__and_module_8_U1 ( .A1(
        n_majority7_module_21__or_module_5_res), .A2(
        n_majority7_module_21__and_module_6_res), .ZN(
        n_majority7_module_21__and_module_8_res) );
  OR2_X1 u_majority7_module_21__or_module_9_U1 ( .A1(
        n_majority7_module_21__and_module_6_res), .A2(
        n_majority7_module_21__or_module_5_res), .ZN(
        n_majority7_module_21__or_module_9_res) );
  OR2_X1 u_majority7_module_21__or_module_10_U1 ( .A1(
        n_majority7_module_21__or_module_7_res), .A2(
        n_majority7_module_21__and_module_7_res), .ZN(
        n_majority7_module_21__or_module_10_res) );
  AND2_X1 u_majority7_module_21__and_module_9_U1 ( .A1(
        n_majority7_module_21__or_module_6_res), .A2(
        n_majority7_module_21__or_module_9_res), .ZN(
        n_majority7_module_21__and_module_9_res) );
  OR2_X1 u_majority7_module_21__or_module_11_U1 ( .A1(
        n_majority7_module_21__or_module_10_res), .A2(
        n_majority7_module_21__and_module_8_res), .ZN(
        n_majority7_module_21__or_module_11_res) );
  AND2_X1 u_majority7_module_21__and_module_10_U1 ( .A1(
        n_majority7_module_21__or_module_8_res), .A2(
        n_majority7_module_21__and_module_9_res), .ZN(
        n_majority7_module_21__and_module_10_res) );
  AND2_X1 u_majority7_module_21__and_module_11_U1 ( .A1(
        n_majority7_module_21__and_module_10_res), .A2(
        n_majority7_module_21__or_module_11_res), .ZN(
        n_majority7_module_21_res) );
  DFF_X1 u_reg_module_22__cini_mul_v000_reg ( .D(n_majority7_module_21_res), 
        .CK(clock_2), .Q(n_reg_module_22_res), .QN() );
  BUF_X1 u_majority7_module_22_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_22_n7) );
  BUF_X1 u_majority7_module_22_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_22_n6) );
  BUF_X1 u_majority7_module_22_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_22_n5) );
  BUF_X1 u_majority7_module_22_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_22_n4) );
  BUF_X1 u_majority7_module_22_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_22_n3) );
  BUF_X1 u_majority7_module_22_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_22_n2) );
  BUF_X1 u_majority7_module_22_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_22_n1) );
  AND2_X1 u_majority7_module_22__and_module_1_U1 ( .A1(
        n_majority7_module_22_n5), .A2(n_majority7_module_22_n4), .ZN(
        n_majority7_module_22__and_module_1_res) );
  OR2_X1 u_majority7_module_22__or_module_1_U1 ( .A1(n_majority7_module_22_n4), 
        .A2(n_majority7_module_22_n5), .ZN(
        n_majority7_module_22__or_module_1_res) );
  AND2_X1 u_majority7_module_22__and_module_2_U1 ( .A1(
        n_majority7_module_22_n7), .A2(n_majority7_module_22_n2), .ZN(
        n_majority7_module_22__and_module_2_res) );
  OR2_X1 u_majority7_module_22__or_module_2_U1 ( .A1(n_majority7_module_22_n2), 
        .A2(n_majority7_module_22_n7), .ZN(
        n_majority7_module_22__or_module_2_res) );
  AND2_X1 u_majority7_module_22__and_module_3_U1 ( .A1(
        n_majority7_module_22_n6), .A2(n_majority7_module_22_n1), .ZN(
        n_majority7_module_22__and_module_3_res) );
  OR2_X1 u_majority7_module_22__or_module_3_U1 ( .A1(n_majority7_module_22_n1), 
        .A2(n_majority7_module_22_n6), .ZN(
        n_majority7_module_22__or_module_3_res) );
  AND2_X1 u_majority7_module_22__and_module_4_U1 ( .A1(
        n_majority7_module_22__and_module_2_res), .A2(
        n_majority7_module_22__and_module_1_res), .ZN(
        n_majority7_module_22__and_module_4_res) );
  OR2_X1 u_majority7_module_22__or_module_4_U1 ( .A1(
        n_majority7_module_22__and_module_1_res), .A2(
        n_majority7_module_22__and_module_2_res), .ZN(
        n_majority7_module_22__or_module_4_res) );
  AND2_X1 u_majority7_module_22__and_module_5_U1 ( .A1(
        n_majority7_module_22__and_module_3_res), .A2(n_majority7_module_22_n3), .ZN(n_majority7_module_22__and_module_5_res) );
  OR2_X1 u_majority7_module_22__or_module_5_U1 ( .A1(n_majority7_module_22_n3), 
        .A2(n_majority7_module_22__and_module_3_res), .ZN(
        n_majority7_module_22__or_module_5_res) );
  AND2_X1 u_majority7_module_22__and_module_6_U1 ( .A1(
        n_majority7_module_22__or_module_1_res), .A2(
        n_majority7_module_22__or_module_2_res), .ZN(
        n_majority7_module_22__and_module_6_res) );
  OR2_X1 u_majority7_module_22__or_module_6_U1 ( .A1(
        n_majority7_module_22__or_module_2_res), .A2(
        n_majority7_module_22__or_module_1_res), .ZN(
        n_majority7_module_22__or_module_6_res) );
  OR2_X1 u_majority7_module_22__or_module_7_U1 ( .A1(
        n_majority7_module_22__and_module_4_res), .A2(
        n_majority7_module_22__and_module_5_res), .ZN(
        n_majority7_module_22__or_module_7_res) );
  AND2_X1 u_majority7_module_22__and_module_7_U1 ( .A1(
        n_majority7_module_22__or_module_3_res), .A2(
        n_majority7_module_22__or_module_4_res), .ZN(
        n_majority7_module_22__and_module_7_res) );
  OR2_X1 u_majority7_module_22__or_module_8_U1 ( .A1(
        n_majority7_module_22__or_module_4_res), .A2(
        n_majority7_module_22__or_module_3_res), .ZN(
        n_majority7_module_22__or_module_8_res) );
  AND2_X1 u_majority7_module_22__and_module_8_U1 ( .A1(
        n_majority7_module_22__or_module_5_res), .A2(
        n_majority7_module_22__and_module_6_res), .ZN(
        n_majority7_module_22__and_module_8_res) );
  OR2_X1 u_majority7_module_22__or_module_9_U1 ( .A1(
        n_majority7_module_22__and_module_6_res), .A2(
        n_majority7_module_22__or_module_5_res), .ZN(
        n_majority7_module_22__or_module_9_res) );
  OR2_X1 u_majority7_module_22__or_module_10_U1 ( .A1(
        n_majority7_module_22__or_module_7_res), .A2(
        n_majority7_module_22__and_module_7_res), .ZN(
        n_majority7_module_22__or_module_10_res) );
  AND2_X1 u_majority7_module_22__and_module_9_U1 ( .A1(
        n_majority7_module_22__or_module_6_res), .A2(
        n_majority7_module_22__or_module_9_res), .ZN(
        n_majority7_module_22__and_module_9_res) );
  OR2_X1 u_majority7_module_22__or_module_11_U1 ( .A1(
        n_majority7_module_22__or_module_10_res), .A2(
        n_majority7_module_22__and_module_8_res), .ZN(
        n_majority7_module_22__or_module_11_res) );
  AND2_X1 u_majority7_module_22__and_module_10_U1 ( .A1(
        n_majority7_module_22__or_module_8_res), .A2(
        n_majority7_module_22__and_module_9_res), .ZN(
        n_majority7_module_22__and_module_10_res) );
  AND2_X1 u_majority7_module_22__and_module_11_U1 ( .A1(
        n_majority7_module_22__and_module_10_res), .A2(
        n_majority7_module_22__or_module_11_res), .ZN(
        n_majority7_module_22_res) );
  DFF_X1 u_reg_module_23__cini_mul_v000_reg ( .D(n_majority7_module_22_res), 
        .CK(clock_2), .Q(n_reg_module_23_res), .QN() );
  BUF_X1 u_majority7_module_23_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_23_n7) );
  BUF_X1 u_majority7_module_23_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_23_n6) );
  BUF_X1 u_majority7_module_23_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_23_n5) );
  BUF_X1 u_majority7_module_23_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_23_n4) );
  BUF_X1 u_majority7_module_23_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_23_n3) );
  BUF_X1 u_majority7_module_23_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_23_n2) );
  BUF_X1 u_majority7_module_23_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_23_n1) );
  AND2_X1 u_majority7_module_23__and_module_1_U1 ( .A1(
        n_majority7_module_23_n5), .A2(n_majority7_module_23_n4), .ZN(
        n_majority7_module_23__and_module_1_res) );
  OR2_X1 u_majority7_module_23__or_module_1_U1 ( .A1(n_majority7_module_23_n4), 
        .A2(n_majority7_module_23_n5), .ZN(
        n_majority7_module_23__or_module_1_res) );
  AND2_X1 u_majority7_module_23__and_module_2_U1 ( .A1(
        n_majority7_module_23_n7), .A2(n_majority7_module_23_n2), .ZN(
        n_majority7_module_23__and_module_2_res) );
  OR2_X1 u_majority7_module_23__or_module_2_U1 ( .A1(n_majority7_module_23_n2), 
        .A2(n_majority7_module_23_n7), .ZN(
        n_majority7_module_23__or_module_2_res) );
  AND2_X1 u_majority7_module_23__and_module_3_U1 ( .A1(
        n_majority7_module_23_n6), .A2(n_majority7_module_23_n1), .ZN(
        n_majority7_module_23__and_module_3_res) );
  OR2_X1 u_majority7_module_23__or_module_3_U1 ( .A1(n_majority7_module_23_n1), 
        .A2(n_majority7_module_23_n6), .ZN(
        n_majority7_module_23__or_module_3_res) );
  AND2_X1 u_majority7_module_23__and_module_4_U1 ( .A1(
        n_majority7_module_23__and_module_2_res), .A2(
        n_majority7_module_23__and_module_1_res), .ZN(
        n_majority7_module_23__and_module_4_res) );
  OR2_X1 u_majority7_module_23__or_module_4_U1 ( .A1(
        n_majority7_module_23__and_module_1_res), .A2(
        n_majority7_module_23__and_module_2_res), .ZN(
        n_majority7_module_23__or_module_4_res) );
  AND2_X1 u_majority7_module_23__and_module_5_U1 ( .A1(
        n_majority7_module_23__and_module_3_res), .A2(n_majority7_module_23_n3), .ZN(n_majority7_module_23__and_module_5_res) );
  OR2_X1 u_majority7_module_23__or_module_5_U1 ( .A1(n_majority7_module_23_n3), 
        .A2(n_majority7_module_23__and_module_3_res), .ZN(
        n_majority7_module_23__or_module_5_res) );
  AND2_X1 u_majority7_module_23__and_module_6_U1 ( .A1(
        n_majority7_module_23__or_module_1_res), .A2(
        n_majority7_module_23__or_module_2_res), .ZN(
        n_majority7_module_23__and_module_6_res) );
  OR2_X1 u_majority7_module_23__or_module_6_U1 ( .A1(
        n_majority7_module_23__or_module_2_res), .A2(
        n_majority7_module_23__or_module_1_res), .ZN(
        n_majority7_module_23__or_module_6_res) );
  OR2_X1 u_majority7_module_23__or_module_7_U1 ( .A1(
        n_majority7_module_23__and_module_4_res), .A2(
        n_majority7_module_23__and_module_5_res), .ZN(
        n_majority7_module_23__or_module_7_res) );
  AND2_X1 u_majority7_module_23__and_module_7_U1 ( .A1(
        n_majority7_module_23__or_module_3_res), .A2(
        n_majority7_module_23__or_module_4_res), .ZN(
        n_majority7_module_23__and_module_7_res) );
  OR2_X1 u_majority7_module_23__or_module_8_U1 ( .A1(
        n_majority7_module_23__or_module_4_res), .A2(
        n_majority7_module_23__or_module_3_res), .ZN(
        n_majority7_module_23__or_module_8_res) );
  AND2_X1 u_majority7_module_23__and_module_8_U1 ( .A1(
        n_majority7_module_23__or_module_5_res), .A2(
        n_majority7_module_23__and_module_6_res), .ZN(
        n_majority7_module_23__and_module_8_res) );
  OR2_X1 u_majority7_module_23__or_module_9_U1 ( .A1(
        n_majority7_module_23__and_module_6_res), .A2(
        n_majority7_module_23__or_module_5_res), .ZN(
        n_majority7_module_23__or_module_9_res) );
  OR2_X1 u_majority7_module_23__or_module_10_U1 ( .A1(
        n_majority7_module_23__or_module_7_res), .A2(
        n_majority7_module_23__and_module_7_res), .ZN(
        n_majority7_module_23__or_module_10_res) );
  AND2_X1 u_majority7_module_23__and_module_9_U1 ( .A1(
        n_majority7_module_23__or_module_6_res), .A2(
        n_majority7_module_23__or_module_9_res), .ZN(
        n_majority7_module_23__and_module_9_res) );
  OR2_X1 u_majority7_module_23__or_module_11_U1 ( .A1(
        n_majority7_module_23__or_module_10_res), .A2(
        n_majority7_module_23__and_module_8_res), .ZN(
        n_majority7_module_23__or_module_11_res) );
  AND2_X1 u_majority7_module_23__and_module_10_U1 ( .A1(
        n_majority7_module_23__or_module_8_res), .A2(
        n_majority7_module_23__and_module_9_res), .ZN(
        n_majority7_module_23__and_module_10_res) );
  AND2_X1 u_majority7_module_23__and_module_11_U1 ( .A1(
        n_majority7_module_23__and_module_10_res), .A2(
        n_majority7_module_23__or_module_11_res), .ZN(
        n_majority7_module_23_res) );
  DFF_X1 u_reg_module_24__cini_mul_v000_reg ( .D(n_majority7_module_23_res), 
        .CK(clock_2), .Q(n_reg_module_24_res), .QN() );
  BUF_X1 u_majority7_module_24_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_24_n7) );
  BUF_X1 u_majority7_module_24_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_24_n6) );
  BUF_X1 u_majority7_module_24_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_24_n5) );
  BUF_X1 u_majority7_module_24_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_24_n4) );
  BUF_X1 u_majority7_module_24_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_24_n3) );
  BUF_X1 u_majority7_module_24_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_24_n2) );
  BUF_X1 u_majority7_module_24_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_24_n1) );
  AND2_X1 u_majority7_module_24__and_module_1_U1 ( .A1(
        n_majority7_module_24_n5), .A2(n_majority7_module_24_n4), .ZN(
        n_majority7_module_24__and_module_1_res) );
  OR2_X1 u_majority7_module_24__or_module_1_U1 ( .A1(n_majority7_module_24_n4), 
        .A2(n_majority7_module_24_n5), .ZN(
        n_majority7_module_24__or_module_1_res) );
  AND2_X1 u_majority7_module_24__and_module_2_U1 ( .A1(
        n_majority7_module_24_n7), .A2(n_majority7_module_24_n2), .ZN(
        n_majority7_module_24__and_module_2_res) );
  OR2_X1 u_majority7_module_24__or_module_2_U1 ( .A1(n_majority7_module_24_n2), 
        .A2(n_majority7_module_24_n7), .ZN(
        n_majority7_module_24__or_module_2_res) );
  AND2_X1 u_majority7_module_24__and_module_3_U1 ( .A1(
        n_majority7_module_24_n6), .A2(n_majority7_module_24_n1), .ZN(
        n_majority7_module_24__and_module_3_res) );
  OR2_X1 u_majority7_module_24__or_module_3_U1 ( .A1(n_majority7_module_24_n1), 
        .A2(n_majority7_module_24_n6), .ZN(
        n_majority7_module_24__or_module_3_res) );
  AND2_X1 u_majority7_module_24__and_module_4_U1 ( .A1(
        n_majority7_module_24__and_module_2_res), .A2(
        n_majority7_module_24__and_module_1_res), .ZN(
        n_majority7_module_24__and_module_4_res) );
  OR2_X1 u_majority7_module_24__or_module_4_U1 ( .A1(
        n_majority7_module_24__and_module_1_res), .A2(
        n_majority7_module_24__and_module_2_res), .ZN(
        n_majority7_module_24__or_module_4_res) );
  AND2_X1 u_majority7_module_24__and_module_5_U1 ( .A1(
        n_majority7_module_24__and_module_3_res), .A2(n_majority7_module_24_n3), .ZN(n_majority7_module_24__and_module_5_res) );
  OR2_X1 u_majority7_module_24__or_module_5_U1 ( .A1(n_majority7_module_24_n3), 
        .A2(n_majority7_module_24__and_module_3_res), .ZN(
        n_majority7_module_24__or_module_5_res) );
  AND2_X1 u_majority7_module_24__and_module_6_U1 ( .A1(
        n_majority7_module_24__or_module_1_res), .A2(
        n_majority7_module_24__or_module_2_res), .ZN(
        n_majority7_module_24__and_module_6_res) );
  OR2_X1 u_majority7_module_24__or_module_6_U1 ( .A1(
        n_majority7_module_24__or_module_2_res), .A2(
        n_majority7_module_24__or_module_1_res), .ZN(
        n_majority7_module_24__or_module_6_res) );
  OR2_X1 u_majority7_module_24__or_module_7_U1 ( .A1(
        n_majority7_module_24__and_module_4_res), .A2(
        n_majority7_module_24__and_module_5_res), .ZN(
        n_majority7_module_24__or_module_7_res) );
  AND2_X1 u_majority7_module_24__and_module_7_U1 ( .A1(
        n_majority7_module_24__or_module_3_res), .A2(
        n_majority7_module_24__or_module_4_res), .ZN(
        n_majority7_module_24__and_module_7_res) );
  OR2_X1 u_majority7_module_24__or_module_8_U1 ( .A1(
        n_majority7_module_24__or_module_4_res), .A2(
        n_majority7_module_24__or_module_3_res), .ZN(
        n_majority7_module_24__or_module_8_res) );
  AND2_X1 u_majority7_module_24__and_module_8_U1 ( .A1(
        n_majority7_module_24__or_module_5_res), .A2(
        n_majority7_module_24__and_module_6_res), .ZN(
        n_majority7_module_24__and_module_8_res) );
  OR2_X1 u_majority7_module_24__or_module_9_U1 ( .A1(
        n_majority7_module_24__and_module_6_res), .A2(
        n_majority7_module_24__or_module_5_res), .ZN(
        n_majority7_module_24__or_module_9_res) );
  OR2_X1 u_majority7_module_24__or_module_10_U1 ( .A1(
        n_majority7_module_24__or_module_7_res), .A2(
        n_majority7_module_24__and_module_7_res), .ZN(
        n_majority7_module_24__or_module_10_res) );
  AND2_X1 u_majority7_module_24__and_module_9_U1 ( .A1(
        n_majority7_module_24__or_module_6_res), .A2(
        n_majority7_module_24__or_module_9_res), .ZN(
        n_majority7_module_24__and_module_9_res) );
  OR2_X1 u_majority7_module_24__or_module_11_U1 ( .A1(
        n_majority7_module_24__or_module_10_res), .A2(
        n_majority7_module_24__and_module_8_res), .ZN(
        n_majority7_module_24__or_module_11_res) );
  AND2_X1 u_majority7_module_24__and_module_10_U1 ( .A1(
        n_majority7_module_24__or_module_8_res), .A2(
        n_majority7_module_24__and_module_9_res), .ZN(
        n_majority7_module_24__and_module_10_res) );
  AND2_X1 u_majority7_module_24__and_module_11_U1 ( .A1(
        n_majority7_module_24__and_module_10_res), .A2(
        n_majority7_module_24__or_module_11_res), .ZN(
        n_majority7_module_24_res) );
  DFF_X1 u_reg_module_25__cini_mul_v000_reg ( .D(n_majority7_module_24_res), 
        .CK(clock_2), .Q(n_reg_module_25_res), .QN() );
  BUF_X1 u_majority7_module_25_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_25_n7) );
  BUF_X1 u_majority7_module_25_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_25_n6) );
  BUF_X1 u_majority7_module_25_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_25_n5) );
  BUF_X1 u_majority7_module_25_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_25_n4) );
  BUF_X1 u_majority7_module_25_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_25_n3) );
  BUF_X1 u_majority7_module_25_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_25_n2) );
  BUF_X1 u_majority7_module_25_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_25_n1) );
  AND2_X1 u_majority7_module_25__and_module_1_U1 ( .A1(
        n_majority7_module_25_n5), .A2(n_majority7_module_25_n4), .ZN(
        n_majority7_module_25__and_module_1_res) );
  OR2_X1 u_majority7_module_25__or_module_1_U1 ( .A1(n_majority7_module_25_n4), 
        .A2(n_majority7_module_25_n5), .ZN(
        n_majority7_module_25__or_module_1_res) );
  AND2_X1 u_majority7_module_25__and_module_2_U1 ( .A1(
        n_majority7_module_25_n7), .A2(n_majority7_module_25_n2), .ZN(
        n_majority7_module_25__and_module_2_res) );
  OR2_X1 u_majority7_module_25__or_module_2_U1 ( .A1(n_majority7_module_25_n2), 
        .A2(n_majority7_module_25_n7), .ZN(
        n_majority7_module_25__or_module_2_res) );
  AND2_X1 u_majority7_module_25__and_module_3_U1 ( .A1(
        n_majority7_module_25_n6), .A2(n_majority7_module_25_n1), .ZN(
        n_majority7_module_25__and_module_3_res) );
  OR2_X1 u_majority7_module_25__or_module_3_U1 ( .A1(n_majority7_module_25_n1), 
        .A2(n_majority7_module_25_n6), .ZN(
        n_majority7_module_25__or_module_3_res) );
  AND2_X1 u_majority7_module_25__and_module_4_U1 ( .A1(
        n_majority7_module_25__and_module_2_res), .A2(
        n_majority7_module_25__and_module_1_res), .ZN(
        n_majority7_module_25__and_module_4_res) );
  OR2_X1 u_majority7_module_25__or_module_4_U1 ( .A1(
        n_majority7_module_25__and_module_1_res), .A2(
        n_majority7_module_25__and_module_2_res), .ZN(
        n_majority7_module_25__or_module_4_res) );
  AND2_X1 u_majority7_module_25__and_module_5_U1 ( .A1(
        n_majority7_module_25__and_module_3_res), .A2(n_majority7_module_25_n3), .ZN(n_majority7_module_25__and_module_5_res) );
  OR2_X1 u_majority7_module_25__or_module_5_U1 ( .A1(n_majority7_module_25_n3), 
        .A2(n_majority7_module_25__and_module_3_res), .ZN(
        n_majority7_module_25__or_module_5_res) );
  AND2_X1 u_majority7_module_25__and_module_6_U1 ( .A1(
        n_majority7_module_25__or_module_1_res), .A2(
        n_majority7_module_25__or_module_2_res), .ZN(
        n_majority7_module_25__and_module_6_res) );
  OR2_X1 u_majority7_module_25__or_module_6_U1 ( .A1(
        n_majority7_module_25__or_module_2_res), .A2(
        n_majority7_module_25__or_module_1_res), .ZN(
        n_majority7_module_25__or_module_6_res) );
  OR2_X1 u_majority7_module_25__or_module_7_U1 ( .A1(
        n_majority7_module_25__and_module_4_res), .A2(
        n_majority7_module_25__and_module_5_res), .ZN(
        n_majority7_module_25__or_module_7_res) );
  AND2_X1 u_majority7_module_25__and_module_7_U1 ( .A1(
        n_majority7_module_25__or_module_3_res), .A2(
        n_majority7_module_25__or_module_4_res), .ZN(
        n_majority7_module_25__and_module_7_res) );
  OR2_X1 u_majority7_module_25__or_module_8_U1 ( .A1(
        n_majority7_module_25__or_module_4_res), .A2(
        n_majority7_module_25__or_module_3_res), .ZN(
        n_majority7_module_25__or_module_8_res) );
  AND2_X1 u_majority7_module_25__and_module_8_U1 ( .A1(
        n_majority7_module_25__or_module_5_res), .A2(
        n_majority7_module_25__and_module_6_res), .ZN(
        n_majority7_module_25__and_module_8_res) );
  OR2_X1 u_majority7_module_25__or_module_9_U1 ( .A1(
        n_majority7_module_25__and_module_6_res), .A2(
        n_majority7_module_25__or_module_5_res), .ZN(
        n_majority7_module_25__or_module_9_res) );
  OR2_X1 u_majority7_module_25__or_module_10_U1 ( .A1(
        n_majority7_module_25__or_module_7_res), .A2(
        n_majority7_module_25__and_module_7_res), .ZN(
        n_majority7_module_25__or_module_10_res) );
  AND2_X1 u_majority7_module_25__and_module_9_U1 ( .A1(
        n_majority7_module_25__or_module_6_res), .A2(
        n_majority7_module_25__or_module_9_res), .ZN(
        n_majority7_module_25__and_module_9_res) );
  OR2_X1 u_majority7_module_25__or_module_11_U1 ( .A1(
        n_majority7_module_25__or_module_10_res), .A2(
        n_majority7_module_25__and_module_8_res), .ZN(
        n_majority7_module_25__or_module_11_res) );
  AND2_X1 u_majority7_module_25__and_module_10_U1 ( .A1(
        n_majority7_module_25__or_module_8_res), .A2(
        n_majority7_module_25__and_module_9_res), .ZN(
        n_majority7_module_25__and_module_10_res) );
  AND2_X1 u_majority7_module_25__and_module_11_U1 ( .A1(
        n_majority7_module_25__and_module_10_res), .A2(
        n_majority7_module_25__or_module_11_res), .ZN(
        n_majority7_module_25_res) );
  DFF_X1 u_reg_module_26__cini_mul_v000_reg ( .D(n_majority7_module_25_res), 
        .CK(clock_2), .Q(n_reg_module_26_res), .QN() );
  BUF_X1 u_majority7_module_26_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_26_n7) );
  BUF_X1 u_majority7_module_26_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_26_n6) );
  BUF_X1 u_majority7_module_26_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_26_n5) );
  BUF_X1 u_majority7_module_26_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_26_n4) );
  BUF_X1 u_majority7_module_26_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_26_n3) );
  BUF_X1 u_majority7_module_26_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_26_n2) );
  BUF_X1 u_majority7_module_26_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_26_n1) );
  AND2_X1 u_majority7_module_26__and_module_1_U1 ( .A1(
        n_majority7_module_26_n5), .A2(n_majority7_module_26_n4), .ZN(
        n_majority7_module_26__and_module_1_res) );
  OR2_X1 u_majority7_module_26__or_module_1_U1 ( .A1(n_majority7_module_26_n4), 
        .A2(n_majority7_module_26_n5), .ZN(
        n_majority7_module_26__or_module_1_res) );
  AND2_X1 u_majority7_module_26__and_module_2_U1 ( .A1(
        n_majority7_module_26_n7), .A2(n_majority7_module_26_n2), .ZN(
        n_majority7_module_26__and_module_2_res) );
  OR2_X1 u_majority7_module_26__or_module_2_U1 ( .A1(n_majority7_module_26_n2), 
        .A2(n_majority7_module_26_n7), .ZN(
        n_majority7_module_26__or_module_2_res) );
  AND2_X1 u_majority7_module_26__and_module_3_U1 ( .A1(
        n_majority7_module_26_n6), .A2(n_majority7_module_26_n1), .ZN(
        n_majority7_module_26__and_module_3_res) );
  OR2_X1 u_majority7_module_26__or_module_3_U1 ( .A1(n_majority7_module_26_n1), 
        .A2(n_majority7_module_26_n6), .ZN(
        n_majority7_module_26__or_module_3_res) );
  AND2_X1 u_majority7_module_26__and_module_4_U1 ( .A1(
        n_majority7_module_26__and_module_2_res), .A2(
        n_majority7_module_26__and_module_1_res), .ZN(
        n_majority7_module_26__and_module_4_res) );
  OR2_X1 u_majority7_module_26__or_module_4_U1 ( .A1(
        n_majority7_module_26__and_module_1_res), .A2(
        n_majority7_module_26__and_module_2_res), .ZN(
        n_majority7_module_26__or_module_4_res) );
  AND2_X1 u_majority7_module_26__and_module_5_U1 ( .A1(
        n_majority7_module_26__and_module_3_res), .A2(n_majority7_module_26_n3), .ZN(n_majority7_module_26__and_module_5_res) );
  OR2_X1 u_majority7_module_26__or_module_5_U1 ( .A1(n_majority7_module_26_n3), 
        .A2(n_majority7_module_26__and_module_3_res), .ZN(
        n_majority7_module_26__or_module_5_res) );
  AND2_X1 u_majority7_module_26__and_module_6_U1 ( .A1(
        n_majority7_module_26__or_module_1_res), .A2(
        n_majority7_module_26__or_module_2_res), .ZN(
        n_majority7_module_26__and_module_6_res) );
  OR2_X1 u_majority7_module_26__or_module_6_U1 ( .A1(
        n_majority7_module_26__or_module_2_res), .A2(
        n_majority7_module_26__or_module_1_res), .ZN(
        n_majority7_module_26__or_module_6_res) );
  OR2_X1 u_majority7_module_26__or_module_7_U1 ( .A1(
        n_majority7_module_26__and_module_4_res), .A2(
        n_majority7_module_26__and_module_5_res), .ZN(
        n_majority7_module_26__or_module_7_res) );
  AND2_X1 u_majority7_module_26__and_module_7_U1 ( .A1(
        n_majority7_module_26__or_module_3_res), .A2(
        n_majority7_module_26__or_module_4_res), .ZN(
        n_majority7_module_26__and_module_7_res) );
  OR2_X1 u_majority7_module_26__or_module_8_U1 ( .A1(
        n_majority7_module_26__or_module_4_res), .A2(
        n_majority7_module_26__or_module_3_res), .ZN(
        n_majority7_module_26__or_module_8_res) );
  AND2_X1 u_majority7_module_26__and_module_8_U1 ( .A1(
        n_majority7_module_26__or_module_5_res), .A2(
        n_majority7_module_26__and_module_6_res), .ZN(
        n_majority7_module_26__and_module_8_res) );
  OR2_X1 u_majority7_module_26__or_module_9_U1 ( .A1(
        n_majority7_module_26__and_module_6_res), .A2(
        n_majority7_module_26__or_module_5_res), .ZN(
        n_majority7_module_26__or_module_9_res) );
  OR2_X1 u_majority7_module_26__or_module_10_U1 ( .A1(
        n_majority7_module_26__or_module_7_res), .A2(
        n_majority7_module_26__and_module_7_res), .ZN(
        n_majority7_module_26__or_module_10_res) );
  AND2_X1 u_majority7_module_26__and_module_9_U1 ( .A1(
        n_majority7_module_26__or_module_6_res), .A2(
        n_majority7_module_26__or_module_9_res), .ZN(
        n_majority7_module_26__and_module_9_res) );
  OR2_X1 u_majority7_module_26__or_module_11_U1 ( .A1(
        n_majority7_module_26__or_module_10_res), .A2(
        n_majority7_module_26__and_module_8_res), .ZN(
        n_majority7_module_26__or_module_11_res) );
  AND2_X1 u_majority7_module_26__and_module_10_U1 ( .A1(
        n_majority7_module_26__or_module_8_res), .A2(
        n_majority7_module_26__and_module_9_res), .ZN(
        n_majority7_module_26__and_module_10_res) );
  AND2_X1 u_majority7_module_26__and_module_11_U1 ( .A1(
        n_majority7_module_26__and_module_10_res), .A2(
        n_majority7_module_26__or_module_11_res), .ZN(
        n_majority7_module_26_res) );
  DFF_X1 u_reg_module_27__cini_mul_v000_reg ( .D(n_majority7_module_26_res), 
        .CK(clock_2), .Q(n_reg_module_27_res), .QN() );
  BUF_X1 u_majority7_module_27_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_27_n7) );
  BUF_X1 u_majority7_module_27_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_27_n6) );
  BUF_X1 u_majority7_module_27_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_27_n5) );
  BUF_X1 u_majority7_module_27_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_27_n4) );
  BUF_X1 u_majority7_module_27_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_27_n3) );
  BUF_X1 u_majority7_module_27_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_27_n2) );
  BUF_X1 u_majority7_module_27_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_27_n1) );
  AND2_X1 u_majority7_module_27__and_module_1_U1 ( .A1(
        n_majority7_module_27_n5), .A2(n_majority7_module_27_n4), .ZN(
        n_majority7_module_27__and_module_1_res) );
  OR2_X1 u_majority7_module_27__or_module_1_U1 ( .A1(n_majority7_module_27_n4), 
        .A2(n_majority7_module_27_n5), .ZN(
        n_majority7_module_27__or_module_1_res) );
  AND2_X1 u_majority7_module_27__and_module_2_U1 ( .A1(
        n_majority7_module_27_n7), .A2(n_majority7_module_27_n2), .ZN(
        n_majority7_module_27__and_module_2_res) );
  OR2_X1 u_majority7_module_27__or_module_2_U1 ( .A1(n_majority7_module_27_n2), 
        .A2(n_majority7_module_27_n7), .ZN(
        n_majority7_module_27__or_module_2_res) );
  AND2_X1 u_majority7_module_27__and_module_3_U1 ( .A1(
        n_majority7_module_27_n6), .A2(n_majority7_module_27_n1), .ZN(
        n_majority7_module_27__and_module_3_res) );
  OR2_X1 u_majority7_module_27__or_module_3_U1 ( .A1(n_majority7_module_27_n1), 
        .A2(n_majority7_module_27_n6), .ZN(
        n_majority7_module_27__or_module_3_res) );
  AND2_X1 u_majority7_module_27__and_module_4_U1 ( .A1(
        n_majority7_module_27__and_module_2_res), .A2(
        n_majority7_module_27__and_module_1_res), .ZN(
        n_majority7_module_27__and_module_4_res) );
  OR2_X1 u_majority7_module_27__or_module_4_U1 ( .A1(
        n_majority7_module_27__and_module_1_res), .A2(
        n_majority7_module_27__and_module_2_res), .ZN(
        n_majority7_module_27__or_module_4_res) );
  AND2_X1 u_majority7_module_27__and_module_5_U1 ( .A1(
        n_majority7_module_27__and_module_3_res), .A2(n_majority7_module_27_n3), .ZN(n_majority7_module_27__and_module_5_res) );
  OR2_X1 u_majority7_module_27__or_module_5_U1 ( .A1(n_majority7_module_27_n3), 
        .A2(n_majority7_module_27__and_module_3_res), .ZN(
        n_majority7_module_27__or_module_5_res) );
  AND2_X1 u_majority7_module_27__and_module_6_U1 ( .A1(
        n_majority7_module_27__or_module_1_res), .A2(
        n_majority7_module_27__or_module_2_res), .ZN(
        n_majority7_module_27__and_module_6_res) );
  OR2_X1 u_majority7_module_27__or_module_6_U1 ( .A1(
        n_majority7_module_27__or_module_2_res), .A2(
        n_majority7_module_27__or_module_1_res), .ZN(
        n_majority7_module_27__or_module_6_res) );
  OR2_X1 u_majority7_module_27__or_module_7_U1 ( .A1(
        n_majority7_module_27__and_module_4_res), .A2(
        n_majority7_module_27__and_module_5_res), .ZN(
        n_majority7_module_27__or_module_7_res) );
  AND2_X1 u_majority7_module_27__and_module_7_U1 ( .A1(
        n_majority7_module_27__or_module_3_res), .A2(
        n_majority7_module_27__or_module_4_res), .ZN(
        n_majority7_module_27__and_module_7_res) );
  OR2_X1 u_majority7_module_27__or_module_8_U1 ( .A1(
        n_majority7_module_27__or_module_4_res), .A2(
        n_majority7_module_27__or_module_3_res), .ZN(
        n_majority7_module_27__or_module_8_res) );
  AND2_X1 u_majority7_module_27__and_module_8_U1 ( .A1(
        n_majority7_module_27__or_module_5_res), .A2(
        n_majority7_module_27__and_module_6_res), .ZN(
        n_majority7_module_27__and_module_8_res) );
  OR2_X1 u_majority7_module_27__or_module_9_U1 ( .A1(
        n_majority7_module_27__and_module_6_res), .A2(
        n_majority7_module_27__or_module_5_res), .ZN(
        n_majority7_module_27__or_module_9_res) );
  OR2_X1 u_majority7_module_27__or_module_10_U1 ( .A1(
        n_majority7_module_27__or_module_7_res), .A2(
        n_majority7_module_27__and_module_7_res), .ZN(
        n_majority7_module_27__or_module_10_res) );
  AND2_X1 u_majority7_module_27__and_module_9_U1 ( .A1(
        n_majority7_module_27__or_module_6_res), .A2(
        n_majority7_module_27__or_module_9_res), .ZN(
        n_majority7_module_27__and_module_9_res) );
  OR2_X1 u_majority7_module_27__or_module_11_U1 ( .A1(
        n_majority7_module_27__or_module_10_res), .A2(
        n_majority7_module_27__and_module_8_res), .ZN(
        n_majority7_module_27__or_module_11_res) );
  AND2_X1 u_majority7_module_27__and_module_10_U1 ( .A1(
        n_majority7_module_27__or_module_8_res), .A2(
        n_majority7_module_27__and_module_9_res), .ZN(
        n_majority7_module_27__and_module_10_res) );
  AND2_X1 u_majority7_module_27__and_module_11_U1 ( .A1(
        n_majority7_module_27__and_module_10_res), .A2(
        n_majority7_module_27__or_module_11_res), .ZN(
        n_majority7_module_27_res) );
  DFF_X1 u_reg_module_28__cini_mul_v000_reg ( .D(n_majority7_module_27_res), 
        .CK(clock_3), .Q(n_reg_module_28_res), .QN() );
  BUF_X1 u_majority7_module_28_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_28_n7) );
  BUF_X1 u_majority7_module_28_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_28_n6) );
  BUF_X1 u_majority7_module_28_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_28_n5) );
  BUF_X1 u_majority7_module_28_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_28_n4) );
  BUF_X1 u_majority7_module_28_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_28_n3) );
  BUF_X1 u_majority7_module_28_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_28_n2) );
  BUF_X1 u_majority7_module_28_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_28_n1) );
  AND2_X1 u_majority7_module_28__and_module_1_U1 ( .A1(
        n_majority7_module_28_n5), .A2(n_majority7_module_28_n4), .ZN(
        n_majority7_module_28__and_module_1_res) );
  OR2_X1 u_majority7_module_28__or_module_1_U1 ( .A1(n_majority7_module_28_n4), 
        .A2(n_majority7_module_28_n5), .ZN(
        n_majority7_module_28__or_module_1_res) );
  AND2_X1 u_majority7_module_28__and_module_2_U1 ( .A1(
        n_majority7_module_28_n7), .A2(n_majority7_module_28_n2), .ZN(
        n_majority7_module_28__and_module_2_res) );
  OR2_X1 u_majority7_module_28__or_module_2_U1 ( .A1(n_majority7_module_28_n2), 
        .A2(n_majority7_module_28_n7), .ZN(
        n_majority7_module_28__or_module_2_res) );
  AND2_X1 u_majority7_module_28__and_module_3_U1 ( .A1(
        n_majority7_module_28_n6), .A2(n_majority7_module_28_n1), .ZN(
        n_majority7_module_28__and_module_3_res) );
  OR2_X1 u_majority7_module_28__or_module_3_U1 ( .A1(n_majority7_module_28_n1), 
        .A2(n_majority7_module_28_n6), .ZN(
        n_majority7_module_28__or_module_3_res) );
  AND2_X1 u_majority7_module_28__and_module_4_U1 ( .A1(
        n_majority7_module_28__and_module_2_res), .A2(
        n_majority7_module_28__and_module_1_res), .ZN(
        n_majority7_module_28__and_module_4_res) );
  OR2_X1 u_majority7_module_28__or_module_4_U1 ( .A1(
        n_majority7_module_28__and_module_1_res), .A2(
        n_majority7_module_28__and_module_2_res), .ZN(
        n_majority7_module_28__or_module_4_res) );
  AND2_X1 u_majority7_module_28__and_module_5_U1 ( .A1(
        n_majority7_module_28__and_module_3_res), .A2(n_majority7_module_28_n3), .ZN(n_majority7_module_28__and_module_5_res) );
  OR2_X1 u_majority7_module_28__or_module_5_U1 ( .A1(n_majority7_module_28_n3), 
        .A2(n_majority7_module_28__and_module_3_res), .ZN(
        n_majority7_module_28__or_module_5_res) );
  AND2_X1 u_majority7_module_28__and_module_6_U1 ( .A1(
        n_majority7_module_28__or_module_1_res), .A2(
        n_majority7_module_28__or_module_2_res), .ZN(
        n_majority7_module_28__and_module_6_res) );
  OR2_X1 u_majority7_module_28__or_module_6_U1 ( .A1(
        n_majority7_module_28__or_module_2_res), .A2(
        n_majority7_module_28__or_module_1_res), .ZN(
        n_majority7_module_28__or_module_6_res) );
  OR2_X1 u_majority7_module_28__or_module_7_U1 ( .A1(
        n_majority7_module_28__and_module_4_res), .A2(
        n_majority7_module_28__and_module_5_res), .ZN(
        n_majority7_module_28__or_module_7_res) );
  AND2_X1 u_majority7_module_28__and_module_7_U1 ( .A1(
        n_majority7_module_28__or_module_3_res), .A2(
        n_majority7_module_28__or_module_4_res), .ZN(
        n_majority7_module_28__and_module_7_res) );
  OR2_X1 u_majority7_module_28__or_module_8_U1 ( .A1(
        n_majority7_module_28__or_module_4_res), .A2(
        n_majority7_module_28__or_module_3_res), .ZN(
        n_majority7_module_28__or_module_8_res) );
  AND2_X1 u_majority7_module_28__and_module_8_U1 ( .A1(
        n_majority7_module_28__or_module_5_res), .A2(
        n_majority7_module_28__and_module_6_res), .ZN(
        n_majority7_module_28__and_module_8_res) );
  OR2_X1 u_majority7_module_28__or_module_9_U1 ( .A1(
        n_majority7_module_28__and_module_6_res), .A2(
        n_majority7_module_28__or_module_5_res), .ZN(
        n_majority7_module_28__or_module_9_res) );
  OR2_X1 u_majority7_module_28__or_module_10_U1 ( .A1(
        n_majority7_module_28__or_module_7_res), .A2(
        n_majority7_module_28__and_module_7_res), .ZN(
        n_majority7_module_28__or_module_10_res) );
  AND2_X1 u_majority7_module_28__and_module_9_U1 ( .A1(
        n_majority7_module_28__or_module_6_res), .A2(
        n_majority7_module_28__or_module_9_res), .ZN(
        n_majority7_module_28__and_module_9_res) );
  OR2_X1 u_majority7_module_28__or_module_11_U1 ( .A1(
        n_majority7_module_28__or_module_10_res), .A2(
        n_majority7_module_28__and_module_8_res), .ZN(
        n_majority7_module_28__or_module_11_res) );
  AND2_X1 u_majority7_module_28__and_module_10_U1 ( .A1(
        n_majority7_module_28__or_module_8_res), .A2(
        n_majority7_module_28__and_module_9_res), .ZN(
        n_majority7_module_28__and_module_10_res) );
  AND2_X1 u_majority7_module_28__and_module_11_U1 ( .A1(
        n_majority7_module_28__and_module_10_res), .A2(
        n_majority7_module_28__or_module_11_res), .ZN(
        n_majority7_module_28_res) );
  DFF_X1 u_reg_module_29__cini_mul_v000_reg ( .D(n_majority7_module_28_res), 
        .CK(clock_3), .Q(n_reg_module_29_res), .QN() );
  BUF_X1 u_majority7_module_29_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_29_n7) );
  BUF_X1 u_majority7_module_29_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_29_n6) );
  BUF_X1 u_majority7_module_29_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_29_n5) );
  BUF_X1 u_majority7_module_29_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_29_n4) );
  BUF_X1 u_majority7_module_29_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_29_n3) );
  BUF_X1 u_majority7_module_29_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_29_n2) );
  BUF_X1 u_majority7_module_29_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_29_n1) );
  AND2_X1 u_majority7_module_29__and_module_1_U1 ( .A1(
        n_majority7_module_29_n5), .A2(n_majority7_module_29_n4), .ZN(
        n_majority7_module_29__and_module_1_res) );
  OR2_X1 u_majority7_module_29__or_module_1_U1 ( .A1(n_majority7_module_29_n4), 
        .A2(n_majority7_module_29_n5), .ZN(
        n_majority7_module_29__or_module_1_res) );
  AND2_X1 u_majority7_module_29__and_module_2_U1 ( .A1(
        n_majority7_module_29_n7), .A2(n_majority7_module_29_n2), .ZN(
        n_majority7_module_29__and_module_2_res) );
  OR2_X1 u_majority7_module_29__or_module_2_U1 ( .A1(n_majority7_module_29_n2), 
        .A2(n_majority7_module_29_n7), .ZN(
        n_majority7_module_29__or_module_2_res) );
  AND2_X1 u_majority7_module_29__and_module_3_U1 ( .A1(
        n_majority7_module_29_n6), .A2(n_majority7_module_29_n1), .ZN(
        n_majority7_module_29__and_module_3_res) );
  OR2_X1 u_majority7_module_29__or_module_3_U1 ( .A1(n_majority7_module_29_n1), 
        .A2(n_majority7_module_29_n6), .ZN(
        n_majority7_module_29__or_module_3_res) );
  AND2_X1 u_majority7_module_29__and_module_4_U1 ( .A1(
        n_majority7_module_29__and_module_2_res), .A2(
        n_majority7_module_29__and_module_1_res), .ZN(
        n_majority7_module_29__and_module_4_res) );
  OR2_X1 u_majority7_module_29__or_module_4_U1 ( .A1(
        n_majority7_module_29__and_module_1_res), .A2(
        n_majority7_module_29__and_module_2_res), .ZN(
        n_majority7_module_29__or_module_4_res) );
  AND2_X1 u_majority7_module_29__and_module_5_U1 ( .A1(
        n_majority7_module_29__and_module_3_res), .A2(n_majority7_module_29_n3), .ZN(n_majority7_module_29__and_module_5_res) );
  OR2_X1 u_majority7_module_29__or_module_5_U1 ( .A1(n_majority7_module_29_n3), 
        .A2(n_majority7_module_29__and_module_3_res), .ZN(
        n_majority7_module_29__or_module_5_res) );
  AND2_X1 u_majority7_module_29__and_module_6_U1 ( .A1(
        n_majority7_module_29__or_module_1_res), .A2(
        n_majority7_module_29__or_module_2_res), .ZN(
        n_majority7_module_29__and_module_6_res) );
  OR2_X1 u_majority7_module_29__or_module_6_U1 ( .A1(
        n_majority7_module_29__or_module_2_res), .A2(
        n_majority7_module_29__or_module_1_res), .ZN(
        n_majority7_module_29__or_module_6_res) );
  OR2_X1 u_majority7_module_29__or_module_7_U1 ( .A1(
        n_majority7_module_29__and_module_4_res), .A2(
        n_majority7_module_29__and_module_5_res), .ZN(
        n_majority7_module_29__or_module_7_res) );
  AND2_X1 u_majority7_module_29__and_module_7_U1 ( .A1(
        n_majority7_module_29__or_module_3_res), .A2(
        n_majority7_module_29__or_module_4_res), .ZN(
        n_majority7_module_29__and_module_7_res) );
  OR2_X1 u_majority7_module_29__or_module_8_U1 ( .A1(
        n_majority7_module_29__or_module_4_res), .A2(
        n_majority7_module_29__or_module_3_res), .ZN(
        n_majority7_module_29__or_module_8_res) );
  AND2_X1 u_majority7_module_29__and_module_8_U1 ( .A1(
        n_majority7_module_29__or_module_5_res), .A2(
        n_majority7_module_29__and_module_6_res), .ZN(
        n_majority7_module_29__and_module_8_res) );
  OR2_X1 u_majority7_module_29__or_module_9_U1 ( .A1(
        n_majority7_module_29__and_module_6_res), .A2(
        n_majority7_module_29__or_module_5_res), .ZN(
        n_majority7_module_29__or_module_9_res) );
  OR2_X1 u_majority7_module_29__or_module_10_U1 ( .A1(
        n_majority7_module_29__or_module_7_res), .A2(
        n_majority7_module_29__and_module_7_res), .ZN(
        n_majority7_module_29__or_module_10_res) );
  AND2_X1 u_majority7_module_29__and_module_9_U1 ( .A1(
        n_majority7_module_29__or_module_6_res), .A2(
        n_majority7_module_29__or_module_9_res), .ZN(
        n_majority7_module_29__and_module_9_res) );
  OR2_X1 u_majority7_module_29__or_module_11_U1 ( .A1(
        n_majority7_module_29__or_module_10_res), .A2(
        n_majority7_module_29__and_module_8_res), .ZN(
        n_majority7_module_29__or_module_11_res) );
  AND2_X1 u_majority7_module_29__and_module_10_U1 ( .A1(
        n_majority7_module_29__or_module_8_res), .A2(
        n_majority7_module_29__and_module_9_res), .ZN(
        n_majority7_module_29__and_module_10_res) );
  AND2_X1 u_majority7_module_29__and_module_11_U1 ( .A1(
        n_majority7_module_29__and_module_10_res), .A2(
        n_majority7_module_29__or_module_11_res), .ZN(
        n_majority7_module_29_res) );
  DFF_X1 u_reg_module_30__cini_mul_v000_reg ( .D(n_majority7_module_29_res), 
        .CK(clock_3), .Q(n_reg_module_30_res), .QN() );
  BUF_X1 u_majority7_module_30_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_30_n7) );
  BUF_X1 u_majority7_module_30_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_30_n6) );
  BUF_X1 u_majority7_module_30_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_30_n5) );
  BUF_X1 u_majority7_module_30_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_30_n4) );
  BUF_X1 u_majority7_module_30_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_30_n3) );
  BUF_X1 u_majority7_module_30_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_30_n2) );
  BUF_X1 u_majority7_module_30_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_30_n1) );
  AND2_X1 u_majority7_module_30__and_module_1_U1 ( .A1(
        n_majority7_module_30_n5), .A2(n_majority7_module_30_n4), .ZN(
        n_majority7_module_30__and_module_1_res) );
  OR2_X1 u_majority7_module_30__or_module_1_U1 ( .A1(n_majority7_module_30_n4), 
        .A2(n_majority7_module_30_n5), .ZN(
        n_majority7_module_30__or_module_1_res) );
  AND2_X1 u_majority7_module_30__and_module_2_U1 ( .A1(
        n_majority7_module_30_n7), .A2(n_majority7_module_30_n2), .ZN(
        n_majority7_module_30__and_module_2_res) );
  OR2_X1 u_majority7_module_30__or_module_2_U1 ( .A1(n_majority7_module_30_n2), 
        .A2(n_majority7_module_30_n7), .ZN(
        n_majority7_module_30__or_module_2_res) );
  AND2_X1 u_majority7_module_30__and_module_3_U1 ( .A1(
        n_majority7_module_30_n6), .A2(n_majority7_module_30_n1), .ZN(
        n_majority7_module_30__and_module_3_res) );
  OR2_X1 u_majority7_module_30__or_module_3_U1 ( .A1(n_majority7_module_30_n1), 
        .A2(n_majority7_module_30_n6), .ZN(
        n_majority7_module_30__or_module_3_res) );
  AND2_X1 u_majority7_module_30__and_module_4_U1 ( .A1(
        n_majority7_module_30__and_module_2_res), .A2(
        n_majority7_module_30__and_module_1_res), .ZN(
        n_majority7_module_30__and_module_4_res) );
  OR2_X1 u_majority7_module_30__or_module_4_U1 ( .A1(
        n_majority7_module_30__and_module_1_res), .A2(
        n_majority7_module_30__and_module_2_res), .ZN(
        n_majority7_module_30__or_module_4_res) );
  AND2_X1 u_majority7_module_30__and_module_5_U1 ( .A1(
        n_majority7_module_30__and_module_3_res), .A2(n_majority7_module_30_n3), .ZN(n_majority7_module_30__and_module_5_res) );
  OR2_X1 u_majority7_module_30__or_module_5_U1 ( .A1(n_majority7_module_30_n3), 
        .A2(n_majority7_module_30__and_module_3_res), .ZN(
        n_majority7_module_30__or_module_5_res) );
  AND2_X1 u_majority7_module_30__and_module_6_U1 ( .A1(
        n_majority7_module_30__or_module_1_res), .A2(
        n_majority7_module_30__or_module_2_res), .ZN(
        n_majority7_module_30__and_module_6_res) );
  OR2_X1 u_majority7_module_30__or_module_6_U1 ( .A1(
        n_majority7_module_30__or_module_2_res), .A2(
        n_majority7_module_30__or_module_1_res), .ZN(
        n_majority7_module_30__or_module_6_res) );
  OR2_X1 u_majority7_module_30__or_module_7_U1 ( .A1(
        n_majority7_module_30__and_module_4_res), .A2(
        n_majority7_module_30__and_module_5_res), .ZN(
        n_majority7_module_30__or_module_7_res) );
  AND2_X1 u_majority7_module_30__and_module_7_U1 ( .A1(
        n_majority7_module_30__or_module_3_res), .A2(
        n_majority7_module_30__or_module_4_res), .ZN(
        n_majority7_module_30__and_module_7_res) );
  OR2_X1 u_majority7_module_30__or_module_8_U1 ( .A1(
        n_majority7_module_30__or_module_4_res), .A2(
        n_majority7_module_30__or_module_3_res), .ZN(
        n_majority7_module_30__or_module_8_res) );
  AND2_X1 u_majority7_module_30__and_module_8_U1 ( .A1(
        n_majority7_module_30__or_module_5_res), .A2(
        n_majority7_module_30__and_module_6_res), .ZN(
        n_majority7_module_30__and_module_8_res) );
  OR2_X1 u_majority7_module_30__or_module_9_U1 ( .A1(
        n_majority7_module_30__and_module_6_res), .A2(
        n_majority7_module_30__or_module_5_res), .ZN(
        n_majority7_module_30__or_module_9_res) );
  OR2_X1 u_majority7_module_30__or_module_10_U1 ( .A1(
        n_majority7_module_30__or_module_7_res), .A2(
        n_majority7_module_30__and_module_7_res), .ZN(
        n_majority7_module_30__or_module_10_res) );
  AND2_X1 u_majority7_module_30__and_module_9_U1 ( .A1(
        n_majority7_module_30__or_module_6_res), .A2(
        n_majority7_module_30__or_module_9_res), .ZN(
        n_majority7_module_30__and_module_9_res) );
  OR2_X1 u_majority7_module_30__or_module_11_U1 ( .A1(
        n_majority7_module_30__or_module_10_res), .A2(
        n_majority7_module_30__and_module_8_res), .ZN(
        n_majority7_module_30__or_module_11_res) );
  AND2_X1 u_majority7_module_30__and_module_10_U1 ( .A1(
        n_majority7_module_30__or_module_8_res), .A2(
        n_majority7_module_30__and_module_9_res), .ZN(
        n_majority7_module_30__and_module_10_res) );
  AND2_X1 u_majority7_module_30__and_module_11_U1 ( .A1(
        n_majority7_module_30__and_module_10_res), .A2(
        n_majority7_module_30__or_module_11_res), .ZN(
        n_majority7_module_30_res) );
  DFF_X1 u_reg_module_31__cini_mul_v000_reg ( .D(n_majority7_module_30_res), 
        .CK(clock_3), .Q(n_reg_module_31_res), .QN() );
  BUF_X1 u_majority7_module_31_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_31_n7) );
  BUF_X1 u_majority7_module_31_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_31_n6) );
  BUF_X1 u_majority7_module_31_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_31_n5) );
  BUF_X1 u_majority7_module_31_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_31_n4) );
  BUF_X1 u_majority7_module_31_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_31_n3) );
  BUF_X1 u_majority7_module_31_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_31_n2) );
  BUF_X1 u_majority7_module_31_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_31_n1) );
  AND2_X1 u_majority7_module_31__and_module_1_U1 ( .A1(
        n_majority7_module_31_n5), .A2(n_majority7_module_31_n4), .ZN(
        n_majority7_module_31__and_module_1_res) );
  OR2_X1 u_majority7_module_31__or_module_1_U1 ( .A1(n_majority7_module_31_n4), 
        .A2(n_majority7_module_31_n5), .ZN(
        n_majority7_module_31__or_module_1_res) );
  AND2_X1 u_majority7_module_31__and_module_2_U1 ( .A1(
        n_majority7_module_31_n7), .A2(n_majority7_module_31_n2), .ZN(
        n_majority7_module_31__and_module_2_res) );
  OR2_X1 u_majority7_module_31__or_module_2_U1 ( .A1(n_majority7_module_31_n2), 
        .A2(n_majority7_module_31_n7), .ZN(
        n_majority7_module_31__or_module_2_res) );
  AND2_X1 u_majority7_module_31__and_module_3_U1 ( .A1(
        n_majority7_module_31_n6), .A2(n_majority7_module_31_n1), .ZN(
        n_majority7_module_31__and_module_3_res) );
  OR2_X1 u_majority7_module_31__or_module_3_U1 ( .A1(n_majority7_module_31_n1), 
        .A2(n_majority7_module_31_n6), .ZN(
        n_majority7_module_31__or_module_3_res) );
  AND2_X1 u_majority7_module_31__and_module_4_U1 ( .A1(
        n_majority7_module_31__and_module_2_res), .A2(
        n_majority7_module_31__and_module_1_res), .ZN(
        n_majority7_module_31__and_module_4_res) );
  OR2_X1 u_majority7_module_31__or_module_4_U1 ( .A1(
        n_majority7_module_31__and_module_1_res), .A2(
        n_majority7_module_31__and_module_2_res), .ZN(
        n_majority7_module_31__or_module_4_res) );
  AND2_X1 u_majority7_module_31__and_module_5_U1 ( .A1(
        n_majority7_module_31__and_module_3_res), .A2(n_majority7_module_31_n3), .ZN(n_majority7_module_31__and_module_5_res) );
  OR2_X1 u_majority7_module_31__or_module_5_U1 ( .A1(n_majority7_module_31_n3), 
        .A2(n_majority7_module_31__and_module_3_res), .ZN(
        n_majority7_module_31__or_module_5_res) );
  AND2_X1 u_majority7_module_31__and_module_6_U1 ( .A1(
        n_majority7_module_31__or_module_1_res), .A2(
        n_majority7_module_31__or_module_2_res), .ZN(
        n_majority7_module_31__and_module_6_res) );
  OR2_X1 u_majority7_module_31__or_module_6_U1 ( .A1(
        n_majority7_module_31__or_module_2_res), .A2(
        n_majority7_module_31__or_module_1_res), .ZN(
        n_majority7_module_31__or_module_6_res) );
  OR2_X1 u_majority7_module_31__or_module_7_U1 ( .A1(
        n_majority7_module_31__and_module_4_res), .A2(
        n_majority7_module_31__and_module_5_res), .ZN(
        n_majority7_module_31__or_module_7_res) );
  AND2_X1 u_majority7_module_31__and_module_7_U1 ( .A1(
        n_majority7_module_31__or_module_3_res), .A2(
        n_majority7_module_31__or_module_4_res), .ZN(
        n_majority7_module_31__and_module_7_res) );
  OR2_X1 u_majority7_module_31__or_module_8_U1 ( .A1(
        n_majority7_module_31__or_module_4_res), .A2(
        n_majority7_module_31__or_module_3_res), .ZN(
        n_majority7_module_31__or_module_8_res) );
  AND2_X1 u_majority7_module_31__and_module_8_U1 ( .A1(
        n_majority7_module_31__or_module_5_res), .A2(
        n_majority7_module_31__and_module_6_res), .ZN(
        n_majority7_module_31__and_module_8_res) );
  OR2_X1 u_majority7_module_31__or_module_9_U1 ( .A1(
        n_majority7_module_31__and_module_6_res), .A2(
        n_majority7_module_31__or_module_5_res), .ZN(
        n_majority7_module_31__or_module_9_res) );
  OR2_X1 u_majority7_module_31__or_module_10_U1 ( .A1(
        n_majority7_module_31__or_module_7_res), .A2(
        n_majority7_module_31__and_module_7_res), .ZN(
        n_majority7_module_31__or_module_10_res) );
  AND2_X1 u_majority7_module_31__and_module_9_U1 ( .A1(
        n_majority7_module_31__or_module_6_res), .A2(
        n_majority7_module_31__or_module_9_res), .ZN(
        n_majority7_module_31__and_module_9_res) );
  OR2_X1 u_majority7_module_31__or_module_11_U1 ( .A1(
        n_majority7_module_31__or_module_10_res), .A2(
        n_majority7_module_31__and_module_8_res), .ZN(
        n_majority7_module_31__or_module_11_res) );
  AND2_X1 u_majority7_module_31__and_module_10_U1 ( .A1(
        n_majority7_module_31__or_module_8_res), .A2(
        n_majority7_module_31__and_module_9_res), .ZN(
        n_majority7_module_31__and_module_10_res) );
  AND2_X1 u_majority7_module_31__and_module_11_U1 ( .A1(
        n_majority7_module_31__and_module_10_res), .A2(
        n_majority7_module_31__or_module_11_res), .ZN(
        n_majority7_module_31_res) );
  DFF_X1 u_reg_module_32__cini_mul_v000_reg ( .D(n_majority7_module_31_res), 
        .CK(clock_3), .Q(n_reg_module_32_res), .QN() );
  BUF_X1 u_majority7_module_32_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_32_n7) );
  BUF_X1 u_majority7_module_32_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_32_n6) );
  BUF_X1 u_majority7_module_32_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_32_n5) );
  BUF_X1 u_majority7_module_32_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_32_n4) );
  BUF_X1 u_majority7_module_32_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_32_n3) );
  BUF_X1 u_majority7_module_32_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_32_n2) );
  BUF_X1 u_majority7_module_32_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_32_n1) );
  AND2_X1 u_majority7_module_32__and_module_1_U1 ( .A1(
        n_majority7_module_32_n5), .A2(n_majority7_module_32_n4), .ZN(
        n_majority7_module_32__and_module_1_res) );
  OR2_X1 u_majority7_module_32__or_module_1_U1 ( .A1(n_majority7_module_32_n4), 
        .A2(n_majority7_module_32_n5), .ZN(
        n_majority7_module_32__or_module_1_res) );
  AND2_X1 u_majority7_module_32__and_module_2_U1 ( .A1(
        n_majority7_module_32_n7), .A2(n_majority7_module_32_n2), .ZN(
        n_majority7_module_32__and_module_2_res) );
  OR2_X1 u_majority7_module_32__or_module_2_U1 ( .A1(n_majority7_module_32_n2), 
        .A2(n_majority7_module_32_n7), .ZN(
        n_majority7_module_32__or_module_2_res) );
  AND2_X1 u_majority7_module_32__and_module_3_U1 ( .A1(
        n_majority7_module_32_n6), .A2(n_majority7_module_32_n1), .ZN(
        n_majority7_module_32__and_module_3_res) );
  OR2_X1 u_majority7_module_32__or_module_3_U1 ( .A1(n_majority7_module_32_n1), 
        .A2(n_majority7_module_32_n6), .ZN(
        n_majority7_module_32__or_module_3_res) );
  AND2_X1 u_majority7_module_32__and_module_4_U1 ( .A1(
        n_majority7_module_32__and_module_2_res), .A2(
        n_majority7_module_32__and_module_1_res), .ZN(
        n_majority7_module_32__and_module_4_res) );
  OR2_X1 u_majority7_module_32__or_module_4_U1 ( .A1(
        n_majority7_module_32__and_module_1_res), .A2(
        n_majority7_module_32__and_module_2_res), .ZN(
        n_majority7_module_32__or_module_4_res) );
  AND2_X1 u_majority7_module_32__and_module_5_U1 ( .A1(
        n_majority7_module_32__and_module_3_res), .A2(n_majority7_module_32_n3), .ZN(n_majority7_module_32__and_module_5_res) );
  OR2_X1 u_majority7_module_32__or_module_5_U1 ( .A1(n_majority7_module_32_n3), 
        .A2(n_majority7_module_32__and_module_3_res), .ZN(
        n_majority7_module_32__or_module_5_res) );
  AND2_X1 u_majority7_module_32__and_module_6_U1 ( .A1(
        n_majority7_module_32__or_module_1_res), .A2(
        n_majority7_module_32__or_module_2_res), .ZN(
        n_majority7_module_32__and_module_6_res) );
  OR2_X1 u_majority7_module_32__or_module_6_U1 ( .A1(
        n_majority7_module_32__or_module_2_res), .A2(
        n_majority7_module_32__or_module_1_res), .ZN(
        n_majority7_module_32__or_module_6_res) );
  OR2_X1 u_majority7_module_32__or_module_7_U1 ( .A1(
        n_majority7_module_32__and_module_4_res), .A2(
        n_majority7_module_32__and_module_5_res), .ZN(
        n_majority7_module_32__or_module_7_res) );
  AND2_X1 u_majority7_module_32__and_module_7_U1 ( .A1(
        n_majority7_module_32__or_module_3_res), .A2(
        n_majority7_module_32__or_module_4_res), .ZN(
        n_majority7_module_32__and_module_7_res) );
  OR2_X1 u_majority7_module_32__or_module_8_U1 ( .A1(
        n_majority7_module_32__or_module_4_res), .A2(
        n_majority7_module_32__or_module_3_res), .ZN(
        n_majority7_module_32__or_module_8_res) );
  AND2_X1 u_majority7_module_32__and_module_8_U1 ( .A1(
        n_majority7_module_32__or_module_5_res), .A2(
        n_majority7_module_32__and_module_6_res), .ZN(
        n_majority7_module_32__and_module_8_res) );
  OR2_X1 u_majority7_module_32__or_module_9_U1 ( .A1(
        n_majority7_module_32__and_module_6_res), .A2(
        n_majority7_module_32__or_module_5_res), .ZN(
        n_majority7_module_32__or_module_9_res) );
  OR2_X1 u_majority7_module_32__or_module_10_U1 ( .A1(
        n_majority7_module_32__or_module_7_res), .A2(
        n_majority7_module_32__and_module_7_res), .ZN(
        n_majority7_module_32__or_module_10_res) );
  AND2_X1 u_majority7_module_32__and_module_9_U1 ( .A1(
        n_majority7_module_32__or_module_6_res), .A2(
        n_majority7_module_32__or_module_9_res), .ZN(
        n_majority7_module_32__and_module_9_res) );
  OR2_X1 u_majority7_module_32__or_module_11_U1 ( .A1(
        n_majority7_module_32__or_module_10_res), .A2(
        n_majority7_module_32__and_module_8_res), .ZN(
        n_majority7_module_32__or_module_11_res) );
  AND2_X1 u_majority7_module_32__and_module_10_U1 ( .A1(
        n_majority7_module_32__or_module_8_res), .A2(
        n_majority7_module_32__and_module_9_res), .ZN(
        n_majority7_module_32__and_module_10_res) );
  AND2_X1 u_majority7_module_32__and_module_11_U1 ( .A1(
        n_majority7_module_32__and_module_10_res), .A2(
        n_majority7_module_32__or_module_11_res), .ZN(
        n_majority7_module_32_res) );
  DFF_X1 u_reg_module_33__cini_mul_v000_reg ( .D(n_majority7_module_32_res), 
        .CK(clock_3), .Q(n_reg_module_33_res), .QN() );
  BUF_X1 u_majority7_module_33_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_33_n7) );
  BUF_X1 u_majority7_module_33_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_33_n6) );
  BUF_X1 u_majority7_module_33_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_33_n5) );
  BUF_X1 u_majority7_module_33_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_33_n4) );
  BUF_X1 u_majority7_module_33_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_33_n3) );
  BUF_X1 u_majority7_module_33_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_33_n2) );
  BUF_X1 u_majority7_module_33_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_33_n1) );
  AND2_X1 u_majority7_module_33__and_module_1_U1 ( .A1(
        n_majority7_module_33_n5), .A2(n_majority7_module_33_n4), .ZN(
        n_majority7_module_33__and_module_1_res) );
  OR2_X1 u_majority7_module_33__or_module_1_U1 ( .A1(n_majority7_module_33_n4), 
        .A2(n_majority7_module_33_n5), .ZN(
        n_majority7_module_33__or_module_1_res) );
  AND2_X1 u_majority7_module_33__and_module_2_U1 ( .A1(
        n_majority7_module_33_n7), .A2(n_majority7_module_33_n2), .ZN(
        n_majority7_module_33__and_module_2_res) );
  OR2_X1 u_majority7_module_33__or_module_2_U1 ( .A1(n_majority7_module_33_n2), 
        .A2(n_majority7_module_33_n7), .ZN(
        n_majority7_module_33__or_module_2_res) );
  AND2_X1 u_majority7_module_33__and_module_3_U1 ( .A1(
        n_majority7_module_33_n6), .A2(n_majority7_module_33_n1), .ZN(
        n_majority7_module_33__and_module_3_res) );
  OR2_X1 u_majority7_module_33__or_module_3_U1 ( .A1(n_majority7_module_33_n1), 
        .A2(n_majority7_module_33_n6), .ZN(
        n_majority7_module_33__or_module_3_res) );
  AND2_X1 u_majority7_module_33__and_module_4_U1 ( .A1(
        n_majority7_module_33__and_module_2_res), .A2(
        n_majority7_module_33__and_module_1_res), .ZN(
        n_majority7_module_33__and_module_4_res) );
  OR2_X1 u_majority7_module_33__or_module_4_U1 ( .A1(
        n_majority7_module_33__and_module_1_res), .A2(
        n_majority7_module_33__and_module_2_res), .ZN(
        n_majority7_module_33__or_module_4_res) );
  AND2_X1 u_majority7_module_33__and_module_5_U1 ( .A1(
        n_majority7_module_33__and_module_3_res), .A2(n_majority7_module_33_n3), .ZN(n_majority7_module_33__and_module_5_res) );
  OR2_X1 u_majority7_module_33__or_module_5_U1 ( .A1(n_majority7_module_33_n3), 
        .A2(n_majority7_module_33__and_module_3_res), .ZN(
        n_majority7_module_33__or_module_5_res) );
  AND2_X1 u_majority7_module_33__and_module_6_U1 ( .A1(
        n_majority7_module_33__or_module_1_res), .A2(
        n_majority7_module_33__or_module_2_res), .ZN(
        n_majority7_module_33__and_module_6_res) );
  OR2_X1 u_majority7_module_33__or_module_6_U1 ( .A1(
        n_majority7_module_33__or_module_2_res), .A2(
        n_majority7_module_33__or_module_1_res), .ZN(
        n_majority7_module_33__or_module_6_res) );
  OR2_X1 u_majority7_module_33__or_module_7_U1 ( .A1(
        n_majority7_module_33__and_module_4_res), .A2(
        n_majority7_module_33__and_module_5_res), .ZN(
        n_majority7_module_33__or_module_7_res) );
  AND2_X1 u_majority7_module_33__and_module_7_U1 ( .A1(
        n_majority7_module_33__or_module_3_res), .A2(
        n_majority7_module_33__or_module_4_res), .ZN(
        n_majority7_module_33__and_module_7_res) );
  OR2_X1 u_majority7_module_33__or_module_8_U1 ( .A1(
        n_majority7_module_33__or_module_4_res), .A2(
        n_majority7_module_33__or_module_3_res), .ZN(
        n_majority7_module_33__or_module_8_res) );
  AND2_X1 u_majority7_module_33__and_module_8_U1 ( .A1(
        n_majority7_module_33__or_module_5_res), .A2(
        n_majority7_module_33__and_module_6_res), .ZN(
        n_majority7_module_33__and_module_8_res) );
  OR2_X1 u_majority7_module_33__or_module_9_U1 ( .A1(
        n_majority7_module_33__and_module_6_res), .A2(
        n_majority7_module_33__or_module_5_res), .ZN(
        n_majority7_module_33__or_module_9_res) );
  OR2_X1 u_majority7_module_33__or_module_10_U1 ( .A1(
        n_majority7_module_33__or_module_7_res), .A2(
        n_majority7_module_33__and_module_7_res), .ZN(
        n_majority7_module_33__or_module_10_res) );
  AND2_X1 u_majority7_module_33__and_module_9_U1 ( .A1(
        n_majority7_module_33__or_module_6_res), .A2(
        n_majority7_module_33__or_module_9_res), .ZN(
        n_majority7_module_33__and_module_9_res) );
  OR2_X1 u_majority7_module_33__or_module_11_U1 ( .A1(
        n_majority7_module_33__or_module_10_res), .A2(
        n_majority7_module_33__and_module_8_res), .ZN(
        n_majority7_module_33__or_module_11_res) );
  AND2_X1 u_majority7_module_33__and_module_10_U1 ( .A1(
        n_majority7_module_33__or_module_8_res), .A2(
        n_majority7_module_33__and_module_9_res), .ZN(
        n_majority7_module_33__and_module_10_res) );
  AND2_X1 u_majority7_module_33__and_module_11_U1 ( .A1(
        n_majority7_module_33__and_module_10_res), .A2(
        n_majority7_module_33__or_module_11_res), .ZN(
        n_majority7_module_33_res) );
  DFF_X1 u_reg_module_34__cini_mul_v000_reg ( .D(n_majority7_module_33_res), 
        .CK(clock_3), .Q(n_reg_module_34_res), .QN() );
  BUF_X1 u_majority7_module_34_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_34_n7) );
  BUF_X1 u_majority7_module_34_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_34_n6) );
  BUF_X1 u_majority7_module_34_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_34_n5) );
  BUF_X1 u_majority7_module_34_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_34_n4) );
  BUF_X1 u_majority7_module_34_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_34_n3) );
  BUF_X1 u_majority7_module_34_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_34_n2) );
  BUF_X1 u_majority7_module_34_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_34_n1) );
  AND2_X1 u_majority7_module_34__and_module_1_U1 ( .A1(
        n_majority7_module_34_n5), .A2(n_majority7_module_34_n4), .ZN(
        n_majority7_module_34__and_module_1_res) );
  OR2_X1 u_majority7_module_34__or_module_1_U1 ( .A1(n_majority7_module_34_n4), 
        .A2(n_majority7_module_34_n5), .ZN(
        n_majority7_module_34__or_module_1_res) );
  AND2_X1 u_majority7_module_34__and_module_2_U1 ( .A1(
        n_majority7_module_34_n7), .A2(n_majority7_module_34_n2), .ZN(
        n_majority7_module_34__and_module_2_res) );
  OR2_X1 u_majority7_module_34__or_module_2_U1 ( .A1(n_majority7_module_34_n2), 
        .A2(n_majority7_module_34_n7), .ZN(
        n_majority7_module_34__or_module_2_res) );
  AND2_X1 u_majority7_module_34__and_module_3_U1 ( .A1(
        n_majority7_module_34_n6), .A2(n_majority7_module_34_n1), .ZN(
        n_majority7_module_34__and_module_3_res) );
  OR2_X1 u_majority7_module_34__or_module_3_U1 ( .A1(n_majority7_module_34_n1), 
        .A2(n_majority7_module_34_n6), .ZN(
        n_majority7_module_34__or_module_3_res) );
  AND2_X1 u_majority7_module_34__and_module_4_U1 ( .A1(
        n_majority7_module_34__and_module_2_res), .A2(
        n_majority7_module_34__and_module_1_res), .ZN(
        n_majority7_module_34__and_module_4_res) );
  OR2_X1 u_majority7_module_34__or_module_4_U1 ( .A1(
        n_majority7_module_34__and_module_1_res), .A2(
        n_majority7_module_34__and_module_2_res), .ZN(
        n_majority7_module_34__or_module_4_res) );
  AND2_X1 u_majority7_module_34__and_module_5_U1 ( .A1(
        n_majority7_module_34__and_module_3_res), .A2(n_majority7_module_34_n3), .ZN(n_majority7_module_34__and_module_5_res) );
  OR2_X1 u_majority7_module_34__or_module_5_U1 ( .A1(n_majority7_module_34_n3), 
        .A2(n_majority7_module_34__and_module_3_res), .ZN(
        n_majority7_module_34__or_module_5_res) );
  AND2_X1 u_majority7_module_34__and_module_6_U1 ( .A1(
        n_majority7_module_34__or_module_1_res), .A2(
        n_majority7_module_34__or_module_2_res), .ZN(
        n_majority7_module_34__and_module_6_res) );
  OR2_X1 u_majority7_module_34__or_module_6_U1 ( .A1(
        n_majority7_module_34__or_module_2_res), .A2(
        n_majority7_module_34__or_module_1_res), .ZN(
        n_majority7_module_34__or_module_6_res) );
  OR2_X1 u_majority7_module_34__or_module_7_U1 ( .A1(
        n_majority7_module_34__and_module_4_res), .A2(
        n_majority7_module_34__and_module_5_res), .ZN(
        n_majority7_module_34__or_module_7_res) );
  AND2_X1 u_majority7_module_34__and_module_7_U1 ( .A1(
        n_majority7_module_34__or_module_3_res), .A2(
        n_majority7_module_34__or_module_4_res), .ZN(
        n_majority7_module_34__and_module_7_res) );
  OR2_X1 u_majority7_module_34__or_module_8_U1 ( .A1(
        n_majority7_module_34__or_module_4_res), .A2(
        n_majority7_module_34__or_module_3_res), .ZN(
        n_majority7_module_34__or_module_8_res) );
  AND2_X1 u_majority7_module_34__and_module_8_U1 ( .A1(
        n_majority7_module_34__or_module_5_res), .A2(
        n_majority7_module_34__and_module_6_res), .ZN(
        n_majority7_module_34__and_module_8_res) );
  OR2_X1 u_majority7_module_34__or_module_9_U1 ( .A1(
        n_majority7_module_34__and_module_6_res), .A2(
        n_majority7_module_34__or_module_5_res), .ZN(
        n_majority7_module_34__or_module_9_res) );
  OR2_X1 u_majority7_module_34__or_module_10_U1 ( .A1(
        n_majority7_module_34__or_module_7_res), .A2(
        n_majority7_module_34__and_module_7_res), .ZN(
        n_majority7_module_34__or_module_10_res) );
  AND2_X1 u_majority7_module_34__and_module_9_U1 ( .A1(
        n_majority7_module_34__or_module_6_res), .A2(
        n_majority7_module_34__or_module_9_res), .ZN(
        n_majority7_module_34__and_module_9_res) );
  OR2_X1 u_majority7_module_34__or_module_11_U1 ( .A1(
        n_majority7_module_34__or_module_10_res), .A2(
        n_majority7_module_34__and_module_8_res), .ZN(
        n_majority7_module_34__or_module_11_res) );
  AND2_X1 u_majority7_module_34__and_module_10_U1 ( .A1(
        n_majority7_module_34__or_module_8_res), .A2(
        n_majority7_module_34__and_module_9_res), .ZN(
        n_majority7_module_34__and_module_10_res) );
  AND2_X1 u_majority7_module_34__and_module_11_U1 ( .A1(
        n_majority7_module_34__and_module_10_res), .A2(
        n_majority7_module_34__or_module_11_res), .ZN(
        n_majority7_module_34_res) );
  DFF_X1 u_reg_module_35__cini_mul_v000_reg ( .D(n_majority7_module_34_res), 
        .CK(clock_3), .Q(n_reg_module_35_res), .QN() );
  BUF_X1 u_majority7_module_35_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_35_n7) );
  BUF_X1 u_majority7_module_35_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_35_n6) );
  BUF_X1 u_majority7_module_35_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_35_n5) );
  BUF_X1 u_majority7_module_35_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_35_n4) );
  BUF_X1 u_majority7_module_35_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_35_n3) );
  BUF_X1 u_majority7_module_35_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_35_n2) );
  BUF_X1 u_majority7_module_35_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_35_n1) );
  AND2_X1 u_majority7_module_35__and_module_1_U1 ( .A1(
        n_majority7_module_35_n5), .A2(n_majority7_module_35_n4), .ZN(
        n_majority7_module_35__and_module_1_res) );
  OR2_X1 u_majority7_module_35__or_module_1_U1 ( .A1(n_majority7_module_35_n4), 
        .A2(n_majority7_module_35_n5), .ZN(
        n_majority7_module_35__or_module_1_res) );
  AND2_X1 u_majority7_module_35__and_module_2_U1 ( .A1(
        n_majority7_module_35_n7), .A2(n_majority7_module_35_n2), .ZN(
        n_majority7_module_35__and_module_2_res) );
  OR2_X1 u_majority7_module_35__or_module_2_U1 ( .A1(n_majority7_module_35_n2), 
        .A2(n_majority7_module_35_n7), .ZN(
        n_majority7_module_35__or_module_2_res) );
  AND2_X1 u_majority7_module_35__and_module_3_U1 ( .A1(
        n_majority7_module_35_n6), .A2(n_majority7_module_35_n1), .ZN(
        n_majority7_module_35__and_module_3_res) );
  OR2_X1 u_majority7_module_35__or_module_3_U1 ( .A1(n_majority7_module_35_n1), 
        .A2(n_majority7_module_35_n6), .ZN(
        n_majority7_module_35__or_module_3_res) );
  AND2_X1 u_majority7_module_35__and_module_4_U1 ( .A1(
        n_majority7_module_35__and_module_2_res), .A2(
        n_majority7_module_35__and_module_1_res), .ZN(
        n_majority7_module_35__and_module_4_res) );
  OR2_X1 u_majority7_module_35__or_module_4_U1 ( .A1(
        n_majority7_module_35__and_module_1_res), .A2(
        n_majority7_module_35__and_module_2_res), .ZN(
        n_majority7_module_35__or_module_4_res) );
  AND2_X1 u_majority7_module_35__and_module_5_U1 ( .A1(
        n_majority7_module_35__and_module_3_res), .A2(n_majority7_module_35_n3), .ZN(n_majority7_module_35__and_module_5_res) );
  OR2_X1 u_majority7_module_35__or_module_5_U1 ( .A1(n_majority7_module_35_n3), 
        .A2(n_majority7_module_35__and_module_3_res), .ZN(
        n_majority7_module_35__or_module_5_res) );
  AND2_X1 u_majority7_module_35__and_module_6_U1 ( .A1(
        n_majority7_module_35__or_module_1_res), .A2(
        n_majority7_module_35__or_module_2_res), .ZN(
        n_majority7_module_35__and_module_6_res) );
  OR2_X1 u_majority7_module_35__or_module_6_U1 ( .A1(
        n_majority7_module_35__or_module_2_res), .A2(
        n_majority7_module_35__or_module_1_res), .ZN(
        n_majority7_module_35__or_module_6_res) );
  OR2_X1 u_majority7_module_35__or_module_7_U1 ( .A1(
        n_majority7_module_35__and_module_4_res), .A2(
        n_majority7_module_35__and_module_5_res), .ZN(
        n_majority7_module_35__or_module_7_res) );
  AND2_X1 u_majority7_module_35__and_module_7_U1 ( .A1(
        n_majority7_module_35__or_module_3_res), .A2(
        n_majority7_module_35__or_module_4_res), .ZN(
        n_majority7_module_35__and_module_7_res) );
  OR2_X1 u_majority7_module_35__or_module_8_U1 ( .A1(
        n_majority7_module_35__or_module_4_res), .A2(
        n_majority7_module_35__or_module_3_res), .ZN(
        n_majority7_module_35__or_module_8_res) );
  AND2_X1 u_majority7_module_35__and_module_8_U1 ( .A1(
        n_majority7_module_35__or_module_5_res), .A2(
        n_majority7_module_35__and_module_6_res), .ZN(
        n_majority7_module_35__and_module_8_res) );
  OR2_X1 u_majority7_module_35__or_module_9_U1 ( .A1(
        n_majority7_module_35__and_module_6_res), .A2(
        n_majority7_module_35__or_module_5_res), .ZN(
        n_majority7_module_35__or_module_9_res) );
  OR2_X1 u_majority7_module_35__or_module_10_U1 ( .A1(
        n_majority7_module_35__or_module_7_res), .A2(
        n_majority7_module_35__and_module_7_res), .ZN(
        n_majority7_module_35__or_module_10_res) );
  AND2_X1 u_majority7_module_35__and_module_9_U1 ( .A1(
        n_majority7_module_35__or_module_6_res), .A2(
        n_majority7_module_35__or_module_9_res), .ZN(
        n_majority7_module_35__and_module_9_res) );
  OR2_X1 u_majority7_module_35__or_module_11_U1 ( .A1(
        n_majority7_module_35__or_module_10_res), .A2(
        n_majority7_module_35__and_module_8_res), .ZN(
        n_majority7_module_35__or_module_11_res) );
  AND2_X1 u_majority7_module_35__and_module_10_U1 ( .A1(
        n_majority7_module_35__or_module_8_res), .A2(
        n_majority7_module_35__and_module_9_res), .ZN(
        n_majority7_module_35__and_module_10_res) );
  AND2_X1 u_majority7_module_35__and_module_11_U1 ( .A1(
        n_majority7_module_35__and_module_10_res), .A2(
        n_majority7_module_35__or_module_11_res), .ZN(
        n_majority7_module_35_res) );
  DFF_X1 u_reg_module_36__cini_mul_v000_reg ( .D(n_majority7_module_35_res), 
        .CK(clock_3), .Q(n_reg_module_36_res), .QN() );
  BUF_X1 u_majority7_module_36_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_36_n7) );
  BUF_X1 u_majority7_module_36_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_36_n6) );
  BUF_X1 u_majority7_module_36_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_36_n5) );
  BUF_X1 u_majority7_module_36_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_36_n4) );
  BUF_X1 u_majority7_module_36_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_36_n3) );
  BUF_X1 u_majority7_module_36_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_36_n2) );
  BUF_X1 u_majority7_module_36_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_36_n1) );
  AND2_X1 u_majority7_module_36__and_module_1_U1 ( .A1(
        n_majority7_module_36_n5), .A2(n_majority7_module_36_n4), .ZN(
        n_majority7_module_36__and_module_1_res) );
  OR2_X1 u_majority7_module_36__or_module_1_U1 ( .A1(n_majority7_module_36_n4), 
        .A2(n_majority7_module_36_n5), .ZN(
        n_majority7_module_36__or_module_1_res) );
  AND2_X1 u_majority7_module_36__and_module_2_U1 ( .A1(
        n_majority7_module_36_n7), .A2(n_majority7_module_36_n2), .ZN(
        n_majority7_module_36__and_module_2_res) );
  OR2_X1 u_majority7_module_36__or_module_2_U1 ( .A1(n_majority7_module_36_n2), 
        .A2(n_majority7_module_36_n7), .ZN(
        n_majority7_module_36__or_module_2_res) );
  AND2_X1 u_majority7_module_36__and_module_3_U1 ( .A1(
        n_majority7_module_36_n6), .A2(n_majority7_module_36_n1), .ZN(
        n_majority7_module_36__and_module_3_res) );
  OR2_X1 u_majority7_module_36__or_module_3_U1 ( .A1(n_majority7_module_36_n1), 
        .A2(n_majority7_module_36_n6), .ZN(
        n_majority7_module_36__or_module_3_res) );
  AND2_X1 u_majority7_module_36__and_module_4_U1 ( .A1(
        n_majority7_module_36__and_module_2_res), .A2(
        n_majority7_module_36__and_module_1_res), .ZN(
        n_majority7_module_36__and_module_4_res) );
  OR2_X1 u_majority7_module_36__or_module_4_U1 ( .A1(
        n_majority7_module_36__and_module_1_res), .A2(
        n_majority7_module_36__and_module_2_res), .ZN(
        n_majority7_module_36__or_module_4_res) );
  AND2_X1 u_majority7_module_36__and_module_5_U1 ( .A1(
        n_majority7_module_36__and_module_3_res), .A2(n_majority7_module_36_n3), .ZN(n_majority7_module_36__and_module_5_res) );
  OR2_X1 u_majority7_module_36__or_module_5_U1 ( .A1(n_majority7_module_36_n3), 
        .A2(n_majority7_module_36__and_module_3_res), .ZN(
        n_majority7_module_36__or_module_5_res) );
  AND2_X1 u_majority7_module_36__and_module_6_U1 ( .A1(
        n_majority7_module_36__or_module_1_res), .A2(
        n_majority7_module_36__or_module_2_res), .ZN(
        n_majority7_module_36__and_module_6_res) );
  OR2_X1 u_majority7_module_36__or_module_6_U1 ( .A1(
        n_majority7_module_36__or_module_2_res), .A2(
        n_majority7_module_36__or_module_1_res), .ZN(
        n_majority7_module_36__or_module_6_res) );
  OR2_X1 u_majority7_module_36__or_module_7_U1 ( .A1(
        n_majority7_module_36__and_module_4_res), .A2(
        n_majority7_module_36__and_module_5_res), .ZN(
        n_majority7_module_36__or_module_7_res) );
  AND2_X1 u_majority7_module_36__and_module_7_U1 ( .A1(
        n_majority7_module_36__or_module_3_res), .A2(
        n_majority7_module_36__or_module_4_res), .ZN(
        n_majority7_module_36__and_module_7_res) );
  OR2_X1 u_majority7_module_36__or_module_8_U1 ( .A1(
        n_majority7_module_36__or_module_4_res), .A2(
        n_majority7_module_36__or_module_3_res), .ZN(
        n_majority7_module_36__or_module_8_res) );
  AND2_X1 u_majority7_module_36__and_module_8_U1 ( .A1(
        n_majority7_module_36__or_module_5_res), .A2(
        n_majority7_module_36__and_module_6_res), .ZN(
        n_majority7_module_36__and_module_8_res) );
  OR2_X1 u_majority7_module_36__or_module_9_U1 ( .A1(
        n_majority7_module_36__and_module_6_res), .A2(
        n_majority7_module_36__or_module_5_res), .ZN(
        n_majority7_module_36__or_module_9_res) );
  OR2_X1 u_majority7_module_36__or_module_10_U1 ( .A1(
        n_majority7_module_36__or_module_7_res), .A2(
        n_majority7_module_36__and_module_7_res), .ZN(
        n_majority7_module_36__or_module_10_res) );
  AND2_X1 u_majority7_module_36__and_module_9_U1 ( .A1(
        n_majority7_module_36__or_module_6_res), .A2(
        n_majority7_module_36__or_module_9_res), .ZN(
        n_majority7_module_36__and_module_9_res) );
  OR2_X1 u_majority7_module_36__or_module_11_U1 ( .A1(
        n_majority7_module_36__or_module_10_res), .A2(
        n_majority7_module_36__and_module_8_res), .ZN(
        n_majority7_module_36__or_module_11_res) );
  AND2_X1 u_majority7_module_36__and_module_10_U1 ( .A1(
        n_majority7_module_36__or_module_8_res), .A2(
        n_majority7_module_36__and_module_9_res), .ZN(
        n_majority7_module_36__and_module_10_res) );
  AND2_X1 u_majority7_module_36__and_module_11_U1 ( .A1(
        n_majority7_module_36__and_module_10_res), .A2(
        n_majority7_module_36__or_module_11_res), .ZN(
        n_majority7_module_36_res) );
  DFF_X1 u_reg_module_37__cini_mul_v000_reg ( .D(n_majority7_module_36_res), 
        .CK(clock_4), .Q(n_reg_module_37_res), .QN() );
  BUF_X1 u_majority7_module_37_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_37_n7) );
  BUF_X1 u_majority7_module_37_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_37_n6) );
  BUF_X1 u_majority7_module_37_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_37_n5) );
  BUF_X1 u_majority7_module_37_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_37_n4) );
  BUF_X1 u_majority7_module_37_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_37_n3) );
  BUF_X1 u_majority7_module_37_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_37_n2) );
  BUF_X1 u_majority7_module_37_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_37_n1) );
  AND2_X1 u_majority7_module_37__and_module_1_U1 ( .A1(
        n_majority7_module_37_n5), .A2(n_majority7_module_37_n4), .ZN(
        n_majority7_module_37__and_module_1_res) );
  OR2_X1 u_majority7_module_37__or_module_1_U1 ( .A1(n_majority7_module_37_n4), 
        .A2(n_majority7_module_37_n5), .ZN(
        n_majority7_module_37__or_module_1_res) );
  AND2_X1 u_majority7_module_37__and_module_2_U1 ( .A1(
        n_majority7_module_37_n7), .A2(n_majority7_module_37_n2), .ZN(
        n_majority7_module_37__and_module_2_res) );
  OR2_X1 u_majority7_module_37__or_module_2_U1 ( .A1(n_majority7_module_37_n2), 
        .A2(n_majority7_module_37_n7), .ZN(
        n_majority7_module_37__or_module_2_res) );
  AND2_X1 u_majority7_module_37__and_module_3_U1 ( .A1(
        n_majority7_module_37_n6), .A2(n_majority7_module_37_n1), .ZN(
        n_majority7_module_37__and_module_3_res) );
  OR2_X1 u_majority7_module_37__or_module_3_U1 ( .A1(n_majority7_module_37_n1), 
        .A2(n_majority7_module_37_n6), .ZN(
        n_majority7_module_37__or_module_3_res) );
  AND2_X1 u_majority7_module_37__and_module_4_U1 ( .A1(
        n_majority7_module_37__and_module_2_res), .A2(
        n_majority7_module_37__and_module_1_res), .ZN(
        n_majority7_module_37__and_module_4_res) );
  OR2_X1 u_majority7_module_37__or_module_4_U1 ( .A1(
        n_majority7_module_37__and_module_1_res), .A2(
        n_majority7_module_37__and_module_2_res), .ZN(
        n_majority7_module_37__or_module_4_res) );
  AND2_X1 u_majority7_module_37__and_module_5_U1 ( .A1(
        n_majority7_module_37__and_module_3_res), .A2(n_majority7_module_37_n3), .ZN(n_majority7_module_37__and_module_5_res) );
  OR2_X1 u_majority7_module_37__or_module_5_U1 ( .A1(n_majority7_module_37_n3), 
        .A2(n_majority7_module_37__and_module_3_res), .ZN(
        n_majority7_module_37__or_module_5_res) );
  AND2_X1 u_majority7_module_37__and_module_6_U1 ( .A1(
        n_majority7_module_37__or_module_1_res), .A2(
        n_majority7_module_37__or_module_2_res), .ZN(
        n_majority7_module_37__and_module_6_res) );
  OR2_X1 u_majority7_module_37__or_module_6_U1 ( .A1(
        n_majority7_module_37__or_module_2_res), .A2(
        n_majority7_module_37__or_module_1_res), .ZN(
        n_majority7_module_37__or_module_6_res) );
  OR2_X1 u_majority7_module_37__or_module_7_U1 ( .A1(
        n_majority7_module_37__and_module_4_res), .A2(
        n_majority7_module_37__and_module_5_res), .ZN(
        n_majority7_module_37__or_module_7_res) );
  AND2_X1 u_majority7_module_37__and_module_7_U1 ( .A1(
        n_majority7_module_37__or_module_3_res), .A2(
        n_majority7_module_37__or_module_4_res), .ZN(
        n_majority7_module_37__and_module_7_res) );
  OR2_X1 u_majority7_module_37__or_module_8_U1 ( .A1(
        n_majority7_module_37__or_module_4_res), .A2(
        n_majority7_module_37__or_module_3_res), .ZN(
        n_majority7_module_37__or_module_8_res) );
  AND2_X1 u_majority7_module_37__and_module_8_U1 ( .A1(
        n_majority7_module_37__or_module_5_res), .A2(
        n_majority7_module_37__and_module_6_res), .ZN(
        n_majority7_module_37__and_module_8_res) );
  OR2_X1 u_majority7_module_37__or_module_9_U1 ( .A1(
        n_majority7_module_37__and_module_6_res), .A2(
        n_majority7_module_37__or_module_5_res), .ZN(
        n_majority7_module_37__or_module_9_res) );
  OR2_X1 u_majority7_module_37__or_module_10_U1 ( .A1(
        n_majority7_module_37__or_module_7_res), .A2(
        n_majority7_module_37__and_module_7_res), .ZN(
        n_majority7_module_37__or_module_10_res) );
  AND2_X1 u_majority7_module_37__and_module_9_U1 ( .A1(
        n_majority7_module_37__or_module_6_res), .A2(
        n_majority7_module_37__or_module_9_res), .ZN(
        n_majority7_module_37__and_module_9_res) );
  OR2_X1 u_majority7_module_37__or_module_11_U1 ( .A1(
        n_majority7_module_37__or_module_10_res), .A2(
        n_majority7_module_37__and_module_8_res), .ZN(
        n_majority7_module_37__or_module_11_res) );
  AND2_X1 u_majority7_module_37__and_module_10_U1 ( .A1(
        n_majority7_module_37__or_module_8_res), .A2(
        n_majority7_module_37__and_module_9_res), .ZN(
        n_majority7_module_37__and_module_10_res) );
  AND2_X1 u_majority7_module_37__and_module_11_U1 ( .A1(
        n_majority7_module_37__and_module_10_res), .A2(
        n_majority7_module_37__or_module_11_res), .ZN(
        n_majority7_module_37_res) );
  DFF_X1 u_reg_module_38__cini_mul_v000_reg ( .D(n_majority7_module_37_res), 
        .CK(clock_4), .Q(n_reg_module_38_res), .QN() );
  BUF_X1 u_majority7_module_38_U7 ( .A(n_xor_module_20_res), .Z(
        n_majority7_module_38_n7) );
  BUF_X1 u_majority7_module_38_U6 ( .A(n_xor_module_32_res), .Z(
        n_majority7_module_38_n6) );
  BUF_X1 u_majority7_module_38_U5 ( .A(n_xor_module_38_res), .Z(
        n_majority7_module_38_n5) );
  BUF_X1 u_majority7_module_38_U4 ( .A(n_xor_module_2_res), .Z(
        n_majority7_module_38_n4) );
  BUF_X1 u_majority7_module_38_U3 ( .A(n_xor_module_8_res), .Z(
        n_majority7_module_38_n3) );
  BUF_X1 u_majority7_module_38_U2 ( .A(n_xor_module_14_res), .Z(
        n_majority7_module_38_n2) );
  BUF_X1 u_majority7_module_38_U1 ( .A(n_xor_module_26_res), .Z(
        n_majority7_module_38_n1) );
  AND2_X1 u_majority7_module_38__and_module_1_U1 ( .A1(
        n_majority7_module_38_n5), .A2(n_majority7_module_38_n4), .ZN(
        n_majority7_module_38__and_module_1_res) );
  OR2_X1 u_majority7_module_38__or_module_1_U1 ( .A1(n_majority7_module_38_n4), 
        .A2(n_majority7_module_38_n5), .ZN(
        n_majority7_module_38__or_module_1_res) );
  AND2_X1 u_majority7_module_38__and_module_2_U1 ( .A1(
        n_majority7_module_38_n7), .A2(n_majority7_module_38_n2), .ZN(
        n_majority7_module_38__and_module_2_res) );
  OR2_X1 u_majority7_module_38__or_module_2_U1 ( .A1(n_majority7_module_38_n2), 
        .A2(n_majority7_module_38_n7), .ZN(
        n_majority7_module_38__or_module_2_res) );
  AND2_X1 u_majority7_module_38__and_module_3_U1 ( .A1(
        n_majority7_module_38_n6), .A2(n_majority7_module_38_n1), .ZN(
        n_majority7_module_38__and_module_3_res) );
  OR2_X1 u_majority7_module_38__or_module_3_U1 ( .A1(n_majority7_module_38_n1), 
        .A2(n_majority7_module_38_n6), .ZN(
        n_majority7_module_38__or_module_3_res) );
  AND2_X1 u_majority7_module_38__and_module_4_U1 ( .A1(
        n_majority7_module_38__and_module_2_res), .A2(
        n_majority7_module_38__and_module_1_res), .ZN(
        n_majority7_module_38__and_module_4_res) );
  OR2_X1 u_majority7_module_38__or_module_4_U1 ( .A1(
        n_majority7_module_38__and_module_1_res), .A2(
        n_majority7_module_38__and_module_2_res), .ZN(
        n_majority7_module_38__or_module_4_res) );
  AND2_X1 u_majority7_module_38__and_module_5_U1 ( .A1(
        n_majority7_module_38__and_module_3_res), .A2(n_majority7_module_38_n3), .ZN(n_majority7_module_38__and_module_5_res) );
  OR2_X1 u_majority7_module_38__or_module_5_U1 ( .A1(n_majority7_module_38_n3), 
        .A2(n_majority7_module_38__and_module_3_res), .ZN(
        n_majority7_module_38__or_module_5_res) );
  AND2_X1 u_majority7_module_38__and_module_6_U1 ( .A1(
        n_majority7_module_38__or_module_1_res), .A2(
        n_majority7_module_38__or_module_2_res), .ZN(
        n_majority7_module_38__and_module_6_res) );
  OR2_X1 u_majority7_module_38__or_module_6_U1 ( .A1(
        n_majority7_module_38__or_module_2_res), .A2(
        n_majority7_module_38__or_module_1_res), .ZN(
        n_majority7_module_38__or_module_6_res) );
  OR2_X1 u_majority7_module_38__or_module_7_U1 ( .A1(
        n_majority7_module_38__and_module_4_res), .A2(
        n_majority7_module_38__and_module_5_res), .ZN(
        n_majority7_module_38__or_module_7_res) );
  AND2_X1 u_majority7_module_38__and_module_7_U1 ( .A1(
        n_majority7_module_38__or_module_3_res), .A2(
        n_majority7_module_38__or_module_4_res), .ZN(
        n_majority7_module_38__and_module_7_res) );
  OR2_X1 u_majority7_module_38__or_module_8_U1 ( .A1(
        n_majority7_module_38__or_module_4_res), .A2(
        n_majority7_module_38__or_module_3_res), .ZN(
        n_majority7_module_38__or_module_8_res) );
  AND2_X1 u_majority7_module_38__and_module_8_U1 ( .A1(
        n_majority7_module_38__or_module_5_res), .A2(
        n_majority7_module_38__and_module_6_res), .ZN(
        n_majority7_module_38__and_module_8_res) );
  OR2_X1 u_majority7_module_38__or_module_9_U1 ( .A1(
        n_majority7_module_38__and_module_6_res), .A2(
        n_majority7_module_38__or_module_5_res), .ZN(
        n_majority7_module_38__or_module_9_res) );
  OR2_X1 u_majority7_module_38__or_module_10_U1 ( .A1(
        n_majority7_module_38__or_module_7_res), .A2(
        n_majority7_module_38__and_module_7_res), .ZN(
        n_majority7_module_38__or_module_10_res) );
  AND2_X1 u_majority7_module_38__and_module_9_U1 ( .A1(
        n_majority7_module_38__or_module_6_res), .A2(
        n_majority7_module_38__or_module_9_res), .ZN(
        n_majority7_module_38__and_module_9_res) );
  OR2_X1 u_majority7_module_38__or_module_11_U1 ( .A1(
        n_majority7_module_38__or_module_10_res), .A2(
        n_majority7_module_38__and_module_8_res), .ZN(
        n_majority7_module_38__or_module_11_res) );
  AND2_X1 u_majority7_module_38__and_module_10_U1 ( .A1(
        n_majority7_module_38__or_module_8_res), .A2(
        n_majority7_module_38__and_module_9_res), .ZN(
        n_majority7_module_38__and_module_10_res) );
  AND2_X1 u_majority7_module_38__and_module_11_U1 ( .A1(
        n_majority7_module_38__and_module_10_res), .A2(
        n_majority7_module_38__or_module_11_res), .ZN(
        n_majority7_module_38_res) );
  DFF_X1 u_reg_module_39__cini_mul_v000_reg ( .D(n_majority7_module_38_res), 
        .CK(clock_4), .Q(n_reg_module_39_res), .QN() );
  BUF_X1 u_majority7_module_39_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_39_n7) );
  BUF_X1 u_majority7_module_39_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_39_n6) );
  BUF_X1 u_majority7_module_39_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_39_n5) );
  BUF_X1 u_majority7_module_39_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_39_n4) );
  BUF_X1 u_majority7_module_39_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_39_n3) );
  BUF_X1 u_majority7_module_39_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_39_n2) );
  BUF_X1 u_majority7_module_39_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_39_n1) );
  AND2_X1 u_majority7_module_39__and_module_1_U1 ( .A1(
        n_majority7_module_39_n5), .A2(n_majority7_module_39_n4), .ZN(
        n_majority7_module_39__and_module_1_res) );
  OR2_X1 u_majority7_module_39__or_module_1_U1 ( .A1(n_majority7_module_39_n4), 
        .A2(n_majority7_module_39_n5), .ZN(
        n_majority7_module_39__or_module_1_res) );
  AND2_X1 u_majority7_module_39__and_module_2_U1 ( .A1(
        n_majority7_module_39_n7), .A2(n_majority7_module_39_n2), .ZN(
        n_majority7_module_39__and_module_2_res) );
  OR2_X1 u_majority7_module_39__or_module_2_U1 ( .A1(n_majority7_module_39_n2), 
        .A2(n_majority7_module_39_n7), .ZN(
        n_majority7_module_39__or_module_2_res) );
  AND2_X1 u_majority7_module_39__and_module_3_U1 ( .A1(
        n_majority7_module_39_n6), .A2(n_majority7_module_39_n1), .ZN(
        n_majority7_module_39__and_module_3_res) );
  OR2_X1 u_majority7_module_39__or_module_3_U1 ( .A1(n_majority7_module_39_n1), 
        .A2(n_majority7_module_39_n6), .ZN(
        n_majority7_module_39__or_module_3_res) );
  AND2_X1 u_majority7_module_39__and_module_4_U1 ( .A1(
        n_majority7_module_39__and_module_2_res), .A2(
        n_majority7_module_39__and_module_1_res), .ZN(
        n_majority7_module_39__and_module_4_res) );
  OR2_X1 u_majority7_module_39__or_module_4_U1 ( .A1(
        n_majority7_module_39__and_module_1_res), .A2(
        n_majority7_module_39__and_module_2_res), .ZN(
        n_majority7_module_39__or_module_4_res) );
  AND2_X1 u_majority7_module_39__and_module_5_U1 ( .A1(
        n_majority7_module_39__and_module_3_res), .A2(n_majority7_module_39_n3), .ZN(n_majority7_module_39__and_module_5_res) );
  OR2_X1 u_majority7_module_39__or_module_5_U1 ( .A1(n_majority7_module_39_n3), 
        .A2(n_majority7_module_39__and_module_3_res), .ZN(
        n_majority7_module_39__or_module_5_res) );
  AND2_X1 u_majority7_module_39__and_module_6_U1 ( .A1(
        n_majority7_module_39__or_module_1_res), .A2(
        n_majority7_module_39__or_module_2_res), .ZN(
        n_majority7_module_39__and_module_6_res) );
  OR2_X1 u_majority7_module_39__or_module_6_U1 ( .A1(
        n_majority7_module_39__or_module_2_res), .A2(
        n_majority7_module_39__or_module_1_res), .ZN(
        n_majority7_module_39__or_module_6_res) );
  OR2_X1 u_majority7_module_39__or_module_7_U1 ( .A1(
        n_majority7_module_39__and_module_4_res), .A2(
        n_majority7_module_39__and_module_5_res), .ZN(
        n_majority7_module_39__or_module_7_res) );
  AND2_X1 u_majority7_module_39__and_module_7_U1 ( .A1(
        n_majority7_module_39__or_module_3_res), .A2(
        n_majority7_module_39__or_module_4_res), .ZN(
        n_majority7_module_39__and_module_7_res) );
  OR2_X1 u_majority7_module_39__or_module_8_U1 ( .A1(
        n_majority7_module_39__or_module_4_res), .A2(
        n_majority7_module_39__or_module_3_res), .ZN(
        n_majority7_module_39__or_module_8_res) );
  AND2_X1 u_majority7_module_39__and_module_8_U1 ( .A1(
        n_majority7_module_39__or_module_5_res), .A2(
        n_majority7_module_39__and_module_6_res), .ZN(
        n_majority7_module_39__and_module_8_res) );
  OR2_X1 u_majority7_module_39__or_module_9_U1 ( .A1(
        n_majority7_module_39__and_module_6_res), .A2(
        n_majority7_module_39__or_module_5_res), .ZN(
        n_majority7_module_39__or_module_9_res) );
  OR2_X1 u_majority7_module_39__or_module_10_U1 ( .A1(
        n_majority7_module_39__or_module_7_res), .A2(
        n_majority7_module_39__and_module_7_res), .ZN(
        n_majority7_module_39__or_module_10_res) );
  AND2_X1 u_majority7_module_39__and_module_9_U1 ( .A1(
        n_majority7_module_39__or_module_6_res), .A2(
        n_majority7_module_39__or_module_9_res), .ZN(
        n_majority7_module_39__and_module_9_res) );
  OR2_X1 u_majority7_module_39__or_module_11_U1 ( .A1(
        n_majority7_module_39__or_module_10_res), .A2(
        n_majority7_module_39__and_module_8_res), .ZN(
        n_majority7_module_39__or_module_11_res) );
  AND2_X1 u_majority7_module_39__and_module_10_U1 ( .A1(
        n_majority7_module_39__or_module_8_res), .A2(
        n_majority7_module_39__and_module_9_res), .ZN(
        n_majority7_module_39__and_module_10_res) );
  AND2_X1 u_majority7_module_39__and_module_11_U1 ( .A1(
        n_majority7_module_39__and_module_10_res), .A2(
        n_majority7_module_39__or_module_11_res), .ZN(
        n_majority7_module_39_res) );
  DFF_X1 u_reg_module_40__cini_mul_v000_reg ( .D(n_majority7_module_39_res), 
        .CK(clock_4), .Q(n_reg_module_40_res), .QN() );
  BUF_X1 u_majority7_module_40_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_40_n7) );
  BUF_X1 u_majority7_module_40_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_40_n6) );
  BUF_X1 u_majority7_module_40_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_40_n5) );
  BUF_X1 u_majority7_module_40_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_40_n4) );
  BUF_X1 u_majority7_module_40_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_40_n3) );
  BUF_X1 u_majority7_module_40_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_40_n2) );
  BUF_X1 u_majority7_module_40_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_40_n1) );
  AND2_X1 u_majority7_module_40__and_module_1_U1 ( .A1(
        n_majority7_module_40_n5), .A2(n_majority7_module_40_n4), .ZN(
        n_majority7_module_40__and_module_1_res) );
  OR2_X1 u_majority7_module_40__or_module_1_U1 ( .A1(n_majority7_module_40_n4), 
        .A2(n_majority7_module_40_n5), .ZN(
        n_majority7_module_40__or_module_1_res) );
  AND2_X1 u_majority7_module_40__and_module_2_U1 ( .A1(
        n_majority7_module_40_n7), .A2(n_majority7_module_40_n2), .ZN(
        n_majority7_module_40__and_module_2_res) );
  OR2_X1 u_majority7_module_40__or_module_2_U1 ( .A1(n_majority7_module_40_n2), 
        .A2(n_majority7_module_40_n7), .ZN(
        n_majority7_module_40__or_module_2_res) );
  AND2_X1 u_majority7_module_40__and_module_3_U1 ( .A1(
        n_majority7_module_40_n6), .A2(n_majority7_module_40_n1), .ZN(
        n_majority7_module_40__and_module_3_res) );
  OR2_X1 u_majority7_module_40__or_module_3_U1 ( .A1(n_majority7_module_40_n1), 
        .A2(n_majority7_module_40_n6), .ZN(
        n_majority7_module_40__or_module_3_res) );
  AND2_X1 u_majority7_module_40__and_module_4_U1 ( .A1(
        n_majority7_module_40__and_module_2_res), .A2(
        n_majority7_module_40__and_module_1_res), .ZN(
        n_majority7_module_40__and_module_4_res) );
  OR2_X1 u_majority7_module_40__or_module_4_U1 ( .A1(
        n_majority7_module_40__and_module_1_res), .A2(
        n_majority7_module_40__and_module_2_res), .ZN(
        n_majority7_module_40__or_module_4_res) );
  AND2_X1 u_majority7_module_40__and_module_5_U1 ( .A1(
        n_majority7_module_40__and_module_3_res), .A2(n_majority7_module_40_n3), .ZN(n_majority7_module_40__and_module_5_res) );
  OR2_X1 u_majority7_module_40__or_module_5_U1 ( .A1(n_majority7_module_40_n3), 
        .A2(n_majority7_module_40__and_module_3_res), .ZN(
        n_majority7_module_40__or_module_5_res) );
  AND2_X1 u_majority7_module_40__and_module_6_U1 ( .A1(
        n_majority7_module_40__or_module_1_res), .A2(
        n_majority7_module_40__or_module_2_res), .ZN(
        n_majority7_module_40__and_module_6_res) );
  OR2_X1 u_majority7_module_40__or_module_6_U1 ( .A1(
        n_majority7_module_40__or_module_2_res), .A2(
        n_majority7_module_40__or_module_1_res), .ZN(
        n_majority7_module_40__or_module_6_res) );
  OR2_X1 u_majority7_module_40__or_module_7_U1 ( .A1(
        n_majority7_module_40__and_module_4_res), .A2(
        n_majority7_module_40__and_module_5_res), .ZN(
        n_majority7_module_40__or_module_7_res) );
  AND2_X1 u_majority7_module_40__and_module_7_U1 ( .A1(
        n_majority7_module_40__or_module_3_res), .A2(
        n_majority7_module_40__or_module_4_res), .ZN(
        n_majority7_module_40__and_module_7_res) );
  OR2_X1 u_majority7_module_40__or_module_8_U1 ( .A1(
        n_majority7_module_40__or_module_4_res), .A2(
        n_majority7_module_40__or_module_3_res), .ZN(
        n_majority7_module_40__or_module_8_res) );
  AND2_X1 u_majority7_module_40__and_module_8_U1 ( .A1(
        n_majority7_module_40__or_module_5_res), .A2(
        n_majority7_module_40__and_module_6_res), .ZN(
        n_majority7_module_40__and_module_8_res) );
  OR2_X1 u_majority7_module_40__or_module_9_U1 ( .A1(
        n_majority7_module_40__and_module_6_res), .A2(
        n_majority7_module_40__or_module_5_res), .ZN(
        n_majority7_module_40__or_module_9_res) );
  OR2_X1 u_majority7_module_40__or_module_10_U1 ( .A1(
        n_majority7_module_40__or_module_7_res), .A2(
        n_majority7_module_40__and_module_7_res), .ZN(
        n_majority7_module_40__or_module_10_res) );
  AND2_X1 u_majority7_module_40__and_module_9_U1 ( .A1(
        n_majority7_module_40__or_module_6_res), .A2(
        n_majority7_module_40__or_module_9_res), .ZN(
        n_majority7_module_40__and_module_9_res) );
  OR2_X1 u_majority7_module_40__or_module_11_U1 ( .A1(
        n_majority7_module_40__or_module_10_res), .A2(
        n_majority7_module_40__and_module_8_res), .ZN(
        n_majority7_module_40__or_module_11_res) );
  AND2_X1 u_majority7_module_40__and_module_10_U1 ( .A1(
        n_majority7_module_40__or_module_8_res), .A2(
        n_majority7_module_40__and_module_9_res), .ZN(
        n_majority7_module_40__and_module_10_res) );
  AND2_X1 u_majority7_module_40__and_module_11_U1 ( .A1(
        n_majority7_module_40__and_module_10_res), .A2(
        n_majority7_module_40__or_module_11_res), .ZN(
        n_majority7_module_40_res) );
  DFF_X1 u_reg_module_41__cini_mul_v000_reg ( .D(n_majority7_module_40_res), 
        .CK(clock_4), .Q(n_reg_module_41_res), .QN() );
  BUF_X1 u_majority7_module_41_U7 ( .A(n_xor_module_22_res), .Z(
        n_majority7_module_41_n7) );
  BUF_X1 u_majority7_module_41_U6 ( .A(n_xor_module_34_res), .Z(
        n_majority7_module_41_n6) );
  BUF_X1 u_majority7_module_41_U5 ( .A(n_xor_module_40_res), .Z(
        n_majority7_module_41_n5) );
  BUF_X1 u_majority7_module_41_U4 ( .A(n_xor_module_4_res), .Z(
        n_majority7_module_41_n4) );
  BUF_X1 u_majority7_module_41_U3 ( .A(n_xor_module_10_res), .Z(
        n_majority7_module_41_n3) );
  BUF_X1 u_majority7_module_41_U2 ( .A(n_xor_module_16_res), .Z(
        n_majority7_module_41_n2) );
  BUF_X1 u_majority7_module_41_U1 ( .A(n_xor_module_28_res), .Z(
        n_majority7_module_41_n1) );
  AND2_X1 u_majority7_module_41__and_module_1_U1 ( .A1(
        n_majority7_module_41_n5), .A2(n_majority7_module_41_n4), .ZN(
        n_majority7_module_41__and_module_1_res) );
  OR2_X1 u_majority7_module_41__or_module_1_U1 ( .A1(n_majority7_module_41_n4), 
        .A2(n_majority7_module_41_n5), .ZN(
        n_majority7_module_41__or_module_1_res) );
  AND2_X1 u_majority7_module_41__and_module_2_U1 ( .A1(
        n_majority7_module_41_n7), .A2(n_majority7_module_41_n2), .ZN(
        n_majority7_module_41__and_module_2_res) );
  OR2_X1 u_majority7_module_41__or_module_2_U1 ( .A1(n_majority7_module_41_n2), 
        .A2(n_majority7_module_41_n7), .ZN(
        n_majority7_module_41__or_module_2_res) );
  AND2_X1 u_majority7_module_41__and_module_3_U1 ( .A1(
        n_majority7_module_41_n6), .A2(n_majority7_module_41_n1), .ZN(
        n_majority7_module_41__and_module_3_res) );
  OR2_X1 u_majority7_module_41__or_module_3_U1 ( .A1(n_majority7_module_41_n1), 
        .A2(n_majority7_module_41_n6), .ZN(
        n_majority7_module_41__or_module_3_res) );
  AND2_X1 u_majority7_module_41__and_module_4_U1 ( .A1(
        n_majority7_module_41__and_module_2_res), .A2(
        n_majority7_module_41__and_module_1_res), .ZN(
        n_majority7_module_41__and_module_4_res) );
  OR2_X1 u_majority7_module_41__or_module_4_U1 ( .A1(
        n_majority7_module_41__and_module_1_res), .A2(
        n_majority7_module_41__and_module_2_res), .ZN(
        n_majority7_module_41__or_module_4_res) );
  AND2_X1 u_majority7_module_41__and_module_5_U1 ( .A1(
        n_majority7_module_41__and_module_3_res), .A2(n_majority7_module_41_n3), .ZN(n_majority7_module_41__and_module_5_res) );
  OR2_X1 u_majority7_module_41__or_module_5_U1 ( .A1(n_majority7_module_41_n3), 
        .A2(n_majority7_module_41__and_module_3_res), .ZN(
        n_majority7_module_41__or_module_5_res) );
  AND2_X1 u_majority7_module_41__and_module_6_U1 ( .A1(
        n_majority7_module_41__or_module_1_res), .A2(
        n_majority7_module_41__or_module_2_res), .ZN(
        n_majority7_module_41__and_module_6_res) );
  OR2_X1 u_majority7_module_41__or_module_6_U1 ( .A1(
        n_majority7_module_41__or_module_2_res), .A2(
        n_majority7_module_41__or_module_1_res), .ZN(
        n_majority7_module_41__or_module_6_res) );
  OR2_X1 u_majority7_module_41__or_module_7_U1 ( .A1(
        n_majority7_module_41__and_module_4_res), .A2(
        n_majority7_module_41__and_module_5_res), .ZN(
        n_majority7_module_41__or_module_7_res) );
  AND2_X1 u_majority7_module_41__and_module_7_U1 ( .A1(
        n_majority7_module_41__or_module_3_res), .A2(
        n_majority7_module_41__or_module_4_res), .ZN(
        n_majority7_module_41__and_module_7_res) );
  OR2_X1 u_majority7_module_41__or_module_8_U1 ( .A1(
        n_majority7_module_41__or_module_4_res), .A2(
        n_majority7_module_41__or_module_3_res), .ZN(
        n_majority7_module_41__or_module_8_res) );
  AND2_X1 u_majority7_module_41__and_module_8_U1 ( .A1(
        n_majority7_module_41__or_module_5_res), .A2(
        n_majority7_module_41__and_module_6_res), .ZN(
        n_majority7_module_41__and_module_8_res) );
  OR2_X1 u_majority7_module_41__or_module_9_U1 ( .A1(
        n_majority7_module_41__and_module_6_res), .A2(
        n_majority7_module_41__or_module_5_res), .ZN(
        n_majority7_module_41__or_module_9_res) );
  OR2_X1 u_majority7_module_41__or_module_10_U1 ( .A1(
        n_majority7_module_41__or_module_7_res), .A2(
        n_majority7_module_41__and_module_7_res), .ZN(
        n_majority7_module_41__or_module_10_res) );
  AND2_X1 u_majority7_module_41__and_module_9_U1 ( .A1(
        n_majority7_module_41__or_module_6_res), .A2(
        n_majority7_module_41__or_module_9_res), .ZN(
        n_majority7_module_41__and_module_9_res) );
  OR2_X1 u_majority7_module_41__or_module_11_U1 ( .A1(
        n_majority7_module_41__or_module_10_res), .A2(
        n_majority7_module_41__and_module_8_res), .ZN(
        n_majority7_module_41__or_module_11_res) );
  AND2_X1 u_majority7_module_41__and_module_10_U1 ( .A1(
        n_majority7_module_41__or_module_8_res), .A2(
        n_majority7_module_41__and_module_9_res), .ZN(
        n_majority7_module_41__and_module_10_res) );
  AND2_X1 u_majority7_module_41__and_module_11_U1 ( .A1(
        n_majority7_module_41__and_module_10_res), .A2(
        n_majority7_module_41__or_module_11_res), .ZN(
        n_majority7_module_41_res) );
  DFF_X1 u_reg_module_42__cini_mul_v000_reg ( .D(n_majority7_module_41_res), 
        .CK(clock_4), .Q(n_reg_module_42_res), .QN() );
  BUF_X1 u_majority7_module_42_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_42_n7) );
  BUF_X1 u_majority7_module_42_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_42_n6) );
  BUF_X1 u_majority7_module_42_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_42_n5) );
  BUF_X1 u_majority7_module_42_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_42_n4) );
  BUF_X1 u_majority7_module_42_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_42_n3) );
  BUF_X1 u_majority7_module_42_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_42_n2) );
  BUF_X1 u_majority7_module_42_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_42_n1) );
  AND2_X1 u_majority7_module_42__and_module_1_U1 ( .A1(
        n_majority7_module_42_n5), .A2(n_majority7_module_42_n4), .ZN(
        n_majority7_module_42__and_module_1_res) );
  OR2_X1 u_majority7_module_42__or_module_1_U1 ( .A1(n_majority7_module_42_n4), 
        .A2(n_majority7_module_42_n5), .ZN(
        n_majority7_module_42__or_module_1_res) );
  AND2_X1 u_majority7_module_42__and_module_2_U1 ( .A1(
        n_majority7_module_42_n7), .A2(n_majority7_module_42_n2), .ZN(
        n_majority7_module_42__and_module_2_res) );
  OR2_X1 u_majority7_module_42__or_module_2_U1 ( .A1(n_majority7_module_42_n2), 
        .A2(n_majority7_module_42_n7), .ZN(
        n_majority7_module_42__or_module_2_res) );
  AND2_X1 u_majority7_module_42__and_module_3_U1 ( .A1(
        n_majority7_module_42_n6), .A2(n_majority7_module_42_n1), .ZN(
        n_majority7_module_42__and_module_3_res) );
  OR2_X1 u_majority7_module_42__or_module_3_U1 ( .A1(n_majority7_module_42_n1), 
        .A2(n_majority7_module_42_n6), .ZN(
        n_majority7_module_42__or_module_3_res) );
  AND2_X1 u_majority7_module_42__and_module_4_U1 ( .A1(
        n_majority7_module_42__and_module_2_res), .A2(
        n_majority7_module_42__and_module_1_res), .ZN(
        n_majority7_module_42__and_module_4_res) );
  OR2_X1 u_majority7_module_42__or_module_4_U1 ( .A1(
        n_majority7_module_42__and_module_1_res), .A2(
        n_majority7_module_42__and_module_2_res), .ZN(
        n_majority7_module_42__or_module_4_res) );
  AND2_X1 u_majority7_module_42__and_module_5_U1 ( .A1(
        n_majority7_module_42__and_module_3_res), .A2(n_majority7_module_42_n3), .ZN(n_majority7_module_42__and_module_5_res) );
  OR2_X1 u_majority7_module_42__or_module_5_U1 ( .A1(n_majority7_module_42_n3), 
        .A2(n_majority7_module_42__and_module_3_res), .ZN(
        n_majority7_module_42__or_module_5_res) );
  AND2_X1 u_majority7_module_42__and_module_6_U1 ( .A1(
        n_majority7_module_42__or_module_1_res), .A2(
        n_majority7_module_42__or_module_2_res), .ZN(
        n_majority7_module_42__and_module_6_res) );
  OR2_X1 u_majority7_module_42__or_module_6_U1 ( .A1(
        n_majority7_module_42__or_module_2_res), .A2(
        n_majority7_module_42__or_module_1_res), .ZN(
        n_majority7_module_42__or_module_6_res) );
  OR2_X1 u_majority7_module_42__or_module_7_U1 ( .A1(
        n_majority7_module_42__and_module_4_res), .A2(
        n_majority7_module_42__and_module_5_res), .ZN(
        n_majority7_module_42__or_module_7_res) );
  AND2_X1 u_majority7_module_42__and_module_7_U1 ( .A1(
        n_majority7_module_42__or_module_3_res), .A2(
        n_majority7_module_42__or_module_4_res), .ZN(
        n_majority7_module_42__and_module_7_res) );
  OR2_X1 u_majority7_module_42__or_module_8_U1 ( .A1(
        n_majority7_module_42__or_module_4_res), .A2(
        n_majority7_module_42__or_module_3_res), .ZN(
        n_majority7_module_42__or_module_8_res) );
  AND2_X1 u_majority7_module_42__and_module_8_U1 ( .A1(
        n_majority7_module_42__or_module_5_res), .A2(
        n_majority7_module_42__and_module_6_res), .ZN(
        n_majority7_module_42__and_module_8_res) );
  OR2_X1 u_majority7_module_42__or_module_9_U1 ( .A1(
        n_majority7_module_42__and_module_6_res), .A2(
        n_majority7_module_42__or_module_5_res), .ZN(
        n_majority7_module_42__or_module_9_res) );
  OR2_X1 u_majority7_module_42__or_module_10_U1 ( .A1(
        n_majority7_module_42__or_module_7_res), .A2(
        n_majority7_module_42__and_module_7_res), .ZN(
        n_majority7_module_42__or_module_10_res) );
  AND2_X1 u_majority7_module_42__and_module_9_U1 ( .A1(
        n_majority7_module_42__or_module_6_res), .A2(
        n_majority7_module_42__or_module_9_res), .ZN(
        n_majority7_module_42__and_module_9_res) );
  OR2_X1 u_majority7_module_42__or_module_11_U1 ( .A1(
        n_majority7_module_42__or_module_10_res), .A2(
        n_majority7_module_42__and_module_8_res), .ZN(
        n_majority7_module_42__or_module_11_res) );
  AND2_X1 u_majority7_module_42__and_module_10_U1 ( .A1(
        n_majority7_module_42__or_module_8_res), .A2(
        n_majority7_module_42__and_module_9_res), .ZN(
        n_majority7_module_42__and_module_10_res) );
  AND2_X1 u_majority7_module_42__and_module_11_U1 ( .A1(
        n_majority7_module_42__and_module_10_res), .A2(
        n_majority7_module_42__or_module_11_res), .ZN(
        n_majority7_module_42_res) );
  DFF_X1 u_reg_module_43__cini_mul_v000_reg ( .D(n_majority7_module_42_res), 
        .CK(clock_4), .Q(n_reg_module_43_res), .QN() );
  BUF_X1 u_majority7_module_43_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_43_n7) );
  BUF_X1 u_majority7_module_43_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_43_n6) );
  BUF_X1 u_majority7_module_43_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_43_n5) );
  BUF_X1 u_majority7_module_43_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_43_n4) );
  BUF_X1 u_majority7_module_43_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_43_n3) );
  BUF_X1 u_majority7_module_43_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_43_n2) );
  BUF_X1 u_majority7_module_43_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_43_n1) );
  AND2_X1 u_majority7_module_43__and_module_1_U1 ( .A1(
        n_majority7_module_43_n5), .A2(n_majority7_module_43_n4), .ZN(
        n_majority7_module_43__and_module_1_res) );
  OR2_X1 u_majority7_module_43__or_module_1_U1 ( .A1(n_majority7_module_43_n4), 
        .A2(n_majority7_module_43_n5), .ZN(
        n_majority7_module_43__or_module_1_res) );
  AND2_X1 u_majority7_module_43__and_module_2_U1 ( .A1(
        n_majority7_module_43_n7), .A2(n_majority7_module_43_n2), .ZN(
        n_majority7_module_43__and_module_2_res) );
  OR2_X1 u_majority7_module_43__or_module_2_U1 ( .A1(n_majority7_module_43_n2), 
        .A2(n_majority7_module_43_n7), .ZN(
        n_majority7_module_43__or_module_2_res) );
  AND2_X1 u_majority7_module_43__and_module_3_U1 ( .A1(
        n_majority7_module_43_n6), .A2(n_majority7_module_43_n1), .ZN(
        n_majority7_module_43__and_module_3_res) );
  OR2_X1 u_majority7_module_43__or_module_3_U1 ( .A1(n_majority7_module_43_n1), 
        .A2(n_majority7_module_43_n6), .ZN(
        n_majority7_module_43__or_module_3_res) );
  AND2_X1 u_majority7_module_43__and_module_4_U1 ( .A1(
        n_majority7_module_43__and_module_2_res), .A2(
        n_majority7_module_43__and_module_1_res), .ZN(
        n_majority7_module_43__and_module_4_res) );
  OR2_X1 u_majority7_module_43__or_module_4_U1 ( .A1(
        n_majority7_module_43__and_module_1_res), .A2(
        n_majority7_module_43__and_module_2_res), .ZN(
        n_majority7_module_43__or_module_4_res) );
  AND2_X1 u_majority7_module_43__and_module_5_U1 ( .A1(
        n_majority7_module_43__and_module_3_res), .A2(n_majority7_module_43_n3), .ZN(n_majority7_module_43__and_module_5_res) );
  OR2_X1 u_majority7_module_43__or_module_5_U1 ( .A1(n_majority7_module_43_n3), 
        .A2(n_majority7_module_43__and_module_3_res), .ZN(
        n_majority7_module_43__or_module_5_res) );
  AND2_X1 u_majority7_module_43__and_module_6_U1 ( .A1(
        n_majority7_module_43__or_module_1_res), .A2(
        n_majority7_module_43__or_module_2_res), .ZN(
        n_majority7_module_43__and_module_6_res) );
  OR2_X1 u_majority7_module_43__or_module_6_U1 ( .A1(
        n_majority7_module_43__or_module_2_res), .A2(
        n_majority7_module_43__or_module_1_res), .ZN(
        n_majority7_module_43__or_module_6_res) );
  OR2_X1 u_majority7_module_43__or_module_7_U1 ( .A1(
        n_majority7_module_43__and_module_4_res), .A2(
        n_majority7_module_43__and_module_5_res), .ZN(
        n_majority7_module_43__or_module_7_res) );
  AND2_X1 u_majority7_module_43__and_module_7_U1 ( .A1(
        n_majority7_module_43__or_module_3_res), .A2(
        n_majority7_module_43__or_module_4_res), .ZN(
        n_majority7_module_43__and_module_7_res) );
  OR2_X1 u_majority7_module_43__or_module_8_U1 ( .A1(
        n_majority7_module_43__or_module_4_res), .A2(
        n_majority7_module_43__or_module_3_res), .ZN(
        n_majority7_module_43__or_module_8_res) );
  AND2_X1 u_majority7_module_43__and_module_8_U1 ( .A1(
        n_majority7_module_43__or_module_5_res), .A2(
        n_majority7_module_43__and_module_6_res), .ZN(
        n_majority7_module_43__and_module_8_res) );
  OR2_X1 u_majority7_module_43__or_module_9_U1 ( .A1(
        n_majority7_module_43__and_module_6_res), .A2(
        n_majority7_module_43__or_module_5_res), .ZN(
        n_majority7_module_43__or_module_9_res) );
  OR2_X1 u_majority7_module_43__or_module_10_U1 ( .A1(
        n_majority7_module_43__or_module_7_res), .A2(
        n_majority7_module_43__and_module_7_res), .ZN(
        n_majority7_module_43__or_module_10_res) );
  AND2_X1 u_majority7_module_43__and_module_9_U1 ( .A1(
        n_majority7_module_43__or_module_6_res), .A2(
        n_majority7_module_43__or_module_9_res), .ZN(
        n_majority7_module_43__and_module_9_res) );
  OR2_X1 u_majority7_module_43__or_module_11_U1 ( .A1(
        n_majority7_module_43__or_module_10_res), .A2(
        n_majority7_module_43__and_module_8_res), .ZN(
        n_majority7_module_43__or_module_11_res) );
  AND2_X1 u_majority7_module_43__and_module_10_U1 ( .A1(
        n_majority7_module_43__or_module_8_res), .A2(
        n_majority7_module_43__and_module_9_res), .ZN(
        n_majority7_module_43__and_module_10_res) );
  AND2_X1 u_majority7_module_43__and_module_11_U1 ( .A1(
        n_majority7_module_43__and_module_10_res), .A2(
        n_majority7_module_43__or_module_11_res), .ZN(
        n_majority7_module_43_res) );
  DFF_X1 u_reg_module_44__cini_mul_v000_reg ( .D(n_majority7_module_43_res), 
        .CK(clock_4), .Q(n_reg_module_44_res), .QN() );
  BUF_X1 u_majority7_module_44_U7 ( .A(n_xor_module_24_res), .Z(
        n_majority7_module_44_n7) );
  BUF_X1 u_majority7_module_44_U6 ( .A(n_xor_module_36_res), .Z(
        n_majority7_module_44_n6) );
  BUF_X1 u_majority7_module_44_U5 ( .A(n_xor_module_42_res), .Z(
        n_majority7_module_44_n5) );
  BUF_X1 u_majority7_module_44_U4 ( .A(n_xor_module_6_res), .Z(
        n_majority7_module_44_n4) );
  BUF_X1 u_majority7_module_44_U3 ( .A(n_xor_module_12_res), .Z(
        n_majority7_module_44_n3) );
  BUF_X1 u_majority7_module_44_U2 ( .A(n_xor_module_18_res), .Z(
        n_majority7_module_44_n2) );
  BUF_X1 u_majority7_module_44_U1 ( .A(n_xor_module_30_res), .Z(
        n_majority7_module_44_n1) );
  AND2_X1 u_majority7_module_44__and_module_1_U1 ( .A1(
        n_majority7_module_44_n5), .A2(n_majority7_module_44_n4), .ZN(
        n_majority7_module_44__and_module_1_res) );
  OR2_X1 u_majority7_module_44__or_module_1_U1 ( .A1(n_majority7_module_44_n4), 
        .A2(n_majority7_module_44_n5), .ZN(
        n_majority7_module_44__or_module_1_res) );
  AND2_X1 u_majority7_module_44__and_module_2_U1 ( .A1(
        n_majority7_module_44_n7), .A2(n_majority7_module_44_n2), .ZN(
        n_majority7_module_44__and_module_2_res) );
  OR2_X1 u_majority7_module_44__or_module_2_U1 ( .A1(n_majority7_module_44_n2), 
        .A2(n_majority7_module_44_n7), .ZN(
        n_majority7_module_44__or_module_2_res) );
  AND2_X1 u_majority7_module_44__and_module_3_U1 ( .A1(
        n_majority7_module_44_n6), .A2(n_majority7_module_44_n1), .ZN(
        n_majority7_module_44__and_module_3_res) );
  OR2_X1 u_majority7_module_44__or_module_3_U1 ( .A1(n_majority7_module_44_n1), 
        .A2(n_majority7_module_44_n6), .ZN(
        n_majority7_module_44__or_module_3_res) );
  AND2_X1 u_majority7_module_44__and_module_4_U1 ( .A1(
        n_majority7_module_44__and_module_2_res), .A2(
        n_majority7_module_44__and_module_1_res), .ZN(
        n_majority7_module_44__and_module_4_res) );
  OR2_X1 u_majority7_module_44__or_module_4_U1 ( .A1(
        n_majority7_module_44__and_module_1_res), .A2(
        n_majority7_module_44__and_module_2_res), .ZN(
        n_majority7_module_44__or_module_4_res) );
  AND2_X1 u_majority7_module_44__and_module_5_U1 ( .A1(
        n_majority7_module_44__and_module_3_res), .A2(n_majority7_module_44_n3), .ZN(n_majority7_module_44__and_module_5_res) );
  OR2_X1 u_majority7_module_44__or_module_5_U1 ( .A1(n_majority7_module_44_n3), 
        .A2(n_majority7_module_44__and_module_3_res), .ZN(
        n_majority7_module_44__or_module_5_res) );
  AND2_X1 u_majority7_module_44__and_module_6_U1 ( .A1(
        n_majority7_module_44__or_module_1_res), .A2(
        n_majority7_module_44__or_module_2_res), .ZN(
        n_majority7_module_44__and_module_6_res) );
  OR2_X1 u_majority7_module_44__or_module_6_U1 ( .A1(
        n_majority7_module_44__or_module_2_res), .A2(
        n_majority7_module_44__or_module_1_res), .ZN(
        n_majority7_module_44__or_module_6_res) );
  OR2_X1 u_majority7_module_44__or_module_7_U1 ( .A1(
        n_majority7_module_44__and_module_4_res), .A2(
        n_majority7_module_44__and_module_5_res), .ZN(
        n_majority7_module_44__or_module_7_res) );
  AND2_X1 u_majority7_module_44__and_module_7_U1 ( .A1(
        n_majority7_module_44__or_module_3_res), .A2(
        n_majority7_module_44__or_module_4_res), .ZN(
        n_majority7_module_44__and_module_7_res) );
  OR2_X1 u_majority7_module_44__or_module_8_U1 ( .A1(
        n_majority7_module_44__or_module_4_res), .A2(
        n_majority7_module_44__or_module_3_res), .ZN(
        n_majority7_module_44__or_module_8_res) );
  AND2_X1 u_majority7_module_44__and_module_8_U1 ( .A1(
        n_majority7_module_44__or_module_5_res), .A2(
        n_majority7_module_44__and_module_6_res), .ZN(
        n_majority7_module_44__and_module_8_res) );
  OR2_X1 u_majority7_module_44__or_module_9_U1 ( .A1(
        n_majority7_module_44__and_module_6_res), .A2(
        n_majority7_module_44__or_module_5_res), .ZN(
        n_majority7_module_44__or_module_9_res) );
  OR2_X1 u_majority7_module_44__or_module_10_U1 ( .A1(
        n_majority7_module_44__or_module_7_res), .A2(
        n_majority7_module_44__and_module_7_res), .ZN(
        n_majority7_module_44__or_module_10_res) );
  AND2_X1 u_majority7_module_44__and_module_9_U1 ( .A1(
        n_majority7_module_44__or_module_6_res), .A2(
        n_majority7_module_44__or_module_9_res), .ZN(
        n_majority7_module_44__and_module_9_res) );
  OR2_X1 u_majority7_module_44__or_module_11_U1 ( .A1(
        n_majority7_module_44__or_module_10_res), .A2(
        n_majority7_module_44__and_module_8_res), .ZN(
        n_majority7_module_44__or_module_11_res) );
  AND2_X1 u_majority7_module_44__and_module_10_U1 ( .A1(
        n_majority7_module_44__or_module_8_res), .A2(
        n_majority7_module_44__and_module_9_res), .ZN(
        n_majority7_module_44__and_module_10_res) );
  AND2_X1 u_majority7_module_44__and_module_11_U1 ( .A1(
        n_majority7_module_44__and_module_10_res), .A2(
        n_majority7_module_44__or_module_11_res), .ZN(
        n_majority7_module_44_res) );
  DFF_X1 u_reg_module_45__cini_mul_v000_reg ( .D(n_majority7_module_44_res), 
        .CK(clock_4), .Q(n_reg_module_45_res), .QN() );
  AND2_X1 u_majority7_module_45__and_module_1_U1 ( .A1(n_xor_module_38_res), 
        .A2(n_xor_module_2_res), .ZN(n_majority7_module_45__and_module_1_res)
         );
  OR2_X1 u_majority7_module_45__or_module_1_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_38_res), .ZN(n_majority7_module_45__or_module_1_res) );
  AND2_X1 u_majority7_module_45__and_module_2_U1 ( .A1(n_xor_module_20_res), 
        .A2(n_xor_module_14_res), .ZN(n_majority7_module_45__and_module_2_res)
         );
  OR2_X1 u_majority7_module_45__or_module_2_U1 ( .A1(n_xor_module_14_res), 
        .A2(n_xor_module_20_res), .ZN(n_majority7_module_45__or_module_2_res)
         );
  AND2_X1 u_majority7_module_45__and_module_3_U1 ( .A1(n_xor_module_32_res), 
        .A2(n_xor_module_26_res), .ZN(n_majority7_module_45__and_module_3_res)
         );
  OR2_X1 u_majority7_module_45__or_module_3_U1 ( .A1(n_xor_module_26_res), 
        .A2(n_xor_module_32_res), .ZN(n_majority7_module_45__or_module_3_res)
         );
  AND2_X1 u_majority7_module_45__and_module_4_U1 ( .A1(
        n_majority7_module_45__and_module_2_res), .A2(
        n_majority7_module_45__and_module_1_res), .ZN(
        n_majority7_module_45__and_module_4_res) );
  OR2_X1 u_majority7_module_45__or_module_4_U1 ( .A1(
        n_majority7_module_45__and_module_1_res), .A2(
        n_majority7_module_45__and_module_2_res), .ZN(
        n_majority7_module_45__or_module_4_res) );
  AND2_X1 u_majority7_module_45__and_module_5_U1 ( .A1(
        n_majority7_module_45__and_module_3_res), .A2(n_xor_module_8_res), 
        .ZN(n_majority7_module_45__and_module_5_res) );
  OR2_X1 u_majority7_module_45__or_module_5_U1 ( .A1(n_xor_module_8_res), .A2(
        n_majority7_module_45__and_module_3_res), .ZN(
        n_majority7_module_45__or_module_5_res) );
  AND2_X1 u_majority7_module_45__and_module_6_U1 ( .A1(
        n_majority7_module_45__or_module_1_res), .A2(
        n_majority7_module_45__or_module_2_res), .ZN(
        n_majority7_module_45__and_module_6_res) );
  OR2_X1 u_majority7_module_45__or_module_6_U1 ( .A1(
        n_majority7_module_45__or_module_2_res), .A2(
        n_majority7_module_45__or_module_1_res), .ZN(
        n_majority7_module_45__or_module_6_res) );
  OR2_X1 u_majority7_module_45__or_module_7_U1 ( .A1(
        n_majority7_module_45__and_module_4_res), .A2(
        n_majority7_module_45__and_module_5_res), .ZN(
        n_majority7_module_45__or_module_7_res) );
  AND2_X1 u_majority7_module_45__and_module_7_U1 ( .A1(
        n_majority7_module_45__or_module_3_res), .A2(
        n_majority7_module_45__or_module_4_res), .ZN(
        n_majority7_module_45__and_module_7_res) );
  OR2_X1 u_majority7_module_45__or_module_8_U1 ( .A1(
        n_majority7_module_45__or_module_4_res), .A2(
        n_majority7_module_45__or_module_3_res), .ZN(
        n_majority7_module_45__or_module_8_res) );
  AND2_X1 u_majority7_module_45__and_module_8_U1 ( .A1(
        n_majority7_module_45__or_module_5_res), .A2(
        n_majority7_module_45__and_module_6_res), .ZN(
        n_majority7_module_45__and_module_8_res) );
  OR2_X1 u_majority7_module_45__or_module_9_U1 ( .A1(
        n_majority7_module_45__and_module_6_res), .A2(
        n_majority7_module_45__or_module_5_res), .ZN(
        n_majority7_module_45__or_module_9_res) );
  OR2_X1 u_majority7_module_45__or_module_10_U1 ( .A1(
        n_majority7_module_45__or_module_7_res), .A2(
        n_majority7_module_45__and_module_7_res), .ZN(
        n_majority7_module_45__or_module_10_res) );
  AND2_X1 u_majority7_module_45__and_module_9_U1 ( .A1(
        n_majority7_module_45__or_module_6_res), .A2(
        n_majority7_module_45__or_module_9_res), .ZN(
        n_majority7_module_45__and_module_9_res) );
  OR2_X1 u_majority7_module_45__or_module_11_U1 ( .A1(
        n_majority7_module_45__or_module_10_res), .A2(
        n_majority7_module_45__and_module_8_res), .ZN(
        n_majority7_module_45__or_module_11_res) );
  AND2_X1 u_majority7_module_45__and_module_10_U1 ( .A1(
        n_majority7_module_45__or_module_8_res), .A2(
        n_majority7_module_45__and_module_9_res), .ZN(
        n_majority7_module_45__and_module_10_res) );
  AND2_X1 u_majority7_module_45__and_module_11_U1 ( .A1(
        n_majority7_module_45__and_module_10_res), .A2(
        n_majority7_module_45__or_module_11_res), .ZN(
        n_majority7_module_45_res) );
  DFF_X1 u_reg_module_46__cini_mul_v000_reg ( .D(n_majority7_module_45_res), 
        .CK(clock_5), .Q(n_reg_module_46_res), .QN() );
  AND2_X1 u_majority7_module_46__and_module_1_U1 ( .A1(n_xor_module_38_res), 
        .A2(n_xor_module_2_res), .ZN(n_majority7_module_46__and_module_1_res)
         );
  OR2_X1 u_majority7_module_46__or_module_1_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_38_res), .ZN(n_majority7_module_46__or_module_1_res) );
  AND2_X1 u_majority7_module_46__and_module_2_U1 ( .A1(n_xor_module_20_res), 
        .A2(n_xor_module_14_res), .ZN(n_majority7_module_46__and_module_2_res)
         );
  OR2_X1 u_majority7_module_46__or_module_2_U1 ( .A1(n_xor_module_14_res), 
        .A2(n_xor_module_20_res), .ZN(n_majority7_module_46__or_module_2_res)
         );
  AND2_X1 u_majority7_module_46__and_module_3_U1 ( .A1(n_xor_module_32_res), 
        .A2(n_xor_module_26_res), .ZN(n_majority7_module_46__and_module_3_res)
         );
  OR2_X1 u_majority7_module_46__or_module_3_U1 ( .A1(n_xor_module_26_res), 
        .A2(n_xor_module_32_res), .ZN(n_majority7_module_46__or_module_3_res)
         );
  AND2_X1 u_majority7_module_46__and_module_4_U1 ( .A1(
        n_majority7_module_46__and_module_2_res), .A2(
        n_majority7_module_46__and_module_1_res), .ZN(
        n_majority7_module_46__and_module_4_res) );
  OR2_X1 u_majority7_module_46__or_module_4_U1 ( .A1(
        n_majority7_module_46__and_module_1_res), .A2(
        n_majority7_module_46__and_module_2_res), .ZN(
        n_majority7_module_46__or_module_4_res) );
  AND2_X1 u_majority7_module_46__and_module_5_U1 ( .A1(
        n_majority7_module_46__and_module_3_res), .A2(n_xor_module_8_res), 
        .ZN(n_majority7_module_46__and_module_5_res) );
  OR2_X1 u_majority7_module_46__or_module_5_U1 ( .A1(n_xor_module_8_res), .A2(
        n_majority7_module_46__and_module_3_res), .ZN(
        n_majority7_module_46__or_module_5_res) );
  AND2_X1 u_majority7_module_46__and_module_6_U1 ( .A1(
        n_majority7_module_46__or_module_1_res), .A2(
        n_majority7_module_46__or_module_2_res), .ZN(
        n_majority7_module_46__and_module_6_res) );
  OR2_X1 u_majority7_module_46__or_module_6_U1 ( .A1(
        n_majority7_module_46__or_module_2_res), .A2(
        n_majority7_module_46__or_module_1_res), .ZN(
        n_majority7_module_46__or_module_6_res) );
  OR2_X1 u_majority7_module_46__or_module_7_U1 ( .A1(
        n_majority7_module_46__and_module_4_res), .A2(
        n_majority7_module_46__and_module_5_res), .ZN(
        n_majority7_module_46__or_module_7_res) );
  AND2_X1 u_majority7_module_46__and_module_7_U1 ( .A1(
        n_majority7_module_46__or_module_3_res), .A2(
        n_majority7_module_46__or_module_4_res), .ZN(
        n_majority7_module_46__and_module_7_res) );
  OR2_X1 u_majority7_module_46__or_module_8_U1 ( .A1(
        n_majority7_module_46__or_module_4_res), .A2(
        n_majority7_module_46__or_module_3_res), .ZN(
        n_majority7_module_46__or_module_8_res) );
  AND2_X1 u_majority7_module_46__and_module_8_U1 ( .A1(
        n_majority7_module_46__or_module_5_res), .A2(
        n_majority7_module_46__and_module_6_res), .ZN(
        n_majority7_module_46__and_module_8_res) );
  OR2_X1 u_majority7_module_46__or_module_9_U1 ( .A1(
        n_majority7_module_46__and_module_6_res), .A2(
        n_majority7_module_46__or_module_5_res), .ZN(
        n_majority7_module_46__or_module_9_res) );
  OR2_X1 u_majority7_module_46__or_module_10_U1 ( .A1(
        n_majority7_module_46__or_module_7_res), .A2(
        n_majority7_module_46__and_module_7_res), .ZN(
        n_majority7_module_46__or_module_10_res) );
  AND2_X1 u_majority7_module_46__and_module_9_U1 ( .A1(
        n_majority7_module_46__or_module_6_res), .A2(
        n_majority7_module_46__or_module_9_res), .ZN(
        n_majority7_module_46__and_module_9_res) );
  OR2_X1 u_majority7_module_46__or_module_11_U1 ( .A1(
        n_majority7_module_46__or_module_10_res), .A2(
        n_majority7_module_46__and_module_8_res), .ZN(
        n_majority7_module_46__or_module_11_res) );
  AND2_X1 u_majority7_module_46__and_module_10_U1 ( .A1(
        n_majority7_module_46__or_module_8_res), .A2(
        n_majority7_module_46__and_module_9_res), .ZN(
        n_majority7_module_46__and_module_10_res) );
  AND2_X1 u_majority7_module_46__and_module_11_U1 ( .A1(
        n_majority7_module_46__and_module_10_res), .A2(
        n_majority7_module_46__or_module_11_res), .ZN(
        n_majority7_module_46_res) );
  DFF_X1 u_reg_module_47__cini_mul_v000_reg ( .D(n_majority7_module_46_res), 
        .CK(clock_5), .Q(n_reg_module_47_res), .QN() );
  AND2_X1 u_majority7_module_47__and_module_1_U1 ( .A1(n_xor_module_38_res), 
        .A2(n_xor_module_2_res), .ZN(n_majority7_module_47__and_module_1_res)
         );
  OR2_X1 u_majority7_module_47__or_module_1_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_38_res), .ZN(n_majority7_module_47__or_module_1_res) );
  AND2_X1 u_majority7_module_47__and_module_2_U1 ( .A1(n_xor_module_20_res), 
        .A2(n_xor_module_14_res), .ZN(n_majority7_module_47__and_module_2_res)
         );
  OR2_X1 u_majority7_module_47__or_module_2_U1 ( .A1(n_xor_module_14_res), 
        .A2(n_xor_module_20_res), .ZN(n_majority7_module_47__or_module_2_res)
         );
  AND2_X1 u_majority7_module_47__and_module_3_U1 ( .A1(n_xor_module_32_res), 
        .A2(n_xor_module_26_res), .ZN(n_majority7_module_47__and_module_3_res)
         );
  OR2_X1 u_majority7_module_47__or_module_3_U1 ( .A1(n_xor_module_26_res), 
        .A2(n_xor_module_32_res), .ZN(n_majority7_module_47__or_module_3_res)
         );
  AND2_X1 u_majority7_module_47__and_module_4_U1 ( .A1(
        n_majority7_module_47__and_module_2_res), .A2(
        n_majority7_module_47__and_module_1_res), .ZN(
        n_majority7_module_47__and_module_4_res) );
  OR2_X1 u_majority7_module_47__or_module_4_U1 ( .A1(
        n_majority7_module_47__and_module_1_res), .A2(
        n_majority7_module_47__and_module_2_res), .ZN(
        n_majority7_module_47__or_module_4_res) );
  AND2_X1 u_majority7_module_47__and_module_5_U1 ( .A1(
        n_majority7_module_47__and_module_3_res), .A2(n_xor_module_8_res), 
        .ZN(n_majority7_module_47__and_module_5_res) );
  OR2_X1 u_majority7_module_47__or_module_5_U1 ( .A1(n_xor_module_8_res), .A2(
        n_majority7_module_47__and_module_3_res), .ZN(
        n_majority7_module_47__or_module_5_res) );
  AND2_X1 u_majority7_module_47__and_module_6_U1 ( .A1(
        n_majority7_module_47__or_module_1_res), .A2(
        n_majority7_module_47__or_module_2_res), .ZN(
        n_majority7_module_47__and_module_6_res) );
  OR2_X1 u_majority7_module_47__or_module_6_U1 ( .A1(
        n_majority7_module_47__or_module_2_res), .A2(
        n_majority7_module_47__or_module_1_res), .ZN(
        n_majority7_module_47__or_module_6_res) );
  OR2_X1 u_majority7_module_47__or_module_7_U1 ( .A1(
        n_majority7_module_47__and_module_4_res), .A2(
        n_majority7_module_47__and_module_5_res), .ZN(
        n_majority7_module_47__or_module_7_res) );
  AND2_X1 u_majority7_module_47__and_module_7_U1 ( .A1(
        n_majority7_module_47__or_module_3_res), .A2(
        n_majority7_module_47__or_module_4_res), .ZN(
        n_majority7_module_47__and_module_7_res) );
  OR2_X1 u_majority7_module_47__or_module_8_U1 ( .A1(
        n_majority7_module_47__or_module_4_res), .A2(
        n_majority7_module_47__or_module_3_res), .ZN(
        n_majority7_module_47__or_module_8_res) );
  AND2_X1 u_majority7_module_47__and_module_8_U1 ( .A1(
        n_majority7_module_47__or_module_5_res), .A2(
        n_majority7_module_47__and_module_6_res), .ZN(
        n_majority7_module_47__and_module_8_res) );
  OR2_X1 u_majority7_module_47__or_module_9_U1 ( .A1(
        n_majority7_module_47__and_module_6_res), .A2(
        n_majority7_module_47__or_module_5_res), .ZN(
        n_majority7_module_47__or_module_9_res) );
  OR2_X1 u_majority7_module_47__or_module_10_U1 ( .A1(
        n_majority7_module_47__or_module_7_res), .A2(
        n_majority7_module_47__and_module_7_res), .ZN(
        n_majority7_module_47__or_module_10_res) );
  AND2_X1 u_majority7_module_47__and_module_9_U1 ( .A1(
        n_majority7_module_47__or_module_6_res), .A2(
        n_majority7_module_47__or_module_9_res), .ZN(
        n_majority7_module_47__and_module_9_res) );
  OR2_X1 u_majority7_module_47__or_module_11_U1 ( .A1(
        n_majority7_module_47__or_module_10_res), .A2(
        n_majority7_module_47__and_module_8_res), .ZN(
        n_majority7_module_47__or_module_11_res) );
  AND2_X1 u_majority7_module_47__and_module_10_U1 ( .A1(
        n_majority7_module_47__or_module_8_res), .A2(
        n_majority7_module_47__and_module_9_res), .ZN(
        n_majority7_module_47__and_module_10_res) );
  AND2_X1 u_majority7_module_47__and_module_11_U1 ( .A1(
        n_majority7_module_47__and_module_10_res), .A2(
        n_majority7_module_47__or_module_11_res), .ZN(
        n_majority7_module_47_res) );
  DFF_X1 u_reg_module_48__cini_mul_v000_reg ( .D(n_majority7_module_47_res), 
        .CK(clock_5), .Q(n_reg_module_48_res), .QN() );
  AND2_X1 u_majority7_module_48__and_module_1_U1 ( .A1(n_xor_module_40_res), 
        .A2(n_xor_module_4_res), .ZN(n_majority7_module_48__and_module_1_res)
         );
  OR2_X1 u_majority7_module_48__or_module_1_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_40_res), .ZN(n_majority7_module_48__or_module_1_res) );
  AND2_X1 u_majority7_module_48__and_module_2_U1 ( .A1(n_xor_module_22_res), 
        .A2(n_xor_module_16_res), .ZN(n_majority7_module_48__and_module_2_res)
         );
  OR2_X1 u_majority7_module_48__or_module_2_U1 ( .A1(n_xor_module_16_res), 
        .A2(n_xor_module_22_res), .ZN(n_majority7_module_48__or_module_2_res)
         );
  AND2_X1 u_majority7_module_48__and_module_3_U1 ( .A1(n_xor_module_34_res), 
        .A2(n_xor_module_28_res), .ZN(n_majority7_module_48__and_module_3_res)
         );
  OR2_X1 u_majority7_module_48__or_module_3_U1 ( .A1(n_xor_module_28_res), 
        .A2(n_xor_module_34_res), .ZN(n_majority7_module_48__or_module_3_res)
         );
  AND2_X1 u_majority7_module_48__and_module_4_U1 ( .A1(
        n_majority7_module_48__and_module_2_res), .A2(
        n_majority7_module_48__and_module_1_res), .ZN(
        n_majority7_module_48__and_module_4_res) );
  OR2_X1 u_majority7_module_48__or_module_4_U1 ( .A1(
        n_majority7_module_48__and_module_1_res), .A2(
        n_majority7_module_48__and_module_2_res), .ZN(
        n_majority7_module_48__or_module_4_res) );
  AND2_X1 u_majority7_module_48__and_module_5_U1 ( .A1(
        n_majority7_module_48__and_module_3_res), .A2(n_xor_module_10_res), 
        .ZN(n_majority7_module_48__and_module_5_res) );
  OR2_X1 u_majority7_module_48__or_module_5_U1 ( .A1(n_xor_module_10_res), 
        .A2(n_majority7_module_48__and_module_3_res), .ZN(
        n_majority7_module_48__or_module_5_res) );
  AND2_X1 u_majority7_module_48__and_module_6_U1 ( .A1(
        n_majority7_module_48__or_module_1_res), .A2(
        n_majority7_module_48__or_module_2_res), .ZN(
        n_majority7_module_48__and_module_6_res) );
  OR2_X1 u_majority7_module_48__or_module_6_U1 ( .A1(
        n_majority7_module_48__or_module_2_res), .A2(
        n_majority7_module_48__or_module_1_res), .ZN(
        n_majority7_module_48__or_module_6_res) );
  OR2_X1 u_majority7_module_48__or_module_7_U1 ( .A1(
        n_majority7_module_48__and_module_4_res), .A2(
        n_majority7_module_48__and_module_5_res), .ZN(
        n_majority7_module_48__or_module_7_res) );
  AND2_X1 u_majority7_module_48__and_module_7_U1 ( .A1(
        n_majority7_module_48__or_module_3_res), .A2(
        n_majority7_module_48__or_module_4_res), .ZN(
        n_majority7_module_48__and_module_7_res) );
  OR2_X1 u_majority7_module_48__or_module_8_U1 ( .A1(
        n_majority7_module_48__or_module_4_res), .A2(
        n_majority7_module_48__or_module_3_res), .ZN(
        n_majority7_module_48__or_module_8_res) );
  AND2_X1 u_majority7_module_48__and_module_8_U1 ( .A1(
        n_majority7_module_48__or_module_5_res), .A2(
        n_majority7_module_48__and_module_6_res), .ZN(
        n_majority7_module_48__and_module_8_res) );
  OR2_X1 u_majority7_module_48__or_module_9_U1 ( .A1(
        n_majority7_module_48__and_module_6_res), .A2(
        n_majority7_module_48__or_module_5_res), .ZN(
        n_majority7_module_48__or_module_9_res) );
  OR2_X1 u_majority7_module_48__or_module_10_U1 ( .A1(
        n_majority7_module_48__or_module_7_res), .A2(
        n_majority7_module_48__and_module_7_res), .ZN(
        n_majority7_module_48__or_module_10_res) );
  AND2_X1 u_majority7_module_48__and_module_9_U1 ( .A1(
        n_majority7_module_48__or_module_6_res), .A2(
        n_majority7_module_48__or_module_9_res), .ZN(
        n_majority7_module_48__and_module_9_res) );
  OR2_X1 u_majority7_module_48__or_module_11_U1 ( .A1(
        n_majority7_module_48__or_module_10_res), .A2(
        n_majority7_module_48__and_module_8_res), .ZN(
        n_majority7_module_48__or_module_11_res) );
  AND2_X1 u_majority7_module_48__and_module_10_U1 ( .A1(
        n_majority7_module_48__or_module_8_res), .A2(
        n_majority7_module_48__and_module_9_res), .ZN(
        n_majority7_module_48__and_module_10_res) );
  AND2_X1 u_majority7_module_48__and_module_11_U1 ( .A1(
        n_majority7_module_48__and_module_10_res), .A2(
        n_majority7_module_48__or_module_11_res), .ZN(
        n_majority7_module_48_res) );
  DFF_X1 u_reg_module_49__cini_mul_v000_reg ( .D(n_majority7_module_48_res), 
        .CK(clock_5), .Q(n_reg_module_49_res), .QN() );
  AND2_X1 u_majority7_module_49__and_module_1_U1 ( .A1(n_xor_module_40_res), 
        .A2(n_xor_module_4_res), .ZN(n_majority7_module_49__and_module_1_res)
         );
  OR2_X1 u_majority7_module_49__or_module_1_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_40_res), .ZN(n_majority7_module_49__or_module_1_res) );
  AND2_X1 u_majority7_module_49__and_module_2_U1 ( .A1(n_xor_module_22_res), 
        .A2(n_xor_module_16_res), .ZN(n_majority7_module_49__and_module_2_res)
         );
  OR2_X1 u_majority7_module_49__or_module_2_U1 ( .A1(n_xor_module_16_res), 
        .A2(n_xor_module_22_res), .ZN(n_majority7_module_49__or_module_2_res)
         );
  AND2_X1 u_majority7_module_49__and_module_3_U1 ( .A1(n_xor_module_34_res), 
        .A2(n_xor_module_28_res), .ZN(n_majority7_module_49__and_module_3_res)
         );
  OR2_X1 u_majority7_module_49__or_module_3_U1 ( .A1(n_xor_module_28_res), 
        .A2(n_xor_module_34_res), .ZN(n_majority7_module_49__or_module_3_res)
         );
  AND2_X1 u_majority7_module_49__and_module_4_U1 ( .A1(
        n_majority7_module_49__and_module_2_res), .A2(
        n_majority7_module_49__and_module_1_res), .ZN(
        n_majority7_module_49__and_module_4_res) );
  OR2_X1 u_majority7_module_49__or_module_4_U1 ( .A1(
        n_majority7_module_49__and_module_1_res), .A2(
        n_majority7_module_49__and_module_2_res), .ZN(
        n_majority7_module_49__or_module_4_res) );
  AND2_X1 u_majority7_module_49__and_module_5_U1 ( .A1(
        n_majority7_module_49__and_module_3_res), .A2(n_xor_module_10_res), 
        .ZN(n_majority7_module_49__and_module_5_res) );
  OR2_X1 u_majority7_module_49__or_module_5_U1 ( .A1(n_xor_module_10_res), 
        .A2(n_majority7_module_49__and_module_3_res), .ZN(
        n_majority7_module_49__or_module_5_res) );
  AND2_X1 u_majority7_module_49__and_module_6_U1 ( .A1(
        n_majority7_module_49__or_module_1_res), .A2(
        n_majority7_module_49__or_module_2_res), .ZN(
        n_majority7_module_49__and_module_6_res) );
  OR2_X1 u_majority7_module_49__or_module_6_U1 ( .A1(
        n_majority7_module_49__or_module_2_res), .A2(
        n_majority7_module_49__or_module_1_res), .ZN(
        n_majority7_module_49__or_module_6_res) );
  OR2_X1 u_majority7_module_49__or_module_7_U1 ( .A1(
        n_majority7_module_49__and_module_4_res), .A2(
        n_majority7_module_49__and_module_5_res), .ZN(
        n_majority7_module_49__or_module_7_res) );
  AND2_X1 u_majority7_module_49__and_module_7_U1 ( .A1(
        n_majority7_module_49__or_module_3_res), .A2(
        n_majority7_module_49__or_module_4_res), .ZN(
        n_majority7_module_49__and_module_7_res) );
  OR2_X1 u_majority7_module_49__or_module_8_U1 ( .A1(
        n_majority7_module_49__or_module_4_res), .A2(
        n_majority7_module_49__or_module_3_res), .ZN(
        n_majority7_module_49__or_module_8_res) );
  AND2_X1 u_majority7_module_49__and_module_8_U1 ( .A1(
        n_majority7_module_49__or_module_5_res), .A2(
        n_majority7_module_49__and_module_6_res), .ZN(
        n_majority7_module_49__and_module_8_res) );
  OR2_X1 u_majority7_module_49__or_module_9_U1 ( .A1(
        n_majority7_module_49__and_module_6_res), .A2(
        n_majority7_module_49__or_module_5_res), .ZN(
        n_majority7_module_49__or_module_9_res) );
  OR2_X1 u_majority7_module_49__or_module_10_U1 ( .A1(
        n_majority7_module_49__or_module_7_res), .A2(
        n_majority7_module_49__and_module_7_res), .ZN(
        n_majority7_module_49__or_module_10_res) );
  AND2_X1 u_majority7_module_49__and_module_9_U1 ( .A1(
        n_majority7_module_49__or_module_6_res), .A2(
        n_majority7_module_49__or_module_9_res), .ZN(
        n_majority7_module_49__and_module_9_res) );
  OR2_X1 u_majority7_module_49__or_module_11_U1 ( .A1(
        n_majority7_module_49__or_module_10_res), .A2(
        n_majority7_module_49__and_module_8_res), .ZN(
        n_majority7_module_49__or_module_11_res) );
  AND2_X1 u_majority7_module_49__and_module_10_U1 ( .A1(
        n_majority7_module_49__or_module_8_res), .A2(
        n_majority7_module_49__and_module_9_res), .ZN(
        n_majority7_module_49__and_module_10_res) );
  AND2_X1 u_majority7_module_49__and_module_11_U1 ( .A1(
        n_majority7_module_49__and_module_10_res), .A2(
        n_majority7_module_49__or_module_11_res), .ZN(
        n_majority7_module_49_res) );
  DFF_X1 u_reg_module_50__cini_mul_v000_reg ( .D(n_majority7_module_49_res), 
        .CK(clock_5), .Q(n_reg_module_50_res), .QN() );
  AND2_X1 u_majority7_module_50__and_module_1_U1 ( .A1(n_xor_module_40_res), 
        .A2(n_xor_module_4_res), .ZN(n_majority7_module_50__and_module_1_res)
         );
  OR2_X1 u_majority7_module_50__or_module_1_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_40_res), .ZN(n_majority7_module_50__or_module_1_res) );
  AND2_X1 u_majority7_module_50__and_module_2_U1 ( .A1(n_xor_module_22_res), 
        .A2(n_xor_module_16_res), .ZN(n_majority7_module_50__and_module_2_res)
         );
  OR2_X1 u_majority7_module_50__or_module_2_U1 ( .A1(n_xor_module_16_res), 
        .A2(n_xor_module_22_res), .ZN(n_majority7_module_50__or_module_2_res)
         );
  AND2_X1 u_majority7_module_50__and_module_3_U1 ( .A1(n_xor_module_34_res), 
        .A2(n_xor_module_28_res), .ZN(n_majority7_module_50__and_module_3_res)
         );
  OR2_X1 u_majority7_module_50__or_module_3_U1 ( .A1(n_xor_module_28_res), 
        .A2(n_xor_module_34_res), .ZN(n_majority7_module_50__or_module_3_res)
         );
  AND2_X1 u_majority7_module_50__and_module_4_U1 ( .A1(
        n_majority7_module_50__and_module_2_res), .A2(
        n_majority7_module_50__and_module_1_res), .ZN(
        n_majority7_module_50__and_module_4_res) );
  OR2_X1 u_majority7_module_50__or_module_4_U1 ( .A1(
        n_majority7_module_50__and_module_1_res), .A2(
        n_majority7_module_50__and_module_2_res), .ZN(
        n_majority7_module_50__or_module_4_res) );
  AND2_X1 u_majority7_module_50__and_module_5_U1 ( .A1(
        n_majority7_module_50__and_module_3_res), .A2(n_xor_module_10_res), 
        .ZN(n_majority7_module_50__and_module_5_res) );
  OR2_X1 u_majority7_module_50__or_module_5_U1 ( .A1(n_xor_module_10_res), 
        .A2(n_majority7_module_50__and_module_3_res), .ZN(
        n_majority7_module_50__or_module_5_res) );
  AND2_X1 u_majority7_module_50__and_module_6_U1 ( .A1(
        n_majority7_module_50__or_module_1_res), .A2(
        n_majority7_module_50__or_module_2_res), .ZN(
        n_majority7_module_50__and_module_6_res) );
  OR2_X1 u_majority7_module_50__or_module_6_U1 ( .A1(
        n_majority7_module_50__or_module_2_res), .A2(
        n_majority7_module_50__or_module_1_res), .ZN(
        n_majority7_module_50__or_module_6_res) );
  OR2_X1 u_majority7_module_50__or_module_7_U1 ( .A1(
        n_majority7_module_50__and_module_4_res), .A2(
        n_majority7_module_50__and_module_5_res), .ZN(
        n_majority7_module_50__or_module_7_res) );
  AND2_X1 u_majority7_module_50__and_module_7_U1 ( .A1(
        n_majority7_module_50__or_module_3_res), .A2(
        n_majority7_module_50__or_module_4_res), .ZN(
        n_majority7_module_50__and_module_7_res) );
  OR2_X1 u_majority7_module_50__or_module_8_U1 ( .A1(
        n_majority7_module_50__or_module_4_res), .A2(
        n_majority7_module_50__or_module_3_res), .ZN(
        n_majority7_module_50__or_module_8_res) );
  AND2_X1 u_majority7_module_50__and_module_8_U1 ( .A1(
        n_majority7_module_50__or_module_5_res), .A2(
        n_majority7_module_50__and_module_6_res), .ZN(
        n_majority7_module_50__and_module_8_res) );
  OR2_X1 u_majority7_module_50__or_module_9_U1 ( .A1(
        n_majority7_module_50__and_module_6_res), .A2(
        n_majority7_module_50__or_module_5_res), .ZN(
        n_majority7_module_50__or_module_9_res) );
  OR2_X1 u_majority7_module_50__or_module_10_U1 ( .A1(
        n_majority7_module_50__or_module_7_res), .A2(
        n_majority7_module_50__and_module_7_res), .ZN(
        n_majority7_module_50__or_module_10_res) );
  AND2_X1 u_majority7_module_50__and_module_9_U1 ( .A1(
        n_majority7_module_50__or_module_6_res), .A2(
        n_majority7_module_50__or_module_9_res), .ZN(
        n_majority7_module_50__and_module_9_res) );
  OR2_X1 u_majority7_module_50__or_module_11_U1 ( .A1(
        n_majority7_module_50__or_module_10_res), .A2(
        n_majority7_module_50__and_module_8_res), .ZN(
        n_majority7_module_50__or_module_11_res) );
  AND2_X1 u_majority7_module_50__and_module_10_U1 ( .A1(
        n_majority7_module_50__or_module_8_res), .A2(
        n_majority7_module_50__and_module_9_res), .ZN(
        n_majority7_module_50__and_module_10_res) );
  AND2_X1 u_majority7_module_50__and_module_11_U1 ( .A1(
        n_majority7_module_50__and_module_10_res), .A2(
        n_majority7_module_50__or_module_11_res), .ZN(
        n_majority7_module_50_res) );
  DFF_X1 u_reg_module_51__cini_mul_v000_reg ( .D(n_majority7_module_50_res), 
        .CK(clock_5), .Q(n_reg_module_51_res), .QN() );
  AND2_X1 u_majority7_module_51__and_module_1_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_51__and_module_1_res)
         );
  OR2_X1 u_majority7_module_51__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_51__or_module_1_res) );
  AND2_X1 u_majority7_module_51__and_module_2_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_xor_module_18_res), .ZN(n_majority7_module_51__and_module_2_res)
         );
  OR2_X1 u_majority7_module_51__or_module_2_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_xor_module_24_res), .ZN(n_majority7_module_51__or_module_2_res)
         );
  AND2_X1 u_majority7_module_51__and_module_3_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_51__and_module_3_res)
         );
  OR2_X1 u_majority7_module_51__or_module_3_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_51__or_module_3_res)
         );
  AND2_X1 u_majority7_module_51__and_module_4_U1 ( .A1(
        n_majority7_module_51__and_module_2_res), .A2(
        n_majority7_module_51__and_module_1_res), .ZN(
        n_majority7_module_51__and_module_4_res) );
  OR2_X1 u_majority7_module_51__or_module_4_U1 ( .A1(
        n_majority7_module_51__and_module_1_res), .A2(
        n_majority7_module_51__and_module_2_res), .ZN(
        n_majority7_module_51__or_module_4_res) );
  AND2_X1 u_majority7_module_51__and_module_5_U1 ( .A1(
        n_majority7_module_51__and_module_3_res), .A2(n_xor_module_12_res), 
        .ZN(n_majority7_module_51__and_module_5_res) );
  OR2_X1 u_majority7_module_51__or_module_5_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_majority7_module_51__and_module_3_res), .ZN(
        n_majority7_module_51__or_module_5_res) );
  AND2_X1 u_majority7_module_51__and_module_6_U1 ( .A1(
        n_majority7_module_51__or_module_1_res), .A2(
        n_majority7_module_51__or_module_2_res), .ZN(
        n_majority7_module_51__and_module_6_res) );
  OR2_X1 u_majority7_module_51__or_module_6_U1 ( .A1(
        n_majority7_module_51__or_module_2_res), .A2(
        n_majority7_module_51__or_module_1_res), .ZN(
        n_majority7_module_51__or_module_6_res) );
  OR2_X1 u_majority7_module_51__or_module_7_U1 ( .A1(
        n_majority7_module_51__and_module_4_res), .A2(
        n_majority7_module_51__and_module_5_res), .ZN(
        n_majority7_module_51__or_module_7_res) );
  AND2_X1 u_majority7_module_51__and_module_7_U1 ( .A1(
        n_majority7_module_51__or_module_3_res), .A2(
        n_majority7_module_51__or_module_4_res), .ZN(
        n_majority7_module_51__and_module_7_res) );
  OR2_X1 u_majority7_module_51__or_module_8_U1 ( .A1(
        n_majority7_module_51__or_module_4_res), .A2(
        n_majority7_module_51__or_module_3_res), .ZN(
        n_majority7_module_51__or_module_8_res) );
  AND2_X1 u_majority7_module_51__and_module_8_U1 ( .A1(
        n_majority7_module_51__or_module_5_res), .A2(
        n_majority7_module_51__and_module_6_res), .ZN(
        n_majority7_module_51__and_module_8_res) );
  OR2_X1 u_majority7_module_51__or_module_9_U1 ( .A1(
        n_majority7_module_51__and_module_6_res), .A2(
        n_majority7_module_51__or_module_5_res), .ZN(
        n_majority7_module_51__or_module_9_res) );
  OR2_X1 u_majority7_module_51__or_module_10_U1 ( .A1(
        n_majority7_module_51__or_module_7_res), .A2(
        n_majority7_module_51__and_module_7_res), .ZN(
        n_majority7_module_51__or_module_10_res) );
  AND2_X1 u_majority7_module_51__and_module_9_U1 ( .A1(
        n_majority7_module_51__or_module_6_res), .A2(
        n_majority7_module_51__or_module_9_res), .ZN(
        n_majority7_module_51__and_module_9_res) );
  OR2_X1 u_majority7_module_51__or_module_11_U1 ( .A1(
        n_majority7_module_51__or_module_10_res), .A2(
        n_majority7_module_51__and_module_8_res), .ZN(
        n_majority7_module_51__or_module_11_res) );
  AND2_X1 u_majority7_module_51__and_module_10_U1 ( .A1(
        n_majority7_module_51__or_module_8_res), .A2(
        n_majority7_module_51__and_module_9_res), .ZN(
        n_majority7_module_51__and_module_10_res) );
  AND2_X1 u_majority7_module_51__and_module_11_U1 ( .A1(
        n_majority7_module_51__and_module_10_res), .A2(
        n_majority7_module_51__or_module_11_res), .ZN(
        n_majority7_module_51_res) );
  DFF_X1 u_reg_module_52__cini_mul_v000_reg ( .D(n_majority7_module_51_res), 
        .CK(clock_5), .Q(n_reg_module_52_res), .QN() );
  AND2_X1 u_majority7_module_52__and_module_1_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_52__and_module_1_res)
         );
  OR2_X1 u_majority7_module_52__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_52__or_module_1_res) );
  AND2_X1 u_majority7_module_52__and_module_2_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_xor_module_18_res), .ZN(n_majority7_module_52__and_module_2_res)
         );
  OR2_X1 u_majority7_module_52__or_module_2_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_xor_module_24_res), .ZN(n_majority7_module_52__or_module_2_res)
         );
  AND2_X1 u_majority7_module_52__and_module_3_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_52__and_module_3_res)
         );
  OR2_X1 u_majority7_module_52__or_module_3_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_52__or_module_3_res)
         );
  AND2_X1 u_majority7_module_52__and_module_4_U1 ( .A1(
        n_majority7_module_52__and_module_2_res), .A2(
        n_majority7_module_52__and_module_1_res), .ZN(
        n_majority7_module_52__and_module_4_res) );
  OR2_X1 u_majority7_module_52__or_module_4_U1 ( .A1(
        n_majority7_module_52__and_module_1_res), .A2(
        n_majority7_module_52__and_module_2_res), .ZN(
        n_majority7_module_52__or_module_4_res) );
  AND2_X1 u_majority7_module_52__and_module_5_U1 ( .A1(
        n_majority7_module_52__and_module_3_res), .A2(n_xor_module_12_res), 
        .ZN(n_majority7_module_52__and_module_5_res) );
  OR2_X1 u_majority7_module_52__or_module_5_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_majority7_module_52__and_module_3_res), .ZN(
        n_majority7_module_52__or_module_5_res) );
  AND2_X1 u_majority7_module_52__and_module_6_U1 ( .A1(
        n_majority7_module_52__or_module_1_res), .A2(
        n_majority7_module_52__or_module_2_res), .ZN(
        n_majority7_module_52__and_module_6_res) );
  OR2_X1 u_majority7_module_52__or_module_6_U1 ( .A1(
        n_majority7_module_52__or_module_2_res), .A2(
        n_majority7_module_52__or_module_1_res), .ZN(
        n_majority7_module_52__or_module_6_res) );
  OR2_X1 u_majority7_module_52__or_module_7_U1 ( .A1(
        n_majority7_module_52__and_module_4_res), .A2(
        n_majority7_module_52__and_module_5_res), .ZN(
        n_majority7_module_52__or_module_7_res) );
  AND2_X1 u_majority7_module_52__and_module_7_U1 ( .A1(
        n_majority7_module_52__or_module_3_res), .A2(
        n_majority7_module_52__or_module_4_res), .ZN(
        n_majority7_module_52__and_module_7_res) );
  OR2_X1 u_majority7_module_52__or_module_8_U1 ( .A1(
        n_majority7_module_52__or_module_4_res), .A2(
        n_majority7_module_52__or_module_3_res), .ZN(
        n_majority7_module_52__or_module_8_res) );
  AND2_X1 u_majority7_module_52__and_module_8_U1 ( .A1(
        n_majority7_module_52__or_module_5_res), .A2(
        n_majority7_module_52__and_module_6_res), .ZN(
        n_majority7_module_52__and_module_8_res) );
  OR2_X1 u_majority7_module_52__or_module_9_U1 ( .A1(
        n_majority7_module_52__and_module_6_res), .A2(
        n_majority7_module_52__or_module_5_res), .ZN(
        n_majority7_module_52__or_module_9_res) );
  OR2_X1 u_majority7_module_52__or_module_10_U1 ( .A1(
        n_majority7_module_52__or_module_7_res), .A2(
        n_majority7_module_52__and_module_7_res), .ZN(
        n_majority7_module_52__or_module_10_res) );
  AND2_X1 u_majority7_module_52__and_module_9_U1 ( .A1(
        n_majority7_module_52__or_module_6_res), .A2(
        n_majority7_module_52__or_module_9_res), .ZN(
        n_majority7_module_52__and_module_9_res) );
  OR2_X1 u_majority7_module_52__or_module_11_U1 ( .A1(
        n_majority7_module_52__or_module_10_res), .A2(
        n_majority7_module_52__and_module_8_res), .ZN(
        n_majority7_module_52__or_module_11_res) );
  AND2_X1 u_majority7_module_52__and_module_10_U1 ( .A1(
        n_majority7_module_52__or_module_8_res), .A2(
        n_majority7_module_52__and_module_9_res), .ZN(
        n_majority7_module_52__and_module_10_res) );
  AND2_X1 u_majority7_module_52__and_module_11_U1 ( .A1(
        n_majority7_module_52__and_module_10_res), .A2(
        n_majority7_module_52__or_module_11_res), .ZN(
        n_majority7_module_52_res) );
  DFF_X1 u_reg_module_53__cini_mul_v000_reg ( .D(n_majority7_module_52_res), 
        .CK(clock_5), .Q(n_reg_module_53_res), .QN() );
  AND2_X1 u_majority7_module_53__and_module_1_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_53__and_module_1_res)
         );
  OR2_X1 u_majority7_module_53__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_53__or_module_1_res) );
  AND2_X1 u_majority7_module_53__and_module_2_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_xor_module_18_res), .ZN(n_majority7_module_53__and_module_2_res)
         );
  OR2_X1 u_majority7_module_53__or_module_2_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_xor_module_24_res), .ZN(n_majority7_module_53__or_module_2_res)
         );
  AND2_X1 u_majority7_module_53__and_module_3_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_53__and_module_3_res)
         );
  OR2_X1 u_majority7_module_53__or_module_3_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_53__or_module_3_res)
         );
  AND2_X1 u_majority7_module_53__and_module_4_U1 ( .A1(
        n_majority7_module_53__and_module_2_res), .A2(
        n_majority7_module_53__and_module_1_res), .ZN(
        n_majority7_module_53__and_module_4_res) );
  OR2_X1 u_majority7_module_53__or_module_4_U1 ( .A1(
        n_majority7_module_53__and_module_1_res), .A2(
        n_majority7_module_53__and_module_2_res), .ZN(
        n_majority7_module_53__or_module_4_res) );
  AND2_X1 u_majority7_module_53__and_module_5_U1 ( .A1(
        n_majority7_module_53__and_module_3_res), .A2(n_xor_module_12_res), 
        .ZN(n_majority7_module_53__and_module_5_res) );
  OR2_X1 u_majority7_module_53__or_module_5_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_majority7_module_53__and_module_3_res), .ZN(
        n_majority7_module_53__or_module_5_res) );
  AND2_X1 u_majority7_module_53__and_module_6_U1 ( .A1(
        n_majority7_module_53__or_module_1_res), .A2(
        n_majority7_module_53__or_module_2_res), .ZN(
        n_majority7_module_53__and_module_6_res) );
  OR2_X1 u_majority7_module_53__or_module_6_U1 ( .A1(
        n_majority7_module_53__or_module_2_res), .A2(
        n_majority7_module_53__or_module_1_res), .ZN(
        n_majority7_module_53__or_module_6_res) );
  OR2_X1 u_majority7_module_53__or_module_7_U1 ( .A1(
        n_majority7_module_53__and_module_4_res), .A2(
        n_majority7_module_53__and_module_5_res), .ZN(
        n_majority7_module_53__or_module_7_res) );
  AND2_X1 u_majority7_module_53__and_module_7_U1 ( .A1(
        n_majority7_module_53__or_module_3_res), .A2(
        n_majority7_module_53__or_module_4_res), .ZN(
        n_majority7_module_53__and_module_7_res) );
  OR2_X1 u_majority7_module_53__or_module_8_U1 ( .A1(
        n_majority7_module_53__or_module_4_res), .A2(
        n_majority7_module_53__or_module_3_res), .ZN(
        n_majority7_module_53__or_module_8_res) );
  AND2_X1 u_majority7_module_53__and_module_8_U1 ( .A1(
        n_majority7_module_53__or_module_5_res), .A2(
        n_majority7_module_53__and_module_6_res), .ZN(
        n_majority7_module_53__and_module_8_res) );
  OR2_X1 u_majority7_module_53__or_module_9_U1 ( .A1(
        n_majority7_module_53__and_module_6_res), .A2(
        n_majority7_module_53__or_module_5_res), .ZN(
        n_majority7_module_53__or_module_9_res) );
  OR2_X1 u_majority7_module_53__or_module_10_U1 ( .A1(
        n_majority7_module_53__or_module_7_res), .A2(
        n_majority7_module_53__and_module_7_res), .ZN(
        n_majority7_module_53__or_module_10_res) );
  AND2_X1 u_majority7_module_53__and_module_9_U1 ( .A1(
        n_majority7_module_53__or_module_6_res), .A2(
        n_majority7_module_53__or_module_9_res), .ZN(
        n_majority7_module_53__and_module_9_res) );
  OR2_X1 u_majority7_module_53__or_module_11_U1 ( .A1(
        n_majority7_module_53__or_module_10_res), .A2(
        n_majority7_module_53__and_module_8_res), .ZN(
        n_majority7_module_53__or_module_11_res) );
  AND2_X1 u_majority7_module_53__and_module_10_U1 ( .A1(
        n_majority7_module_53__or_module_8_res), .A2(
        n_majority7_module_53__and_module_9_res), .ZN(
        n_majority7_module_53__and_module_10_res) );
  AND2_X1 u_majority7_module_53__and_module_11_U1 ( .A1(
        n_majority7_module_53__and_module_10_res), .A2(
        n_majority7_module_53__or_module_11_res), .ZN(
        n_majority7_module_53_res) );
  DFF_X1 u_reg_module_54__cini_mul_v000_reg ( .D(n_majority7_module_53_res), 
        .CK(clock_5), .Q(n_reg_module_54_res), .QN() );
  AND2_X1 u_majority7_module_54__and_module_1_U1 ( .A1(n_xor_module_38_res), 
        .A2(n_xor_module_2_res), .ZN(n_majority7_module_54__and_module_1_res)
         );
  OR2_X1 u_majority7_module_54__or_module_1_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_38_res), .ZN(n_majority7_module_54__or_module_1_res) );
  AND2_X1 u_majority7_module_54__and_module_2_U1 ( .A1(n_xor_module_20_res), 
        .A2(n_xor_module_14_res), .ZN(n_majority7_module_54__and_module_2_res)
         );
  OR2_X1 u_majority7_module_54__or_module_2_U1 ( .A1(n_xor_module_14_res), 
        .A2(n_xor_module_20_res), .ZN(n_majority7_module_54__or_module_2_res)
         );
  AND2_X1 u_majority7_module_54__and_module_3_U1 ( .A1(n_xor_module_32_res), 
        .A2(n_xor_module_26_res), .ZN(n_majority7_module_54__and_module_3_res)
         );
  OR2_X1 u_majority7_module_54__or_module_3_U1 ( .A1(n_xor_module_26_res), 
        .A2(n_xor_module_32_res), .ZN(n_majority7_module_54__or_module_3_res)
         );
  AND2_X1 u_majority7_module_54__and_module_4_U1 ( .A1(
        n_majority7_module_54__and_module_2_res), .A2(
        n_majority7_module_54__and_module_1_res), .ZN(
        n_majority7_module_54__and_module_4_res) );
  OR2_X1 u_majority7_module_54__or_module_4_U1 ( .A1(
        n_majority7_module_54__and_module_1_res), .A2(
        n_majority7_module_54__and_module_2_res), .ZN(
        n_majority7_module_54__or_module_4_res) );
  AND2_X1 u_majority7_module_54__and_module_5_U1 ( .A1(
        n_majority7_module_54__and_module_3_res), .A2(n_xor_module_8_res), 
        .ZN(n_majority7_module_54__and_module_5_res) );
  OR2_X1 u_majority7_module_54__or_module_5_U1 ( .A1(n_xor_module_8_res), .A2(
        n_majority7_module_54__and_module_3_res), .ZN(
        n_majority7_module_54__or_module_5_res) );
  AND2_X1 u_majority7_module_54__and_module_6_U1 ( .A1(
        n_majority7_module_54__or_module_1_res), .A2(
        n_majority7_module_54__or_module_2_res), .ZN(
        n_majority7_module_54__and_module_6_res) );
  OR2_X1 u_majority7_module_54__or_module_6_U1 ( .A1(
        n_majority7_module_54__or_module_2_res), .A2(
        n_majority7_module_54__or_module_1_res), .ZN(
        n_majority7_module_54__or_module_6_res) );
  OR2_X1 u_majority7_module_54__or_module_7_U1 ( .A1(
        n_majority7_module_54__and_module_4_res), .A2(
        n_majority7_module_54__and_module_5_res), .ZN(
        n_majority7_module_54__or_module_7_res) );
  AND2_X1 u_majority7_module_54__and_module_7_U1 ( .A1(
        n_majority7_module_54__or_module_3_res), .A2(
        n_majority7_module_54__or_module_4_res), .ZN(
        n_majority7_module_54__and_module_7_res) );
  OR2_X1 u_majority7_module_54__or_module_8_U1 ( .A1(
        n_majority7_module_54__or_module_4_res), .A2(
        n_majority7_module_54__or_module_3_res), .ZN(
        n_majority7_module_54__or_module_8_res) );
  AND2_X1 u_majority7_module_54__and_module_8_U1 ( .A1(
        n_majority7_module_54__or_module_5_res), .A2(
        n_majority7_module_54__and_module_6_res), .ZN(
        n_majority7_module_54__and_module_8_res) );
  OR2_X1 u_majority7_module_54__or_module_9_U1 ( .A1(
        n_majority7_module_54__and_module_6_res), .A2(
        n_majority7_module_54__or_module_5_res), .ZN(
        n_majority7_module_54__or_module_9_res) );
  OR2_X1 u_majority7_module_54__or_module_10_U1 ( .A1(
        n_majority7_module_54__or_module_7_res), .A2(
        n_majority7_module_54__and_module_7_res), .ZN(
        n_majority7_module_54__or_module_10_res) );
  AND2_X1 u_majority7_module_54__and_module_9_U1 ( .A1(
        n_majority7_module_54__or_module_6_res), .A2(
        n_majority7_module_54__or_module_9_res), .ZN(
        n_majority7_module_54__and_module_9_res) );
  OR2_X1 u_majority7_module_54__or_module_11_U1 ( .A1(
        n_majority7_module_54__or_module_10_res), .A2(
        n_majority7_module_54__and_module_8_res), .ZN(
        n_majority7_module_54__or_module_11_res) );
  AND2_X1 u_majority7_module_54__and_module_10_U1 ( .A1(
        n_majority7_module_54__or_module_8_res), .A2(
        n_majority7_module_54__and_module_9_res), .ZN(
        n_majority7_module_54__and_module_10_res) );
  AND2_X1 u_majority7_module_54__and_module_11_U1 ( .A1(
        n_majority7_module_54__and_module_10_res), .A2(
        n_majority7_module_54__or_module_11_res), .ZN(
        n_majority7_module_54_res) );
  DFF_X1 u_reg_module_55__cini_mul_v000_reg ( .D(n_majority7_module_54_res), 
        .CK(clock_6), .Q(n_reg_module_55_res), .QN() );
  AND2_X1 u_majority7_module_55__and_module_1_U1 ( .A1(n_xor_module_38_res), 
        .A2(n_xor_module_2_res), .ZN(n_majority7_module_55__and_module_1_res)
         );
  OR2_X1 u_majority7_module_55__or_module_1_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_38_res), .ZN(n_majority7_module_55__or_module_1_res) );
  AND2_X1 u_majority7_module_55__and_module_2_U1 ( .A1(n_xor_module_20_res), 
        .A2(n_xor_module_14_res), .ZN(n_majority7_module_55__and_module_2_res)
         );
  OR2_X1 u_majority7_module_55__or_module_2_U1 ( .A1(n_xor_module_14_res), 
        .A2(n_xor_module_20_res), .ZN(n_majority7_module_55__or_module_2_res)
         );
  AND2_X1 u_majority7_module_55__and_module_3_U1 ( .A1(n_xor_module_32_res), 
        .A2(n_xor_module_26_res), .ZN(n_majority7_module_55__and_module_3_res)
         );
  OR2_X1 u_majority7_module_55__or_module_3_U1 ( .A1(n_xor_module_26_res), 
        .A2(n_xor_module_32_res), .ZN(n_majority7_module_55__or_module_3_res)
         );
  AND2_X1 u_majority7_module_55__and_module_4_U1 ( .A1(
        n_majority7_module_55__and_module_2_res), .A2(
        n_majority7_module_55__and_module_1_res), .ZN(
        n_majority7_module_55__and_module_4_res) );
  OR2_X1 u_majority7_module_55__or_module_4_U1 ( .A1(
        n_majority7_module_55__and_module_1_res), .A2(
        n_majority7_module_55__and_module_2_res), .ZN(
        n_majority7_module_55__or_module_4_res) );
  AND2_X1 u_majority7_module_55__and_module_5_U1 ( .A1(
        n_majority7_module_55__and_module_3_res), .A2(n_xor_module_8_res), 
        .ZN(n_majority7_module_55__and_module_5_res) );
  OR2_X1 u_majority7_module_55__or_module_5_U1 ( .A1(n_xor_module_8_res), .A2(
        n_majority7_module_55__and_module_3_res), .ZN(
        n_majority7_module_55__or_module_5_res) );
  AND2_X1 u_majority7_module_55__and_module_6_U1 ( .A1(
        n_majority7_module_55__or_module_1_res), .A2(
        n_majority7_module_55__or_module_2_res), .ZN(
        n_majority7_module_55__and_module_6_res) );
  OR2_X1 u_majority7_module_55__or_module_6_U1 ( .A1(
        n_majority7_module_55__or_module_2_res), .A2(
        n_majority7_module_55__or_module_1_res), .ZN(
        n_majority7_module_55__or_module_6_res) );
  OR2_X1 u_majority7_module_55__or_module_7_U1 ( .A1(
        n_majority7_module_55__and_module_4_res), .A2(
        n_majority7_module_55__and_module_5_res), .ZN(
        n_majority7_module_55__or_module_7_res) );
  AND2_X1 u_majority7_module_55__and_module_7_U1 ( .A1(
        n_majority7_module_55__or_module_3_res), .A2(
        n_majority7_module_55__or_module_4_res), .ZN(
        n_majority7_module_55__and_module_7_res) );
  OR2_X1 u_majority7_module_55__or_module_8_U1 ( .A1(
        n_majority7_module_55__or_module_4_res), .A2(
        n_majority7_module_55__or_module_3_res), .ZN(
        n_majority7_module_55__or_module_8_res) );
  AND2_X1 u_majority7_module_55__and_module_8_U1 ( .A1(
        n_majority7_module_55__or_module_5_res), .A2(
        n_majority7_module_55__and_module_6_res), .ZN(
        n_majority7_module_55__and_module_8_res) );
  OR2_X1 u_majority7_module_55__or_module_9_U1 ( .A1(
        n_majority7_module_55__and_module_6_res), .A2(
        n_majority7_module_55__or_module_5_res), .ZN(
        n_majority7_module_55__or_module_9_res) );
  OR2_X1 u_majority7_module_55__or_module_10_U1 ( .A1(
        n_majority7_module_55__or_module_7_res), .A2(
        n_majority7_module_55__and_module_7_res), .ZN(
        n_majority7_module_55__or_module_10_res) );
  AND2_X1 u_majority7_module_55__and_module_9_U1 ( .A1(
        n_majority7_module_55__or_module_6_res), .A2(
        n_majority7_module_55__or_module_9_res), .ZN(
        n_majority7_module_55__and_module_9_res) );
  OR2_X1 u_majority7_module_55__or_module_11_U1 ( .A1(
        n_majority7_module_55__or_module_10_res), .A2(
        n_majority7_module_55__and_module_8_res), .ZN(
        n_majority7_module_55__or_module_11_res) );
  AND2_X1 u_majority7_module_55__and_module_10_U1 ( .A1(
        n_majority7_module_55__or_module_8_res), .A2(
        n_majority7_module_55__and_module_9_res), .ZN(
        n_majority7_module_55__and_module_10_res) );
  AND2_X1 u_majority7_module_55__and_module_11_U1 ( .A1(
        n_majority7_module_55__and_module_10_res), .A2(
        n_majority7_module_55__or_module_11_res), .ZN(
        n_majority7_module_55_res) );
  DFF_X1 u_reg_module_56__cini_mul_v000_reg ( .D(n_majority7_module_55_res), 
        .CK(clock_6), .Q(n_reg_module_56_res), .QN() );
  AND2_X1 u_majority7_module_56__and_module_1_U1 ( .A1(n_xor_module_38_res), 
        .A2(n_xor_module_2_res), .ZN(n_majority7_module_56__and_module_1_res)
         );
  OR2_X1 u_majority7_module_56__or_module_1_U1 ( .A1(n_xor_module_2_res), .A2(
        n_xor_module_38_res), .ZN(n_majority7_module_56__or_module_1_res) );
  AND2_X1 u_majority7_module_56__and_module_2_U1 ( .A1(n_xor_module_20_res), 
        .A2(n_xor_module_14_res), .ZN(n_majority7_module_56__and_module_2_res)
         );
  OR2_X1 u_majority7_module_56__or_module_2_U1 ( .A1(n_xor_module_14_res), 
        .A2(n_xor_module_20_res), .ZN(n_majority7_module_56__or_module_2_res)
         );
  AND2_X1 u_majority7_module_56__and_module_3_U1 ( .A1(n_xor_module_32_res), 
        .A2(n_xor_module_26_res), .ZN(n_majority7_module_56__and_module_3_res)
         );
  OR2_X1 u_majority7_module_56__or_module_3_U1 ( .A1(n_xor_module_26_res), 
        .A2(n_xor_module_32_res), .ZN(n_majority7_module_56__or_module_3_res)
         );
  AND2_X1 u_majority7_module_56__and_module_4_U1 ( .A1(
        n_majority7_module_56__and_module_2_res), .A2(
        n_majority7_module_56__and_module_1_res), .ZN(
        n_majority7_module_56__and_module_4_res) );
  OR2_X1 u_majority7_module_56__or_module_4_U1 ( .A1(
        n_majority7_module_56__and_module_1_res), .A2(
        n_majority7_module_56__and_module_2_res), .ZN(
        n_majority7_module_56__or_module_4_res) );
  AND2_X1 u_majority7_module_56__and_module_5_U1 ( .A1(
        n_majority7_module_56__and_module_3_res), .A2(n_xor_module_8_res), 
        .ZN(n_majority7_module_56__and_module_5_res) );
  OR2_X1 u_majority7_module_56__or_module_5_U1 ( .A1(n_xor_module_8_res), .A2(
        n_majority7_module_56__and_module_3_res), .ZN(
        n_majority7_module_56__or_module_5_res) );
  AND2_X1 u_majority7_module_56__and_module_6_U1 ( .A1(
        n_majority7_module_56__or_module_1_res), .A2(
        n_majority7_module_56__or_module_2_res), .ZN(
        n_majority7_module_56__and_module_6_res) );
  OR2_X1 u_majority7_module_56__or_module_6_U1 ( .A1(
        n_majority7_module_56__or_module_2_res), .A2(
        n_majority7_module_56__or_module_1_res), .ZN(
        n_majority7_module_56__or_module_6_res) );
  OR2_X1 u_majority7_module_56__or_module_7_U1 ( .A1(
        n_majority7_module_56__and_module_4_res), .A2(
        n_majority7_module_56__and_module_5_res), .ZN(
        n_majority7_module_56__or_module_7_res) );
  AND2_X1 u_majority7_module_56__and_module_7_U1 ( .A1(
        n_majority7_module_56__or_module_3_res), .A2(
        n_majority7_module_56__or_module_4_res), .ZN(
        n_majority7_module_56__and_module_7_res) );
  OR2_X1 u_majority7_module_56__or_module_8_U1 ( .A1(
        n_majority7_module_56__or_module_4_res), .A2(
        n_majority7_module_56__or_module_3_res), .ZN(
        n_majority7_module_56__or_module_8_res) );
  AND2_X1 u_majority7_module_56__and_module_8_U1 ( .A1(
        n_majority7_module_56__or_module_5_res), .A2(
        n_majority7_module_56__and_module_6_res), .ZN(
        n_majority7_module_56__and_module_8_res) );
  OR2_X1 u_majority7_module_56__or_module_9_U1 ( .A1(
        n_majority7_module_56__and_module_6_res), .A2(
        n_majority7_module_56__or_module_5_res), .ZN(
        n_majority7_module_56__or_module_9_res) );
  OR2_X1 u_majority7_module_56__or_module_10_U1 ( .A1(
        n_majority7_module_56__or_module_7_res), .A2(
        n_majority7_module_56__and_module_7_res), .ZN(
        n_majority7_module_56__or_module_10_res) );
  AND2_X1 u_majority7_module_56__and_module_9_U1 ( .A1(
        n_majority7_module_56__or_module_6_res), .A2(
        n_majority7_module_56__or_module_9_res), .ZN(
        n_majority7_module_56__and_module_9_res) );
  OR2_X1 u_majority7_module_56__or_module_11_U1 ( .A1(
        n_majority7_module_56__or_module_10_res), .A2(
        n_majority7_module_56__and_module_8_res), .ZN(
        n_majority7_module_56__or_module_11_res) );
  AND2_X1 u_majority7_module_56__and_module_10_U1 ( .A1(
        n_majority7_module_56__or_module_8_res), .A2(
        n_majority7_module_56__and_module_9_res), .ZN(
        n_majority7_module_56__and_module_10_res) );
  AND2_X1 u_majority7_module_56__and_module_11_U1 ( .A1(
        n_majority7_module_56__and_module_10_res), .A2(
        n_majority7_module_56__or_module_11_res), .ZN(
        n_majority7_module_56_res) );
  DFF_X1 u_reg_module_57__cini_mul_v000_reg ( .D(n_majority7_module_56_res), 
        .CK(clock_6), .Q(n_reg_module_57_res), .QN() );
  AND2_X1 u_majority7_module_57__and_module_1_U1 ( .A1(n_xor_module_40_res), 
        .A2(n_xor_module_4_res), .ZN(n_majority7_module_57__and_module_1_res)
         );
  OR2_X1 u_majority7_module_57__or_module_1_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_40_res), .ZN(n_majority7_module_57__or_module_1_res) );
  AND2_X1 u_majority7_module_57__and_module_2_U1 ( .A1(n_xor_module_22_res), 
        .A2(n_xor_module_16_res), .ZN(n_majority7_module_57__and_module_2_res)
         );
  OR2_X1 u_majority7_module_57__or_module_2_U1 ( .A1(n_xor_module_16_res), 
        .A2(n_xor_module_22_res), .ZN(n_majority7_module_57__or_module_2_res)
         );
  AND2_X1 u_majority7_module_57__and_module_3_U1 ( .A1(n_xor_module_34_res), 
        .A2(n_xor_module_28_res), .ZN(n_majority7_module_57__and_module_3_res)
         );
  OR2_X1 u_majority7_module_57__or_module_3_U1 ( .A1(n_xor_module_28_res), 
        .A2(n_xor_module_34_res), .ZN(n_majority7_module_57__or_module_3_res)
         );
  AND2_X1 u_majority7_module_57__and_module_4_U1 ( .A1(
        n_majority7_module_57__and_module_2_res), .A2(
        n_majority7_module_57__and_module_1_res), .ZN(
        n_majority7_module_57__and_module_4_res) );
  OR2_X1 u_majority7_module_57__or_module_4_U1 ( .A1(
        n_majority7_module_57__and_module_1_res), .A2(
        n_majority7_module_57__and_module_2_res), .ZN(
        n_majority7_module_57__or_module_4_res) );
  AND2_X1 u_majority7_module_57__and_module_5_U1 ( .A1(
        n_majority7_module_57__and_module_3_res), .A2(n_xor_module_10_res), 
        .ZN(n_majority7_module_57__and_module_5_res) );
  OR2_X1 u_majority7_module_57__or_module_5_U1 ( .A1(n_xor_module_10_res), 
        .A2(n_majority7_module_57__and_module_3_res), .ZN(
        n_majority7_module_57__or_module_5_res) );
  AND2_X1 u_majority7_module_57__and_module_6_U1 ( .A1(
        n_majority7_module_57__or_module_1_res), .A2(
        n_majority7_module_57__or_module_2_res), .ZN(
        n_majority7_module_57__and_module_6_res) );
  OR2_X1 u_majority7_module_57__or_module_6_U1 ( .A1(
        n_majority7_module_57__or_module_2_res), .A2(
        n_majority7_module_57__or_module_1_res), .ZN(
        n_majority7_module_57__or_module_6_res) );
  OR2_X1 u_majority7_module_57__or_module_7_U1 ( .A1(
        n_majority7_module_57__and_module_4_res), .A2(
        n_majority7_module_57__and_module_5_res), .ZN(
        n_majority7_module_57__or_module_7_res) );
  AND2_X1 u_majority7_module_57__and_module_7_U1 ( .A1(
        n_majority7_module_57__or_module_3_res), .A2(
        n_majority7_module_57__or_module_4_res), .ZN(
        n_majority7_module_57__and_module_7_res) );
  OR2_X1 u_majority7_module_57__or_module_8_U1 ( .A1(
        n_majority7_module_57__or_module_4_res), .A2(
        n_majority7_module_57__or_module_3_res), .ZN(
        n_majority7_module_57__or_module_8_res) );
  AND2_X1 u_majority7_module_57__and_module_8_U1 ( .A1(
        n_majority7_module_57__or_module_5_res), .A2(
        n_majority7_module_57__and_module_6_res), .ZN(
        n_majority7_module_57__and_module_8_res) );
  OR2_X1 u_majority7_module_57__or_module_9_U1 ( .A1(
        n_majority7_module_57__and_module_6_res), .A2(
        n_majority7_module_57__or_module_5_res), .ZN(
        n_majority7_module_57__or_module_9_res) );
  OR2_X1 u_majority7_module_57__or_module_10_U1 ( .A1(
        n_majority7_module_57__or_module_7_res), .A2(
        n_majority7_module_57__and_module_7_res), .ZN(
        n_majority7_module_57__or_module_10_res) );
  AND2_X1 u_majority7_module_57__and_module_9_U1 ( .A1(
        n_majority7_module_57__or_module_6_res), .A2(
        n_majority7_module_57__or_module_9_res), .ZN(
        n_majority7_module_57__and_module_9_res) );
  OR2_X1 u_majority7_module_57__or_module_11_U1 ( .A1(
        n_majority7_module_57__or_module_10_res), .A2(
        n_majority7_module_57__and_module_8_res), .ZN(
        n_majority7_module_57__or_module_11_res) );
  AND2_X1 u_majority7_module_57__and_module_10_U1 ( .A1(
        n_majority7_module_57__or_module_8_res), .A2(
        n_majority7_module_57__and_module_9_res), .ZN(
        n_majority7_module_57__and_module_10_res) );
  AND2_X1 u_majority7_module_57__and_module_11_U1 ( .A1(
        n_majority7_module_57__and_module_10_res), .A2(
        n_majority7_module_57__or_module_11_res), .ZN(
        n_majority7_module_57_res) );
  DFF_X1 u_reg_module_58__cini_mul_v000_reg ( .D(n_majority7_module_57_res), 
        .CK(clock_6), .Q(n_reg_module_58_res), .QN() );
  AND2_X1 u_majority7_module_58__and_module_1_U1 ( .A1(n_xor_module_40_res), 
        .A2(n_xor_module_4_res), .ZN(n_majority7_module_58__and_module_1_res)
         );
  OR2_X1 u_majority7_module_58__or_module_1_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_40_res), .ZN(n_majority7_module_58__or_module_1_res) );
  AND2_X1 u_majority7_module_58__and_module_2_U1 ( .A1(n_xor_module_22_res), 
        .A2(n_xor_module_16_res), .ZN(n_majority7_module_58__and_module_2_res)
         );
  OR2_X1 u_majority7_module_58__or_module_2_U1 ( .A1(n_xor_module_16_res), 
        .A2(n_xor_module_22_res), .ZN(n_majority7_module_58__or_module_2_res)
         );
  AND2_X1 u_majority7_module_58__and_module_3_U1 ( .A1(n_xor_module_34_res), 
        .A2(n_xor_module_28_res), .ZN(n_majority7_module_58__and_module_3_res)
         );
  OR2_X1 u_majority7_module_58__or_module_3_U1 ( .A1(n_xor_module_28_res), 
        .A2(n_xor_module_34_res), .ZN(n_majority7_module_58__or_module_3_res)
         );
  AND2_X1 u_majority7_module_58__and_module_4_U1 ( .A1(
        n_majority7_module_58__and_module_2_res), .A2(
        n_majority7_module_58__and_module_1_res), .ZN(
        n_majority7_module_58__and_module_4_res) );
  OR2_X1 u_majority7_module_58__or_module_4_U1 ( .A1(
        n_majority7_module_58__and_module_1_res), .A2(
        n_majority7_module_58__and_module_2_res), .ZN(
        n_majority7_module_58__or_module_4_res) );
  AND2_X1 u_majority7_module_58__and_module_5_U1 ( .A1(
        n_majority7_module_58__and_module_3_res), .A2(n_xor_module_10_res), 
        .ZN(n_majority7_module_58__and_module_5_res) );
  OR2_X1 u_majority7_module_58__or_module_5_U1 ( .A1(n_xor_module_10_res), 
        .A2(n_majority7_module_58__and_module_3_res), .ZN(
        n_majority7_module_58__or_module_5_res) );
  AND2_X1 u_majority7_module_58__and_module_6_U1 ( .A1(
        n_majority7_module_58__or_module_1_res), .A2(
        n_majority7_module_58__or_module_2_res), .ZN(
        n_majority7_module_58__and_module_6_res) );
  OR2_X1 u_majority7_module_58__or_module_6_U1 ( .A1(
        n_majority7_module_58__or_module_2_res), .A2(
        n_majority7_module_58__or_module_1_res), .ZN(
        n_majority7_module_58__or_module_6_res) );
  OR2_X1 u_majority7_module_58__or_module_7_U1 ( .A1(
        n_majority7_module_58__and_module_4_res), .A2(
        n_majority7_module_58__and_module_5_res), .ZN(
        n_majority7_module_58__or_module_7_res) );
  AND2_X1 u_majority7_module_58__and_module_7_U1 ( .A1(
        n_majority7_module_58__or_module_3_res), .A2(
        n_majority7_module_58__or_module_4_res), .ZN(
        n_majority7_module_58__and_module_7_res) );
  OR2_X1 u_majority7_module_58__or_module_8_U1 ( .A1(
        n_majority7_module_58__or_module_4_res), .A2(
        n_majority7_module_58__or_module_3_res), .ZN(
        n_majority7_module_58__or_module_8_res) );
  AND2_X1 u_majority7_module_58__and_module_8_U1 ( .A1(
        n_majority7_module_58__or_module_5_res), .A2(
        n_majority7_module_58__and_module_6_res), .ZN(
        n_majority7_module_58__and_module_8_res) );
  OR2_X1 u_majority7_module_58__or_module_9_U1 ( .A1(
        n_majority7_module_58__and_module_6_res), .A2(
        n_majority7_module_58__or_module_5_res), .ZN(
        n_majority7_module_58__or_module_9_res) );
  OR2_X1 u_majority7_module_58__or_module_10_U1 ( .A1(
        n_majority7_module_58__or_module_7_res), .A2(
        n_majority7_module_58__and_module_7_res), .ZN(
        n_majority7_module_58__or_module_10_res) );
  AND2_X1 u_majority7_module_58__and_module_9_U1 ( .A1(
        n_majority7_module_58__or_module_6_res), .A2(
        n_majority7_module_58__or_module_9_res), .ZN(
        n_majority7_module_58__and_module_9_res) );
  OR2_X1 u_majority7_module_58__or_module_11_U1 ( .A1(
        n_majority7_module_58__or_module_10_res), .A2(
        n_majority7_module_58__and_module_8_res), .ZN(
        n_majority7_module_58__or_module_11_res) );
  AND2_X1 u_majority7_module_58__and_module_10_U1 ( .A1(
        n_majority7_module_58__or_module_8_res), .A2(
        n_majority7_module_58__and_module_9_res), .ZN(
        n_majority7_module_58__and_module_10_res) );
  AND2_X1 u_majority7_module_58__and_module_11_U1 ( .A1(
        n_majority7_module_58__and_module_10_res), .A2(
        n_majority7_module_58__or_module_11_res), .ZN(
        n_majority7_module_58_res) );
  DFF_X1 u_reg_module_59__cini_mul_v000_reg ( .D(n_majority7_module_58_res), 
        .CK(clock_6), .Q(n_reg_module_59_res), .QN() );
  AND2_X1 u_majority7_module_59__and_module_1_U1 ( .A1(n_xor_module_40_res), 
        .A2(n_xor_module_4_res), .ZN(n_majority7_module_59__and_module_1_res)
         );
  OR2_X1 u_majority7_module_59__or_module_1_U1 ( .A1(n_xor_module_4_res), .A2(
        n_xor_module_40_res), .ZN(n_majority7_module_59__or_module_1_res) );
  AND2_X1 u_majority7_module_59__and_module_2_U1 ( .A1(n_xor_module_22_res), 
        .A2(n_xor_module_16_res), .ZN(n_majority7_module_59__and_module_2_res)
         );
  OR2_X1 u_majority7_module_59__or_module_2_U1 ( .A1(n_xor_module_16_res), 
        .A2(n_xor_module_22_res), .ZN(n_majority7_module_59__or_module_2_res)
         );
  AND2_X1 u_majority7_module_59__and_module_3_U1 ( .A1(n_xor_module_34_res), 
        .A2(n_xor_module_28_res), .ZN(n_majority7_module_59__and_module_3_res)
         );
  OR2_X1 u_majority7_module_59__or_module_3_U1 ( .A1(n_xor_module_28_res), 
        .A2(n_xor_module_34_res), .ZN(n_majority7_module_59__or_module_3_res)
         );
  AND2_X1 u_majority7_module_59__and_module_4_U1 ( .A1(
        n_majority7_module_59__and_module_2_res), .A2(
        n_majority7_module_59__and_module_1_res), .ZN(
        n_majority7_module_59__and_module_4_res) );
  OR2_X1 u_majority7_module_59__or_module_4_U1 ( .A1(
        n_majority7_module_59__and_module_1_res), .A2(
        n_majority7_module_59__and_module_2_res), .ZN(
        n_majority7_module_59__or_module_4_res) );
  AND2_X1 u_majority7_module_59__and_module_5_U1 ( .A1(
        n_majority7_module_59__and_module_3_res), .A2(n_xor_module_10_res), 
        .ZN(n_majority7_module_59__and_module_5_res) );
  OR2_X1 u_majority7_module_59__or_module_5_U1 ( .A1(n_xor_module_10_res), 
        .A2(n_majority7_module_59__and_module_3_res), .ZN(
        n_majority7_module_59__or_module_5_res) );
  AND2_X1 u_majority7_module_59__and_module_6_U1 ( .A1(
        n_majority7_module_59__or_module_1_res), .A2(
        n_majority7_module_59__or_module_2_res), .ZN(
        n_majority7_module_59__and_module_6_res) );
  OR2_X1 u_majority7_module_59__or_module_6_U1 ( .A1(
        n_majority7_module_59__or_module_2_res), .A2(
        n_majority7_module_59__or_module_1_res), .ZN(
        n_majority7_module_59__or_module_6_res) );
  OR2_X1 u_majority7_module_59__or_module_7_U1 ( .A1(
        n_majority7_module_59__and_module_4_res), .A2(
        n_majority7_module_59__and_module_5_res), .ZN(
        n_majority7_module_59__or_module_7_res) );
  AND2_X1 u_majority7_module_59__and_module_7_U1 ( .A1(
        n_majority7_module_59__or_module_3_res), .A2(
        n_majority7_module_59__or_module_4_res), .ZN(
        n_majority7_module_59__and_module_7_res) );
  OR2_X1 u_majority7_module_59__or_module_8_U1 ( .A1(
        n_majority7_module_59__or_module_4_res), .A2(
        n_majority7_module_59__or_module_3_res), .ZN(
        n_majority7_module_59__or_module_8_res) );
  AND2_X1 u_majority7_module_59__and_module_8_U1 ( .A1(
        n_majority7_module_59__or_module_5_res), .A2(
        n_majority7_module_59__and_module_6_res), .ZN(
        n_majority7_module_59__and_module_8_res) );
  OR2_X1 u_majority7_module_59__or_module_9_U1 ( .A1(
        n_majority7_module_59__and_module_6_res), .A2(
        n_majority7_module_59__or_module_5_res), .ZN(
        n_majority7_module_59__or_module_9_res) );
  OR2_X1 u_majority7_module_59__or_module_10_U1 ( .A1(
        n_majority7_module_59__or_module_7_res), .A2(
        n_majority7_module_59__and_module_7_res), .ZN(
        n_majority7_module_59__or_module_10_res) );
  AND2_X1 u_majority7_module_59__and_module_9_U1 ( .A1(
        n_majority7_module_59__or_module_6_res), .A2(
        n_majority7_module_59__or_module_9_res), .ZN(
        n_majority7_module_59__and_module_9_res) );
  OR2_X1 u_majority7_module_59__or_module_11_U1 ( .A1(
        n_majority7_module_59__or_module_10_res), .A2(
        n_majority7_module_59__and_module_8_res), .ZN(
        n_majority7_module_59__or_module_11_res) );
  AND2_X1 u_majority7_module_59__and_module_10_U1 ( .A1(
        n_majority7_module_59__or_module_8_res), .A2(
        n_majority7_module_59__and_module_9_res), .ZN(
        n_majority7_module_59__and_module_10_res) );
  AND2_X1 u_majority7_module_59__and_module_11_U1 ( .A1(
        n_majority7_module_59__and_module_10_res), .A2(
        n_majority7_module_59__or_module_11_res), .ZN(
        n_majority7_module_59_res) );
  DFF_X1 u_reg_module_60__cini_mul_v000_reg ( .D(n_majority7_module_59_res), 
        .CK(clock_6), .Q(n_reg_module_60_res), .QN() );
  AND2_X1 u_majority7_module_60__and_module_1_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_60__and_module_1_res)
         );
  OR2_X1 u_majority7_module_60__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_60__or_module_1_res) );
  AND2_X1 u_majority7_module_60__and_module_2_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_xor_module_18_res), .ZN(n_majority7_module_60__and_module_2_res)
         );
  OR2_X1 u_majority7_module_60__or_module_2_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_xor_module_24_res), .ZN(n_majority7_module_60__or_module_2_res)
         );
  AND2_X1 u_majority7_module_60__and_module_3_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_60__and_module_3_res)
         );
  OR2_X1 u_majority7_module_60__or_module_3_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_60__or_module_3_res)
         );
  AND2_X1 u_majority7_module_60__and_module_4_U1 ( .A1(
        n_majority7_module_60__and_module_2_res), .A2(
        n_majority7_module_60__and_module_1_res), .ZN(
        n_majority7_module_60__and_module_4_res) );
  OR2_X1 u_majority7_module_60__or_module_4_U1 ( .A1(
        n_majority7_module_60__and_module_1_res), .A2(
        n_majority7_module_60__and_module_2_res), .ZN(
        n_majority7_module_60__or_module_4_res) );
  AND2_X1 u_majority7_module_60__and_module_5_U1 ( .A1(
        n_majority7_module_60__and_module_3_res), .A2(n_xor_module_12_res), 
        .ZN(n_majority7_module_60__and_module_5_res) );
  OR2_X1 u_majority7_module_60__or_module_5_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_majority7_module_60__and_module_3_res), .ZN(
        n_majority7_module_60__or_module_5_res) );
  AND2_X1 u_majority7_module_60__and_module_6_U1 ( .A1(
        n_majority7_module_60__or_module_1_res), .A2(
        n_majority7_module_60__or_module_2_res), .ZN(
        n_majority7_module_60__and_module_6_res) );
  OR2_X1 u_majority7_module_60__or_module_6_U1 ( .A1(
        n_majority7_module_60__or_module_2_res), .A2(
        n_majority7_module_60__or_module_1_res), .ZN(
        n_majority7_module_60__or_module_6_res) );
  OR2_X1 u_majority7_module_60__or_module_7_U1 ( .A1(
        n_majority7_module_60__and_module_4_res), .A2(
        n_majority7_module_60__and_module_5_res), .ZN(
        n_majority7_module_60__or_module_7_res) );
  AND2_X1 u_majority7_module_60__and_module_7_U1 ( .A1(
        n_majority7_module_60__or_module_3_res), .A2(
        n_majority7_module_60__or_module_4_res), .ZN(
        n_majority7_module_60__and_module_7_res) );
  OR2_X1 u_majority7_module_60__or_module_8_U1 ( .A1(
        n_majority7_module_60__or_module_4_res), .A2(
        n_majority7_module_60__or_module_3_res), .ZN(
        n_majority7_module_60__or_module_8_res) );
  AND2_X1 u_majority7_module_60__and_module_8_U1 ( .A1(
        n_majority7_module_60__or_module_5_res), .A2(
        n_majority7_module_60__and_module_6_res), .ZN(
        n_majority7_module_60__and_module_8_res) );
  OR2_X1 u_majority7_module_60__or_module_9_U1 ( .A1(
        n_majority7_module_60__and_module_6_res), .A2(
        n_majority7_module_60__or_module_5_res), .ZN(
        n_majority7_module_60__or_module_9_res) );
  OR2_X1 u_majority7_module_60__or_module_10_U1 ( .A1(
        n_majority7_module_60__or_module_7_res), .A2(
        n_majority7_module_60__and_module_7_res), .ZN(
        n_majority7_module_60__or_module_10_res) );
  AND2_X1 u_majority7_module_60__and_module_9_U1 ( .A1(
        n_majority7_module_60__or_module_6_res), .A2(
        n_majority7_module_60__or_module_9_res), .ZN(
        n_majority7_module_60__and_module_9_res) );
  OR2_X1 u_majority7_module_60__or_module_11_U1 ( .A1(
        n_majority7_module_60__or_module_10_res), .A2(
        n_majority7_module_60__and_module_8_res), .ZN(
        n_majority7_module_60__or_module_11_res) );
  AND2_X1 u_majority7_module_60__and_module_10_U1 ( .A1(
        n_majority7_module_60__or_module_8_res), .A2(
        n_majority7_module_60__and_module_9_res), .ZN(
        n_majority7_module_60__and_module_10_res) );
  AND2_X1 u_majority7_module_60__and_module_11_U1 ( .A1(
        n_majority7_module_60__and_module_10_res), .A2(
        n_majority7_module_60__or_module_11_res), .ZN(
        n_majority7_module_60_res) );
  DFF_X1 u_reg_module_61__cini_mul_v000_reg ( .D(n_majority7_module_60_res), 
        .CK(clock_6), .Q(n_reg_module_61_res), .QN() );
  AND2_X1 u_majority7_module_61__and_module_1_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_61__and_module_1_res)
         );
  OR2_X1 u_majority7_module_61__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_61__or_module_1_res) );
  AND2_X1 u_majority7_module_61__and_module_2_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_xor_module_18_res), .ZN(n_majority7_module_61__and_module_2_res)
         );
  OR2_X1 u_majority7_module_61__or_module_2_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_xor_module_24_res), .ZN(n_majority7_module_61__or_module_2_res)
         );
  AND2_X1 u_majority7_module_61__and_module_3_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_61__and_module_3_res)
         );
  OR2_X1 u_majority7_module_61__or_module_3_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_61__or_module_3_res)
         );
  AND2_X1 u_majority7_module_61__and_module_4_U1 ( .A1(
        n_majority7_module_61__and_module_2_res), .A2(
        n_majority7_module_61__and_module_1_res), .ZN(
        n_majority7_module_61__and_module_4_res) );
  OR2_X1 u_majority7_module_61__or_module_4_U1 ( .A1(
        n_majority7_module_61__and_module_1_res), .A2(
        n_majority7_module_61__and_module_2_res), .ZN(
        n_majority7_module_61__or_module_4_res) );
  AND2_X1 u_majority7_module_61__and_module_5_U1 ( .A1(
        n_majority7_module_61__and_module_3_res), .A2(n_xor_module_12_res), 
        .ZN(n_majority7_module_61__and_module_5_res) );
  OR2_X1 u_majority7_module_61__or_module_5_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_majority7_module_61__and_module_3_res), .ZN(
        n_majority7_module_61__or_module_5_res) );
  AND2_X1 u_majority7_module_61__and_module_6_U1 ( .A1(
        n_majority7_module_61__or_module_1_res), .A2(
        n_majority7_module_61__or_module_2_res), .ZN(
        n_majority7_module_61__and_module_6_res) );
  OR2_X1 u_majority7_module_61__or_module_6_U1 ( .A1(
        n_majority7_module_61__or_module_2_res), .A2(
        n_majority7_module_61__or_module_1_res), .ZN(
        n_majority7_module_61__or_module_6_res) );
  OR2_X1 u_majority7_module_61__or_module_7_U1 ( .A1(
        n_majority7_module_61__and_module_4_res), .A2(
        n_majority7_module_61__and_module_5_res), .ZN(
        n_majority7_module_61__or_module_7_res) );
  AND2_X1 u_majority7_module_61__and_module_7_U1 ( .A1(
        n_majority7_module_61__or_module_3_res), .A2(
        n_majority7_module_61__or_module_4_res), .ZN(
        n_majority7_module_61__and_module_7_res) );
  OR2_X1 u_majority7_module_61__or_module_8_U1 ( .A1(
        n_majority7_module_61__or_module_4_res), .A2(
        n_majority7_module_61__or_module_3_res), .ZN(
        n_majority7_module_61__or_module_8_res) );
  AND2_X1 u_majority7_module_61__and_module_8_U1 ( .A1(
        n_majority7_module_61__or_module_5_res), .A2(
        n_majority7_module_61__and_module_6_res), .ZN(
        n_majority7_module_61__and_module_8_res) );
  OR2_X1 u_majority7_module_61__or_module_9_U1 ( .A1(
        n_majority7_module_61__and_module_6_res), .A2(
        n_majority7_module_61__or_module_5_res), .ZN(
        n_majority7_module_61__or_module_9_res) );
  OR2_X1 u_majority7_module_61__or_module_10_U1 ( .A1(
        n_majority7_module_61__or_module_7_res), .A2(
        n_majority7_module_61__and_module_7_res), .ZN(
        n_majority7_module_61__or_module_10_res) );
  AND2_X1 u_majority7_module_61__and_module_9_U1 ( .A1(
        n_majority7_module_61__or_module_6_res), .A2(
        n_majority7_module_61__or_module_9_res), .ZN(
        n_majority7_module_61__and_module_9_res) );
  OR2_X1 u_majority7_module_61__or_module_11_U1 ( .A1(
        n_majority7_module_61__or_module_10_res), .A2(
        n_majority7_module_61__and_module_8_res), .ZN(
        n_majority7_module_61__or_module_11_res) );
  AND2_X1 u_majority7_module_61__and_module_10_U1 ( .A1(
        n_majority7_module_61__or_module_8_res), .A2(
        n_majority7_module_61__and_module_9_res), .ZN(
        n_majority7_module_61__and_module_10_res) );
  AND2_X1 u_majority7_module_61__and_module_11_U1 ( .A1(
        n_majority7_module_61__and_module_10_res), .A2(
        n_majority7_module_61__or_module_11_res), .ZN(
        n_majority7_module_61_res) );
  DFF_X1 u_reg_module_62__cini_mul_v000_reg ( .D(n_majority7_module_61_res), 
        .CK(clock_6), .Q(n_reg_module_62_res), .QN() );
  AND2_X1 u_majority7_module_62__and_module_1_U1 ( .A1(n_xor_module_42_res), 
        .A2(n_xor_module_6_res), .ZN(n_majority7_module_62__and_module_1_res)
         );
  OR2_X1 u_majority7_module_62__or_module_1_U1 ( .A1(n_xor_module_6_res), .A2(
        n_xor_module_42_res), .ZN(n_majority7_module_62__or_module_1_res) );
  AND2_X1 u_majority7_module_62__and_module_2_U1 ( .A1(n_xor_module_24_res), 
        .A2(n_xor_module_18_res), .ZN(n_majority7_module_62__and_module_2_res)
         );
  OR2_X1 u_majority7_module_62__or_module_2_U1 ( .A1(n_xor_module_18_res), 
        .A2(n_xor_module_24_res), .ZN(n_majority7_module_62__or_module_2_res)
         );
  AND2_X1 u_majority7_module_62__and_module_3_U1 ( .A1(n_xor_module_36_res), 
        .A2(n_xor_module_30_res), .ZN(n_majority7_module_62__and_module_3_res)
         );
  OR2_X1 u_majority7_module_62__or_module_3_U1 ( .A1(n_xor_module_30_res), 
        .A2(n_xor_module_36_res), .ZN(n_majority7_module_62__or_module_3_res)
         );
  AND2_X1 u_majority7_module_62__and_module_4_U1 ( .A1(
        n_majority7_module_62__and_module_2_res), .A2(
        n_majority7_module_62__and_module_1_res), .ZN(
        n_majority7_module_62__and_module_4_res) );
  OR2_X1 u_majority7_module_62__or_module_4_U1 ( .A1(
        n_majority7_module_62__and_module_1_res), .A2(
        n_majority7_module_62__and_module_2_res), .ZN(
        n_majority7_module_62__or_module_4_res) );
  AND2_X1 u_majority7_module_62__and_module_5_U1 ( .A1(
        n_majority7_module_62__and_module_3_res), .A2(n_xor_module_12_res), 
        .ZN(n_majority7_module_62__and_module_5_res) );
  OR2_X1 u_majority7_module_62__or_module_5_U1 ( .A1(n_xor_module_12_res), 
        .A2(n_majority7_module_62__and_module_3_res), .ZN(
        n_majority7_module_62__or_module_5_res) );
  AND2_X1 u_majority7_module_62__and_module_6_U1 ( .A1(
        n_majority7_module_62__or_module_1_res), .A2(
        n_majority7_module_62__or_module_2_res), .ZN(
        n_majority7_module_62__and_module_6_res) );
  OR2_X1 u_majority7_module_62__or_module_6_U1 ( .A1(
        n_majority7_module_62__or_module_2_res), .A2(
        n_majority7_module_62__or_module_1_res), .ZN(
        n_majority7_module_62__or_module_6_res) );
  OR2_X1 u_majority7_module_62__or_module_7_U1 ( .A1(
        n_majority7_module_62__and_module_4_res), .A2(
        n_majority7_module_62__and_module_5_res), .ZN(
        n_majority7_module_62__or_module_7_res) );
  AND2_X1 u_majority7_module_62__and_module_7_U1 ( .A1(
        n_majority7_module_62__or_module_3_res), .A2(
        n_majority7_module_62__or_module_4_res), .ZN(
        n_majority7_module_62__and_module_7_res) );
  OR2_X1 u_majority7_module_62__or_module_8_U1 ( .A1(
        n_majority7_module_62__or_module_4_res), .A2(
        n_majority7_module_62__or_module_3_res), .ZN(
        n_majority7_module_62__or_module_8_res) );
  AND2_X1 u_majority7_module_62__and_module_8_U1 ( .A1(
        n_majority7_module_62__or_module_5_res), .A2(
        n_majority7_module_62__and_module_6_res), .ZN(
        n_majority7_module_62__and_module_8_res) );
  OR2_X1 u_majority7_module_62__or_module_9_U1 ( .A1(
        n_majority7_module_62__and_module_6_res), .A2(
        n_majority7_module_62__or_module_5_res), .ZN(
        n_majority7_module_62__or_module_9_res) );
  OR2_X1 u_majority7_module_62__or_module_10_U1 ( .A1(
        n_majority7_module_62__or_module_7_res), .A2(
        n_majority7_module_62__and_module_7_res), .ZN(
        n_majority7_module_62__or_module_10_res) );
  AND2_X1 u_majority7_module_62__and_module_9_U1 ( .A1(
        n_majority7_module_62__or_module_6_res), .A2(
        n_majority7_module_62__or_module_9_res), .ZN(
        n_majority7_module_62__and_module_9_res) );
  OR2_X1 u_majority7_module_62__or_module_11_U1 ( .A1(
        n_majority7_module_62__or_module_10_res), .A2(
        n_majority7_module_62__and_module_8_res), .ZN(
        n_majority7_module_62__or_module_11_res) );
  AND2_X1 u_majority7_module_62__and_module_10_U1 ( .A1(
        n_majority7_module_62__or_module_8_res), .A2(
        n_majority7_module_62__and_module_9_res), .ZN(
        n_majority7_module_62__and_module_10_res) );
  AND2_X1 u_majority7_module_62__and_module_11_U1 ( .A1(
        n_majority7_module_62__and_module_10_res), .A2(
        n_majority7_module_62__or_module_11_res), .ZN(
        n_majority7_module_62_res) );
  DFF_X1 u_reg_module_63__cini_mul_v000_reg ( .D(n_majority7_module_62_res), 
        .CK(clock_6), .Q(n_reg_module_63_res), .QN() );
  AND2_X1 u_and_module_1_U1 ( .A1(n_reg_module_1_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_1_res) );
  DFF_X1 u_reg_module_64__cini_mul_v000_reg ( .D(n_and_module_1_res), .CK(
        clock_0), .Q(n_reg_module_64_res), .QN() );
  AND2_X1 u_and_module_2_U1 ( .A1(n_reg_module_4_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_2_res) );
  XOR2_X1 u_xor_module_43_U1 ( .A(p_rand_3), .B(n_and_module_2_res), .Z(
        n_xor_module_43_res) );
  DFF_X1 u_reg_module_65__cini_mul_v000_reg ( .D(n_xor_module_43_res), .CK(
        clock_0), .Q(n_reg_module_65_res), .QN() );
  AND2_X1 u_and_module_3_U1 ( .A1(n_reg_module_7_res), .A2(io_i0_s0_d0), .ZN(
        n_and_module_3_res) );
  XOR2_X1 u_xor_module_44_U1 ( .A(p_rand_4), .B(n_and_module_3_res), .Z(
        n_xor_module_44_res) );
  DFF_X1 u_reg_module_66__cini_mul_v000_reg ( .D(n_xor_module_44_res), .CK(
        clock_0), .Q(n_reg_module_66_res), .QN() );
  AND2_X1 u_and_module_4_U1 ( .A1(n_reg_module_2_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_4_res) );
  XOR2_X1 u_xor_module_45_U1 ( .A(p_rand_3), .B(n_and_module_4_res), .Z(
        n_xor_module_45_res) );
  DFF_X1 u_reg_module_67__cini_mul_v000_reg ( .D(n_xor_module_45_res), .CK(
        clock_0), .Q(n_reg_module_67_res), .QN() );
  AND2_X1 u_and_module_5_U1 ( .A1(n_reg_module_5_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_5_res) );
  DFF_X1 u_reg_module_68__cini_mul_v000_reg ( .D(n_and_module_5_res), .CK(
        clock_0), .Q(n_reg_module_68_res), .QN() );
  AND2_X1 u_and_module_6_U1 ( .A1(n_reg_module_8_res), .A2(io_i0_s1_d0), .ZN(
        n_and_module_6_res) );
  XOR2_X1 u_xor_module_46_U1 ( .A(p_rand_5), .B(n_and_module_6_res), .Z(
        n_xor_module_46_res) );
  DFF_X1 u_reg_module_69__cini_mul_v000_reg ( .D(n_xor_module_46_res), .CK(
        clock_0), .Q(n_reg_module_69_res), .QN() );
  AND2_X1 u_and_module_7_U1 ( .A1(n_reg_module_3_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_7_res) );
  XOR2_X1 u_xor_module_47_U1 ( .A(p_rand_4), .B(n_and_module_7_res), .Z(
        n_xor_module_47_res) );
  DFF_X1 u_reg_module_70__cini_mul_v000_reg ( .D(n_xor_module_47_res), .CK(
        clock_0), .Q(n_reg_module_70_res), .QN() );
  AND2_X1 u_and_module_8_U1 ( .A1(n_reg_module_6_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_8_res) );
  XOR2_X1 u_xor_module_48_U1 ( .A(p_rand_5), .B(n_and_module_8_res), .Z(
        n_xor_module_48_res) );
  DFF_X1 u_reg_module_71__cini_mul_v000_reg ( .D(n_xor_module_48_res), .CK(
        clock_0), .Q(n_reg_module_71_res), .QN() );
  AND2_X1 u_and_module_9_U1 ( .A1(n_reg_module_9_res), .A2(io_i0_s2_d0), .ZN(
        n_and_module_9_res) );
  DFF_X1 u_reg_module_72__cini_mul_v000_reg ( .D(n_and_module_9_res), .CK(
        clock_0), .Q(n_reg_module_72_res), .QN() );
  AND2_X1 u_and_module_10_U1 ( .A1(n_reg_module_10_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_10_res) );
  DFF_X1 u_reg_module_73__cini_mul_v000_reg ( .D(n_and_module_10_res), .CK(
        clock_1), .Q(n_reg_module_73_res), .QN() );
  AND2_X1 u_and_module_11_U1 ( .A1(n_reg_module_13_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_11_res) );
  XOR2_X1 u_xor_module_49_U1 ( .A(p_rand_3), .B(n_and_module_11_res), .Z(
        n_xor_module_49_res) );
  DFF_X1 u_reg_module_74__cini_mul_v000_reg ( .D(n_xor_module_49_res), .CK(
        clock_1), .Q(n_reg_module_74_res), .QN() );
  AND2_X1 u_and_module_12_U1 ( .A1(n_reg_module_16_res), .A2(io_i0_s0_d1), 
        .ZN(n_and_module_12_res) );
  XOR2_X1 u_xor_module_50_U1 ( .A(p_rand_4), .B(n_and_module_12_res), .Z(
        n_xor_module_50_res) );
  DFF_X1 u_reg_module_75__cini_mul_v000_reg ( .D(n_xor_module_50_res), .CK(
        clock_1), .Q(n_reg_module_75_res), .QN() );
  AND2_X1 u_and_module_13_U1 ( .A1(n_reg_module_11_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_13_res) );
  XOR2_X1 u_xor_module_51_U1 ( .A(p_rand_3), .B(n_and_module_13_res), .Z(
        n_xor_module_51_res) );
  DFF_X1 u_reg_module_76__cini_mul_v000_reg ( .D(n_xor_module_51_res), .CK(
        clock_1), .Q(n_reg_module_76_res), .QN() );
  AND2_X1 u_and_module_14_U1 ( .A1(n_reg_module_14_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_14_res) );
  DFF_X1 u_reg_module_77__cini_mul_v000_reg ( .D(n_and_module_14_res), .CK(
        clock_1), .Q(n_reg_module_77_res), .QN() );
  AND2_X1 u_and_module_15_U1 ( .A1(n_reg_module_17_res), .A2(io_i0_s1_d1), 
        .ZN(n_and_module_15_res) );
  XOR2_X1 u_xor_module_52_U1 ( .A(p_rand_5), .B(n_and_module_15_res), .Z(
        n_xor_module_52_res) );
  DFF_X1 u_reg_module_78__cini_mul_v000_reg ( .D(n_xor_module_52_res), .CK(
        clock_1), .Q(n_reg_module_78_res), .QN() );
  AND2_X1 u_and_module_16_U1 ( .A1(n_reg_module_12_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_16_res) );
  XOR2_X1 u_xor_module_53_U1 ( .A(p_rand_4), .B(n_and_module_16_res), .Z(
        n_xor_module_53_res) );
  DFF_X1 u_reg_module_79__cini_mul_v000_reg ( .D(n_xor_module_53_res), .CK(
        clock_1), .Q(n_reg_module_79_res), .QN() );
  AND2_X1 u_and_module_17_U1 ( .A1(n_reg_module_15_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_17_res) );
  XOR2_X1 u_xor_module_54_U1 ( .A(p_rand_5), .B(n_and_module_17_res), .Z(
        n_xor_module_54_res) );
  DFF_X1 u_reg_module_80__cini_mul_v000_reg ( .D(n_xor_module_54_res), .CK(
        clock_1), .Q(n_reg_module_80_res), .QN() );
  AND2_X1 u_and_module_18_U1 ( .A1(n_reg_module_18_res), .A2(io_i0_s2_d1), 
        .ZN(n_and_module_18_res) );
  DFF_X1 u_reg_module_81__cini_mul_v000_reg ( .D(n_and_module_18_res), .CK(
        clock_1), .Q(n_reg_module_81_res), .QN() );
  AND2_X1 u_and_module_19_U1 ( .A1(n_reg_module_19_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_19_res) );
  DFF_X1 u_reg_module_82__cini_mul_v000_reg ( .D(n_and_module_19_res), .CK(
        clock_2), .Q(n_reg_module_82_res), .QN() );
  AND2_X1 u_and_module_20_U1 ( .A1(n_reg_module_22_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_20_res) );
  XOR2_X1 u_xor_module_55_U1 ( .A(p_rand_3), .B(n_and_module_20_res), .Z(
        n_xor_module_55_res) );
  DFF_X1 u_reg_module_83__cini_mul_v000_reg ( .D(n_xor_module_55_res), .CK(
        clock_2), .Q(n_reg_module_83_res), .QN() );
  AND2_X1 u_and_module_21_U1 ( .A1(n_reg_module_25_res), .A2(io_i0_s0_d2), 
        .ZN(n_and_module_21_res) );
  XOR2_X1 u_xor_module_56_U1 ( .A(p_rand_4), .B(n_and_module_21_res), .Z(
        n_xor_module_56_res) );
  DFF_X1 u_reg_module_84__cini_mul_v000_reg ( .D(n_xor_module_56_res), .CK(
        clock_2), .Q(n_reg_module_84_res), .QN() );
  AND2_X1 u_and_module_22_U1 ( .A1(n_reg_module_20_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_22_res) );
  XOR2_X1 u_xor_module_57_U1 ( .A(p_rand_3), .B(n_and_module_22_res), .Z(
        n_xor_module_57_res) );
  DFF_X1 u_reg_module_85__cini_mul_v000_reg ( .D(n_xor_module_57_res), .CK(
        clock_2), .Q(n_reg_module_85_res), .QN() );
  AND2_X1 u_and_module_23_U1 ( .A1(n_reg_module_23_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_23_res) );
  DFF_X1 u_reg_module_86__cini_mul_v000_reg ( .D(n_and_module_23_res), .CK(
        clock_2), .Q(n_reg_module_86_res), .QN() );
  AND2_X1 u_and_module_24_U1 ( .A1(n_reg_module_26_res), .A2(io_i0_s1_d2), 
        .ZN(n_and_module_24_res) );
  XOR2_X1 u_xor_module_58_U1 ( .A(p_rand_5), .B(n_and_module_24_res), .Z(
        n_xor_module_58_res) );
  DFF_X1 u_reg_module_87__cini_mul_v000_reg ( .D(n_xor_module_58_res), .CK(
        clock_2), .Q(n_reg_module_87_res), .QN() );
  AND2_X1 u_and_module_25_U1 ( .A1(n_reg_module_21_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_25_res) );
  XOR2_X1 u_xor_module_59_U1 ( .A(p_rand_4), .B(n_and_module_25_res), .Z(
        n_xor_module_59_res) );
  DFF_X1 u_reg_module_88__cini_mul_v000_reg ( .D(n_xor_module_59_res), .CK(
        clock_2), .Q(n_reg_module_88_res), .QN() );
  AND2_X1 u_and_module_26_U1 ( .A1(n_reg_module_24_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_26_res) );
  XOR2_X1 u_xor_module_60_U1 ( .A(p_rand_5), .B(n_and_module_26_res), .Z(
        n_xor_module_60_res) );
  DFF_X1 u_reg_module_89__cini_mul_v000_reg ( .D(n_xor_module_60_res), .CK(
        clock_2), .Q(n_reg_module_89_res), .QN() );
  AND2_X1 u_and_module_27_U1 ( .A1(n_reg_module_27_res), .A2(io_i0_s2_d2), 
        .ZN(n_and_module_27_res) );
  DFF_X1 u_reg_module_90__cini_mul_v000_reg ( .D(n_and_module_27_res), .CK(
        clock_2), .Q(n_reg_module_90_res), .QN() );
  AND2_X1 u_and_module_28_U1 ( .A1(n_reg_module_28_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_28_res) );
  DFF_X1 u_reg_module_91__cini_mul_v000_reg ( .D(n_and_module_28_res), .CK(
        clock_3), .Q(n_reg_module_91_res), .QN() );
  AND2_X1 u_and_module_29_U1 ( .A1(n_reg_module_31_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_29_res) );
  XOR2_X1 u_xor_module_61_U1 ( .A(p_rand_3), .B(n_and_module_29_res), .Z(
        n_xor_module_61_res) );
  DFF_X1 u_reg_module_92__cini_mul_v000_reg ( .D(n_xor_module_61_res), .CK(
        clock_3), .Q(n_reg_module_92_res), .QN() );
  AND2_X1 u_and_module_30_U1 ( .A1(n_reg_module_34_res), .A2(io_i0_s0_d3), 
        .ZN(n_and_module_30_res) );
  XOR2_X1 u_xor_module_62_U1 ( .A(p_rand_4), .B(n_and_module_30_res), .Z(
        n_xor_module_62_res) );
  DFF_X1 u_reg_module_93__cini_mul_v000_reg ( .D(n_xor_module_62_res), .CK(
        clock_3), .Q(n_reg_module_93_res), .QN() );
  AND2_X1 u_and_module_31_U1 ( .A1(n_reg_module_29_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_31_res) );
  XOR2_X1 u_xor_module_63_U1 ( .A(p_rand_3), .B(n_and_module_31_res), .Z(
        n_xor_module_63_res) );
  DFF_X1 u_reg_module_94__cini_mul_v000_reg ( .D(n_xor_module_63_res), .CK(
        clock_3), .Q(n_reg_module_94_res), .QN() );
  AND2_X1 u_and_module_32_U1 ( .A1(n_reg_module_32_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_32_res) );
  DFF_X1 u_reg_module_95__cini_mul_v000_reg ( .D(n_and_module_32_res), .CK(
        clock_3), .Q(n_reg_module_95_res), .QN() );
  AND2_X1 u_and_module_33_U1 ( .A1(n_reg_module_35_res), .A2(io_i0_s1_d3), 
        .ZN(n_and_module_33_res) );
  XOR2_X1 u_xor_module_64_U1 ( .A(p_rand_5), .B(n_and_module_33_res), .Z(
        n_xor_module_64_res) );
  DFF_X1 u_reg_module_96__cini_mul_v000_reg ( .D(n_xor_module_64_res), .CK(
        clock_3), .Q(n_reg_module_96_res), .QN() );
  AND2_X1 u_and_module_34_U1 ( .A1(n_reg_module_30_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_34_res) );
  XOR2_X1 u_xor_module_65_U1 ( .A(p_rand_4), .B(n_and_module_34_res), .Z(
        n_xor_module_65_res) );
  DFF_X1 u_reg_module_97__cini_mul_v000_reg ( .D(n_xor_module_65_res), .CK(
        clock_3), .Q(n_reg_module_97_res), .QN() );
  AND2_X1 u_and_module_35_U1 ( .A1(n_reg_module_33_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_35_res) );
  XOR2_X1 u_xor_module_66_U1 ( .A(p_rand_5), .B(n_and_module_35_res), .Z(
        n_xor_module_66_res) );
  DFF_X1 u_reg_module_98__cini_mul_v000_reg ( .D(n_xor_module_66_res), .CK(
        clock_3), .Q(n_reg_module_98_res), .QN() );
  AND2_X1 u_and_module_36_U1 ( .A1(n_reg_module_36_res), .A2(io_i0_s2_d3), 
        .ZN(n_and_module_36_res) );
  DFF_X1 u_reg_module_99__cini_mul_v000_reg ( .D(n_and_module_36_res), .CK(
        clock_3), .Q(n_reg_module_99_res), .QN() );
  AND2_X1 u_and_module_37_U1 ( .A1(n_reg_module_37_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_37_res) );
  DFF_X1 u_reg_module_100__cini_mul_v000_reg ( .D(n_and_module_37_res), .CK(
        clock_4), .Q(n_reg_module_100_res), .QN() );
  AND2_X1 u_and_module_38_U1 ( .A1(n_reg_module_40_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_38_res) );
  XOR2_X1 u_xor_module_67_U1 ( .A(p_rand_3), .B(n_and_module_38_res), .Z(
        n_xor_module_67_res) );
  DFF_X1 u_reg_module_101__cini_mul_v000_reg ( .D(n_xor_module_67_res), .CK(
        clock_4), .Q(n_reg_module_101_res), .QN() );
  AND2_X1 u_and_module_39_U1 ( .A1(n_reg_module_43_res), .A2(io_i0_s0_d4), 
        .ZN(n_and_module_39_res) );
  XOR2_X1 u_xor_module_68_U1 ( .A(p_rand_4), .B(n_and_module_39_res), .Z(
        n_xor_module_68_res) );
  DFF_X1 u_reg_module_102__cini_mul_v000_reg ( .D(n_xor_module_68_res), .CK(
        clock_4), .Q(n_reg_module_102_res), .QN() );
  AND2_X1 u_and_module_40_U1 ( .A1(n_reg_module_38_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_40_res) );
  XOR2_X1 u_xor_module_69_U1 ( .A(p_rand_3), .B(n_and_module_40_res), .Z(
        n_xor_module_69_res) );
  DFF_X1 u_reg_module_103__cini_mul_v000_reg ( .D(n_xor_module_69_res), .CK(
        clock_4), .Q(n_reg_module_103_res), .QN() );
  AND2_X1 u_and_module_41_U1 ( .A1(n_reg_module_41_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_41_res) );
  DFF_X1 u_reg_module_104__cini_mul_v000_reg ( .D(n_and_module_41_res), .CK(
        clock_4), .Q(n_reg_module_104_res), .QN() );
  AND2_X1 u_and_module_42_U1 ( .A1(n_reg_module_44_res), .A2(io_i0_s1_d4), 
        .ZN(n_and_module_42_res) );
  XOR2_X1 u_xor_module_70_U1 ( .A(p_rand_5), .B(n_and_module_42_res), .Z(
        n_xor_module_70_res) );
  DFF_X1 u_reg_module_105__cini_mul_v000_reg ( .D(n_xor_module_70_res), .CK(
        clock_4), .Q(n_reg_module_105_res), .QN() );
  AND2_X1 u_and_module_43_U1 ( .A1(n_reg_module_39_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_43_res) );
  XOR2_X1 u_xor_module_71_U1 ( .A(p_rand_4), .B(n_and_module_43_res), .Z(
        n_xor_module_71_res) );
  DFF_X1 u_reg_module_106__cini_mul_v000_reg ( .D(n_xor_module_71_res), .CK(
        clock_4), .Q(n_reg_module_106_res), .QN() );
  AND2_X1 u_and_module_44_U1 ( .A1(n_reg_module_42_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_44_res) );
  XOR2_X1 u_xor_module_72_U1 ( .A(p_rand_5), .B(n_and_module_44_res), .Z(
        n_xor_module_72_res) );
  DFF_X1 u_reg_module_107__cini_mul_v000_reg ( .D(n_xor_module_72_res), .CK(
        clock_4), .Q(n_reg_module_107_res), .QN() );
  AND2_X1 u_and_module_45_U1 ( .A1(n_reg_module_45_res), .A2(io_i0_s2_d4), 
        .ZN(n_and_module_45_res) );
  DFF_X1 u_reg_module_108__cini_mul_v000_reg ( .D(n_and_module_45_res), .CK(
        clock_4), .Q(n_reg_module_108_res), .QN() );
  AND2_X1 u_and_module_46_U1 ( .A1(n_reg_module_46_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_46_res) );
  DFF_X1 u_reg_module_109__cini_mul_v000_reg ( .D(n_and_module_46_res), .CK(
        clock_5), .Q(n_reg_module_109_res), .QN() );
  AND2_X1 u_and_module_47_U1 ( .A1(n_reg_module_49_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_47_res) );
  XOR2_X1 u_xor_module_73_U1 ( .A(p_rand_3), .B(n_and_module_47_res), .Z(
        n_xor_module_73_res) );
  DFF_X1 u_reg_module_110__cini_mul_v000_reg ( .D(n_xor_module_73_res), .CK(
        clock_5), .Q(n_reg_module_110_res), .QN() );
  AND2_X1 u_and_module_48_U1 ( .A1(n_reg_module_52_res), .A2(io_i0_s0_d5), 
        .ZN(n_and_module_48_res) );
  XOR2_X1 u_xor_module_74_U1 ( .A(p_rand_4), .B(n_and_module_48_res), .Z(
        n_xor_module_74_res) );
  DFF_X1 u_reg_module_111__cini_mul_v000_reg ( .D(n_xor_module_74_res), .CK(
        clock_5), .Q(n_reg_module_111_res), .QN() );
  AND2_X1 u_and_module_49_U1 ( .A1(n_reg_module_47_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_49_res) );
  XOR2_X1 u_xor_module_75_U1 ( .A(p_rand_3), .B(n_and_module_49_res), .Z(
        n_xor_module_75_res) );
  DFF_X1 u_reg_module_112__cini_mul_v000_reg ( .D(n_xor_module_75_res), .CK(
        clock_5), .Q(n_reg_module_112_res), .QN() );
  AND2_X1 u_and_module_50_U1 ( .A1(n_reg_module_50_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_50_res) );
  DFF_X1 u_reg_module_113__cini_mul_v000_reg ( .D(n_and_module_50_res), .CK(
        clock_5), .Q(n_reg_module_113_res), .QN() );
  AND2_X1 u_and_module_51_U1 ( .A1(n_reg_module_53_res), .A2(io_i0_s1_d5), 
        .ZN(n_and_module_51_res) );
  XOR2_X1 u_xor_module_76_U1 ( .A(p_rand_5), .B(n_and_module_51_res), .Z(
        n_xor_module_76_res) );
  DFF_X1 u_reg_module_114__cini_mul_v000_reg ( .D(n_xor_module_76_res), .CK(
        clock_5), .Q(n_reg_module_114_res), .QN() );
  AND2_X1 u_and_module_52_U1 ( .A1(n_reg_module_48_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_52_res) );
  XOR2_X1 u_xor_module_77_U1 ( .A(p_rand_4), .B(n_and_module_52_res), .Z(
        n_xor_module_77_res) );
  DFF_X1 u_reg_module_115__cini_mul_v000_reg ( .D(n_xor_module_77_res), .CK(
        clock_5), .Q(n_reg_module_115_res), .QN() );
  AND2_X1 u_and_module_53_U1 ( .A1(n_reg_module_51_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_53_res) );
  XOR2_X1 u_xor_module_78_U1 ( .A(p_rand_5), .B(n_and_module_53_res), .Z(
        n_xor_module_78_res) );
  DFF_X1 u_reg_module_116__cini_mul_v000_reg ( .D(n_xor_module_78_res), .CK(
        clock_5), .Q(n_reg_module_116_res), .QN() );
  AND2_X1 u_and_module_54_U1 ( .A1(n_reg_module_54_res), .A2(io_i0_s2_d5), 
        .ZN(n_and_module_54_res) );
  DFF_X1 u_reg_module_117__cini_mul_v000_reg ( .D(n_and_module_54_res), .CK(
        clock_5), .Q(n_reg_module_117_res), .QN() );
  AND2_X1 u_and_module_55_U1 ( .A1(n_reg_module_55_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_55_res) );
  DFF_X1 u_reg_module_118__cini_mul_v000_reg ( .D(n_and_module_55_res), .CK(
        clock_6), .Q(n_reg_module_118_res), .QN() );
  AND2_X1 u_and_module_56_U1 ( .A1(n_reg_module_58_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_56_res) );
  XOR2_X1 u_xor_module_79_U1 ( .A(p_rand_3), .B(n_and_module_56_res), .Z(
        n_xor_module_79_res) );
  DFF_X1 u_reg_module_119__cini_mul_v000_reg ( .D(n_xor_module_79_res), .CK(
        clock_6), .Q(n_reg_module_119_res), .QN() );
  AND2_X1 u_and_module_57_U1 ( .A1(n_reg_module_61_res), .A2(io_i0_s0_d6), 
        .ZN(n_and_module_57_res) );
  XOR2_X1 u_xor_module_80_U1 ( .A(p_rand_4), .B(n_and_module_57_res), .Z(
        n_xor_module_80_res) );
  DFF_X1 u_reg_module_120__cini_mul_v000_reg ( .D(n_xor_module_80_res), .CK(
        clock_6), .Q(n_reg_module_120_res), .QN() );
  AND2_X1 u_and_module_58_U1 ( .A1(n_reg_module_56_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_58_res) );
  XOR2_X1 u_xor_module_81_U1 ( .A(p_rand_3), .B(n_and_module_58_res), .Z(
        n_xor_module_81_res) );
  DFF_X1 u_reg_module_121__cini_mul_v000_reg ( .D(n_xor_module_81_res), .CK(
        clock_6), .Q(n_reg_module_121_res), .QN() );
  AND2_X1 u_and_module_59_U1 ( .A1(n_reg_module_59_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_59_res) );
  DFF_X1 u_reg_module_122__cini_mul_v000_reg ( .D(n_and_module_59_res), .CK(
        clock_6), .Q(n_reg_module_122_res), .QN() );
  AND2_X1 u_and_module_60_U1 ( .A1(n_reg_module_62_res), .A2(io_i0_s1_d6), 
        .ZN(n_and_module_60_res) );
  XOR2_X1 u_xor_module_82_U1 ( .A(p_rand_5), .B(n_and_module_60_res), .Z(
        n_xor_module_82_res) );
  DFF_X1 u_reg_module_123__cini_mul_v000_reg ( .D(n_xor_module_82_res), .CK(
        clock_6), .Q(n_reg_module_123_res), .QN() );
  AND2_X1 u_and_module_61_U1 ( .A1(n_reg_module_57_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_61_res) );
  XOR2_X1 u_xor_module_83_U1 ( .A(p_rand_4), .B(n_and_module_61_res), .Z(
        n_xor_module_83_res) );
  DFF_X1 u_reg_module_124__cini_mul_v000_reg ( .D(n_xor_module_83_res), .CK(
        clock_6), .Q(n_reg_module_124_res), .QN() );
  AND2_X1 u_and_module_62_U1 ( .A1(n_reg_module_60_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_62_res) );
  XOR2_X1 u_xor_module_84_U1 ( .A(p_rand_5), .B(n_and_module_62_res), .Z(
        n_xor_module_84_res) );
  DFF_X1 u_reg_module_125__cini_mul_v000_reg ( .D(n_xor_module_84_res), .CK(
        clock_6), .Q(n_reg_module_125_res), .QN() );
  AND2_X1 u_and_module_63_U1 ( .A1(n_reg_module_63_res), .A2(io_i0_s2_d6), 
        .ZN(n_and_module_63_res) );
  DFF_X1 u_reg_module_126__cini_mul_v000_reg ( .D(n_and_module_63_res), .CK(
        clock_6), .Q(n_reg_module_126_res), .QN() );
  XOR2_X1 u_xor_module_85_U1 ( .A(n_reg_module_65_res), .B(n_reg_module_64_res), .Z(n_xor_module_85_res) );
  XOR2_X1 u_xor_module_86_U1 ( .A(n_reg_module_66_res), .B(n_xor_module_85_res), .Z(io_o0_s0_d0) );
  XOR2_X1 u_xor_module_87_U1 ( .A(n_reg_module_67_res), .B(n_reg_module_68_res), .Z(n_xor_module_87_res) );
  XOR2_X1 u_xor_module_88_U1 ( .A(n_reg_module_69_res), .B(n_xor_module_87_res), .Z(io_o0_s1_d0) );
  XOR2_X1 u_xor_module_89_U1 ( .A(n_reg_module_70_res), .B(n_reg_module_72_res), .Z(n_xor_module_89_res) );
  XOR2_X1 u_xor_module_90_U1 ( .A(n_reg_module_71_res), .B(n_xor_module_89_res), .Z(io_o0_s2_d0) );
  XOR2_X1 u_xor_module_91_U1 ( .A(n_reg_module_74_res), .B(n_reg_module_73_res), .Z(n_xor_module_91_res) );
  XOR2_X1 u_xor_module_92_U1 ( .A(n_reg_module_75_res), .B(n_xor_module_91_res), .Z(io_o0_s0_d1) );
  XOR2_X1 u_xor_module_93_U1 ( .A(n_reg_module_76_res), .B(n_reg_module_77_res), .Z(n_xor_module_93_res) );
  XOR2_X1 u_xor_module_94_U1 ( .A(n_reg_module_78_res), .B(n_xor_module_93_res), .Z(io_o0_s1_d1) );
  XOR2_X1 u_xor_module_95_U1 ( .A(n_reg_module_79_res), .B(n_reg_module_81_res), .Z(n_xor_module_95_res) );
  XOR2_X1 u_xor_module_96_U1 ( .A(n_reg_module_80_res), .B(n_xor_module_95_res), .Z(io_o0_s2_d1) );
  XOR2_X1 u_xor_module_97_U1 ( .A(n_reg_module_83_res), .B(n_reg_module_82_res), .Z(n_xor_module_97_res) );
  XOR2_X1 u_xor_module_98_U1 ( .A(n_reg_module_84_res), .B(n_xor_module_97_res), .Z(io_o0_s0_d2) );
  XOR2_X1 u_xor_module_99_U1 ( .A(n_reg_module_85_res), .B(n_reg_module_86_res), .Z(n_xor_module_99_res) );
  XOR2_X1 u_xor_module_100_U1 ( .A(n_reg_module_87_res), .B(
        n_xor_module_99_res), .Z(io_o0_s1_d2) );
  XOR2_X1 u_xor_module_101_U1 ( .A(n_reg_module_88_res), .B(
        n_reg_module_90_res), .Z(n_xor_module_101_res) );
  XOR2_X1 u_xor_module_102_U1 ( .A(n_reg_module_89_res), .B(
        n_xor_module_101_res), .Z(io_o0_s2_d2) );
  XOR2_X1 u_xor_module_103_U1 ( .A(n_reg_module_92_res), .B(
        n_reg_module_91_res), .Z(n_xor_module_103_res) );
  XOR2_X1 u_xor_module_104_U1 ( .A(n_reg_module_93_res), .B(
        n_xor_module_103_res), .Z(io_o0_s0_d3) );
  XOR2_X1 u_xor_module_105_U1 ( .A(n_reg_module_94_res), .B(
        n_reg_module_95_res), .Z(n_xor_module_105_res) );
  XOR2_X1 u_xor_module_106_U1 ( .A(n_reg_module_96_res), .B(
        n_xor_module_105_res), .Z(io_o0_s1_d3) );
  XOR2_X1 u_xor_module_107_U1 ( .A(n_reg_module_97_res), .B(
        n_reg_module_99_res), .Z(n_xor_module_107_res) );
  XOR2_X1 u_xor_module_108_U1 ( .A(n_reg_module_98_res), .B(
        n_xor_module_107_res), .Z(io_o0_s2_d3) );
  XOR2_X1 u_xor_module_109_U1 ( .A(n_reg_module_101_res), .B(
        n_reg_module_100_res), .Z(n_xor_module_109_res) );
  XOR2_X1 u_xor_module_110_U1 ( .A(n_reg_module_102_res), .B(
        n_xor_module_109_res), .Z(io_o0_s0_d4) );
  XOR2_X1 u_xor_module_111_U1 ( .A(n_reg_module_103_res), .B(
        n_reg_module_104_res), .Z(n_xor_module_111_res) );
  XOR2_X1 u_xor_module_112_U1 ( .A(n_reg_module_105_res), .B(
        n_xor_module_111_res), .Z(io_o0_s1_d4) );
  XOR2_X1 u_xor_module_113_U1 ( .A(n_reg_module_106_res), .B(
        n_reg_module_108_res), .Z(n_xor_module_113_res) );
  XOR2_X1 u_xor_module_114_U1 ( .A(n_reg_module_107_res), .B(
        n_xor_module_113_res), .Z(io_o0_s2_d4) );
  XOR2_X1 u_xor_module_115_U1 ( .A(n_reg_module_110_res), .B(
        n_reg_module_109_res), .Z(n_xor_module_115_res) );
  XOR2_X1 u_xor_module_116_U1 ( .A(n_reg_module_111_res), .B(
        n_xor_module_115_res), .Z(io_o0_s0_d5) );
  XOR2_X1 u_xor_module_117_U1 ( .A(n_reg_module_112_res), .B(
        n_reg_module_113_res), .Z(n_xor_module_117_res) );
  XOR2_X1 u_xor_module_118_U1 ( .A(n_reg_module_114_res), .B(
        n_xor_module_117_res), .Z(io_o0_s1_d5) );
  XOR2_X1 u_xor_module_119_U1 ( .A(n_reg_module_115_res), .B(
        n_reg_module_117_res), .Z(n_xor_module_119_res) );
  XOR2_X1 u_xor_module_120_U1 ( .A(n_reg_module_116_res), .B(
        n_xor_module_119_res), .Z(io_o0_s2_d5) );
  XOR2_X1 u_xor_module_121_U1 ( .A(n_reg_module_119_res), .B(
        n_reg_module_118_res), .Z(n_xor_module_121_res) );
  XOR2_X1 u_xor_module_122_U1 ( .A(n_reg_module_120_res), .B(
        n_xor_module_121_res), .Z(io_o0_s0_d6) );
  XOR2_X1 u_xor_module_123_U1 ( .A(n_reg_module_121_res), .B(
        n_reg_module_122_res), .Z(n_xor_module_123_res) );
  XOR2_X1 u_xor_module_124_U1 ( .A(n_reg_module_123_res), .B(
        n_xor_module_123_res), .Z(io_o0_s1_d6) );
  XOR2_X1 u_xor_module_125_U1 ( .A(n_reg_module_124_res), .B(
        n_reg_module_126_res), .Z(n_xor_module_125_res) );
  XOR2_X1 u_xor_module_126_U1 ( .A(n_reg_module_125_res), .B(
        n_xor_module_125_res), .Z(io_o0_s2_d6) );
endmodule

