
module DefaultSbox_keyAdd ( clock, reset, io_state, io_key, io_out );
  input [3:0] io_state;
  input [3:0] io_key;
  output [3:0] io_out;
  input clock, reset;
  wire   sbox_io_o0, sbox_io_o1, sbox_io_o2, sbox_io_o3, sbox_n38, sbox_n37,
         sbox_n36, sbox_n35, sbox_n34, sbox_n33, sbox_n32, sbox_n31, sbox_n30,
         sbox_n29, sbox_n28, sbox_n27, sbox_n26, sbox_n25, sbox_n24, sbox_n23,
         sbox_n22, sbox_n21, sbox_n20, sbox_n19, sbox_n18, sbox_n17, sbox_n16,
         sbox_n15, sbox_n14, sbox_n13, sbox_n12, sbox_n11, sbox_n10, sbox_n9,
         sbox_n8, sbox_n7, sbox_n6, sbox_n5, sbox_n4, sbox_n3, sbox_n2,
         sbox_n1;

  XOR2_X1 U5 ( .A(sbox_io_o3), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 U6 ( .A(sbox_io_o2), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 U7 ( .A(sbox_io_o1), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 U8 ( .A(sbox_io_o0), .B(io_key[0]), .Z(io_out[0]) );
  INV_X1 sbox_U42 ( .A(io_state[3]), .ZN(sbox_n13) );
  INV_X1 sbox_U41 ( .A(io_state[0]), .ZN(sbox_n31) );
  NAND2_X1 sbox_U40 ( .A1(sbox_n13), .A2(sbox_n31), .ZN(sbox_n38) );
  INV_X1 sbox_U39 ( .A(io_state[1]), .ZN(sbox_n18) );
  NAND2_X1 sbox_U38 ( .A1(io_state[2]), .A2(sbox_n18), .ZN(sbox_n14) );
  NOR2_X1 sbox_U37 ( .A1(sbox_n38), .A2(sbox_n14), .ZN(sbox_n20) );
  NOR2_X1 sbox_U36 ( .A1(io_state[0]), .A2(sbox_n14), .ZN(sbox_n37) );
  AND2_X1 sbox_U35 ( .A1(sbox_n37), .A2(io_state[3]), .ZN(sbox_n3) );
  NOR2_X1 sbox_U34 ( .A1(io_state[3]), .A2(io_state[2]), .ZN(sbox_n36) );
  AND2_X1 sbox_U33 ( .A1(sbox_n36), .A2(io_state[1]), .ZN(sbox_n24) );
  AND2_X1 sbox_U32 ( .A1(sbox_n24), .A2(sbox_n31), .ZN(sbox_n15) );
  NOR2_X1 sbox_U31 ( .A1(sbox_n3), .A2(sbox_n15), .ZN(sbox_n33) );
  NOR2_X1 sbox_U30 ( .A1(io_state[2]), .A2(io_state[1]), .ZN(sbox_n35) );
  NAND2_X1 sbox_U29 ( .A1(sbox_n35), .A2(io_state[0]), .ZN(sbox_n34) );
  NAND2_X1 sbox_U28 ( .A1(sbox_n33), .A2(sbox_n34), .ZN(sbox_n26) );
  NOR2_X1 sbox_U27 ( .A1(sbox_n20), .A2(sbox_n26), .ZN(sbox_n27) );
  NOR2_X1 sbox_U26 ( .A1(sbox_n13), .A2(io_state[2]), .ZN(sbox_n5) );
  NAND2_X1 sbox_U25 ( .A1(sbox_n5), .A2(io_state[1]), .ZN(sbox_n32) );
  NOR2_X1 sbox_U24 ( .A1(io_state[0]), .A2(sbox_n32), .ZN(sbox_n29) );
  NAND2_X1 sbox_U23 ( .A1(io_state[1]), .A2(io_state[2]), .ZN(sbox_n8) );
  NOR2_X1 sbox_U22 ( .A1(sbox_n31), .A2(sbox_n8), .ZN(sbox_n30) );
  NOR2_X1 sbox_U21 ( .A1(sbox_n29), .A2(sbox_n30), .ZN(sbox_n28) );
  NAND2_X1 sbox_U20 ( .A1(sbox_n27), .A2(sbox_n28), .ZN(sbox_io_o0) );
  NOR2_X1 sbox_U19 ( .A1(io_state[0]), .A2(sbox_n8), .ZN(sbox_n25) );
  NOR2_X1 sbox_U18 ( .A1(sbox_n25), .A2(sbox_n26), .ZN(sbox_n21) );
  AND2_X1 sbox_U17 ( .A1(io_state[0]), .A2(sbox_n24), .ZN(sbox_n19) );
  NOR2_X1 sbox_U16 ( .A1(sbox_n14), .A2(sbox_n13), .ZN(sbox_n23) );
  NOR2_X1 sbox_U15 ( .A1(sbox_n19), .A2(sbox_n23), .ZN(sbox_n22) );
  NAND2_X1 sbox_U14 ( .A1(sbox_n21), .A2(sbox_n22), .ZN(sbox_io_o1) );
  NOR2_X1 sbox_U13 ( .A1(sbox_n19), .A2(sbox_n20), .ZN(sbox_n16) );
  NAND2_X1 sbox_U12 ( .A1(sbox_n5), .A2(sbox_n18), .ZN(sbox_n17) );
  NAND2_X1 sbox_U11 ( .A1(sbox_n16), .A2(sbox_n17), .ZN(sbox_n7) );
  NOR2_X1 sbox_U10 ( .A1(sbox_n15), .A2(sbox_n7), .ZN(sbox_n9) );
  NOR2_X1 sbox_U9 ( .A1(io_state[3]), .A2(sbox_n14), .ZN(sbox_n11) );
  NOR2_X1 sbox_U8 ( .A1(sbox_n13), .A2(sbox_n8), .ZN(sbox_n12) );
  NOR2_X1 sbox_U7 ( .A1(sbox_n11), .A2(sbox_n12), .ZN(sbox_n10) );
  NAND2_X1 sbox_U6 ( .A1(sbox_n9), .A2(sbox_n10), .ZN(sbox_io_o2) );
  NOR2_X1 sbox_U5 ( .A1(io_state[3]), .A2(sbox_n8), .ZN(sbox_n6) );
  NOR2_X1 sbox_U4 ( .A1(sbox_n6), .A2(sbox_n7), .ZN(sbox_n1) );
  AND2_X1 sbox_U3 ( .A1(io_state[0]), .A2(sbox_n5), .ZN(sbox_n4) );
  NOR2_X1 sbox_U2 ( .A1(sbox_n3), .A2(sbox_n4), .ZN(sbox_n2) );
  NAND2_X1 sbox_U1 ( .A1(sbox_n1), .A2(sbox_n2), .ZN(sbox_io_o3) );
endmodule

