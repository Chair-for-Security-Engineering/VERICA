
module PresentSbox_keyAdd_detection_sifaTest ( clock, reset, io_state, io_key, 
        io_error );
  input [3:0] io_state;
  input [3:0] io_key;
  input clock, reset;
  output io_error;
  wire   n7, n8, n9, n10, n11, n12, PresentSbox_keyAdd_sbox_io_o3,
         PresentSbox_keyAdd_sbox_io_o2, PresentSbox_keyAdd_sbox_io_o1,
         PresentSbox_keyAdd_sbox_io_o0, PresentSbox_keyAdd_sbox_n18,
         PresentSbox_keyAdd_sbox_n17, PresentSbox_keyAdd_sbox_n16,
         PresentSbox_keyAdd_sbox_n15, PresentSbox_keyAdd_sbox_n14,
         PresentSbox_keyAdd_sbox_n13, PresentSbox_keyAdd_sbox_n12,
         PresentSbox_keyAdd_sbox_n11, PresentSbox_keyAdd_sbox_n10,
         PresentSbox_keyAdd_sbox_n9, PresentSbox_keyAdd_sbox_n8,
         PresentSbox_keyAdd_sbox_n7, PresentSbox_keyAdd_sbox_n6,
         PresentSbox_keyAdd_sbox_n5, PresentSbox_keyAdd_sbox_n4,
         PresentSbox_keyAdd_sbox_n3, PresentSbox_keyAdd_sbox_n2,
         PresentSbox_keyAdd_sbox_n1, PresentSbox_keyAdd_1_sbox_io_o3,
         PresentSbox_keyAdd_1_sbox_io_o2, PresentSbox_keyAdd_1_sbox_io_o1,
         PresentSbox_keyAdd_1_sbox_io_o0, PresentSbox_keyAdd_1_sbox_n18,
         PresentSbox_keyAdd_1_sbox_n17, PresentSbox_keyAdd_1_sbox_n16,
         PresentSbox_keyAdd_1_sbox_n15, PresentSbox_keyAdd_1_sbox_n14,
         PresentSbox_keyAdd_1_sbox_n13, PresentSbox_keyAdd_1_sbox_n12,
         PresentSbox_keyAdd_1_sbox_n11, PresentSbox_keyAdd_1_sbox_n10,
         PresentSbox_keyAdd_1_sbox_n9, PresentSbox_keyAdd_1_sbox_n8,
         PresentSbox_keyAdd_1_sbox_n7, PresentSbox_keyAdd_1_sbox_n6,
         PresentSbox_keyAdd_1_sbox_n5, PresentSbox_keyAdd_1_sbox_n4,
         PresentSbox_keyAdd_1_sbox_n3, PresentSbox_keyAdd_1_sbox_n2,
         PresentSbox_keyAdd_1_sbox_n1;
  wire   [3:0] output_sbox_0;
  wire   [3:0] output_sbox_1;
  wire io_state0, io_state1, io_state2, io_state3;

  BUF_X1 B00 ( .A(io_state[0]), .Z(io_state0) );
  BUF_X1 B01 ( .A(io_state[1]), .Z(io_state1) );
  BUF_X1 B02 ( .A(io_state[2]), .Z(io_state2) );
  BUF_X1 B03 ( .A(io_state[3]), .Z(io_state3) );

  NAND2_X1 det_U8 ( .A1(n7), .A2(n8), .ZN(io_error) );
  NOR2_X1 det_U9 ( .A1(n9), .A2(n10), .ZN(n8) );
  XOR2_X1 det_U10 ( .A(output_sbox_1[1]), .B(output_sbox_0[1]), .Z(n10) );
  XOR2_X1 det_U11 ( .A(output_sbox_1[0]), .B(output_sbox_0[0]), .Z(n9) );
  NOR2_X1 det_U12 ( .A1(n11), .A2(n12), .ZN(n7) );
  XOR2_X1 det_U13 ( .A(output_sbox_1[3]), .B(output_sbox_0[3]), .Z(n12) );
  XOR2_X1 det_U14 ( .A(output_sbox_1[2]), .B(output_sbox_0[2]), .Z(n11) );
  XOR2_X1 PresentSbox_keyAdd_U4 ( .A(PresentSbox_keyAdd_sbox_io_o0), .B(
        io_key[0]), .Z(output_sbox_0[0]) );
  XOR2_X1 PresentSbox_keyAdd_U3 ( .A(PresentSbox_keyAdd_sbox_io_o1), .B(
        io_key[1]), .Z(output_sbox_0[1]) );
  XOR2_X1 PresentSbox_keyAdd_U2 ( .A(PresentSbox_keyAdd_sbox_io_o2), .B(
        io_key[2]), .Z(output_sbox_0[2]) );
  XOR2_X1 PresentSbox_keyAdd_U1 ( .A(PresentSbox_keyAdd_sbox_io_o3), .B(
        io_key[3]), .Z(output_sbox_0[3]) );
  INV_X1 PresentSbox_keyAdd_sbox_U022 ( .A(io_state[1]), .ZN(
        PresentSbox_keyAdd_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U021 ( .A1(PresentSbox_keyAdd_sbox_n18), .A2(
        io_state[2]), .ZN(PresentSbox_keyAdd_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_sbox_U020 ( .A1(io_state[2]), .A2(
        PresentSbox_keyAdd_sbox_n18), .ZN(PresentSbox_keyAdd_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_sbox_U019 ( .A1(PresentSbox_keyAdd_sbox_n1), .A2(
        PresentSbox_keyAdd_sbox_n17), .ZN(PresentSbox_keyAdd_sbox_n13) );
  INV_X1 PresentSbox_keyAdd_sbox_U018 ( .A(io_state[3]), .ZN(
        PresentSbox_keyAdd_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U017 ( .A(PresentSbox_keyAdd_sbox_n13), .B(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n15) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U016 ( .A1(PresentSbox_keyAdd_sbox_n13), .A2(
        io_state[0]), .ZN(PresentSbox_keyAdd_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_sbox_U015 ( .A1(PresentSbox_keyAdd_sbox_n11), .A2(
        PresentSbox_keyAdd_sbox_n1), .ZN(PresentSbox_keyAdd_sbox_n14) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U014 ( .A(io_state[0]), .B(io_state[2]), 
        .ZN(PresentSbox_keyAdd_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U013 ( .A(PresentSbox_keyAdd_sbox_n14), .B(
        PresentSbox_keyAdd_sbox_n4), .Z(PresentSbox_keyAdd_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_sbox_U012 ( .A1(PresentSbox_keyAdd_sbox_n15), 
        .A2(PresentSbox_keyAdd_sbox_n16), .ZN(PresentSbox_keyAdd_sbox_n3) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U011 ( .A(PresentSbox_keyAdd_sbox_n14), .B(
        io_state[3]), .ZN(PresentSbox_keyAdd_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U010 ( .A(PresentSbox_keyAdd_sbox_n3), .B(
        PresentSbox_keyAdd_sbox_n6), .Z(PresentSbox_keyAdd_sbox_io_o0) );
  XNOR2_X1 PresentSbox_keyAdd_sbox_U009 ( .A(io_state[0]), .B(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U008 ( .A(PresentSbox_keyAdd_sbox_n13), .B(
        PresentSbox_keyAdd_sbox_n2), .Z(PresentSbox_keyAdd_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_sbox_U007 ( .A1(PresentSbox_keyAdd_sbox_n11), .A2(
        PresentSbox_keyAdd_sbox_n12), .ZN(PresentSbox_keyAdd_sbox_n10) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U006 ( .A(PresentSbox_keyAdd_sbox_n4), .B(
        PresentSbox_keyAdd_sbox_n10), .Z(PresentSbox_keyAdd_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_sbox_U005 ( .A1(PresentSbox_keyAdd_sbox_n8), .A2(
        PresentSbox_keyAdd_sbox_n9), .ZN(PresentSbox_keyAdd_sbox_n7) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U004 ( .A(PresentSbox_keyAdd_sbox_n7), .B(
        io_state[2]), .Z(PresentSbox_keyAdd_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U003 ( .A(PresentSbox_keyAdd_sbox_n5), .B(
        PresentSbox_keyAdd_sbox_n6), .Z(PresentSbox_keyAdd_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U002 ( .A(PresentSbox_keyAdd_sbox_n3), .B(
        PresentSbox_keyAdd_sbox_n4), .Z(PresentSbox_keyAdd_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_sbox_U001 ( .A(PresentSbox_keyAdd_sbox_n1), .B(
        PresentSbox_keyAdd_sbox_n2), .Z(PresentSbox_keyAdd_sbox_io_o3) );
  XOR2_X1 PresentSbox_keyAdd_1_U4 ( .A(PresentSbox_keyAdd_1_sbox_io_o0), .B(
        io_key[0]), .Z(output_sbox_1[0]) );
  XOR2_X1 PresentSbox_keyAdd_1_U3 ( .A(PresentSbox_keyAdd_1_sbox_io_o1), .B(
        io_key[1]), .Z(output_sbox_1[1]) );
  XOR2_X1 PresentSbox_keyAdd_1_U2 ( .A(PresentSbox_keyAdd_1_sbox_io_o2), .B(
        io_key[2]), .Z(output_sbox_1[2]) );
  XOR2_X1 PresentSbox_keyAdd_1_U1 ( .A(PresentSbox_keyAdd_1_sbox_io_o3), .B(
        io_key[3]), .Z(output_sbox_1[3]) );
  INV_X1 PresentSbox_keyAdd_1_sbox_U022 ( .A(io_state1), .ZN(
        PresentSbox_keyAdd_1_sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U021 ( .A1(PresentSbox_keyAdd_1_sbox_n18), 
        .A2(io_state2), .ZN(PresentSbox_keyAdd_1_sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_1_sbox_U020 ( .A1(io_state2), .A2(
        PresentSbox_keyAdd_1_sbox_n18), .ZN(PresentSbox_keyAdd_1_sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U019 ( .A1(PresentSbox_keyAdd_1_sbox_n1), 
        .A2(PresentSbox_keyAdd_1_sbox_n17), .ZN(PresentSbox_keyAdd_1_sbox_n13)
         );
  INV_X1 PresentSbox_keyAdd_1_sbox_U018 ( .A(io_state3), .ZN(
        PresentSbox_keyAdd_1_sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U017 ( .A(PresentSbox_keyAdd_1_sbox_n13), 
        .B(PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n15)
         );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U016 ( .A1(PresentSbox_keyAdd_1_sbox_n13), 
        .A2(io_state0), .ZN(PresentSbox_keyAdd_1_sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U015 ( .A1(PresentSbox_keyAdd_1_sbox_n11), 
        .A2(PresentSbox_keyAdd_1_sbox_n1), .ZN(PresentSbox_keyAdd_1_sbox_n14)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U014 ( .A(io_state0), .B(io_state2), 
        .ZN(PresentSbox_keyAdd_1_sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U013 ( .A(PresentSbox_keyAdd_1_sbox_n14), 
        .B(PresentSbox_keyAdd_1_sbox_n4), .Z(PresentSbox_keyAdd_1_sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U012 ( .A1(PresentSbox_keyAdd_1_sbox_n15), 
        .A2(PresentSbox_keyAdd_1_sbox_n16), .ZN(PresentSbox_keyAdd_1_sbox_n3)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U011 ( .A(PresentSbox_keyAdd_1_sbox_n14), 
        .B(io_state3), .ZN(PresentSbox_keyAdd_1_sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U010 ( .A(PresentSbox_keyAdd_1_sbox_n3), 
        .B(PresentSbox_keyAdd_1_sbox_n6), .Z(PresentSbox_keyAdd_1_sbox_io_o0)
         );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U009 ( .A(io_state0), .B(
        PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U008 ( .A(PresentSbox_keyAdd_1_sbox_n13), 
        .B(PresentSbox_keyAdd_1_sbox_n2), .Z(PresentSbox_keyAdd_1_sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U007 ( .A1(PresentSbox_keyAdd_1_sbox_n11), 
        .A2(PresentSbox_keyAdd_1_sbox_n12), .ZN(PresentSbox_keyAdd_1_sbox_n10)
         );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U006 ( .A(PresentSbox_keyAdd_1_sbox_n4), .B(
        PresentSbox_keyAdd_1_sbox_n10), .Z(PresentSbox_keyAdd_1_sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U005 ( .A1(PresentSbox_keyAdd_1_sbox_n8), 
        .A2(PresentSbox_keyAdd_1_sbox_n9), .ZN(PresentSbox_keyAdd_1_sbox_n7)
         );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U004 ( .A(PresentSbox_keyAdd_1_sbox_n7), .B(
        io_state2), .Z(PresentSbox_keyAdd_1_sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U003 ( .A(PresentSbox_keyAdd_1_sbox_n5), .B(
        PresentSbox_keyAdd_1_sbox_n6), .Z(PresentSbox_keyAdd_1_sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U002 ( .A(PresentSbox_keyAdd_1_sbox_n3), .B(
        PresentSbox_keyAdd_1_sbox_n4), .Z(PresentSbox_keyAdd_1_sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U001 ( .A(PresentSbox_keyAdd_1_sbox_n1), .B(
        PresentSbox_keyAdd_1_sbox_n2), .Z(PresentSbox_keyAdd_1_sbox_io_o3) );
endmodule

