
module andSININA ( port_a_0, port_a_1, port_b_0, port_b_1, port_c_0, port_c_1, 
        port_r, clk, reset );
  input [2:0] port_a_0;
  input [2:0] port_a_1;
  input [2:0] port_b_0;
  input [2:0] port_b_1;
  output [2:0] port_c_0;
  output [2:0] port_c_1;
  input [1:0] port_r;
  input clk, reset;
  wire   mul_n12, mul_n11, mul_n10, mul_n9, mul_n8, mul_n7, mul_n6, mul_n5,
         mul_n4, mul_n3, mul_n2, mul_n1, mul_N13, mul_N12, mul_N11, mul_N10,
         mul_N9, mul_N8, cor_maj_23_port_o, cor_maj_22_port_o,
         cor_maj_21_port_o, cor_maj_20_port_o, cor_maj_19_port_o,
         cor_maj_18_port_o, cor_maj_17_port_o, cor_maj_16_port_o,
         cor_maj_15_port_o, cor_maj_14_port_o, cor_maj_13_port_o,
         cor_maj_12_port_o, cor_maj_12_n3, cor_maj_12_n2, cor_maj_12_n1,
         cor_maj_13_n6, cor_maj_13_n5, cor_maj_13_n4, cor_maj_14_n6,
         cor_maj_14_n5, cor_maj_14_n4, cor_maj_15_n6, cor_maj_15_n5,
         cor_maj_15_n4, cor_maj_16_n6, cor_maj_16_n5, cor_maj_16_n4,
         cor_maj_17_n6, cor_maj_17_n5, cor_maj_17_n4, cor_maj_18_n6,
         cor_maj_18_n5, cor_maj_18_n4, cor_maj_19_n6, cor_maj_19_n5,
         cor_maj_19_n4, cor_maj_20_n6, cor_maj_20_n5, cor_maj_20_n4,
         cor_maj_21_n6, cor_maj_21_n5, cor_maj_21_n4, cor_maj_22_n6,
         cor_maj_22_n5, cor_maj_22_n4, cor_maj_23_n6, cor_maj_23_n5,
         cor_maj_23_n4;
  wire   [2:0] mul_port_c_0_0;
  wire   [2:0] mul_port_c_0_1;
  wire   [2:0] mul_port_c_1_0;
  wire   [2:0] mul_port_c_1_1;
  wire   [2:0] cor_port_v_0_0;
  wire   [2:0] cor_port_v_0_1;
  wire   [2:0] cor_port_v_1_0;
  wire   [2:0] cor_port_v_1_1;
  wire   [2:0] comp_port_c_0;
  wire   [2:0] comp_port_c_1;
  wire   [2:0] mul_xor2_7_port_z;
  wire   [2:0] mul_xor2_6_port_z;
  wire   [2:0] mul_xor2_6_port_a0;
  wire   [2:0] mul_xor2_5_port_z;
  wire   [2:0] mul_xor2_4_port_z;
  wire   [2:0] mul_xor2_4_port_a0;
  wire wire0, wire1, wire2, wire3, wire4, wire5, wire6, wire7, wire8, wire9, wire10, wire11, wire12, wire13, wire14, wire15, wire16, wire17, wire18, wire19, wire20, wire21, wire22, wire23, wire24, wire25, wire26, wire27, wire28, wire29, wire30, wire31, wire32, wire33, wire34, wire35, wire36, wire37, wire38, wire39, wire40, wire41, wire42, wire43, wire44, wire45, wire46, wire47, wire48, wire49, wire50, wire51, wire52, wire53, wire54, wire55, wire56, wire57, wire58, wire59, wire60, wire61, wire62, wire63, wire64, wire65, wire66, wire67, wire68, wire69, wire70, wire71, wire72, wire73, wire74, wire75, wire76, wire77, wire78, wire79, wire80, wire81, wire82, wire83, wire84, wire85, wire86, wire87, wire88, wire89, wire90, wire91, wire92, wire93, wire94, wire95;

  DFF_X1 result_0_reg_2_ ( .D(comp_port_c_0[2]), .CK(clk), .Q(port_c_0[2]), .QN() );
  DFF_X1 result_0_reg_1_ ( .D(comp_port_c_0[1]), .CK(clk), .Q(port_c_0[1]), .QN() );
  DFF_X1 result_0_reg_0_ ( .D(comp_port_c_0[0]), .CK(clk), .Q(port_c_0[0]), .QN() );
  DFF_X1 result_1_reg_2_ ( .D(comp_port_c_1[2]), .CK(clk), .Q(port_c_1[2]), .QN() );
  DFF_X1 result_1_reg_1_ ( .D(comp_port_c_1[1]), .CK(clk), .Q(port_c_1[1]), .QN() );
  DFF_X1 result_1_reg_0_ ( .D(comp_port_c_1[0]), .CK(clk), .Q(port_c_1[0]), .QN() );
  INV_X1 mul_U26 ( .A(port_a_1[2]), .ZN(mul_n4) );
  INV_X1 mul_U25 ( .A(port_a_1[1]), .ZN(mul_n5) );
  INV_X1 mul_U24 ( .A(port_a_1[0]), .ZN(mul_n6) );
  INV_X1 mul_U23 ( .A(port_a_0[2]), .ZN(mul_n1) );
  INV_X1 mul_U22 ( .A(port_a_0[1]), .ZN(mul_n2) );
  INV_X1 mul_U21 ( .A(port_a_0[0]), .ZN(mul_n3) );
  INV_X1 mul_U20 ( .A(port_b_0[2]), .ZN(mul_n7) );
  INV_X1 mul_U19 ( .A(port_b_0[1]), .ZN(mul_n8) );
  INV_X1 mul_U18 ( .A(port_b_0[0]), .ZN(mul_n9) );
  INV_X1 mul_U17 ( .A(port_b_1[2]), .ZN(mul_n10) );
  INV_X1 mul_U16 ( .A(port_b_1[1]), .ZN(mul_n11) );
  INV_X1 mul_U15 ( .A(port_b_1[0]), .ZN(mul_n12) );
  INV_X1 mul_U14_0 (.A(mul_n1), .ZN(wire0)); 
  INV_X1 mul_U14_1 (.A(mul_n10), .ZN(wire1)); 
  AND2_X1 mul_U14_2 ( .A1(wire0), .A2(wire1), .ZN(mul_xor2_4_port_a0[2]) ); 
  INV_X1 mul_U13_3 (.A(mul_n2), .ZN(wire2)); 
  INV_X1 mul_U13_4 (.A(mul_n11), .ZN(wire3)); 
  AND2_X1 mul_U13_5 ( .A1(wire2), .A2(wire3), .ZN(mul_xor2_4_port_a0[1]) ); 
  INV_X1 mul_U12_6 (.A(mul_n3), .ZN(wire4)); 
  INV_X1 mul_U12_7 (.A(mul_n12), .ZN(wire5)); 
  AND2_X1 mul_U12_8 ( .A1(wire4), .A2(wire5), .ZN(mul_xor2_4_port_a0[0]) ); 
  INV_X1 mul_U11_9 (.A(mul_n4), .ZN(wire6)); 
  INV_X1 mul_U11_10 (.A(mul_n7), .ZN(wire7)); 
  AND2_X1 mul_U11_11 ( .A1(wire6), .A2(wire7), .ZN(mul_xor2_6_port_a0[2]) ); 
  INV_X1 mul_U10_12 (.A(mul_n5), .ZN(wire8)); 
  INV_X1 mul_U10_13 (.A(mul_n8), .ZN(wire9)); 
  AND2_X1 mul_U10_14 ( .A1(wire8), .A2(wire9), .ZN(mul_xor2_6_port_a0[1]) ); 
  INV_X1 mul_U9_15 (.A(mul_n6), .ZN(wire10)); 
  INV_X1 mul_U9_16 (.A(mul_n9), .ZN(wire11)); 
  AND2_X1 mul_U9_17 ( .A1(wire10), .A2(wire11), .ZN(mul_xor2_6_port_a0[0]) ); 
  INV_X1 mul_U8_18 (.A(mul_n7), .ZN(wire12)); 
  INV_X1 mul_U8_19 (.A(mul_n1), .ZN(wire13)); 
  AND2_X1 mul_U8_20 ( .A1(wire12), .A2(wire13), .ZN(mul_N8) ); 
  INV_X1 mul_U7_21 (.A(mul_n8), .ZN(wire14)); 
  INV_X1 mul_U7_22 (.A(mul_n2), .ZN(wire15)); 
  AND2_X1 mul_U7_23 ( .A1(wire14), .A2(wire15), .ZN(mul_N9) ); 
  INV_X1 mul_U6_24 (.A(mul_n9), .ZN(wire16)); 
  INV_X1 mul_U6_25 (.A(mul_n3), .ZN(wire17)); 
  AND2_X1 mul_U6_26 ( .A1(wire16), .A2(wire17), .ZN(mul_N10) ); 
  INV_X1 mul_U5_27 (.A(mul_n4), .ZN(wire18)); 
  INV_X1 mul_U5_28 (.A(mul_n10), .ZN(wire19)); 
  AND2_X1 mul_U5_29 ( .A1(wire18), .A2(wire19), .ZN(mul_N11) ); 
  INV_X1 mul_U4_30 (.A(mul_n5), .ZN(wire20)); 
  INV_X1 mul_U4_31 (.A(mul_n11), .ZN(wire21)); 
  AND2_X1 mul_U4_32 ( .A1(wire20), .A2(wire21), .ZN(mul_N12) ); 
  INV_X1 mul_U3_33 (.A(mul_n6), .ZN(wire22)); 
  INV_X1 mul_U3_34 (.A(mul_n12), .ZN(wire23)); 
  AND2_X1 mul_U3_35 ( .A1(wire22), .A2(wire23), .ZN(mul_N13) ); 
  DFF_X1 mul_u_1_1_reg_0_ ( .D(mul_N13), .CK(clk), .Q(mul_port_c_1_1[0]), .QN() );
  DFF_X1 mul_u_1_1_reg_1_ ( .D(mul_N12), .CK(clk), .Q(mul_port_c_1_1[1]), .QN() );
  DFF_X1 mul_u_1_1_reg_2_ ( .D(mul_N11), .CK(clk), .Q(mul_port_c_1_1[2]), .QN() );
  DFF_X1 mul_u_1_0_reg_0_ ( .D(mul_xor2_7_port_z[0]), .CK(clk), .Q(mul_port_c_1_0[0]), .QN() );
  DFF_X1 mul_u_1_0_reg_1_ ( .D(mul_xor2_7_port_z[1]), .CK(clk), .Q(mul_port_c_1_0[1]), .QN() );
  DFF_X1 mul_u_1_0_reg_2_ ( .D(mul_xor2_7_port_z[2]), .CK(clk), .Q(mul_port_c_1_0[2]), .QN() );
  DFF_X1 mul_u_0_1_reg_0_ ( .D(mul_xor2_5_port_z[0]), .CK(clk), .Q(mul_port_c_0_1[0]), .QN() );
  DFF_X1 mul_u_0_1_reg_1_ ( .D(mul_xor2_5_port_z[1]), .CK(clk), .Q(mul_port_c_0_1[1]), .QN() );
  DFF_X1 mul_u_0_1_reg_2_ ( .D(mul_xor2_5_port_z[2]), .CK(clk), .Q(mul_port_c_0_1[2]), .QN() );
  DFF_X1 mul_u_0_0_reg_0_ ( .D(mul_N10), .CK(clk), .Q(mul_port_c_0_0[0]), .QN() );
  DFF_X1 mul_u_0_0_reg_1_ ( .D(mul_N9), .CK(clk), .Q(mul_port_c_0_0[1]), .QN());
  DFF_X1 mul_u_0_0_reg_2_ ( .D(mul_N8), .CK(clk), .Q(mul_port_c_0_0[2]), .QN());
  XOR2_X1 mul_xor2_4_U3 ( .A(port_r[0]), .B(mul_xor2_4_port_a0[2]), .Z(mul_xor2_4_port_z[2]) );
  XOR2_X1 mul_xor2_4_U2 ( .A(port_r[0]), .B(mul_xor2_4_port_a0[1]), .Z(mul_xor2_4_port_z[1]) );
  XOR2_X1 mul_xor2_4_U1 ( .A(port_r[0]), .B(mul_xor2_4_port_a0[0]), .Z(mul_xor2_4_port_z[0]) );
  XOR2_X1 mul_xor2_5_U3 ( .A(port_r[1]), .B(mul_xor2_4_port_z[2]), .Z(mul_xor2_5_port_z[2]) );
  XOR2_X1 mul_xor2_5_U2 ( .A(port_r[1]), .B(mul_xor2_4_port_z[1]), .Z(mul_xor2_5_port_z[1]) );
  XOR2_X1 mul_xor2_5_U1 ( .A(port_r[1]), .B(mul_xor2_4_port_z[0]), .Z(mul_xor2_5_port_z[0]) );
  XOR2_X1 mul_xor2_6_U3 ( .A(port_r[0]), .B(mul_xor2_6_port_a0[2]), .Z(mul_xor2_6_port_z[2]) );
  XOR2_X1 mul_xor2_6_U2 ( .A(port_r[0]), .B(mul_xor2_6_port_a0[1]), .Z(mul_xor2_6_port_z[1]) );
  XOR2_X1 mul_xor2_6_U1 ( .A(port_r[0]), .B(mul_xor2_6_port_a0[0]), .Z(mul_xor2_6_port_z[0]) );
  XOR2_X1 mul_xor2_7_U3 ( .A(port_r[1]), .B(mul_xor2_6_port_z[2]), .Z(mul_xor2_7_port_z[2]) );
  XOR2_X1 mul_xor2_7_U2 ( .A(port_r[1]), .B(mul_xor2_6_port_z[1]), .Z(mul_xor2_7_port_z[1]) );
  XOR2_X1 mul_xor2_7_U1 ( .A(port_r[1]), .B(mul_xor2_6_port_z[0]), .Z(mul_xor2_7_port_z[0]) );
  DFF_X1 cor_m_1_1_reg_0_ ( .D(cor_maj_21_port_o), .CK(clk), .Q(cor_port_v_1_1[0]), .QN() );
  DFF_X1 cor_m_1_1_reg_1_ ( .D(cor_maj_22_port_o), .CK(clk), .Q(cor_port_v_1_1[1]), .QN() );
  DFF_X1 cor_m_1_1_reg_2_ ( .D(cor_maj_23_port_o), .CK(clk), .Q(cor_port_v_1_1[2]), .QN() );
  DFF_X1 cor_m_1_0_reg_0_ ( .D(cor_maj_18_port_o), .CK(clk), .Q(cor_port_v_1_0[0]), .QN() );
  DFF_X1 cor_m_1_0_reg_1_ ( .D(cor_maj_19_port_o), .CK(clk), .Q(cor_port_v_1_0[1]), .QN() );
  DFF_X1 cor_m_1_0_reg_2_ ( .D(cor_maj_20_port_o), .CK(clk), .Q(cor_port_v_1_0[2]), .QN() );
  DFF_X1 cor_m_0_1_reg_0_ ( .D(cor_maj_15_port_o), .CK(clk), .Q(cor_port_v_0_1[0]), .QN() );
  DFF_X1 cor_m_0_1_reg_1_ ( .D(cor_maj_16_port_o), .CK(clk), .Q(cor_port_v_0_1[1]), .QN() );
  DFF_X1 cor_m_0_1_reg_2_ ( .D(cor_maj_17_port_o), .CK(clk), .Q(cor_port_v_0_1[2]), .QN() );
  DFF_X1 cor_m_0_0_reg_0_ ( .D(cor_maj_12_port_o), .CK(clk), .Q(cor_port_v_0_0[0]), .QN() );
  DFF_X1 cor_m_0_0_reg_1_ ( .D(cor_maj_13_port_o), .CK(clk), .Q(cor_port_v_0_0[1]), .QN() );
  DFF_X1 cor_m_0_0_reg_2_ ( .D(cor_maj_14_port_o), .CK(clk), .Q(cor_port_v_0_0[2]), .QN() );
  INV_X1 cor_maj_12_U4_36 (.A(mul_port_c_0_0[1]), .ZN(wire24)); 
  INV_X1 cor_maj_12_U4_37 (.A(mul_port_c_0_0[0]), .ZN(wire25)); 
  AND2_X1 cor_maj_12_U4_38 ( .A1(wire24), .A2(wire25), .ZN(wire26) ); 
  INV_X1 cor_maj_12_U4_39 (.A(wire26), .ZN(cor_maj_12_n3)); 
  AND2_X1 cor_maj_12_U3_40 ( .A1(mul_port_c_0_0[2]), .A2(cor_maj_12_n3), .ZN(wire27) ); 
  INV_X1 cor_maj_12_U3_41 (.A(wire27), .ZN(cor_maj_12_n2)); 
  AND2_X1 cor_maj_12_U2_42 ( .A1(mul_port_c_0_0[1]), .A2(mul_port_c_0_0[0]), .ZN(wire28) ); 
  INV_X1 cor_maj_12_U2_43 (.A(wire28), .ZN(cor_maj_12_n1)); 
  AND2_X1 cor_maj_12_U1_44 ( .A1(cor_maj_12_n1), .A2(cor_maj_12_n2), .ZN(wire29) ); 
  INV_X1 cor_maj_12_U1_45 (.A(wire29), .ZN(cor_maj_12_port_o)); 
  INV_X1 cor_maj_13_U4_46 (.A(mul_port_c_0_0[1]), .ZN(wire30)); 
  INV_X1 cor_maj_13_U4_47 (.A(mul_port_c_0_0[0]), .ZN(wire31)); 
  AND2_X1 cor_maj_13_U4_48 ( .A1(wire30), .A2(wire31), .ZN(wire32) ); 
  INV_X1 cor_maj_13_U4_49 (.A(wire32), .ZN(cor_maj_13_n4)); 
  AND2_X1 cor_maj_13_U3_50 ( .A1(mul_port_c_0_0[2]), .A2(cor_maj_13_n4), .ZN(wire33) ); 
  INV_X1 cor_maj_13_U3_51 (.A(wire33), .ZN(cor_maj_13_n5)); 
  AND2_X1 cor_maj_13_U2_52 ( .A1(mul_port_c_0_0[1]), .A2(mul_port_c_0_0[0]), .ZN(wire34) ); 
  INV_X1 cor_maj_13_U2_53 (.A(wire34), .ZN(cor_maj_13_n6)); 
  AND2_X1 cor_maj_13_U1_54 ( .A1(cor_maj_13_n6), .A2(cor_maj_13_n5), .ZN(wire35) ); 
  INV_X1 cor_maj_13_U1_55 (.A(wire35), .ZN(cor_maj_13_port_o)); 
  INV_X1 cor_maj_14_U4_56 (.A(mul_port_c_0_0[1]), .ZN(wire36)); 
  INV_X1 cor_maj_14_U4_57 (.A(mul_port_c_0_0[0]), .ZN(wire37)); 
  AND2_X1 cor_maj_14_U4_58 ( .A1(wire36), .A2(wire37), .ZN(wire38) ); 
  INV_X1 cor_maj_14_U4_59 (.A(wire38), .ZN(cor_maj_14_n4)); 
  AND2_X1 cor_maj_14_U3_60 ( .A1(mul_port_c_0_0[2]), .A2(cor_maj_14_n4), .ZN(wire39) ); 
  INV_X1 cor_maj_14_U3_61 (.A(wire39), .ZN(cor_maj_14_n5)); 
  AND2_X1 cor_maj_14_U2_62 ( .A1(mul_port_c_0_0[1]), .A2(mul_port_c_0_0[0]), .ZN(wire40) ); 
  INV_X1 cor_maj_14_U2_63 (.A(wire40), .ZN(cor_maj_14_n6)); 
  AND2_X1 cor_maj_14_U1_64 ( .A1(cor_maj_14_n6), .A2(cor_maj_14_n5), .ZN(wire41) ); 
  INV_X1 cor_maj_14_U1_65 (.A(wire41), .ZN(cor_maj_14_port_o)); 
  INV_X1 cor_maj_15_U4_66 (.A(mul_port_c_0_1[1]), .ZN(wire42)); 
  INV_X1 cor_maj_15_U4_67 (.A(mul_port_c_0_1[0]), .ZN(wire43)); 
  AND2_X1 cor_maj_15_U4_68 ( .A1(wire42), .A2(wire43), .ZN(wire44) ); 
  INV_X1 cor_maj_15_U4_69 (.A(wire44), .ZN(cor_maj_15_n4)); 
  AND2_X1 cor_maj_15_U3_70 ( .A1(mul_port_c_0_1[2]), .A2(cor_maj_15_n4), .ZN(wire45) ); 
  INV_X1 cor_maj_15_U3_71 (.A(wire45), .ZN(cor_maj_15_n5)); 
  AND2_X1 cor_maj_15_U2_72 ( .A1(mul_port_c_0_1[1]), .A2(mul_port_c_0_1[0]), .ZN(wire46) ); 
  INV_X1 cor_maj_15_U2_73 (.A(wire46), .ZN(cor_maj_15_n6)); 
  AND2_X1 cor_maj_15_U1_74 ( .A1(cor_maj_15_n6), .A2(cor_maj_15_n5), .ZN(wire47) ); 
  INV_X1 cor_maj_15_U1_75 (.A(wire47), .ZN(cor_maj_15_port_o)); 
  INV_X1 cor_maj_16_U4_76 (.A(mul_port_c_0_1[1]), .ZN(wire48)); 
  INV_X1 cor_maj_16_U4_77 (.A(mul_port_c_0_1[0]), .ZN(wire49)); 
  AND2_X1 cor_maj_16_U4_78 ( .A1(wire48), .A2(wire49), .ZN(wire50) ); 
  INV_X1 cor_maj_16_U4_79 (.A(wire50), .ZN(cor_maj_16_n4)); 
  AND2_X1 cor_maj_16_U3_80 ( .A1(mul_port_c_0_1[2]), .A2(cor_maj_16_n4), .ZN(wire51) ); 
  INV_X1 cor_maj_16_U3_81 (.A(wire51), .ZN(cor_maj_16_n5)); 
  AND2_X1 cor_maj_16_U2_82 ( .A1(mul_port_c_0_1[1]), .A2(mul_port_c_0_1[0]), .ZN(wire52) ); 
  INV_X1 cor_maj_16_U2_83 (.A(wire52), .ZN(cor_maj_16_n6)); 
  AND2_X1 cor_maj_16_U1_84 ( .A1(cor_maj_16_n6), .A2(cor_maj_16_n5), .ZN(wire53) ); 
  INV_X1 cor_maj_16_U1_85 (.A(wire53), .ZN(cor_maj_16_port_o)); 
  INV_X1 cor_maj_17_U4_86 (.A(mul_port_c_0_1[1]), .ZN(wire54)); 
  INV_X1 cor_maj_17_U4_87 (.A(mul_port_c_0_1[0]), .ZN(wire55)); 
  AND2_X1 cor_maj_17_U4_88 ( .A1(wire54), .A2(wire55), .ZN(wire56) ); 
  INV_X1 cor_maj_17_U4_89 (.A(wire56), .ZN(cor_maj_17_n4)); 
  AND2_X1 cor_maj_17_U3_90 ( .A1(mul_port_c_0_1[2]), .A2(cor_maj_17_n4), .ZN(wire57) ); 
  INV_X1 cor_maj_17_U3_91 (.A(wire57), .ZN(cor_maj_17_n5)); 
  AND2_X1 cor_maj_17_U2_92 ( .A1(mul_port_c_0_1[1]), .A2(mul_port_c_0_1[0]), .ZN(wire58) ); 
  INV_X1 cor_maj_17_U2_93 (.A(wire58), .ZN(cor_maj_17_n6)); 
  AND2_X1 cor_maj_17_U1_94 ( .A1(cor_maj_17_n6), .A2(cor_maj_17_n5), .ZN(wire59) ); 
  INV_X1 cor_maj_17_U1_95 (.A(wire59), .ZN(cor_maj_17_port_o)); 
  INV_X1 cor_maj_18_U4_96 (.A(mul_port_c_1_0[1]), .ZN(wire60)); 
  INV_X1 cor_maj_18_U4_97 (.A(mul_port_c_1_0[0]), .ZN(wire61)); 
  AND2_X1 cor_maj_18_U4_98 ( .A1(wire60), .A2(wire61), .ZN(wire62) ); 
  INV_X1 cor_maj_18_U4_99 (.A(wire62), .ZN(cor_maj_18_n4)); 
  AND2_X1 cor_maj_18_U3_100 ( .A1(mul_port_c_1_0[2]), .A2(cor_maj_18_n4), .ZN(wire63) ); 
  INV_X1 cor_maj_18_U3_101 (.A(wire63), .ZN(cor_maj_18_n5)); 
  AND2_X1 cor_maj_18_U2_102 ( .A1(mul_port_c_1_0[1]), .A2(mul_port_c_1_0[0]), .ZN(wire64) ); 
  INV_X1 cor_maj_18_U2_103 (.A(wire64), .ZN(cor_maj_18_n6)); 
  AND2_X1 cor_maj_18_U1_104 ( .A1(cor_maj_18_n6), .A2(cor_maj_18_n5), .ZN(wire65) ); 
  INV_X1 cor_maj_18_U1_105 (.A(wire65), .ZN(cor_maj_18_port_o)); 
  INV_X1 cor_maj_19_U4_106 (.A(mul_port_c_1_0[1]), .ZN(wire66)); 
  INV_X1 cor_maj_19_U4_107 (.A(mul_port_c_1_0[0]), .ZN(wire67)); 
  AND2_X1 cor_maj_19_U4_108 ( .A1(wire66), .A2(wire67), .ZN(wire68) ); 
  INV_X1 cor_maj_19_U4_109 (.A(wire68), .ZN(cor_maj_19_n4)); 
  AND2_X1 cor_maj_19_U3_110 ( .A1(mul_port_c_1_0[2]), .A2(cor_maj_19_n4), .ZN(wire69) ); 
  INV_X1 cor_maj_19_U3_111 (.A(wire69), .ZN(cor_maj_19_n5)); 
  AND2_X1 cor_maj_19_U2_112 ( .A1(mul_port_c_1_0[1]), .A2(mul_port_c_1_0[0]), .ZN(wire70) ); 
  INV_X1 cor_maj_19_U2_113 (.A(wire70), .ZN(cor_maj_19_n6)); 
  AND2_X1 cor_maj_19_U1_114 ( .A1(cor_maj_19_n6), .A2(cor_maj_19_n5), .ZN(wire71) ); 
  INV_X1 cor_maj_19_U1_115 (.A(wire71), .ZN(cor_maj_19_port_o)); 
  INV_X1 cor_maj_20_U4_116 (.A(mul_port_c_1_0[1]), .ZN(wire72)); 
  INV_X1 cor_maj_20_U4_117 (.A(mul_port_c_1_0[0]), .ZN(wire73)); 
  AND2_X1 cor_maj_20_U4_118 ( .A1(wire72), .A2(wire73), .ZN(wire74) ); 
  INV_X1 cor_maj_20_U4_119 (.A(wire74), .ZN(cor_maj_20_n4)); 
  AND2_X1 cor_maj_20_U3_120 ( .A1(mul_port_c_1_0[2]), .A2(cor_maj_20_n4), .ZN(wire75) ); 
  INV_X1 cor_maj_20_U3_121 (.A(wire75), .ZN(cor_maj_20_n5)); 
  AND2_X1 cor_maj_20_U2_122 ( .A1(mul_port_c_1_0[1]), .A2(mul_port_c_1_0[0]), .ZN(wire76) ); 
  INV_X1 cor_maj_20_U2_123 (.A(wire76), .ZN(cor_maj_20_n6)); 
  AND2_X1 cor_maj_20_U1_124 ( .A1(cor_maj_20_n6), .A2(cor_maj_20_n5), .ZN(wire77) ); 
  INV_X1 cor_maj_20_U1_125 (.A(wire77), .ZN(cor_maj_20_port_o)); 
  INV_X1 cor_maj_21_U4_126 (.A(mul_port_c_1_1[1]), .ZN(wire78)); 
  INV_X1 cor_maj_21_U4_127 (.A(mul_port_c_1_1[0]), .ZN(wire79)); 
  AND2_X1 cor_maj_21_U4_128 ( .A1(wire78), .A2(wire79), .ZN(wire80) ); 
  INV_X1 cor_maj_21_U4_129 (.A(wire80), .ZN(cor_maj_21_n4)); 
  AND2_X1 cor_maj_21_U3_130 ( .A1(mul_port_c_1_1[2]), .A2(cor_maj_21_n4), .ZN(wire81) ); 
  INV_X1 cor_maj_21_U3_131 (.A(wire81), .ZN(cor_maj_21_n5)); 
  AND2_X1 cor_maj_21_U2_132 ( .A1(mul_port_c_1_1[1]), .A2(mul_port_c_1_1[0]), .ZN(wire82) ); 
  INV_X1 cor_maj_21_U2_133 (.A(wire82), .ZN(cor_maj_21_n6)); 
  AND2_X1 cor_maj_21_U1_134 ( .A1(cor_maj_21_n6), .A2(cor_maj_21_n5), .ZN(wire83) ); 
  INV_X1 cor_maj_21_U1_135 (.A(wire83), .ZN(cor_maj_21_port_o)); 
  INV_X1 cor_maj_22_U4_136 (.A(mul_port_c_1_1[1]), .ZN(wire84)); 
  INV_X1 cor_maj_22_U4_137 (.A(mul_port_c_1_1[0]), .ZN(wire85)); 
  AND2_X1 cor_maj_22_U4_138 ( .A1(wire84), .A2(wire85), .ZN(wire86) ); 
  INV_X1 cor_maj_22_U4_139 (.A(wire86), .ZN(cor_maj_22_n4)); 
  AND2_X1 cor_maj_22_U3_140 ( .A1(mul_port_c_1_1[2]), .A2(cor_maj_22_n4), .ZN(wire87) ); 
  INV_X1 cor_maj_22_U3_141 (.A(wire87), .ZN(cor_maj_22_n5)); 
  AND2_X1 cor_maj_22_U2_142 ( .A1(mul_port_c_1_1[1]), .A2(mul_port_c_1_1[0]), .ZN(wire88) ); 
  INV_X1 cor_maj_22_U2_143 (.A(wire88), .ZN(cor_maj_22_n6)); 
  AND2_X1 cor_maj_22_U1_144 ( .A1(cor_maj_22_n6), .A2(cor_maj_22_n5), .ZN(wire89) ); 
  INV_X1 cor_maj_22_U1_145 (.A(wire89), .ZN(cor_maj_22_port_o)); 
  INV_X1 cor_maj_23_U4_146 (.A(mul_port_c_1_1[1]), .ZN(wire90)); 
  INV_X1 cor_maj_23_U4_147 (.A(mul_port_c_1_1[0]), .ZN(wire91)); 
  AND2_X1 cor_maj_23_U4_148 ( .A1(wire90), .A2(wire91), .ZN(wire92) ); 
  INV_X1 cor_maj_23_U4_149 (.A(wire92), .ZN(cor_maj_23_n4)); 
  AND2_X1 cor_maj_23_U3_150 ( .A1(mul_port_c_1_1[2]), .A2(cor_maj_23_n4), .ZN(wire93) ); 
  INV_X1 cor_maj_23_U3_151 (.A(wire93), .ZN(cor_maj_23_n5)); 
  AND2_X1 cor_maj_23_U2_152 ( .A1(mul_port_c_1_1[1]), .A2(mul_port_c_1_1[0]), .ZN(wire94) ); 
  INV_X1 cor_maj_23_U2_153 (.A(wire94), .ZN(cor_maj_23_n6)); 
  AND2_X1 cor_maj_23_U1_154 ( .A1(cor_maj_23_n6), .A2(cor_maj_23_n5), .ZN(wire95) ); 
  INV_X1 cor_maj_23_U1_155 (.A(wire95), .ZN(cor_maj_23_port_o)); 
  XOR2_X1 comp_U6 ( .A(cor_port_v_0_1[2]), .B(cor_port_v_0_0[2]), .Z(comp_port_c_0[2]) );
  XOR2_X1 comp_U5 ( .A(cor_port_v_0_1[1]), .B(cor_port_v_0_0[1]), .Z(comp_port_c_0[1]) );
  XOR2_X1 comp_U4 ( .A(cor_port_v_0_1[0]), .B(cor_port_v_0_0[0]), .Z(comp_port_c_0[0]) );
  XOR2_X1 comp_U3 ( .A(cor_port_v_1_1[2]), .B(cor_port_v_1_0[2]), .Z(comp_port_c_1[2]) );
  XOR2_X1 comp_U2 ( .A(cor_port_v_1_1[1]), .B(cor_port_v_1_0[1]), .Z(comp_port_c_1[1]) );
  XOR2_X1 comp_U1 ( .A(cor_port_v_1_1[0]), .B(cor_port_v_1_0[0]), .Z(comp_port_c_1[0]) );
endmodule

