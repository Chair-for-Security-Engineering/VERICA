module PresentSbox_keyAdd ( clock, reset, io_state, io_key, io_out );
  input [3:0] io_state;
  input [3:0] io_key;
  output [3:0] io_out;
  input clock, reset;
  wire   sbox_io_o0, sbox_io_o1, sbox_io_o2, sbox_io_o3, sbox_n18, sbox_n17,
         sbox_n16, sbox_n15, sbox_n14, sbox_n13, sbox_n12, sbox_n11, sbox_n10,
         sbox_n9, sbox_n8, sbox_n7, sbox_n6, sbox_n5, sbox_n4, sbox_n3,
         sbox_n2, sbox_n1;
  wire io_state0, io_state1, io_state2, io_state3;

  BUF_X1 B00 ( .A(io_state[0]), .Z(io_state0) );
  BUF_X1 B01 ( .A(io_state[1]), .Z(io_state1) );
  BUF_X1 B02 ( .A(io_state[2]), .Z(io_state2) );
  BUF_X1 B03 ( .A(io_state[3]), .Z(io_state3) );

  XOR2_X1 PresentSbox_keyAdd_U1 ( .A(sbox_io_o3), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 PresentSbox_keyAdd_U2 ( .A(sbox_io_o2), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 PresentSbox_keyAdd_U3 ( .A(sbox_io_o1), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 PresentSbox_keyAdd_U4 ( .A(sbox_io_o0), .B(io_key[0]), .Z(io_out[0]) );
  INV_X1 PresentSbox_keyAdd_1_sbox_U022 ( .A(io_state1), .ZN(sbox_n18) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U021 ( .A1(sbox_n18), .A2(io_state2), .ZN(sbox_n1) );
  AND2_X1 PresentSbox_keyAdd_1_sbox_U020 ( .A1(io_state2), .A2(sbox_n18), .ZN(sbox_n17) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U019 ( .A1(sbox_n1), .A2(sbox_n17), .ZN(sbox_n13) );
  INV_X1 PresentSbox_keyAdd_1_sbox_U018 ( .A(io_state3), .ZN(sbox_n12) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U017 ( .A(sbox_n13), .B(sbox_n12), .ZN(sbox_n15) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U016 ( .A1(sbox_n13), .A2(io_state0), .ZN(sbox_n11) );
  OR2_X1 PresentSbox_keyAdd_1_sbox_U015 ( .A1(sbox_n11), .A2(sbox_n1), .ZN(sbox_n14) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U014 ( .A(io_state0), .B(io_state2), .ZN(sbox_n4) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U013 ( .A(sbox_n14), .B(sbox_n4), .Z(sbox_n16) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U012 ( .A1(sbox_n15), .A2(sbox_n16), .ZN(sbox_n3) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U011 ( .A(sbox_n14), .B(io_state3), .ZN(sbox_n6) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U010 ( .A(sbox_n3), .B(sbox_n6), .Z(sbox_io_o0) );
  XNOR2_X1 PresentSbox_keyAdd_1_sbox_U009 ( .A(io_state0), .B(sbox_n12), .ZN(sbox_n2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U008 ( .A(sbox_n13), .B(sbox_n2), .Z(sbox_n8) );
  NOR2_X1 PresentSbox_keyAdd_1_sbox_U007 ( .A1(sbox_n11), .A2(sbox_n12), .ZN(sbox_n10) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U006 ( .A(sbox_n4), .B(sbox_n10), .Z(sbox_n9) );
  NAND2_X1 PresentSbox_keyAdd_1_sbox_U005 ( .A1(sbox_n8), .A2(sbox_n9), .ZN(sbox_n7) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U004 ( .A(sbox_n7), .B(io_state2), .Z(sbox_n5) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U003 ( .A(sbox_n5), .B(sbox_n6), .Z(sbox_io_o1) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U002 ( .A(sbox_n3), .B(sbox_n4), .Z(sbox_io_o2) );
  XOR2_X1 PresentSbox_keyAdd_1_sbox_U00PresentSbox_keyAdd_1_sbox_U0221 ( .A(sbox_n1), .B(sbox_n2), .Z(sbox_io_o3) );
endmodule