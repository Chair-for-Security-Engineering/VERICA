
module AesSbox_keyAdd_detection ( clock, reset, io_state, io_key, io_out, 
        io_error );
  input [7:0] io_state;
  input [7:0] io_key;
  output [7:0] io_out;
  input clock, reset;
  output io_error;
  wire   n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, AesSbox_keyAdd_sbox_io_o7,
         AesSbox_keyAdd_sbox_io_o6, AesSbox_keyAdd_sbox_io_o5,
         AesSbox_keyAdd_sbox_io_o4, AesSbox_keyAdd_sbox_io_o3,
         AesSbox_keyAdd_sbox_io_o2, AesSbox_keyAdd_sbox_io_o1,
         AesSbox_keyAdd_sbox_io_o0, AesSbox_keyAdd_sbox_n128,
         AesSbox_keyAdd_sbox_n127, AesSbox_keyAdd_sbox_n126,
         AesSbox_keyAdd_sbox_n125, AesSbox_keyAdd_sbox_n124,
         AesSbox_keyAdd_sbox_n123, AesSbox_keyAdd_sbox_n122,
         AesSbox_keyAdd_sbox_n121, AesSbox_keyAdd_sbox_n120,
         AesSbox_keyAdd_sbox_n119, AesSbox_keyAdd_sbox_n118,
         AesSbox_keyAdd_sbox_n117, AesSbox_keyAdd_sbox_n116,
         AesSbox_keyAdd_sbox_n115, AesSbox_keyAdd_sbox_n114,
         AesSbox_keyAdd_sbox_n113, AesSbox_keyAdd_sbox_n112,
         AesSbox_keyAdd_sbox_n111, AesSbox_keyAdd_sbox_n110,
         AesSbox_keyAdd_sbox_n109, AesSbox_keyAdd_sbox_n108,
         AesSbox_keyAdd_sbox_n107, AesSbox_keyAdd_sbox_n106,
         AesSbox_keyAdd_sbox_n105, AesSbox_keyAdd_sbox_n104,
         AesSbox_keyAdd_sbox_n103, AesSbox_keyAdd_sbox_n102,
         AesSbox_keyAdd_sbox_n101, AesSbox_keyAdd_sbox_n100,
         AesSbox_keyAdd_sbox_n99, AesSbox_keyAdd_sbox_n98,
         AesSbox_keyAdd_sbox_n97, AesSbox_keyAdd_sbox_n96,
         AesSbox_keyAdd_sbox_n95, AesSbox_keyAdd_sbox_n94,
         AesSbox_keyAdd_sbox_n93, AesSbox_keyAdd_sbox_n92,
         AesSbox_keyAdd_sbox_n91, AesSbox_keyAdd_sbox_n90,
         AesSbox_keyAdd_sbox_n89, AesSbox_keyAdd_sbox_n88,
         AesSbox_keyAdd_sbox_n87, AesSbox_keyAdd_sbox_n86,
         AesSbox_keyAdd_sbox_n85, AesSbox_keyAdd_sbox_n84,
         AesSbox_keyAdd_sbox_n83, AesSbox_keyAdd_sbox_n82,
         AesSbox_keyAdd_sbox_n81, AesSbox_keyAdd_sbox_n80,
         AesSbox_keyAdd_sbox_n79, AesSbox_keyAdd_sbox_n78,
         AesSbox_keyAdd_sbox_n77, AesSbox_keyAdd_sbox_n76,
         AesSbox_keyAdd_sbox_n75, AesSbox_keyAdd_sbox_n74,
         AesSbox_keyAdd_sbox_n73, AesSbox_keyAdd_sbox_n72,
         AesSbox_keyAdd_sbox_n71, AesSbox_keyAdd_sbox_n70,
         AesSbox_keyAdd_sbox_n69, AesSbox_keyAdd_sbox_n68,
         AesSbox_keyAdd_sbox_n67, AesSbox_keyAdd_sbox_n66,
         AesSbox_keyAdd_sbox_n65, AesSbox_keyAdd_sbox_n64,
         AesSbox_keyAdd_sbox_n63, AesSbox_keyAdd_sbox_n62,
         AesSbox_keyAdd_sbox_n61, AesSbox_keyAdd_sbox_n60,
         AesSbox_keyAdd_sbox_n59, AesSbox_keyAdd_sbox_n58,
         AesSbox_keyAdd_sbox_n57, AesSbox_keyAdd_sbox_n56,
         AesSbox_keyAdd_sbox_n55, AesSbox_keyAdd_sbox_n54,
         AesSbox_keyAdd_sbox_n53, AesSbox_keyAdd_sbox_n52,
         AesSbox_keyAdd_sbox_n51, AesSbox_keyAdd_sbox_n50,
         AesSbox_keyAdd_sbox_n49, AesSbox_keyAdd_sbox_n48,
         AesSbox_keyAdd_sbox_n47, AesSbox_keyAdd_sbox_n46,
         AesSbox_keyAdd_sbox_n45, AesSbox_keyAdd_sbox_n44,
         AesSbox_keyAdd_sbox_n43, AesSbox_keyAdd_sbox_n42,
         AesSbox_keyAdd_sbox_n41, AesSbox_keyAdd_sbox_n40,
         AesSbox_keyAdd_sbox_n39, AesSbox_keyAdd_sbox_n38,
         AesSbox_keyAdd_sbox_n37, AesSbox_keyAdd_sbox_n36,
         AesSbox_keyAdd_sbox_n35, AesSbox_keyAdd_sbox_n34,
         AesSbox_keyAdd_sbox_n33, AesSbox_keyAdd_sbox_n32,
         AesSbox_keyAdd_sbox_n31, AesSbox_keyAdd_sbox_n30,
         AesSbox_keyAdd_sbox_n29, AesSbox_keyAdd_sbox_n28,
         AesSbox_keyAdd_sbox_n27, AesSbox_keyAdd_sbox_n26,
         AesSbox_keyAdd_sbox_n25, AesSbox_keyAdd_sbox_n24,
         AesSbox_keyAdd_sbox_n23, AesSbox_keyAdd_sbox_n22,
         AesSbox_keyAdd_sbox_n21, AesSbox_keyAdd_sbox_n20,
         AesSbox_keyAdd_sbox_n19, AesSbox_keyAdd_sbox_n18,
         AesSbox_keyAdd_sbox_n17, AesSbox_keyAdd_sbox_n16,
         AesSbox_keyAdd_sbox_n15, AesSbox_keyAdd_sbox_n14,
         AesSbox_keyAdd_sbox_n13, AesSbox_keyAdd_sbox_n12,
         AesSbox_keyAdd_sbox_n11, AesSbox_keyAdd_sbox_n10,
         AesSbox_keyAdd_sbox_n9, AesSbox_keyAdd_sbox_n8,
         AesSbox_keyAdd_sbox_n7, AesSbox_keyAdd_sbox_n6,
         AesSbox_keyAdd_sbox_n5, AesSbox_keyAdd_sbox_n4,
         AesSbox_keyAdd_sbox_n3, AesSbox_keyAdd_sbox_n2,
         AesSbox_keyAdd_sbox_n1, AesSbox_keyAdd_1_sbox_io_o7,
         AesSbox_keyAdd_1_sbox_io_o6, AesSbox_keyAdd_1_sbox_io_o5,
         AesSbox_keyAdd_1_sbox_io_o4, AesSbox_keyAdd_1_sbox_io_o3,
         AesSbox_keyAdd_1_sbox_io_o2, AesSbox_keyAdd_1_sbox_io_o1,
         AesSbox_keyAdd_1_sbox_io_o0, AesSbox_keyAdd_1_sbox_n128,
         AesSbox_keyAdd_1_sbox_n127, AesSbox_keyAdd_1_sbox_n126,
         AesSbox_keyAdd_1_sbox_n125, AesSbox_keyAdd_1_sbox_n124,
         AesSbox_keyAdd_1_sbox_n123, AesSbox_keyAdd_1_sbox_n122,
         AesSbox_keyAdd_1_sbox_n121, AesSbox_keyAdd_1_sbox_n120,
         AesSbox_keyAdd_1_sbox_n119, AesSbox_keyAdd_1_sbox_n118,
         AesSbox_keyAdd_1_sbox_n117, AesSbox_keyAdd_1_sbox_n116,
         AesSbox_keyAdd_1_sbox_n115, AesSbox_keyAdd_1_sbox_n114,
         AesSbox_keyAdd_1_sbox_n113, AesSbox_keyAdd_1_sbox_n112,
         AesSbox_keyAdd_1_sbox_n111, AesSbox_keyAdd_1_sbox_n110,
         AesSbox_keyAdd_1_sbox_n109, AesSbox_keyAdd_1_sbox_n108,
         AesSbox_keyAdd_1_sbox_n107, AesSbox_keyAdd_1_sbox_n106,
         AesSbox_keyAdd_1_sbox_n105, AesSbox_keyAdd_1_sbox_n104,
         AesSbox_keyAdd_1_sbox_n103, AesSbox_keyAdd_1_sbox_n102,
         AesSbox_keyAdd_1_sbox_n101, AesSbox_keyAdd_1_sbox_n100,
         AesSbox_keyAdd_1_sbox_n99, AesSbox_keyAdd_1_sbox_n98,
         AesSbox_keyAdd_1_sbox_n97, AesSbox_keyAdd_1_sbox_n96,
         AesSbox_keyAdd_1_sbox_n95, AesSbox_keyAdd_1_sbox_n94,
         AesSbox_keyAdd_1_sbox_n93, AesSbox_keyAdd_1_sbox_n92,
         AesSbox_keyAdd_1_sbox_n91, AesSbox_keyAdd_1_sbox_n90,
         AesSbox_keyAdd_1_sbox_n89, AesSbox_keyAdd_1_sbox_n88,
         AesSbox_keyAdd_1_sbox_n87, AesSbox_keyAdd_1_sbox_n86,
         AesSbox_keyAdd_1_sbox_n85, AesSbox_keyAdd_1_sbox_n84,
         AesSbox_keyAdd_1_sbox_n83, AesSbox_keyAdd_1_sbox_n82,
         AesSbox_keyAdd_1_sbox_n81, AesSbox_keyAdd_1_sbox_n80,
         AesSbox_keyAdd_1_sbox_n79, AesSbox_keyAdd_1_sbox_n78,
         AesSbox_keyAdd_1_sbox_n77, AesSbox_keyAdd_1_sbox_n76,
         AesSbox_keyAdd_1_sbox_n75, AesSbox_keyAdd_1_sbox_n74,
         AesSbox_keyAdd_1_sbox_n73, AesSbox_keyAdd_1_sbox_n72,
         AesSbox_keyAdd_1_sbox_n71, AesSbox_keyAdd_1_sbox_n70,
         AesSbox_keyAdd_1_sbox_n69, AesSbox_keyAdd_1_sbox_n68,
         AesSbox_keyAdd_1_sbox_n67, AesSbox_keyAdd_1_sbox_n66,
         AesSbox_keyAdd_1_sbox_n65, AesSbox_keyAdd_1_sbox_n64,
         AesSbox_keyAdd_1_sbox_n63, AesSbox_keyAdd_1_sbox_n62,
         AesSbox_keyAdd_1_sbox_n61, AesSbox_keyAdd_1_sbox_n60,
         AesSbox_keyAdd_1_sbox_n59, AesSbox_keyAdd_1_sbox_n58,
         AesSbox_keyAdd_1_sbox_n57, AesSbox_keyAdd_1_sbox_n56,
         AesSbox_keyAdd_1_sbox_n55, AesSbox_keyAdd_1_sbox_n54,
         AesSbox_keyAdd_1_sbox_n53, AesSbox_keyAdd_1_sbox_n52,
         AesSbox_keyAdd_1_sbox_n51, AesSbox_keyAdd_1_sbox_n50,
         AesSbox_keyAdd_1_sbox_n49, AesSbox_keyAdd_1_sbox_n48,
         AesSbox_keyAdd_1_sbox_n47, AesSbox_keyAdd_1_sbox_n46,
         AesSbox_keyAdd_1_sbox_n45, AesSbox_keyAdd_1_sbox_n44,
         AesSbox_keyAdd_1_sbox_n43, AesSbox_keyAdd_1_sbox_n42,
         AesSbox_keyAdd_1_sbox_n41, AesSbox_keyAdd_1_sbox_n40,
         AesSbox_keyAdd_1_sbox_n39, AesSbox_keyAdd_1_sbox_n38,
         AesSbox_keyAdd_1_sbox_n37, AesSbox_keyAdd_1_sbox_n36,
         AesSbox_keyAdd_1_sbox_n35, AesSbox_keyAdd_1_sbox_n34,
         AesSbox_keyAdd_1_sbox_n33, AesSbox_keyAdd_1_sbox_n32,
         AesSbox_keyAdd_1_sbox_n31, AesSbox_keyAdd_1_sbox_n30,
         AesSbox_keyAdd_1_sbox_n29, AesSbox_keyAdd_1_sbox_n28,
         AesSbox_keyAdd_1_sbox_n27, AesSbox_keyAdd_1_sbox_n26,
         AesSbox_keyAdd_1_sbox_n25, AesSbox_keyAdd_1_sbox_n24,
         AesSbox_keyAdd_1_sbox_n23, AesSbox_keyAdd_1_sbox_n22,
         AesSbox_keyAdd_1_sbox_n21, AesSbox_keyAdd_1_sbox_n20,
         AesSbox_keyAdd_1_sbox_n19, AesSbox_keyAdd_1_sbox_n18,
         AesSbox_keyAdd_1_sbox_n17, AesSbox_keyAdd_1_sbox_n16,
         AesSbox_keyAdd_1_sbox_n15, AesSbox_keyAdd_1_sbox_n14,
         AesSbox_keyAdd_1_sbox_n13, AesSbox_keyAdd_1_sbox_n12,
         AesSbox_keyAdd_1_sbox_n11, AesSbox_keyAdd_1_sbox_n10,
         AesSbox_keyAdd_1_sbox_n9, AesSbox_keyAdd_1_sbox_n8,
         AesSbox_keyAdd_1_sbox_n7, AesSbox_keyAdd_1_sbox_n6,
         AesSbox_keyAdd_1_sbox_n5, AesSbox_keyAdd_1_sbox_n4,
         AesSbox_keyAdd_1_sbox_n3, AesSbox_keyAdd_1_sbox_n2,
         AesSbox_keyAdd_1_sbox_n1;
  wire   [7:0] output_sbox_0;
  wire   [7:0] output_sbox_1;

  NOR2_X1 det_U0032 ( .A1(io_error), .A2(n23), .ZN(io_out[7]) );
  NOR2_X1 det_U0033 ( .A1(io_error), .A2(n24), .ZN(io_out[6]) );
  NOR2_X1 det_U0034 ( .A1(io_error), .A2(n25), .ZN(io_out[5]) );
  NOR2_X1 det_U0035 ( .A1(io_error), .A2(n26), .ZN(io_out[4]) );
  NOR2_X1 det_U0036 ( .A1(io_error), .A2(n27), .ZN(io_out[3]) );
  NOR2_X1 det_U0037 ( .A1(io_error), .A2(n28), .ZN(io_out[2]) );
  NOR2_X1 det_U0038 ( .A1(io_error), .A2(n29), .ZN(io_out[1]) );
  NOR2_X1 det_U0039 ( .A1(io_error), .A2(n30), .ZN(io_out[0]) );
  NAND2_X1 det_U0040 ( .A1(n31), .A2(n32), .ZN(io_error) );
  NOR2_X1 det_U0041 ( .A1(n33), .A2(n34), .ZN(n32) );
  NAND2_X1 det_U0042 ( .A1(n35), .A2(n36), .ZN(n34) );
  XOR2_X1 det_U0043 ( .A(n28), .B(output_sbox_1[2]), .Z(n36) );
  INV_X1 det_U0044 ( .A(output_sbox_0[2]), .ZN(n28) );
  XOR2_X1 det_U0045 ( .A(n27), .B(output_sbox_1[3]), .Z(n35) );
  INV_X1 det_U0046 ( .A(output_sbox_0[3]), .ZN(n27) );
  NAND2_X1 det_U0047 ( .A1(n37), .A2(n38), .ZN(n33) );
  XOR2_X1 det_U0048 ( .A(n30), .B(output_sbox_1[0]), .Z(n38) );
  INV_X1 det_U0049 ( .A(output_sbox_0[0]), .ZN(n30) );
  XOR2_X1 det_U0050 ( .A(n29), .B(output_sbox_1[1]), .Z(n37) );
  INV_X1 det_U0051 ( .A(output_sbox_0[1]), .ZN(n29) );
  NOR2_X1 det_U0052 ( .A1(n39), .A2(n40), .ZN(n31) );
  NAND2_X1 det_U0053 ( .A1(n41), .A2(n42), .ZN(n40) );
  XOR2_X1 det_U0054 ( .A(n24), .B(output_sbox_1[6]), .Z(n42) );
  INV_X1 det_U0055 ( .A(output_sbox_0[6]), .ZN(n24) );
  XOR2_X1 det_U0056 ( .A(n23), .B(output_sbox_1[7]), .Z(n41) );
  INV_X1 det_U0057 ( .A(output_sbox_0[7]), .ZN(n23) );
  NAND2_X1 det_U0058 ( .A1(n43), .A2(n44), .ZN(n39) );
  XOR2_X1 det_U0059 ( .A(n26), .B(output_sbox_1[4]), .Z(n44) );
  INV_X1 det_U0060 ( .A(output_sbox_0[4]), .ZN(n26) );
  XOR2_X1 det_U0061 ( .A(n25), .B(output_sbox_1[5]), .Z(n43) );
  INV_X1 det_U0062 ( .A(output_sbox_0[5]), .ZN(n25) );
  XOR2_X1 AesSbox_keyAdd_U0008 ( .A(AesSbox_keyAdd_sbox_io_o0), .B(io_key[0]), 
        .Z(output_sbox_0[0]) );
  XOR2_X1 AesSbox_keyAdd_U0007 ( .A(AesSbox_keyAdd_sbox_io_o1), .B(io_key[1]), 
        .Z(output_sbox_0[1]) );
  XOR2_X1 AesSbox_keyAdd_U0006 ( .A(AesSbox_keyAdd_sbox_io_o2), .B(io_key[2]), 
        .Z(output_sbox_0[2]) );
  XOR2_X1 AesSbox_keyAdd_U0005 ( .A(AesSbox_keyAdd_sbox_io_o3), .B(io_key[3]), 
        .Z(output_sbox_0[3]) );
  XOR2_X1 AesSbox_keyAdd_U0004 ( .A(AesSbox_keyAdd_sbox_io_o4), .B(io_key[4]), 
        .Z(output_sbox_0[4]) );
  XOR2_X1 AesSbox_keyAdd_U0003 ( .A(AesSbox_keyAdd_sbox_io_o5), .B(io_key[5]), 
        .Z(output_sbox_0[5]) );
  XOR2_X1 AesSbox_keyAdd_U0002 ( .A(AesSbox_keyAdd_sbox_io_o6), .B(io_key[6]), 
        .Z(output_sbox_0[6]) );
  XOR2_X1 AesSbox_keyAdd_U0001 ( .A(AesSbox_keyAdd_sbox_io_o7), .B(io_key[7]), 
        .Z(output_sbox_0[7]) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0136 ( .A(io_state[0]), .B(io_state[3]), .Z(
        AesSbox_keyAdd_sbox_n71) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0135 ( .A(io_state[2]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_sbox_n107) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0134 ( .A(AesSbox_keyAdd_sbox_n71), .B(
        AesSbox_keyAdd_sbox_n107), .Z(AesSbox_keyAdd_sbox_n75) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0133 ( .A(io_state[1]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_sbox_n126) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0132 ( .A(io_state[6]), .B(io_state[4]), .ZN(
        AesSbox_keyAdd_sbox_n125) );
  INV_X1 AesSbox_keyAdd_sbox_U0131 ( .A(AesSbox_keyAdd_sbox_n125), .ZN(
        AesSbox_keyAdd_sbox_n108) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0130 ( .A(AesSbox_keyAdd_sbox_n108), .B(
        AesSbox_keyAdd_sbox_n126), .Z(AesSbox_keyAdd_sbox_n74) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0129 ( .A1(AesSbox_keyAdd_sbox_n74), .A2(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n117) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0128 ( .A(io_state[3]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_sbox_n124) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0127 ( .A(AesSbox_keyAdd_sbox_n107), .B(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n128) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0126 ( .A1(AesSbox_keyAdd_sbox_n124), .A2(
        AesSbox_keyAdd_sbox_n128), .ZN(AesSbox_keyAdd_sbox_n127) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0125 ( .A(AesSbox_keyAdd_sbox_n117), .B(
        AesSbox_keyAdd_sbox_n127), .ZN(AesSbox_keyAdd_sbox_n100) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0124 ( .A(AesSbox_keyAdd_sbox_n126), .B(
        AesSbox_keyAdd_sbox_n100), .ZN(AesSbox_keyAdd_sbox_n120) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0123 ( .A(AesSbox_keyAdd_sbox_n125), .B(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n61) );
  INV_X1 AesSbox_keyAdd_sbox_U0122 ( .A(AesSbox_keyAdd_sbox_n124), .ZN(
        AesSbox_keyAdd_sbox_n73) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0121 ( .A(io_state[0]), .B(io_state[6]), .Z(
        AesSbox_keyAdd_sbox_n48) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0120 ( .A(AesSbox_keyAdd_sbox_n73), .B(
        AesSbox_keyAdd_sbox_n48), .Z(AesSbox_keyAdd_sbox_n64) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0119 ( .A1(AesSbox_keyAdd_sbox_n64), .A2(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n113) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0118 ( .A(io_state[1]), .B(io_state[2]), .Z(
        AesSbox_keyAdd_sbox_n119) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0117 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_sbox_n119), .Z(AesSbox_keyAdd_sbox_n66) );
  INV_X1 AesSbox_keyAdd_sbox_U0116 ( .A(AesSbox_keyAdd_sbox_n66), .ZN(
        AesSbox_keyAdd_sbox_n115) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0115 ( .A(AesSbox_keyAdd_sbox_n115), .B(
        io_state[6]), .ZN(AesSbox_keyAdd_sbox_n14) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0114 ( .A(io_state[0]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_sbox_n116) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0113 ( .A(AesSbox_keyAdd_sbox_n14), .B(
        AesSbox_keyAdd_sbox_n116), .Z(AesSbox_keyAdd_sbox_n65) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0112 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n58) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0111 ( .A1(AesSbox_keyAdd_sbox_n65), .A2(
        AesSbox_keyAdd_sbox_n58), .ZN(AesSbox_keyAdd_sbox_n123) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0110 ( .A(AesSbox_keyAdd_sbox_n113), .B(
        AesSbox_keyAdd_sbox_n123), .Z(AesSbox_keyAdd_sbox_n122) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0109 ( .A(AesSbox_keyAdd_sbox_n61), .B(
        AesSbox_keyAdd_sbox_n122), .ZN(AesSbox_keyAdd_sbox_n121) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0108 ( .A(AesSbox_keyAdd_sbox_n120), .B(
        AesSbox_keyAdd_sbox_n121), .Z(AesSbox_keyAdd_sbox_n109) );
  INV_X1 AesSbox_keyAdd_sbox_U0107 ( .A(AesSbox_keyAdd_sbox_n109), .ZN(
        AesSbox_keyAdd_sbox_n94) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0106 ( .A(AesSbox_keyAdd_sbox_n119), .B(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n45) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0105 ( .A1(AesSbox_keyAdd_sbox_n45), .A2(
        AesSbox_keyAdd_sbox_n116), .ZN(AesSbox_keyAdd_sbox_n118) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0104 ( .A(AesSbox_keyAdd_sbox_n117), .B(
        AesSbox_keyAdd_sbox_n118), .Z(AesSbox_keyAdd_sbox_n104) );
  INV_X1 AesSbox_keyAdd_sbox_U0103 ( .A(AesSbox_keyAdd_sbox_n116), .ZN(
        AesSbox_keyAdd_sbox_n43) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0102 ( .A(AesSbox_keyAdd_sbox_n104), .B(
        AesSbox_keyAdd_sbox_n43), .Z(AesSbox_keyAdd_sbox_n110) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0101 ( .A(AesSbox_keyAdd_sbox_n115), .B(
        io_state[3]), .ZN(AesSbox_keyAdd_sbox_n25) );
  AND2_X1 AesSbox_keyAdd_sbox_U0100 ( .A1(AesSbox_keyAdd_sbox_n25), .A2(
        io_state[7]), .ZN(AesSbox_keyAdd_sbox_n114) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0099 ( .A(AesSbox_keyAdd_sbox_n113), .B(
        AesSbox_keyAdd_sbox_n114), .ZN(AesSbox_keyAdd_sbox_n112) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0098 ( .A(AesSbox_keyAdd_sbox_n45), .B(
        AesSbox_keyAdd_sbox_n112), .ZN(AesSbox_keyAdd_sbox_n111) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0097 ( .A(AesSbox_keyAdd_sbox_n110), .B(
        AesSbox_keyAdd_sbox_n111), .Z(AesSbox_keyAdd_sbox_n81) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0096 ( .A(AesSbox_keyAdd_sbox_n109), .B(
        AesSbox_keyAdd_sbox_n81), .Z(AesSbox_keyAdd_sbox_n84) );
  AND2_X1 AesSbox_keyAdd_sbox_U0095 ( .A1(AesSbox_keyAdd_sbox_n94), .A2(
        AesSbox_keyAdd_sbox_n84), .ZN(AesSbox_keyAdd_sbox_n101) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0094 ( .A(AesSbox_keyAdd_sbox_n25), .B(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n50) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0093 ( .A(AesSbox_keyAdd_sbox_n107), .B(
        AesSbox_keyAdd_sbox_n108), .Z(AesSbox_keyAdd_sbox_n68) );
  AND2_X1 AesSbox_keyAdd_sbox_U0092 ( .A1(AesSbox_keyAdd_sbox_n68), .A2(
        AesSbox_keyAdd_sbox_n48), .ZN(AesSbox_keyAdd_sbox_n98) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0091 ( .A(AesSbox_keyAdd_sbox_n66), .B(
        AesSbox_keyAdd_sbox_n68), .ZN(AesSbox_keyAdd_sbox_n33) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0090 ( .A1(AesSbox_keyAdd_sbox_n50), .A2(
        AesSbox_keyAdd_sbox_n33), .ZN(AesSbox_keyAdd_sbox_n106) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0089 ( .A(AesSbox_keyAdd_sbox_n98), .B(
        AesSbox_keyAdd_sbox_n106), .Z(AesSbox_keyAdd_sbox_n105) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0088 ( .A(AesSbox_keyAdd_sbox_n50), .B(
        AesSbox_keyAdd_sbox_n105), .Z(AesSbox_keyAdd_sbox_n102) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0087 ( .A(AesSbox_keyAdd_sbox_n33), .B(
        AesSbox_keyAdd_sbox_n104), .Z(AesSbox_keyAdd_sbox_n103) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0086 ( .A(AesSbox_keyAdd_sbox_n102), .B(
        AesSbox_keyAdd_sbox_n103), .Z(AesSbox_keyAdd_sbox_n85) );
  INV_X1 AesSbox_keyAdd_sbox_U0085 ( .A(AesSbox_keyAdd_sbox_n85), .ZN(
        AesSbox_keyAdd_sbox_n77) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0084 ( .A1(AesSbox_keyAdd_sbox_n101), .A2(
        AesSbox_keyAdd_sbox_n77), .ZN(AesSbox_keyAdd_sbox_n93) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0083 ( .A(AesSbox_keyAdd_sbox_n48), .B(
        AesSbox_keyAdd_sbox_n100), .ZN(AesSbox_keyAdd_sbox_n95) );
  AND2_X1 AesSbox_keyAdd_sbox_U0082 ( .A1(AesSbox_keyAdd_sbox_n66), .A2(
        AesSbox_keyAdd_sbox_n14), .ZN(AesSbox_keyAdd_sbox_n99) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0081 ( .A(AesSbox_keyAdd_sbox_n98), .B(
        AesSbox_keyAdd_sbox_n99), .Z(AesSbox_keyAdd_sbox_n97) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0080 ( .A(AesSbox_keyAdd_sbox_n68), .B(
        AesSbox_keyAdd_sbox_n97), .Z(AesSbox_keyAdd_sbox_n96) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0079 ( .A(AesSbox_keyAdd_sbox_n95), .B(
        AesSbox_keyAdd_sbox_n96), .Z(AesSbox_keyAdd_sbox_n91) );
  INV_X1 AesSbox_keyAdd_sbox_U0078 ( .A(AesSbox_keyAdd_sbox_n91), .ZN(
        AesSbox_keyAdd_sbox_n90) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0077 ( .A1(AesSbox_keyAdd_sbox_n90), .A2(
        AesSbox_keyAdd_sbox_n94), .ZN(AesSbox_keyAdd_sbox_n80) );
  INV_X1 AesSbox_keyAdd_sbox_U0076 ( .A(AesSbox_keyAdd_sbox_n80), .ZN(
        AesSbox_keyAdd_sbox_n88) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0075 ( .A(AesSbox_keyAdd_sbox_n93), .B(
        AesSbox_keyAdd_sbox_n88), .Z(AesSbox_keyAdd_sbox_n92) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0074 ( .A(AesSbox_keyAdd_sbox_n92), .B(
        AesSbox_keyAdd_sbox_n84), .ZN(AesSbox_keyAdd_sbox_n13) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0073 ( .A1(AesSbox_keyAdd_sbox_n81), .A2(
        AesSbox_keyAdd_sbox_n91), .ZN(AesSbox_keyAdd_sbox_n89) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0072 ( .A(AesSbox_keyAdd_sbox_n77), .B(
        AesSbox_keyAdd_sbox_n90), .Z(AesSbox_keyAdd_sbox_n79) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0071 ( .A1(AesSbox_keyAdd_sbox_n89), .A2(
        AesSbox_keyAdd_sbox_n79), .ZN(AesSbox_keyAdd_sbox_n87) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0070 ( .A(AesSbox_keyAdd_sbox_n87), .B(
        AesSbox_keyAdd_sbox_n88), .Z(AesSbox_keyAdd_sbox_n86) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0069 ( .A(AesSbox_keyAdd_sbox_n86), .B(
        AesSbox_keyAdd_sbox_n79), .Z(AesSbox_keyAdd_sbox_n59) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0068 ( .A(AesSbox_keyAdd_sbox_n13), .B(
        AesSbox_keyAdd_sbox_n59), .Z(AesSbox_keyAdd_sbox_n46) );
  INV_X1 AesSbox_keyAdd_sbox_U0067 ( .A(AesSbox_keyAdd_sbox_n46), .ZN(
        AesSbox_keyAdd_sbox_n42) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0066 ( .A(AesSbox_keyAdd_sbox_n80), .B(
        AesSbox_keyAdd_sbox_n85), .Z(AesSbox_keyAdd_sbox_n83) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0065 ( .A1(AesSbox_keyAdd_sbox_n83), .A2(
        AesSbox_keyAdd_sbox_n84), .ZN(AesSbox_keyAdd_sbox_n82) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0064 ( .A(AesSbox_keyAdd_sbox_n82), .B(
        AesSbox_keyAdd_sbox_n81), .ZN(AesSbox_keyAdd_sbox_n32) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0063 ( .A(AesSbox_keyAdd_sbox_n80), .B(
        AesSbox_keyAdd_sbox_n81), .Z(AesSbox_keyAdd_sbox_n78) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0062 ( .A1(AesSbox_keyAdd_sbox_n78), .A2(
        AesSbox_keyAdd_sbox_n79), .ZN(AesSbox_keyAdd_sbox_n76) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0061 ( .A(AesSbox_keyAdd_sbox_n76), .B(
        AesSbox_keyAdd_sbox_n77), .ZN(AesSbox_keyAdd_sbox_n24) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0060 ( .A(AesSbox_keyAdd_sbox_n32), .B(
        AesSbox_keyAdd_sbox_n24), .ZN(AesSbox_keyAdd_sbox_n70) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0059 ( .A(AesSbox_keyAdd_sbox_n42), .B(
        AesSbox_keyAdd_sbox_n70), .Z(AesSbox_keyAdd_sbox_n72) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0058 ( .A1(AesSbox_keyAdd_sbox_n75), .A2(
        AesSbox_keyAdd_sbox_n72), .ZN(AesSbox_keyAdd_sbox_n22) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0057 ( .A1(AesSbox_keyAdd_sbox_n74), .A2(
        AesSbox_keyAdd_sbox_n70), .ZN(AesSbox_keyAdd_sbox_n40) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0056 ( .A(AesSbox_keyAdd_sbox_n22), .B(
        AesSbox_keyAdd_sbox_n40), .ZN(AesSbox_keyAdd_sbox_n55) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0055 ( .A1(AesSbox_keyAdd_sbox_n72), .A2(
        AesSbox_keyAdd_sbox_n73), .ZN(AesSbox_keyAdd_sbox_n69) );
  AND2_X1 AesSbox_keyAdd_sbox_U0054 ( .A1(AesSbox_keyAdd_sbox_n70), .A2(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n41) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0053 ( .A(AesSbox_keyAdd_sbox_n69), .B(
        AesSbox_keyAdd_sbox_n41), .Z(AesSbox_keyAdd_sbox_n15) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0052 ( .A(AesSbox_keyAdd_sbox_n13), .B(
        AesSbox_keyAdd_sbox_n32), .ZN(AesSbox_keyAdd_sbox_n47) );
  AND2_X1 AesSbox_keyAdd_sbox_U0051 ( .A1(AesSbox_keyAdd_sbox_n68), .A2(
        AesSbox_keyAdd_sbox_n47), .ZN(AesSbox_keyAdd_sbox_n67) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0050 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n67), .Z(AesSbox_keyAdd_sbox_n4) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0049 ( .A1(AesSbox_keyAdd_sbox_n13), .A2(
        AesSbox_keyAdd_sbox_n66), .ZN(AesSbox_keyAdd_sbox_n16) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0048 ( .A1(AesSbox_keyAdd_sbox_n59), .A2(
        AesSbox_keyAdd_sbox_n65), .ZN(AesSbox_keyAdd_sbox_n62) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0047 ( .A(AesSbox_keyAdd_sbox_n16), .B(
        AesSbox_keyAdd_sbox_n62), .Z(AesSbox_keyAdd_sbox_n28) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0046 ( .A(AesSbox_keyAdd_sbox_n4), .B(
        AesSbox_keyAdd_sbox_n28), .ZN(AesSbox_keyAdd_sbox_n35) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0045 ( .A(AesSbox_keyAdd_sbox_n24), .B(
        AesSbox_keyAdd_sbox_n59), .ZN(AesSbox_keyAdd_sbox_n60) );
  AND2_X1 AesSbox_keyAdd_sbox_U0044 ( .A1(AesSbox_keyAdd_sbox_n60), .A2(
        AesSbox_keyAdd_sbox_n64), .ZN(AesSbox_keyAdd_sbox_n56) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0043 ( .A(AesSbox_keyAdd_sbox_n35), .B(
        AesSbox_keyAdd_sbox_n56), .Z(AesSbox_keyAdd_sbox_n63) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0042 ( .A(AesSbox_keyAdd_sbox_n55), .B(
        AesSbox_keyAdd_sbox_n63), .Z(AesSbox_keyAdd_sbox_io_o0) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0041 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n62), .Z(AesSbox_keyAdd_sbox_n52) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0040 ( .A1(AesSbox_keyAdd_sbox_n60), .A2(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n51) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0039 ( .A1(AesSbox_keyAdd_sbox_n58), .A2(
        AesSbox_keyAdd_sbox_n59), .ZN(AesSbox_keyAdd_sbox_n57) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0038 ( .A(AesSbox_keyAdd_sbox_n56), .B(
        AesSbox_keyAdd_sbox_n57), .Z(AesSbox_keyAdd_sbox_n29) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0037 ( .A(AesSbox_keyAdd_sbox_n51), .B(
        AesSbox_keyAdd_sbox_n29), .ZN(AesSbox_keyAdd_sbox_n34) );
  INV_X1 AesSbox_keyAdd_sbox_U0036 ( .A(AesSbox_keyAdd_sbox_n55), .ZN(
        AesSbox_keyAdd_sbox_n54) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0035 ( .A(AesSbox_keyAdd_sbox_n34), .B(
        AesSbox_keyAdd_sbox_n54), .Z(AesSbox_keyAdd_sbox_n53) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0034 ( .A(AesSbox_keyAdd_sbox_n52), .B(
        AesSbox_keyAdd_sbox_n53), .Z(AesSbox_keyAdd_sbox_io_o1) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0033 ( .A1(io_state[7]), .A2(
        AesSbox_keyAdd_sbox_n24), .ZN(AesSbox_keyAdd_sbox_n31) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0032 ( .A(AesSbox_keyAdd_sbox_n51), .B(
        AesSbox_keyAdd_sbox_n31), .ZN(AesSbox_keyAdd_sbox_n5) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0031 ( .A1(AesSbox_keyAdd_sbox_n50), .A2(
        AesSbox_keyAdd_sbox_n32), .ZN(AesSbox_keyAdd_sbox_n49) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0030 ( .A(AesSbox_keyAdd_sbox_n5), .B(
        AesSbox_keyAdd_sbox_n49), .ZN(AesSbox_keyAdd_sbox_n20) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0029 ( .A1(AesSbox_keyAdd_sbox_n47), .A2(
        AesSbox_keyAdd_sbox_n48), .ZN(AesSbox_keyAdd_sbox_n3) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0028 ( .A1(AesSbox_keyAdd_sbox_n45), .A2(
        AesSbox_keyAdd_sbox_n46), .ZN(AesSbox_keyAdd_sbox_n44) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0027 ( .A(AesSbox_keyAdd_sbox_n3), .B(
        AesSbox_keyAdd_sbox_n44), .ZN(AesSbox_keyAdd_sbox_n23) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0026 ( .A(AesSbox_keyAdd_sbox_n20), .B(
        AesSbox_keyAdd_sbox_n23), .ZN(AesSbox_keyAdd_sbox_n36) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0025 ( .A1(AesSbox_keyAdd_sbox_n42), .A2(
        AesSbox_keyAdd_sbox_n43), .ZN(AesSbox_keyAdd_sbox_n38) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0024 ( .A(AesSbox_keyAdd_sbox_n40), .B(
        AesSbox_keyAdd_sbox_n41), .Z(AesSbox_keyAdd_sbox_n39) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0023 ( .A(AesSbox_keyAdd_sbox_n38), .B(
        AesSbox_keyAdd_sbox_n39), .Z(AesSbox_keyAdd_sbox_n37) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0022 ( .A(AesSbox_keyAdd_sbox_n36), .B(
        AesSbox_keyAdd_sbox_n37), .Z(AesSbox_keyAdd_sbox_io_o2) );
  INV_X1 AesSbox_keyAdd_sbox_U0021 ( .A(AesSbox_keyAdd_sbox_n35), .ZN(
        AesSbox_keyAdd_sbox_n19) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0020 ( .A(AesSbox_keyAdd_sbox_n19), .B(
        AesSbox_keyAdd_sbox_n34), .Z(AesSbox_keyAdd_sbox_io_o3) );
  NOR2_X1 AesSbox_keyAdd_sbox_U0019 ( .A1(AesSbox_keyAdd_sbox_n32), .A2(
        AesSbox_keyAdd_sbox_n33), .ZN(AesSbox_keyAdd_sbox_n12) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0018 ( .A(AesSbox_keyAdd_sbox_n31), .B(
        AesSbox_keyAdd_sbox_n12), .Z(AesSbox_keyAdd_sbox_n30) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0017 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n30), .Z(AesSbox_keyAdd_sbox_n26) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0016 ( .A(AesSbox_keyAdd_sbox_n28), .B(
        AesSbox_keyAdd_sbox_n29), .ZN(AesSbox_keyAdd_sbox_n27) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0015 ( .A(AesSbox_keyAdd_sbox_n26), .B(
        AesSbox_keyAdd_sbox_n27), .Z(AesSbox_keyAdd_sbox_io_o4) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0014 ( .A1(AesSbox_keyAdd_sbox_n24), .A2(
        AesSbox_keyAdd_sbox_n25), .ZN(AesSbox_keyAdd_sbox_n21) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0013 ( .A(AesSbox_keyAdd_sbox_n22), .B(
        AesSbox_keyAdd_sbox_n23), .Z(AesSbox_keyAdd_sbox_n10) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0012 ( .A(AesSbox_keyAdd_sbox_n21), .B(
        AesSbox_keyAdd_sbox_n10), .Z(AesSbox_keyAdd_sbox_n17) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0011 ( .A(AesSbox_keyAdd_sbox_n19), .B(
        AesSbox_keyAdd_sbox_n20), .Z(AesSbox_keyAdd_sbox_n18) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0010 ( .A(AesSbox_keyAdd_sbox_n17), .B(
        AesSbox_keyAdd_sbox_n18), .Z(AesSbox_keyAdd_sbox_io_o5) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U0009 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n16), .ZN(AesSbox_keyAdd_sbox_n8) );
  NAND2_X1 AesSbox_keyAdd_sbox_U0008 ( .A1(AesSbox_keyAdd_sbox_n13), .A2(
        AesSbox_keyAdd_sbox_n14), .ZN(AesSbox_keyAdd_sbox_n11) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0007 ( .A(AesSbox_keyAdd_sbox_n11), .B(
        AesSbox_keyAdd_sbox_n12), .Z(AesSbox_keyAdd_sbox_n7) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0006 ( .A(AesSbox_keyAdd_sbox_n7), .B(
        AesSbox_keyAdd_sbox_n10), .Z(AesSbox_keyAdd_sbox_n9) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0005 ( .A(AesSbox_keyAdd_sbox_n8), .B(
        AesSbox_keyAdd_sbox_n9), .Z(AesSbox_keyAdd_sbox_io_o6) );
  INV_X1 AesSbox_keyAdd_sbox_U0004 ( .A(AesSbox_keyAdd_sbox_n7), .ZN(
        AesSbox_keyAdd_sbox_n6) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0003 ( .A(AesSbox_keyAdd_sbox_n5), .B(
        AesSbox_keyAdd_sbox_n6), .Z(AesSbox_keyAdd_sbox_n1) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0002 ( .A(AesSbox_keyAdd_sbox_n3), .B(
        AesSbox_keyAdd_sbox_n4), .Z(AesSbox_keyAdd_sbox_n2) );
  XOR2_X1 AesSbox_keyAdd_sbox_U0001 ( .A(AesSbox_keyAdd_sbox_n1), .B(
        AesSbox_keyAdd_sbox_n2), .Z(AesSbox_keyAdd_sbox_io_o7) );
  XOR2_X1 AesSbox_keyAdd_1_U0008 ( .A(AesSbox_keyAdd_1_sbox_io_o0), .B(io_key[0]), 
        .Z(output_sbox_1[0]) );
  XOR2_X1 AesSbox_keyAdd_1_U0007 ( .A(AesSbox_keyAdd_1_sbox_io_o1), .B(io_key[1]), 
        .Z(output_sbox_1[1]) );
  XOR2_X1 AesSbox_keyAdd_1_U0006 ( .A(AesSbox_keyAdd_1_sbox_io_o2), .B(io_key[2]), 
        .Z(output_sbox_1[2]) );
  XOR2_X1 AesSbox_keyAdd_1_U0005 ( .A(AesSbox_keyAdd_1_sbox_io_o3), .B(io_key[3]), 
        .Z(output_sbox_1[3]) );
  XOR2_X1 AesSbox_keyAdd_1_U0004 ( .A(AesSbox_keyAdd_1_sbox_io_o4), .B(io_key[4]), 
        .Z(output_sbox_1[4]) );
  XOR2_X1 AesSbox_keyAdd_1_U0003 ( .A(AesSbox_keyAdd_1_sbox_io_o5), .B(io_key[5]), 
        .Z(output_sbox_1[5]) );
  XOR2_X1 AesSbox_keyAdd_1_U0002 ( .A(AesSbox_keyAdd_1_sbox_io_o6), .B(io_key[6]), 
        .Z(output_sbox_1[6]) );
  XOR2_X1 AesSbox_keyAdd_1_U0001 ( .A(AesSbox_keyAdd_1_sbox_io_o7), .B(io_key[7]), 
        .Z(output_sbox_1[7]) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0136 ( .A(io_state[0]), .B(io_state[3]), .Z(
        AesSbox_keyAdd_1_sbox_n71) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0135 ( .A(io_state[2]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_1_sbox_n107) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0134 ( .A(AesSbox_keyAdd_1_sbox_n71), .B(
        AesSbox_keyAdd_1_sbox_n107), .Z(AesSbox_keyAdd_1_sbox_n75) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0133 ( .A(io_state[1]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_1_sbox_n126) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0132 ( .A(io_state[6]), .B(io_state[4]), .ZN(
        AesSbox_keyAdd_1_sbox_n125) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0131 ( .A(AesSbox_keyAdd_1_sbox_n125), .ZN(
        AesSbox_keyAdd_1_sbox_n108) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0130 ( .A(AesSbox_keyAdd_1_sbox_n108), .B(
        AesSbox_keyAdd_1_sbox_n126), .Z(AesSbox_keyAdd_1_sbox_n74) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0129 ( .A1(AesSbox_keyAdd_1_sbox_n74), .A2(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n117) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0128 ( .A(io_state[3]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_1_sbox_n124) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0127 ( .A(AesSbox_keyAdd_1_sbox_n107), .B(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n128) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0126 ( .A1(AesSbox_keyAdd_1_sbox_n124), .A2(
        AesSbox_keyAdd_1_sbox_n128), .ZN(AesSbox_keyAdd_1_sbox_n127) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0125 ( .A(AesSbox_keyAdd_1_sbox_n117), .B(
        AesSbox_keyAdd_1_sbox_n127), .ZN(AesSbox_keyAdd_1_sbox_n100) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0124 ( .A(AesSbox_keyAdd_1_sbox_n126), .B(
        AesSbox_keyAdd_1_sbox_n100), .ZN(AesSbox_keyAdd_1_sbox_n120) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0123 ( .A(AesSbox_keyAdd_1_sbox_n125), .B(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n61) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0122 ( .A(AesSbox_keyAdd_1_sbox_n124), .ZN(
        AesSbox_keyAdd_1_sbox_n73) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0121 ( .A(io_state[0]), .B(io_state[6]), .Z(
        AesSbox_keyAdd_1_sbox_n48) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0120 ( .A(AesSbox_keyAdd_1_sbox_n73), .B(
        AesSbox_keyAdd_1_sbox_n48), .Z(AesSbox_keyAdd_1_sbox_n64) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0119 ( .A1(AesSbox_keyAdd_1_sbox_n64), .A2(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n113) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0118 ( .A(io_state[1]), .B(io_state[2]), .Z(
        AesSbox_keyAdd_1_sbox_n119) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0117 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_1_sbox_n119), .Z(AesSbox_keyAdd_1_sbox_n66) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0116 ( .A(AesSbox_keyAdd_1_sbox_n66), .ZN(
        AesSbox_keyAdd_1_sbox_n115) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0115 ( .A(AesSbox_keyAdd_1_sbox_n115), .B(
        io_state[6]), .ZN(AesSbox_keyAdd_1_sbox_n14) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0114 ( .A(io_state[0]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_1_sbox_n116) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0113 ( .A(AesSbox_keyAdd_1_sbox_n14), .B(
        AesSbox_keyAdd_1_sbox_n116), .Z(AesSbox_keyAdd_1_sbox_n65) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0112 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n58) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0111 ( .A1(AesSbox_keyAdd_1_sbox_n65), .A2(
        AesSbox_keyAdd_1_sbox_n58), .ZN(AesSbox_keyAdd_1_sbox_n123) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0110 ( .A(AesSbox_keyAdd_1_sbox_n113), .B(
        AesSbox_keyAdd_1_sbox_n123), .Z(AesSbox_keyAdd_1_sbox_n122) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0109 ( .A(AesSbox_keyAdd_1_sbox_n61), .B(
        AesSbox_keyAdd_1_sbox_n122), .ZN(AesSbox_keyAdd_1_sbox_n121) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0108 ( .A(AesSbox_keyAdd_1_sbox_n120), .B(
        AesSbox_keyAdd_1_sbox_n121), .Z(AesSbox_keyAdd_1_sbox_n109) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0107 ( .A(AesSbox_keyAdd_1_sbox_n109), .ZN(
        AesSbox_keyAdd_1_sbox_n94) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0106 ( .A(AesSbox_keyAdd_1_sbox_n119), .B(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n45) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0105 ( .A1(AesSbox_keyAdd_1_sbox_n45), .A2(
        AesSbox_keyAdd_1_sbox_n116), .ZN(AesSbox_keyAdd_1_sbox_n118) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0104 ( .A(AesSbox_keyAdd_1_sbox_n117), .B(
        AesSbox_keyAdd_1_sbox_n118), .Z(AesSbox_keyAdd_1_sbox_n104) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0103 ( .A(AesSbox_keyAdd_1_sbox_n116), .ZN(
        AesSbox_keyAdd_1_sbox_n43) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0102 ( .A(AesSbox_keyAdd_1_sbox_n104), .B(
        AesSbox_keyAdd_1_sbox_n43), .Z(AesSbox_keyAdd_1_sbox_n110) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0101 ( .A(AesSbox_keyAdd_1_sbox_n115), .B(
        io_state[3]), .ZN(AesSbox_keyAdd_1_sbox_n25) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0100 ( .A1(AesSbox_keyAdd_1_sbox_n25), .A2(
        io_state[7]), .ZN(AesSbox_keyAdd_1_sbox_n114) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0099 ( .A(AesSbox_keyAdd_1_sbox_n113), .B(
        AesSbox_keyAdd_1_sbox_n114), .ZN(AesSbox_keyAdd_1_sbox_n112) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0098 ( .A(AesSbox_keyAdd_1_sbox_n45), .B(
        AesSbox_keyAdd_1_sbox_n112), .ZN(AesSbox_keyAdd_1_sbox_n111) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0097 ( .A(AesSbox_keyAdd_1_sbox_n110), .B(
        AesSbox_keyAdd_1_sbox_n111), .Z(AesSbox_keyAdd_1_sbox_n81) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0096 ( .A(AesSbox_keyAdd_1_sbox_n109), .B(
        AesSbox_keyAdd_1_sbox_n81), .Z(AesSbox_keyAdd_1_sbox_n84) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0095 ( .A1(AesSbox_keyAdd_1_sbox_n94), .A2(
        AesSbox_keyAdd_1_sbox_n84), .ZN(AesSbox_keyAdd_1_sbox_n101) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0094 ( .A(AesSbox_keyAdd_1_sbox_n25), .B(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n50) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0093 ( .A(AesSbox_keyAdd_1_sbox_n107), .B(
        AesSbox_keyAdd_1_sbox_n108), .Z(AesSbox_keyAdd_1_sbox_n68) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0092 ( .A1(AesSbox_keyAdd_1_sbox_n68), .A2(
        AesSbox_keyAdd_1_sbox_n48), .ZN(AesSbox_keyAdd_1_sbox_n98) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0091 ( .A(AesSbox_keyAdd_1_sbox_n66), .B(
        AesSbox_keyAdd_1_sbox_n68), .ZN(AesSbox_keyAdd_1_sbox_n33) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0090 ( .A1(AesSbox_keyAdd_1_sbox_n50), .A2(
        AesSbox_keyAdd_1_sbox_n33), .ZN(AesSbox_keyAdd_1_sbox_n106) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0089 ( .A(AesSbox_keyAdd_1_sbox_n98), .B(
        AesSbox_keyAdd_1_sbox_n106), .Z(AesSbox_keyAdd_1_sbox_n105) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0088 ( .A(AesSbox_keyAdd_1_sbox_n50), .B(
        AesSbox_keyAdd_1_sbox_n105), .Z(AesSbox_keyAdd_1_sbox_n102) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0087 ( .A(AesSbox_keyAdd_1_sbox_n33), .B(
        AesSbox_keyAdd_1_sbox_n104), .Z(AesSbox_keyAdd_1_sbox_n103) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0086 ( .A(AesSbox_keyAdd_1_sbox_n102), .B(
        AesSbox_keyAdd_1_sbox_n103), .Z(AesSbox_keyAdd_1_sbox_n85) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0085 ( .A(AesSbox_keyAdd_1_sbox_n85), .ZN(
        AesSbox_keyAdd_1_sbox_n77) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0084 ( .A1(AesSbox_keyAdd_1_sbox_n101), .A2(
        AesSbox_keyAdd_1_sbox_n77), .ZN(AesSbox_keyAdd_1_sbox_n93) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0083 ( .A(AesSbox_keyAdd_1_sbox_n48), .B(
        AesSbox_keyAdd_1_sbox_n100), .ZN(AesSbox_keyAdd_1_sbox_n95) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0082 ( .A1(AesSbox_keyAdd_1_sbox_n66), .A2(
        AesSbox_keyAdd_1_sbox_n14), .ZN(AesSbox_keyAdd_1_sbox_n99) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0081 ( .A(AesSbox_keyAdd_1_sbox_n98), .B(
        AesSbox_keyAdd_1_sbox_n99), .Z(AesSbox_keyAdd_1_sbox_n97) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0080 ( .A(AesSbox_keyAdd_1_sbox_n68), .B(
        AesSbox_keyAdd_1_sbox_n97), .Z(AesSbox_keyAdd_1_sbox_n96) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0079 ( .A(AesSbox_keyAdd_1_sbox_n95), .B(
        AesSbox_keyAdd_1_sbox_n96), .Z(AesSbox_keyAdd_1_sbox_n91) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0078 ( .A(AesSbox_keyAdd_1_sbox_n91), .ZN(
        AesSbox_keyAdd_1_sbox_n90) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0077 ( .A1(AesSbox_keyAdd_1_sbox_n90), .A2(
        AesSbox_keyAdd_1_sbox_n94), .ZN(AesSbox_keyAdd_1_sbox_n80) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0076 ( .A(AesSbox_keyAdd_1_sbox_n80), .ZN(
        AesSbox_keyAdd_1_sbox_n88) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0075 ( .A(AesSbox_keyAdd_1_sbox_n93), .B(
        AesSbox_keyAdd_1_sbox_n88), .Z(AesSbox_keyAdd_1_sbox_n92) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0074 ( .A(AesSbox_keyAdd_1_sbox_n92), .B(
        AesSbox_keyAdd_1_sbox_n84), .ZN(AesSbox_keyAdd_1_sbox_n13) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0073 ( .A1(AesSbox_keyAdd_1_sbox_n81), .A2(
        AesSbox_keyAdd_1_sbox_n91), .ZN(AesSbox_keyAdd_1_sbox_n89) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0072 ( .A(AesSbox_keyAdd_1_sbox_n77), .B(
        AesSbox_keyAdd_1_sbox_n90), .Z(AesSbox_keyAdd_1_sbox_n79) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0071 ( .A1(AesSbox_keyAdd_1_sbox_n89), .A2(
        AesSbox_keyAdd_1_sbox_n79), .ZN(AesSbox_keyAdd_1_sbox_n87) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0070 ( .A(AesSbox_keyAdd_1_sbox_n87), .B(
        AesSbox_keyAdd_1_sbox_n88), .Z(AesSbox_keyAdd_1_sbox_n86) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0069 ( .A(AesSbox_keyAdd_1_sbox_n86), .B(
        AesSbox_keyAdd_1_sbox_n79), .Z(AesSbox_keyAdd_1_sbox_n59) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0068 ( .A(AesSbox_keyAdd_1_sbox_n13), .B(
        AesSbox_keyAdd_1_sbox_n59), .Z(AesSbox_keyAdd_1_sbox_n46) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0067 ( .A(AesSbox_keyAdd_1_sbox_n46), .ZN(
        AesSbox_keyAdd_1_sbox_n42) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0066 ( .A(AesSbox_keyAdd_1_sbox_n80), .B(
        AesSbox_keyAdd_1_sbox_n85), .Z(AesSbox_keyAdd_1_sbox_n83) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0065 ( .A1(AesSbox_keyAdd_1_sbox_n83), .A2(
        AesSbox_keyAdd_1_sbox_n84), .ZN(AesSbox_keyAdd_1_sbox_n82) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0064 ( .A(AesSbox_keyAdd_1_sbox_n82), .B(
        AesSbox_keyAdd_1_sbox_n81), .ZN(AesSbox_keyAdd_1_sbox_n32) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0063 ( .A(AesSbox_keyAdd_1_sbox_n80), .B(
        AesSbox_keyAdd_1_sbox_n81), .Z(AesSbox_keyAdd_1_sbox_n78) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0062 ( .A1(AesSbox_keyAdd_1_sbox_n78), .A2(
        AesSbox_keyAdd_1_sbox_n79), .ZN(AesSbox_keyAdd_1_sbox_n76) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0061 ( .A(AesSbox_keyAdd_1_sbox_n76), .B(
        AesSbox_keyAdd_1_sbox_n77), .ZN(AesSbox_keyAdd_1_sbox_n24) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U060 ( .A(AesSbox_keyAdd_1_sbox_n32), .B(
        AesSbox_keyAdd_1_sbox_n24), .ZN(AesSbox_keyAdd_1_sbox_n70) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0059 ( .A(AesSbox_keyAdd_1_sbox_n42), .B(
        AesSbox_keyAdd_1_sbox_n70), .Z(AesSbox_keyAdd_1_sbox_n72) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0058 ( .A1(AesSbox_keyAdd_1_sbox_n75), .A2(
        AesSbox_keyAdd_1_sbox_n72), .ZN(AesSbox_keyAdd_1_sbox_n22) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0057 ( .A1(AesSbox_keyAdd_1_sbox_n74), .A2(
        AesSbox_keyAdd_1_sbox_n70), .ZN(AesSbox_keyAdd_1_sbox_n40) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0056 ( .A(AesSbox_keyAdd_1_sbox_n22), .B(
        AesSbox_keyAdd_1_sbox_n40), .ZN(AesSbox_keyAdd_1_sbox_n55) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0055 ( .A1(AesSbox_keyAdd_1_sbox_n72), .A2(
        AesSbox_keyAdd_1_sbox_n73), .ZN(AesSbox_keyAdd_1_sbox_n69) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0054 ( .A1(AesSbox_keyAdd_1_sbox_n70), .A2(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n41) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0053 ( .A(AesSbox_keyAdd_1_sbox_n69), .B(
        AesSbox_keyAdd_1_sbox_n41), .Z(AesSbox_keyAdd_1_sbox_n15) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0052 ( .A(AesSbox_keyAdd_1_sbox_n13), .B(
        AesSbox_keyAdd_1_sbox_n32), .ZN(AesSbox_keyAdd_1_sbox_n47) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0051 ( .A1(AesSbox_keyAdd_1_sbox_n68), .A2(
        AesSbox_keyAdd_1_sbox_n47), .ZN(AesSbox_keyAdd_1_sbox_n67) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0050 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n67), .Z(AesSbox_keyAdd_1_sbox_n4) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0049 ( .A1(AesSbox_keyAdd_1_sbox_n13), .A2(
        AesSbox_keyAdd_1_sbox_n66), .ZN(AesSbox_keyAdd_1_sbox_n16) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0048 ( .A1(AesSbox_keyAdd_1_sbox_n59), .A2(
        AesSbox_keyAdd_1_sbox_n65), .ZN(AesSbox_keyAdd_1_sbox_n62) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0047 ( .A(AesSbox_keyAdd_1_sbox_n16), .B(
        AesSbox_keyAdd_1_sbox_n62), .Z(AesSbox_keyAdd_1_sbox_n28) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0046 ( .A(AesSbox_keyAdd_1_sbox_n4), .B(
        AesSbox_keyAdd_1_sbox_n28), .ZN(AesSbox_keyAdd_1_sbox_n35) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0045 ( .A(AesSbox_keyAdd_1_sbox_n24), .B(
        AesSbox_keyAdd_1_sbox_n59), .ZN(AesSbox_keyAdd_1_sbox_n60) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U0044 ( .A1(AesSbox_keyAdd_1_sbox_n60), .A2(
        AesSbox_keyAdd_1_sbox_n64), .ZN(AesSbox_keyAdd_1_sbox_n56) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0043 ( .A(AesSbox_keyAdd_1_sbox_n35), .B(
        AesSbox_keyAdd_1_sbox_n56), .Z(AesSbox_keyAdd_1_sbox_n63) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0042 ( .A(AesSbox_keyAdd_1_sbox_n55), .B(
        AesSbox_keyAdd_1_sbox_n63), .Z(AesSbox_keyAdd_1_sbox_io_o0) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0041 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n62), .Z(AesSbox_keyAdd_1_sbox_n52) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0040 ( .A1(AesSbox_keyAdd_1_sbox_n60), .A2(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n51) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0039 ( .A1(AesSbox_keyAdd_1_sbox_n58), .A2(
        AesSbox_keyAdd_1_sbox_n59), .ZN(AesSbox_keyAdd_1_sbox_n57) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0038 ( .A(AesSbox_keyAdd_1_sbox_n56), .B(
        AesSbox_keyAdd_1_sbox_n57), .Z(AesSbox_keyAdd_1_sbox_n29) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0037 ( .A(AesSbox_keyAdd_1_sbox_n51), .B(
        AesSbox_keyAdd_1_sbox_n29), .ZN(AesSbox_keyAdd_1_sbox_n34) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0036 ( .A(AesSbox_keyAdd_1_sbox_n55), .ZN(
        AesSbox_keyAdd_1_sbox_n54) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0035 ( .A(AesSbox_keyAdd_1_sbox_n34), .B(
        AesSbox_keyAdd_1_sbox_n54), .Z(AesSbox_keyAdd_1_sbox_n53) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0034 ( .A(AesSbox_keyAdd_1_sbox_n52), .B(
        AesSbox_keyAdd_1_sbox_n53), .Z(AesSbox_keyAdd_1_sbox_io_o1) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0033 ( .A1(io_state[7]), .A2(
        AesSbox_keyAdd_1_sbox_n24), .ZN(AesSbox_keyAdd_1_sbox_n31) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0032 ( .A(AesSbox_keyAdd_1_sbox_n51), .B(
        AesSbox_keyAdd_1_sbox_n31), .ZN(AesSbox_keyAdd_1_sbox_n5) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0031 ( .A1(AesSbox_keyAdd_1_sbox_n50), .A2(
        AesSbox_keyAdd_1_sbox_n32), .ZN(AesSbox_keyAdd_1_sbox_n49) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0030 ( .A(AesSbox_keyAdd_1_sbox_n5), .B(
        AesSbox_keyAdd_1_sbox_n49), .ZN(AesSbox_keyAdd_1_sbox_n20) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0029 ( .A1(AesSbox_keyAdd_1_sbox_n47), .A2(
        AesSbox_keyAdd_1_sbox_n48), .ZN(AesSbox_keyAdd_1_sbox_n3) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0028 ( .A1(AesSbox_keyAdd_1_sbox_n45), .A2(
        AesSbox_keyAdd_1_sbox_n46), .ZN(AesSbox_keyAdd_1_sbox_n44) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0027 ( .A(AesSbox_keyAdd_1_sbox_n3), .B(
        AesSbox_keyAdd_1_sbox_n44), .ZN(AesSbox_keyAdd_1_sbox_n23) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0026 ( .A(AesSbox_keyAdd_1_sbox_n20), .B(
        AesSbox_keyAdd_1_sbox_n23), .ZN(AesSbox_keyAdd_1_sbox_n36) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0025 ( .A1(AesSbox_keyAdd_1_sbox_n42), .A2(
        AesSbox_keyAdd_1_sbox_n43), .ZN(AesSbox_keyAdd_1_sbox_n38) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0024 ( .A(AesSbox_keyAdd_1_sbox_n40), .B(
        AesSbox_keyAdd_1_sbox_n41), .Z(AesSbox_keyAdd_1_sbox_n39) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0023 ( .A(AesSbox_keyAdd_1_sbox_n38), .B(
        AesSbox_keyAdd_1_sbox_n39), .Z(AesSbox_keyAdd_1_sbox_n37) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0022 ( .A(AesSbox_keyAdd_1_sbox_n36), .B(
        AesSbox_keyAdd_1_sbox_n37), .Z(AesSbox_keyAdd_1_sbox_io_o2) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0021 ( .A(AesSbox_keyAdd_1_sbox_n35), .ZN(
        AesSbox_keyAdd_1_sbox_n19) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0020 ( .A(AesSbox_keyAdd_1_sbox_n19), .B(
        AesSbox_keyAdd_1_sbox_n34), .Z(AesSbox_keyAdd_1_sbox_io_o3) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U0019 ( .A1(AesSbox_keyAdd_1_sbox_n32), .A2(
        AesSbox_keyAdd_1_sbox_n33), .ZN(AesSbox_keyAdd_1_sbox_n12) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0018 ( .A(AesSbox_keyAdd_1_sbox_n31), .B(
        AesSbox_keyAdd_1_sbox_n12), .Z(AesSbox_keyAdd_1_sbox_n30) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0017 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n30), .Z(AesSbox_keyAdd_1_sbox_n26) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0016 ( .A(AesSbox_keyAdd_1_sbox_n28), .B(
        AesSbox_keyAdd_1_sbox_n29), .ZN(AesSbox_keyAdd_1_sbox_n27) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0015 ( .A(AesSbox_keyAdd_1_sbox_n26), .B(
        AesSbox_keyAdd_1_sbox_n27), .Z(AesSbox_keyAdd_1_sbox_io_o4) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0014 ( .A1(AesSbox_keyAdd_1_sbox_n24), .A2(
        AesSbox_keyAdd_1_sbox_n25), .ZN(AesSbox_keyAdd_1_sbox_n21) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0013 ( .A(AesSbox_keyAdd_1_sbox_n22), .B(
        AesSbox_keyAdd_1_sbox_n23), .Z(AesSbox_keyAdd_1_sbox_n10) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0012 ( .A(AesSbox_keyAdd_1_sbox_n21), .B(
        AesSbox_keyAdd_1_sbox_n10), .Z(AesSbox_keyAdd_1_sbox_n17) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0011 ( .A(AesSbox_keyAdd_1_sbox_n19), .B(
        AesSbox_keyAdd_1_sbox_n20), .Z(AesSbox_keyAdd_1_sbox_n18) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0010 ( .A(AesSbox_keyAdd_1_sbox_n17), .B(
        AesSbox_keyAdd_1_sbox_n18), .Z(AesSbox_keyAdd_1_sbox_io_o5) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U0009 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n16), .ZN(AesSbox_keyAdd_1_sbox_n8) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U0008 ( .A1(AesSbox_keyAdd_1_sbox_n13), .A2(
        AesSbox_keyAdd_1_sbox_n14), .ZN(AesSbox_keyAdd_1_sbox_n11) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0007 ( .A(AesSbox_keyAdd_1_sbox_n11), .B(
        AesSbox_keyAdd_1_sbox_n12), .Z(AesSbox_keyAdd_1_sbox_n7) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0006 ( .A(AesSbox_keyAdd_1_sbox_n7), .B(
        AesSbox_keyAdd_1_sbox_n10), .Z(AesSbox_keyAdd_1_sbox_n9) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0005 ( .A(AesSbox_keyAdd_1_sbox_n8), .B(
        AesSbox_keyAdd_1_sbox_n9), .Z(AesSbox_keyAdd_1_sbox_io_o6) );
  INV_X1 AesSbox_keyAdd_1_sbox_U0004 ( .A(AesSbox_keyAdd_1_sbox_n7), .ZN(
        AesSbox_keyAdd_1_sbox_n6) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0003 ( .A(AesSbox_keyAdd_1_sbox_n5), .B(
        AesSbox_keyAdd_1_sbox_n6), .Z(AesSbox_keyAdd_1_sbox_n1) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0002 ( .A(AesSbox_keyAdd_1_sbox_n3), .B(
        AesSbox_keyAdd_1_sbox_n4), .Z(AesSbox_keyAdd_1_sbox_n2) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U0001 ( .A(AesSbox_keyAdd_1_sbox_n1), .B(
        AesSbox_keyAdd_1_sbox_n2), .Z(AesSbox_keyAdd_1_sbox_io_o7) );
endmodule

