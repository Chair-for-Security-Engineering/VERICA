
module Sbox_andOptimized ( clock_0, reset_0, io_i0_s0, io_i0_s1, io_i1_s0, 
        io_i1_s1, io_i2_s0, io_i2_s1, io_i3_s0, io_i3_s1, io_k0_s0, io_k0_s1, 
        io_k1_s0, io_k1_s1, io_k2_s0, io_k2_s1, io_k3_s0, io_k3_s1, p_rand_0, 
        p_rand_1, p_rand_2, p_rand_3, io_o0_s0, io_o0_s1, io_o1_s0, io_o1_s1, 
        io_o2_s0, io_o2_s1, io_o3_s0, io_o3_s1 );
  input clock_0, reset_0, io_i0_s0, io_i0_s1, io_i1_s0, io_i1_s1, io_i2_s0,
         io_i2_s1, io_i3_s0, io_i3_s1, io_k0_s0, io_k0_s1, io_k1_s0, io_k1_s1,
         io_k2_s0, io_k2_s1, io_k3_s0, io_k3_s1, p_rand_0, p_rand_1, p_rand_2,
         p_rand_3;
  output io_o0_s0, io_o0_s1, io_o1_s0, io_o1_s1, io_o2_s0, io_o2_s1, io_o3_s0,
         io_o3_s1;
  wire   n_xor_module_1_res, n_xor_module_2_res, n_not_module_1_res,
         n_not_module_2_res, n_reg_module_1_res, n_not_module_3_res,
         n_and_module_1_res, n_xor_module_3_res, n_not_module_4_res,
         n_and_module_2_res, n_xor_module_4_res, n_reg_module_2_res,
         n_and_module_3_res, n_reg_module_3_res, n_reg_module_4_res,
         n_and_module_4_res, n_reg_module_5_res, n_reg_module_6_res,
         n_xor_module_5_res, n_xor_module_6_res, n_reg_module_7_res,
         n_and_module_5_res, n_reg_module_8_res, n_reg_module_9_res,
         n_and_module_6_res, n_reg_module_10_res, n_reg_module_11_res,
         n_xor_module_7_res, n_xor_module_8_res, n_xor_module_9_res,
         n_xor_module_10_res, n_xor_module_11_res, n_xor_module_12_res,
         n_xor_module_13_res, n_xor_module_14_res, n_not_module_5_res,
         n_xor_module_15_res, n_xor_module_16_res, n_xor_module_17_res,
         n_xor_module_18_res, n_xor_module_19_res, n_xor_module_20_res,
         n_not_module_6_res, n_reg_module_12_res, n_not_module_7_res,
         n_and_module_7_res, n_xor_module_21_res, n_not_module_8_res,
         n_and_module_8_res, n_xor_module_22_res, n_reg_module_13_res,
         n_and_module_9_res, n_reg_module_14_res, n_reg_module_15_res,
         n_and_module_10_res, n_reg_module_16_res, n_reg_module_17_res,
         n_xor_module_23_res, n_xor_module_24_res, n_reg_module_18_res,
         n_and_module_11_res, n_reg_module_19_res, n_reg_module_20_res,
         n_and_module_12_res, n_reg_module_21_res, n_reg_module_22_res,
         n_xor_module_25_res, n_xor_module_26_res, n_xor_module_27_res,
         n_xor_module_28_res, n_xor_module_29_res, n_xor_module_30_res,
         n_xor_module_31_res, n_xor_module_32_res, n_not_module_9_res,
         n_xor_module_33_res, n_xor_module_34_res, n_xor_module_35_res,
         n_xor_module_36_res, n_reg_module_23_res, n_not_module_10_res,
         n_and_module_13_res, n_xor_module_37_res, n_not_module_11_res,
         n_and_module_14_res, n_xor_module_38_res, n_reg_module_24_res,
         n_and_module_15_res, n_reg_module_25_res, n_reg_module_26_res,
         n_and_module_16_res, n_reg_module_27_res, n_reg_module_28_res,
         n_xor_module_39_res, n_xor_module_40_res, n_reg_module_29_res,
         n_and_module_17_res, n_reg_module_30_res, n_reg_module_31_res,
         n_and_module_18_res, n_reg_module_32_res, n_reg_module_33_res,
         n_xor_module_41_res, n_xor_module_42_res, n_reg_module_34_res,
         n_not_module_12_res, n_and_module_19_res, n_xor_module_43_res,
         n_not_module_13_res, n_and_module_20_res, n_xor_module_44_res,
         n_reg_module_35_res, n_and_module_21_res, n_reg_module_36_res,
         n_reg_module_37_res, n_and_module_22_res, n_reg_module_38_res,
         n_reg_module_39_res, n_xor_module_45_res, n_xor_module_46_res,
         n_reg_module_40_res, n_and_module_23_res, n_reg_module_41_res,
         n_reg_module_42_res, n_and_module_24_res, n_reg_module_43_res,
         n_reg_module_44_res, n_xor_module_47_res, n_xor_module_48_res,
         n_xor_module_49_res, n_xor_module_50_res, n_xor_module_51_res,
         n_xor_module_52_res, n_xor_module_53_res, n_xor_module_54_res,
         n_xor_module_55_res, n_xor_module_56_res, n_xor_module_57_res,
         n_xor_module_58_res, n_xor_module_59_res, n_xor_module_60_res,
         n_xor_module_61_res, n_xor_module_62_res, n_xor_module_63_res,
         n_xor_module_64_res, n_xor_module_65_res, n_xor_module_66_res,
         n_xor_module_67_res, n_xor_module_68_res, n_xor_module_69_res,
         n_xor_module_70_res;

  XOR2_X1 u_xor_module_1_U1 ( .A(io_i2_s0), .B(io_i1_s0), .Z(
        n_xor_module_1_res) );
  XOR2_X1 u_xor_module_2_U1 ( .A(io_i2_s1), .B(io_i1_s1), .Z(
        n_xor_module_2_res) );
  INV_X1 u_not_module_1_U1 ( .A(n_xor_module_1_res), .ZN(n_not_module_1_res)
         );
  INV_X1 u_not_module_2_U1 ( .A(io_i0_s0), .ZN(n_not_module_2_res) );
  DFF_X1 u_reg_module_1__hpc_r0_reg ( .D(p_rand_0), .CK(clock_0), .Q(
        n_reg_module_1_res), .QN() );
  INV_X1 u_not_module_3_U1 ( .A(n_not_module_1_res), .ZN(n_not_module_3_res)
         );
  AND2_X1 u_and_module_1_U1 ( .A1(n_not_module_3_res), .A2(n_reg_module_1_res), 
        .ZN(n_and_module_1_res) );
  XOR2_X1 u_xor_module_3_U1 ( .A(p_rand_0), .B(io_i0_s1), .Z(
        n_xor_module_3_res) );
  INV_X1 u_not_module_4_U1 ( .A(n_xor_module_2_res), .ZN(n_not_module_4_res)
         );
  AND2_X1 u_and_module_2_U1 ( .A1(n_not_module_4_res), .A2(n_reg_module_1_res), 
        .ZN(n_and_module_2_res) );
  XOR2_X1 u_xor_module_4_U1 ( .A(p_rand_0), .B(n_not_module_2_res), .Z(
        n_xor_module_4_res) );
  DFF_X1 u_reg_module_2__hpc_r0_reg ( .D(n_not_module_2_res), .CK(clock_0), 
        .Q(n_reg_module_2_res), .QN() );
  AND2_X1 u_and_module_3_U1 ( .A1(n_reg_module_2_res), .A2(n_not_module_1_res), 
        .ZN(n_and_module_3_res) );
  DFF_X1 u_reg_module_3__hpc_r0_reg ( .D(n_and_module_3_res), .CK(clock_0), 
        .Q(n_reg_module_3_res), .QN() );
  DFF_X1 u_reg_module_4__hpc_r0_reg ( .D(n_xor_module_3_res), .CK(clock_0), 
        .Q(n_reg_module_4_res), .QN() );
  AND2_X1 u_and_module_4_U1 ( .A1(n_reg_module_4_res), .A2(n_not_module_1_res), 
        .ZN(n_and_module_4_res) );
  DFF_X1 u_reg_module_5__hpc_r0_reg ( .D(n_and_module_4_res), .CK(clock_0), 
        .Q(n_reg_module_5_res), .QN() );
  DFF_X1 u_reg_module_6__hpc_r0_reg ( .D(n_and_module_1_res), .CK(clock_0), 
        .Q(n_reg_module_6_res), .QN() );
  XOR2_X1 u_xor_module_5_U1 ( .A(n_reg_module_6_res), .B(n_reg_module_5_res), 
        .Z(n_xor_module_5_res) );
  XOR2_X1 u_xor_module_6_U1 ( .A(n_xor_module_5_res), .B(n_reg_module_3_res), 
        .Z(n_xor_module_6_res) );
  DFF_X1 u_reg_module_7__hpc_r0_reg ( .D(io_i0_s1), .CK(clock_0), .Q(
        n_reg_module_7_res), .QN() );
  AND2_X1 u_and_module_5_U1 ( .A1(n_reg_module_7_res), .A2(n_xor_module_2_res), 
        .ZN(n_and_module_5_res) );
  DFF_X1 u_reg_module_8__hpc_r0_reg ( .D(n_and_module_5_res), .CK(clock_0), 
        .Q(n_reg_module_8_res), .QN() );
  DFF_X1 u_reg_module_9__hpc_r0_reg ( .D(n_xor_module_4_res), .CK(clock_0), 
        .Q(n_reg_module_9_res), .QN() );
  AND2_X1 u_and_module_6_U1 ( .A1(n_reg_module_9_res), .A2(n_xor_module_2_res), 
        .ZN(n_and_module_6_res) );
  DFF_X1 u_reg_module_10__hpc_r0_reg ( .D(n_and_module_6_res), .CK(clock_0), 
        .Q(n_reg_module_10_res), .QN() );
  DFF_X1 u_reg_module_11__hpc_r0_reg ( .D(n_and_module_2_res), .CK(clock_0), 
        .Q(n_reg_module_11_res), .QN() );
  XOR2_X1 u_xor_module_7_U1 ( .A(n_reg_module_11_res), .B(n_reg_module_10_res), 
        .Z(n_xor_module_7_res) );
  XOR2_X1 u_xor_module_8_U1 ( .A(n_xor_module_7_res), .B(n_reg_module_8_res), 
        .Z(n_xor_module_8_res) );
  XOR2_X1 u_xor_module_9_U1 ( .A(io_i2_s0), .B(io_i0_s0), .Z(
        n_xor_module_9_res) );
  XOR2_X1 u_xor_module_10_U1 ( .A(io_i2_s1), .B(io_i0_s1), .Z(
        n_xor_module_10_res) );
  XOR2_X1 u_xor_module_11_U1 ( .A(io_i3_s0), .B(n_xor_module_9_res), .Z(
        n_xor_module_11_res) );
  XOR2_X1 u_xor_module_12_U1 ( .A(io_i3_s1), .B(n_xor_module_10_res), .Z(
        n_xor_module_12_res) );
  XOR2_X1 u_xor_module_13_U1 ( .A(n_xor_module_6_res), .B(n_xor_module_11_res), 
        .Z(n_xor_module_13_res) );
  XOR2_X1 u_xor_module_14_U1 ( .A(n_xor_module_8_res), .B(n_xor_module_12_res), 
        .Z(n_xor_module_14_res) );
  INV_X1 u_not_module_5_U1 ( .A(n_xor_module_13_res), .ZN(n_not_module_5_res)
         );
  XOR2_X1 u_xor_module_15_U1 ( .A(io_i1_s0), .B(io_i0_s0), .Z(
        n_xor_module_15_res) );
  XOR2_X1 u_xor_module_16_U1 ( .A(io_i1_s1), .B(io_i0_s1), .Z(
        n_xor_module_16_res) );
  XOR2_X1 u_xor_module_17_U1 ( .A(io_i2_s0), .B(n_xor_module_15_res), .Z(
        n_xor_module_17_res) );
  XOR2_X1 u_xor_module_18_U1 ( .A(io_i2_s1), .B(n_xor_module_16_res), .Z(
        n_xor_module_18_res) );
  XOR2_X1 u_xor_module_19_U1 ( .A(io_i3_s0), .B(n_xor_module_17_res), .Z(
        n_xor_module_19_res) );
  XOR2_X1 u_xor_module_20_U1 ( .A(io_i3_s1), .B(n_xor_module_18_res), .Z(
        n_xor_module_20_res) );
  INV_X1 u_not_module_6_U1 ( .A(io_i2_s0), .ZN(n_not_module_6_res) );
  DFF_X1 u_reg_module_12__hpc_r0_reg ( .D(p_rand_1), .CK(clock_0), .Q(
        n_reg_module_12_res), .QN() );
  INV_X1 u_not_module_7_U1 ( .A(n_not_module_6_res), .ZN(n_not_module_7_res)
         );
  AND2_X1 u_and_module_7_U1 ( .A1(n_not_module_7_res), .A2(n_reg_module_12_res), .ZN(n_and_module_7_res) );
  XOR2_X1 u_xor_module_21_U1 ( .A(p_rand_1), .B(io_i1_s1), .Z(
        n_xor_module_21_res) );
  INV_X1 u_not_module_8_U1 ( .A(io_i2_s1), .ZN(n_not_module_8_res) );
  AND2_X1 u_and_module_8_U1 ( .A1(n_not_module_8_res), .A2(n_reg_module_12_res), .ZN(n_and_module_8_res) );
  XOR2_X1 u_xor_module_22_U1 ( .A(p_rand_1), .B(io_i1_s0), .Z(
        n_xor_module_22_res) );
  DFF_X1 u_reg_module_13__hpc_r0_reg ( .D(io_i1_s0), .CK(clock_0), .Q(
        n_reg_module_13_res), .QN() );
  AND2_X1 u_and_module_9_U1 ( .A1(n_reg_module_13_res), .A2(n_not_module_6_res), .ZN(n_and_module_9_res) );
  DFF_X1 u_reg_module_14__hpc_r0_reg ( .D(n_and_module_9_res), .CK(clock_0), 
        .Q(n_reg_module_14_res), .QN() );
  DFF_X1 u_reg_module_15__hpc_r0_reg ( .D(n_xor_module_21_res), .CK(clock_0), 
        .Q(n_reg_module_15_res), .QN() );
  AND2_X1 u_and_module_10_U1 ( .A1(n_reg_module_15_res), .A2(
        n_not_module_6_res), .ZN(n_and_module_10_res) );
  DFF_X1 u_reg_module_16__hpc_r0_reg ( .D(n_and_module_10_res), .CK(clock_0), 
        .Q(n_reg_module_16_res), .QN() );
  DFF_X1 u_reg_module_17__hpc_r0_reg ( .D(n_and_module_7_res), .CK(clock_0), 
        .Q(n_reg_module_17_res), .QN() );
  XOR2_X1 u_xor_module_23_U1 ( .A(n_reg_module_17_res), .B(n_reg_module_16_res), .Z(n_xor_module_23_res) );
  XOR2_X1 u_xor_module_24_U1 ( .A(n_xor_module_23_res), .B(n_reg_module_14_res), .Z(n_xor_module_24_res) );
  DFF_X1 u_reg_module_18__hpc_r0_reg ( .D(io_i1_s1), .CK(clock_0), .Q(
        n_reg_module_18_res), .QN() );
  AND2_X1 u_and_module_11_U1 ( .A1(n_reg_module_18_res), .A2(io_i2_s1), .ZN(
        n_and_module_11_res) );
  DFF_X1 u_reg_module_19__hpc_r0_reg ( .D(n_and_module_11_res), .CK(clock_0), 
        .Q(n_reg_module_19_res), .QN() );
  DFF_X1 u_reg_module_20__hpc_r0_reg ( .D(n_xor_module_22_res), .CK(clock_0), 
        .Q(n_reg_module_20_res), .QN() );
  AND2_X1 u_and_module_12_U1 ( .A1(n_reg_module_20_res), .A2(io_i2_s1), .ZN(
        n_and_module_12_res) );
  DFF_X1 u_reg_module_21__hpc_r0_reg ( .D(n_and_module_12_res), .CK(clock_0), 
        .Q(n_reg_module_21_res), .QN() );
  DFF_X1 u_reg_module_22__hpc_r0_reg ( .D(n_and_module_8_res), .CK(clock_0), 
        .Q(n_reg_module_22_res), .QN() );
  XOR2_X1 u_xor_module_25_U1 ( .A(n_reg_module_22_res), .B(n_reg_module_21_res), .Z(n_xor_module_25_res) );
  XOR2_X1 u_xor_module_26_U1 ( .A(n_xor_module_25_res), .B(n_reg_module_19_res), .Z(n_xor_module_26_res) );
  XOR2_X1 u_xor_module_27_U1 ( .A(io_i2_s0), .B(io_i0_s0), .Z(
        n_xor_module_27_res) );
  XOR2_X1 u_xor_module_28_U1 ( .A(io_i2_s1), .B(io_i0_s1), .Z(
        n_xor_module_28_res) );
  XOR2_X1 u_xor_module_29_U1 ( .A(n_xor_module_6_res), .B(n_xor_module_27_res), 
        .Z(n_xor_module_29_res) );
  XOR2_X1 u_xor_module_30_U1 ( .A(n_xor_module_8_res), .B(n_xor_module_28_res), 
        .Z(n_xor_module_30_res) );
  XOR2_X1 u_xor_module_31_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_29_res), .Z(n_xor_module_31_res) );
  XOR2_X1 u_xor_module_32_U1 ( .A(n_xor_module_26_res), .B(n_xor_module_30_res), .Z(n_xor_module_32_res) );
  INV_X1 u_not_module_9_U1 ( .A(n_xor_module_31_res), .ZN(n_not_module_9_res)
         );
  XOR2_X1 u_xor_module_33_U1 ( .A(io_i2_s0), .B(io_i1_s0), .Z(
        n_xor_module_33_res) );
  XOR2_X1 u_xor_module_34_U1 ( .A(io_i2_s1), .B(io_i1_s1), .Z(
        n_xor_module_34_res) );
  XOR2_X1 u_xor_module_35_U1 ( .A(io_i3_s0), .B(n_xor_module_33_res), .Z(
        n_xor_module_35_res) );
  XOR2_X1 u_xor_module_36_U1 ( .A(io_i3_s1), .B(n_xor_module_34_res), .Z(
        n_xor_module_36_res) );
  DFF_X1 u_reg_module_23__hpc_r0_reg ( .D(p_rand_2), .CK(clock_0), .Q(
        n_reg_module_23_res), .QN() );
  INV_X1 u_not_module_10_U1 ( .A(n_not_module_5_res), .ZN(n_not_module_10_res)
         );
  AND2_X1 u_and_module_13_U1 ( .A1(n_not_module_10_res), .A2(
        n_reg_module_23_res), .ZN(n_and_module_13_res) );
  XOR2_X1 u_xor_module_37_U1 ( .A(p_rand_2), .B(n_xor_module_20_res), .Z(
        n_xor_module_37_res) );
  INV_X1 u_not_module_11_U1 ( .A(n_xor_module_14_res), .ZN(n_not_module_11_res) );
  AND2_X1 u_and_module_14_U1 ( .A1(n_not_module_11_res), .A2(
        n_reg_module_23_res), .ZN(n_and_module_14_res) );
  XOR2_X1 u_xor_module_38_U1 ( .A(p_rand_2), .B(n_xor_module_19_res), .Z(
        n_xor_module_38_res) );
  DFF_X1 u_reg_module_24__hpc_r0_reg ( .D(n_xor_module_19_res), .CK(clock_0), 
        .Q(n_reg_module_24_res), .QN() );
  AND2_X1 u_and_module_15_U1 ( .A1(n_reg_module_24_res), .A2(
        n_not_module_5_res), .ZN(n_and_module_15_res) );
  DFF_X1 u_reg_module_25__hpc_r0_reg ( .D(n_and_module_15_res), .CK(clock_0), 
        .Q(n_reg_module_25_res), .QN() );
  DFF_X1 u_reg_module_26__hpc_r0_reg ( .D(n_xor_module_37_res), .CK(clock_0), 
        .Q(n_reg_module_26_res), .QN() );
  AND2_X1 u_and_module_16_U1 ( .A1(n_reg_module_26_res), .A2(
        n_not_module_5_res), .ZN(n_and_module_16_res) );
  DFF_X1 u_reg_module_27__hpc_r0_reg ( .D(n_and_module_16_res), .CK(clock_0), 
        .Q(n_reg_module_27_res), .QN() );
  DFF_X1 u_reg_module_28__hpc_r0_reg ( .D(n_and_module_13_res), .CK(clock_0), 
        .Q(n_reg_module_28_res), .QN() );
  XOR2_X1 u_xor_module_39_U1 ( .A(n_reg_module_28_res), .B(n_reg_module_27_res), .Z(n_xor_module_39_res) );
  XOR2_X1 u_xor_module_40_U1 ( .A(n_xor_module_39_res), .B(n_reg_module_25_res), .Z(n_xor_module_40_res) );
  DFF_X1 u_reg_module_29__hpc_r0_reg ( .D(n_xor_module_20_res), .CK(clock_0), 
        .Q(n_reg_module_29_res), .QN() );
  AND2_X1 u_and_module_17_U1 ( .A1(n_reg_module_29_res), .A2(
        n_xor_module_14_res), .ZN(n_and_module_17_res) );
  DFF_X1 u_reg_module_30__hpc_r0_reg ( .D(n_and_module_17_res), .CK(clock_0), 
        .Q(n_reg_module_30_res), .QN() );
  DFF_X1 u_reg_module_31__hpc_r0_reg ( .D(n_xor_module_38_res), .CK(clock_0), 
        .Q(n_reg_module_31_res), .QN() );
  AND2_X1 u_and_module_18_U1 ( .A1(n_reg_module_31_res), .A2(
        n_xor_module_14_res), .ZN(n_and_module_18_res) );
  DFF_X1 u_reg_module_32__hpc_r0_reg ( .D(n_and_module_18_res), .CK(clock_0), 
        .Q(n_reg_module_32_res), .QN() );
  DFF_X1 u_reg_module_33__hpc_r0_reg ( .D(n_and_module_14_res), .CK(clock_0), 
        .Q(n_reg_module_33_res), .QN() );
  XOR2_X1 u_xor_module_41_U1 ( .A(n_reg_module_33_res), .B(n_reg_module_32_res), .Z(n_xor_module_41_res) );
  XOR2_X1 u_xor_module_42_U1 ( .A(n_xor_module_41_res), .B(n_reg_module_30_res), .Z(n_xor_module_42_res) );
  DFF_X1 u_reg_module_34__hpc_r0_reg ( .D(p_rand_3), .CK(clock_0), .Q(
        n_reg_module_34_res), .QN() );
  INV_X1 u_not_module_12_U1 ( .A(n_not_module_9_res), .ZN(n_not_module_12_res)
         );
  AND2_X1 u_and_module_19_U1 ( .A1(n_not_module_12_res), .A2(
        n_reg_module_34_res), .ZN(n_and_module_19_res) );
  XOR2_X1 u_xor_module_43_U1 ( .A(p_rand_3), .B(n_xor_module_36_res), .Z(
        n_xor_module_43_res) );
  INV_X1 u_not_module_13_U1 ( .A(n_xor_module_32_res), .ZN(n_not_module_13_res) );
  AND2_X1 u_and_module_20_U1 ( .A1(n_not_module_13_res), .A2(
        n_reg_module_34_res), .ZN(n_and_module_20_res) );
  XOR2_X1 u_xor_module_44_U1 ( .A(p_rand_3), .B(n_xor_module_35_res), .Z(
        n_xor_module_44_res) );
  DFF_X1 u_reg_module_35__hpc_r0_reg ( .D(n_xor_module_35_res), .CK(clock_0), 
        .Q(n_reg_module_35_res), .QN() );
  AND2_X1 u_and_module_21_U1 ( .A1(n_reg_module_35_res), .A2(
        n_not_module_9_res), .ZN(n_and_module_21_res) );
  DFF_X1 u_reg_module_36__hpc_r0_reg ( .D(n_and_module_21_res), .CK(clock_0), 
        .Q(n_reg_module_36_res), .QN() );
  DFF_X1 u_reg_module_37__hpc_r0_reg ( .D(n_xor_module_43_res), .CK(clock_0), 
        .Q(n_reg_module_37_res), .QN() );
  AND2_X1 u_and_module_22_U1 ( .A1(n_reg_module_37_res), .A2(
        n_not_module_9_res), .ZN(n_and_module_22_res) );
  DFF_X1 u_reg_module_38__hpc_r0_reg ( .D(n_and_module_22_res), .CK(clock_0), 
        .Q(n_reg_module_38_res), .QN() );
  DFF_X1 u_reg_module_39__hpc_r0_reg ( .D(n_and_module_19_res), .CK(clock_0), 
        .Q(n_reg_module_39_res), .QN() );
  XOR2_X1 u_xor_module_45_U1 ( .A(n_reg_module_39_res), .B(n_reg_module_38_res), .Z(n_xor_module_45_res) );
  XOR2_X1 u_xor_module_46_U1 ( .A(n_xor_module_45_res), .B(n_reg_module_36_res), .Z(n_xor_module_46_res) );
  DFF_X1 u_reg_module_40__hpc_r0_reg ( .D(n_xor_module_36_res), .CK(clock_0), 
        .Q(n_reg_module_40_res), .QN() );
  AND2_X1 u_and_module_23_U1 ( .A1(n_reg_module_40_res), .A2(
        n_xor_module_32_res), .ZN(n_and_module_23_res) );
  DFF_X1 u_reg_module_41__hpc_r0_reg ( .D(n_and_module_23_res), .CK(clock_0), 
        .Q(n_reg_module_41_res), .QN() );
  DFF_X1 u_reg_module_42__hpc_r0_reg ( .D(n_xor_module_44_res), .CK(clock_0), 
        .Q(n_reg_module_42_res), .QN() );
  AND2_X1 u_and_module_24_U1 ( .A1(n_reg_module_42_res), .A2(
        n_xor_module_32_res), .ZN(n_and_module_24_res) );
  DFF_X1 u_reg_module_43__hpc_r0_reg ( .D(n_and_module_24_res), .CK(clock_0), 
        .Q(n_reg_module_43_res), .QN() );
  DFF_X1 u_reg_module_44__hpc_r0_reg ( .D(n_and_module_20_res), .CK(clock_0), 
        .Q(n_reg_module_44_res), .QN() );
  XOR2_X1 u_xor_module_47_U1 ( .A(n_reg_module_44_res), .B(n_reg_module_43_res), .Z(n_xor_module_47_res) );
  XOR2_X1 u_xor_module_48_U1 ( .A(n_xor_module_47_res), .B(n_reg_module_41_res), .Z(n_xor_module_48_res) );
  XOR2_X1 u_xor_module_49_U1 ( .A(n_xor_module_6_res), .B(io_i3_s0), .Z(
        n_xor_module_49_res) );
  XOR2_X1 u_xor_module_50_U1 ( .A(n_xor_module_8_res), .B(io_i3_s1), .Z(
        n_xor_module_50_res) );
  XOR2_X1 u_xor_module_51_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_49_res), .Z(n_xor_module_51_res) );
  XOR2_X1 u_xor_module_52_U1 ( .A(n_xor_module_26_res), .B(n_xor_module_50_res), .Z(n_xor_module_52_res) );
  XOR2_X1 u_xor_module_53_U1 ( .A(n_xor_module_46_res), .B(n_xor_module_51_res), .Z(n_xor_module_53_res) );
  XOR2_X1 u_xor_module_54_U1 ( .A(n_xor_module_48_res), .B(n_xor_module_52_res), .Z(n_xor_module_54_res) );
  XOR2_X1 u_xor_module_55_U1 ( .A(io_i3_s0), .B(io_i2_s0), .Z(
        n_xor_module_55_res) );
  XOR2_X1 u_xor_module_56_U1 ( .A(io_i3_s1), .B(io_i2_s1), .Z(
        n_xor_module_56_res) );
  XOR2_X1 u_xor_module_57_U1 ( .A(n_xor_module_6_res), .B(n_xor_module_55_res), 
        .Z(n_xor_module_57_res) );
  XOR2_X1 u_xor_module_58_U1 ( .A(n_xor_module_8_res), .B(n_xor_module_56_res), 
        .Z(n_xor_module_58_res) );
  XOR2_X1 u_xor_module_59_U1 ( .A(n_xor_module_40_res), .B(n_xor_module_57_res), .Z(n_xor_module_59_res) );
  XOR2_X1 u_xor_module_60_U1 ( .A(n_xor_module_42_res), .B(n_xor_module_58_res), .Z(n_xor_module_60_res) );
  XOR2_X1 u_xor_module_61_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_59_res), .Z(n_xor_module_61_res) );
  XOR2_X1 u_xor_module_62_U1 ( .A(n_xor_module_26_res), .B(n_xor_module_60_res), .Z(n_xor_module_62_res) );
  XOR2_X1 u_xor_module_63_U1 ( .A(io_i2_s0), .B(io_i0_s0), .Z(
        n_xor_module_63_res) );
  XOR2_X1 u_xor_module_64_U1 ( .A(io_i2_s1), .B(io_i0_s1), .Z(
        n_xor_module_64_res) );
  XOR2_X1 u_xor_module_65_U1 ( .A(n_xor_module_46_res), .B(n_xor_module_63_res), .Z(n_xor_module_65_res) );
  XOR2_X1 u_xor_module_66_U1 ( .A(n_xor_module_48_res), .B(n_xor_module_64_res), .Z(n_xor_module_66_res) );
  XOR2_X1 u_xor_module_67_U1 ( .A(io_i3_s0), .B(io_i0_s0), .Z(
        n_xor_module_67_res) );
  XOR2_X1 u_xor_module_68_U1 ( .A(io_i3_s1), .B(io_i0_s1), .Z(
        n_xor_module_68_res) );
  XOR2_X1 u_xor_module_69_U1 ( .A(n_xor_module_24_res), .B(n_xor_module_67_res), .Z(n_xor_module_69_res) );
  XOR2_X1 u_xor_module_70_U1 ( .A(n_xor_module_26_res), .B(n_xor_module_68_res), .Z(n_xor_module_70_res) );
  XOR2_X1 u_xor_module_71_U1 ( .A(io_k0_s0), .B(n_xor_module_53_res), .Z(
        io_o0_s0) );
  XOR2_X1 u_xor_module_72_U1 ( .A(io_k0_s1), .B(n_xor_module_54_res), .Z(
        io_o0_s1) );
  XOR2_X1 u_xor_module_73_U1 ( .A(io_k1_s0), .B(n_xor_module_61_res), .Z(
        io_o1_s0) );
  XOR2_X1 u_xor_module_74_U1 ( .A(io_k1_s1), .B(n_xor_module_62_res), .Z(
        io_o1_s1) );
  XOR2_X1 u_xor_module_75_U1 ( .A(io_k2_s0), .B(n_xor_module_65_res), .Z(
        io_o2_s0) );
  XOR2_X1 u_xor_module_76_U1 ( .A(io_k2_s1), .B(n_xor_module_66_res), .Z(
        io_o2_s1) );
  XOR2_X1 u_xor_module_77_U1 ( .A(io_k3_s0), .B(n_xor_module_69_res), .Z(
        io_o3_s0) );
  XOR2_X1 u_xor_module_78_U1 ( .A(io_k3_s1), .B(n_xor_module_70_res), .Z(
        io_o3_s1) );
endmodule

