module KeyAddition ( clock, reset, io_state, io_key, io_out );
  input [15:0] io_state;
  input [15:0] io_key;
  output [15:0] io_out;
  input clock, reset;


  XOR2_X1 U17 ( .A(io_state[9]), .B(io_key[9]), .Z(io_out[9]) );
  XOR2_X1 U18 ( .A(io_state[8]), .B(io_key[8]), .Z(io_out[8]) );
  XOR2_X1 U19 ( .A(io_state[7]), .B(io_key[7]), .Z(io_out[7]) );
  XOR2_X1 U20 ( .A(io_state[6]), .B(io_key[6]), .Z(io_out[6]) );
  XOR2_X1 U21 ( .A(io_state[5]), .B(io_key[5]), .Z(io_out[5]) );
  XOR2_X1 U22 ( .A(io_state[4]), .B(io_key[4]), .Z(io_out[4]) );
  XOR2_X1 U23 ( .A(io_state[3]), .B(io_key[3]), .Z(io_out[3]) );
  XOR2_X1 U24 ( .A(io_state[2]), .B(io_key[2]), .Z(io_out[2]) );
  XOR2_X1 U25 ( .A(io_state[1]), .B(io_key[1]), .Z(io_out[1]) );
  XOR2_X1 U26 ( .A(io_state[15]), .B(io_key[15]), .Z(io_out[15]) );
  XOR2_X1 U27 ( .A(io_state[14]), .B(io_key[14]), .Z(io_out[14]) );
  XOR2_X1 U28 ( .A(io_state[13]), .B(io_key[13]), .Z(io_out[13]) );
  XOR2_X1 U29 ( .A(io_state[12]), .B(io_key[12]), .Z(io_out[12]) );
  XOR2_X1 U30 ( .A(io_state[11]), .B(io_key[11]), .Z(io_out[11]) );
  XOR2_X1 U31 ( .A(io_state[10]), .B(io_key[10]), .Z(io_out[10]) );
  XOR2_X1 U32 ( .A(io_state[0]), .B(io_key[0]), .Z(io_out[0]) );
endmodule
