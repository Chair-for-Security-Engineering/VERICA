
module CINI ( io_a_0, io_a_1, io_b_0, io_b_1, io_c_0, io_c_1, io_rand, clk, 
        reset );
  input [4:0] io_a_0;
  input [4:0] io_a_1;
  input [4:0] io_b_0;
  input [4:0] io_b_1;
  output [4:0] io_c_0;
  output [4:0] io_c_1;
  input [0:0] io_rand;
  input clk, reset;
  wire   simpleNot_10_port_z, simpleNot_11_port_z, simpleNot_12_port_z,
         simpleNot_13_port_z, simpleNot_14_port_z, simpleNot_15_port_z,
         simpleNot_16_port_z, simpleNot_17_port_z, simpleNot_18_port_z,
         simpleNot_19_port_z, simpleXor_10_port_z, simpleXor_11_port_z,
         simpleXor_12_port_z, simpleXor_13_port_z, simpleXor_14_port_z,
         simpleXor_15_port_z, simpleXor_16_port_z, simpleXor_17_port_z,
         simpleXor_18_port_z, simpleXor_19_port_z, n_zz_io_c_0_2_1_,
         n_zz_io_c_0_0_, n_zz_io_c_1_2_1_, n_zz_io_c_1_0_, n_zz_io_c_0_5_1_,
         n_zz_io_c_0_3_0_, n_zz_io_c_1_5_1_, n_zz_io_c_1_3_0_,
         n_zz_io_c_0_8_1_, n_zz_io_c_0_6_0_, n_zz_io_c_1_8_1_,
         n_zz_io_c_1_6_0_, n_zz_io_c_0_11_1_, n_zz_io_c_0_9_0_,
         n_zz_io_c_1_11_1_, n_zz_io_c_1_9_0_, n_zz_io_c_0_14_1_,
         n_zz_io_c_0_12_0_, n_zz_io_c_1_14_1_, n_zz_io_c_1_12_0_, N0, N1, N2,
         N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         cor_maj_19_port_o, cor_maj_18_port_o, cor_maj_17_port_o,
         cor_maj_16_port_o, cor_maj_15_port_o, cor_maj_14_port_o,
         cor_maj_13_port_o, cor_maj_12_port_o, cor_maj_11_port_o,
         cor_maj_10_port_o, cor_maj_10_n13, cor_maj_10_n12, cor_maj_10_n11,
         cor_maj_10_n10, cor_maj_10_n9, cor_maj_10_n8, cor_maj_10_n7,
         cor_maj_10_n6, cor_maj_10_n5, cor_maj_10_n4, cor_maj_10_n3,
         cor_maj_10_n2, cor_maj_10_n1, cor_maj_11_n26, cor_maj_11_n25,
         cor_maj_11_n24, cor_maj_11_n23, cor_maj_11_n22, cor_maj_11_n21,
         cor_maj_11_n20, cor_maj_11_n19, cor_maj_11_n18, cor_maj_11_n17,
         cor_maj_11_n16, cor_maj_11_n15, cor_maj_11_n14, cor_maj_12_n26,
         cor_maj_12_n25, cor_maj_12_n24, cor_maj_12_n23, cor_maj_12_n22,
         cor_maj_12_n21, cor_maj_12_n20, cor_maj_12_n19, cor_maj_12_n18,
         cor_maj_12_n17, cor_maj_12_n16, cor_maj_12_n15, cor_maj_12_n14,
         cor_maj_13_n26, cor_maj_13_n25, cor_maj_13_n24, cor_maj_13_n23,
         cor_maj_13_n22, cor_maj_13_n21, cor_maj_13_n20, cor_maj_13_n19,
         cor_maj_13_n18, cor_maj_13_n17, cor_maj_13_n16, cor_maj_13_n15,
         cor_maj_13_n14, cor_maj_14_n26, cor_maj_14_n25, cor_maj_14_n24,
         cor_maj_14_n23, cor_maj_14_n22, cor_maj_14_n21, cor_maj_14_n20,
         cor_maj_14_n19, cor_maj_14_n18, cor_maj_14_n17, cor_maj_14_n16,
         cor_maj_14_n15, cor_maj_14_n14, cor_maj_15_n26, cor_maj_15_n25,
         cor_maj_15_n24, cor_maj_15_n23, cor_maj_15_n22, cor_maj_15_n21,
         cor_maj_15_n20, cor_maj_15_n19, cor_maj_15_n18, cor_maj_15_n17,
         cor_maj_15_n16, cor_maj_15_n15, cor_maj_15_n14, cor_maj_16_n26,
         cor_maj_16_n25, cor_maj_16_n24, cor_maj_16_n23, cor_maj_16_n22,
         cor_maj_16_n21, cor_maj_16_n20, cor_maj_16_n19, cor_maj_16_n18,
         cor_maj_16_n17, cor_maj_16_n16, cor_maj_16_n15, cor_maj_16_n14,
         cor_maj_17_n26, cor_maj_17_n25, cor_maj_17_n24, cor_maj_17_n23,
         cor_maj_17_n22, cor_maj_17_n21, cor_maj_17_n20, cor_maj_17_n19,
         cor_maj_17_n18, cor_maj_17_n17, cor_maj_17_n16, cor_maj_17_n15,
         cor_maj_17_n14, cor_maj_18_n26, cor_maj_18_n25, cor_maj_18_n24,
         cor_maj_18_n23, cor_maj_18_n22, cor_maj_18_n21, cor_maj_18_n20,
         cor_maj_18_n19, cor_maj_18_n18, cor_maj_18_n17, cor_maj_18_n16,
         cor_maj_18_n15, cor_maj_18_n14, cor_maj_19_n26, cor_maj_19_n25,
         cor_maj_19_n24, cor_maj_19_n23, cor_maj_19_n22, cor_maj_19_n21,
         cor_maj_19_n20, cor_maj_19_n19, cor_maj_19_n18, cor_maj_19_n17,
         cor_maj_19_n16, cor_maj_19_n15, cor_maj_19_n14;
  wire   [4:0] v_1_0_1;
  wire   [4:0] v_1_1_0;
  wire   [4:0] cor_port_v_0_1;
  wire   [4:0] cor_port_v_1_0;
  wire   [4:0] u_0_1;
  wire   [4:0] u_1_0;
  wire   [4:0] rand_reg_0;
  wire   [4:0] rand_reg_1;
  wire   [4:0] b_reg_0;
  wire   [4:0] b_reg_1;

  DFF_X1 b_reg_1_reg_4_ ( .D(io_b_1[4]), .CK(clk), .Q(b_reg_1[4]), .QN() );
  DFF_X1 b_reg_1_reg_3_ ( .D(io_b_1[3]), .CK(clk), .Q(b_reg_1[3]), .QN() );
  DFF_X1 b_reg_1_reg_2_ ( .D(io_b_1[2]), .CK(clk), .Q(b_reg_1[2]), .QN() );
  DFF_X1 b_reg_1_reg_1_ ( .D(io_b_1[1]), .CK(clk), .Q(b_reg_1[1]), .QN() );
  DFF_X1 b_reg_1_reg_0_ ( .D(io_b_1[0]), .CK(clk), .Q(b_reg_1[0]), .QN() );
  DFF_X1 u_zz_io_c_0_2_reg_1_ ( .D(N11), .CK(clk), .Q(n_zz_io_c_0_2_1_), .QN()
         );
  DFF_X1 b_reg_0_reg_4_ ( .D(io_b_0[4]), .CK(clk), .Q(b_reg_0[4]), .QN() );
  DFF_X1 b_reg_0_reg_3_ ( .D(io_b_0[3]), .CK(clk), .Q(b_reg_0[3]), .QN() );
  DFF_X1 b_reg_0_reg_2_ ( .D(io_b_0[2]), .CK(clk), .Q(b_reg_0[2]), .QN() );
  DFF_X1 b_reg_0_reg_1_ ( .D(io_b_0[1]), .CK(clk), .Q(b_reg_0[1]), .QN() );
  DFF_X1 b_reg_0_reg_0_ ( .D(io_b_0[0]), .CK(clk), .Q(b_reg_0[0]), .QN() );
  DFF_X1 u_zz_io_c_0_2_reg_0_ ( .D(N10), .CK(clk), .Q(n_zz_io_c_0_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_14_reg_1_ ( .D(N29), .CK(clk), .Q(n_zz_io_c_1_14_1_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_14_reg_0_ ( .D(N28), .CK(clk), .Q(n_zz_io_c_1_12_0_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_1_ ( .D(N27), .CK(clk), .Q(n_zz_io_c_0_14_1_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_14_reg_0_ ( .D(N26), .CK(clk), .Q(n_zz_io_c_0_12_0_), 
        .QN() );
  DFF_X1 rand_reg_0_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[4]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[3]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[2]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[1]), 
        .QN() );
  DFF_X1 rand_reg_0_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_0[0]), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_1_ ( .D(N25), .CK(clk), .Q(n_zz_io_c_1_11_1_), 
        .QN() );
  DFF_X1 u_zz_io_c_1_11_reg_0_ ( .D(N24), .CK(clk), .Q(n_zz_io_c_1_9_0_), 
        .QN() );
  DFF_X1 u_0_1_reg_4_ ( .D(N8), .CK(clk), .Q(u_0_1[4]), .QN() );
  DFF_X1 u_0_1_reg_3_ ( .D(N6), .CK(clk), .Q(u_0_1[3]), .QN() );
  DFF_X1 u_0_1_reg_2_ ( .D(N4), .CK(clk), .Q(u_0_1[2]), .QN() );
  DFF_X1 u_0_1_reg_1_ ( .D(N2), .CK(clk), .Q(u_0_1[1]), .QN() );
  DFF_X1 u_0_1_reg_0_ ( .D(N0), .CK(clk), .Q(u_0_1[0]), .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_1_ ( .D(N23), .CK(clk), .Q(n_zz_io_c_0_11_1_), 
        .QN() );
  DFF_X1 u_zz_io_c_0_11_reg_0_ ( .D(N22), .CK(clk), .Q(n_zz_io_c_0_9_0_), 
        .QN() );
  DFF_X1 rand_reg_1_reg_4_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_1[4]), 
        .QN() );
  DFF_X1 u_1_0_reg_4_ ( .D(N9), .CK(clk), .Q(u_1_0[4]), .QN() );
  DFF_X1 rand_reg_1_reg_3_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_1[3]), 
        .QN() );
  DFF_X1 u_1_0_reg_3_ ( .D(N7), .CK(clk), .Q(u_1_0[3]), .QN() );
  DFF_X1 rand_reg_1_reg_2_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_1[2]), 
        .QN() );
  DFF_X1 u_1_0_reg_2_ ( .D(N5), .CK(clk), .Q(u_1_0[2]), .QN() );
  DFF_X1 rand_reg_1_reg_1_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_1[1]), 
        .QN() );
  DFF_X1 u_1_0_reg_1_ ( .D(N3), .CK(clk), .Q(u_1_0[1]), .QN() );
  DFF_X1 rand_reg_1_reg_0_ ( .D(io_rand[0]), .CK(clk), .Q(rand_reg_1[0]), 
        .QN() );
  DFF_X1 u_1_0_reg_0_ ( .D(N1), .CK(clk), .Q(u_1_0[0]), .QN() );
  DFF_X1 u_zz_io_c_1_8_reg_1_ ( .D(N21), .CK(clk), .Q(n_zz_io_c_1_8_1_), .QN()
         );
  DFF_X1 u_zz_io_c_1_8_reg_0_ ( .D(N20), .CK(clk), .Q(n_zz_io_c_1_6_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_8_reg_1_ ( .D(N19), .CK(clk), .Q(n_zz_io_c_0_8_1_), .QN()
         );
  DFF_X1 u_zz_io_c_0_8_reg_0_ ( .D(N18), .CK(clk), .Q(n_zz_io_c_0_6_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_5_reg_1_ ( .D(N17), .CK(clk), .Q(n_zz_io_c_1_5_1_), .QN()
         );
  DFF_X1 u_zz_io_c_1_5_reg_0_ ( .D(N16), .CK(clk), .Q(n_zz_io_c_1_3_0_), .QN()
         );
  DFF_X1 u_zz_io_c_0_5_reg_1_ ( .D(N15), .CK(clk), .Q(n_zz_io_c_0_5_1_), .QN()
         );
  DFF_X1 u_zz_io_c_0_5_reg_0_ ( .D(N14), .CK(clk), .Q(n_zz_io_c_0_3_0_), .QN()
         );
  DFF_X1 u_zz_io_c_1_2_reg_1_ ( .D(N13), .CK(clk), .Q(n_zz_io_c_1_2_1_), .QN()
         );
  DFF_X1 u_zz_io_c_1_2_reg_0_ ( .D(N12), .CK(clk), .Q(n_zz_io_c_1_0_), .QN()
         );
  XOR2_X2 U3 ( .A(io_rand[0]), .B(io_b_0[4]), .Z(v_1_1_0[4]) );
  XOR2_X2 U4 ( .A(io_rand[0]), .B(io_b_0[3]), .Z(v_1_1_0[3]) );
  XOR2_X2 U5 ( .A(io_rand[0]), .B(io_b_0[2]), .Z(v_1_1_0[2]) );
  XOR2_X2 U6 ( .A(io_rand[0]), .B(io_b_0[1]), .Z(v_1_1_0[1]) );
  XOR2_X2 U7 ( .A(io_rand[0]), .B(io_b_0[0]), .Z(v_1_1_0[0]) );
  XOR2_X2 U8 ( .A(io_rand[0]), .B(io_b_1[4]), .Z(v_1_0_1[4]) );
  XOR2_X2 U9 ( .A(io_rand[0]), .B(io_b_1[3]), .Z(v_1_0_1[3]) );
  XOR2_X2 U10 ( .A(io_rand[0]), .B(io_b_1[2]), .Z(v_1_0_1[2]) );
  XOR2_X2 U11 ( .A(io_rand[0]), .B(io_b_1[1]), .Z(v_1_0_1[1]) );
  XOR2_X2 U12 ( .A(io_rand[0]), .B(io_b_1[0]), .Z(v_1_0_1[0]) );
  AND2_X1 U53 ( .A1(b_reg_1[0]), .A2(io_a_1[0]), .ZN(N12) );
  AND2_X1 U54 ( .A1(b_reg_0[1]), .A2(io_a_0[1]), .ZN(N14) );
  AND2_X1 U55 ( .A1(b_reg_1[1]), .A2(io_a_1[1]), .ZN(N16) );
  AND2_X1 U56 ( .A1(b_reg_0[2]), .A2(io_a_0[2]), .ZN(N18) );
  AND2_X1 U57 ( .A1(b_reg_1[2]), .A2(io_a_1[2]), .ZN(N20) );
  AND2_X1 U58 ( .A1(b_reg_0[3]), .A2(io_a_0[3]), .ZN(N22) );
  AND2_X1 U59 ( .A1(b_reg_1[3]), .A2(io_a_1[3]), .ZN(N24) );
  AND2_X1 U60 ( .A1(b_reg_0[4]), .A2(io_a_0[4]), .ZN(N26) );
  AND2_X1 U61 ( .A1(b_reg_1[4]), .A2(io_a_1[4]), .ZN(N28) );
  AND2_X1 U62 ( .A1(b_reg_0[0]), .A2(io_a_0[0]), .ZN(N10) );
  AND2_X1 U63 ( .A1(io_a_1[0]), .A2(cor_port_v_1_0[0]), .ZN(N13) );
  AND2_X1 U64 ( .A1(io_a_0[1]), .A2(cor_port_v_0_1[1]), .ZN(N15) );
  AND2_X1 U65 ( .A1(io_a_1[1]), .A2(cor_port_v_1_0[1]), .ZN(N17) );
  AND2_X1 U66 ( .A1(io_a_0[2]), .A2(cor_port_v_0_1[2]), .ZN(N19) );
  AND2_X1 U67 ( .A1(io_a_1[2]), .A2(cor_port_v_1_0[2]), .ZN(N21) );
  AND2_X1 U68 ( .A1(simpleNot_11_port_z), .A2(rand_reg_1[0]), .ZN(N1) );
  AND2_X1 U69 ( .A1(simpleNot_13_port_z), .A2(rand_reg_1[1]), .ZN(N3) );
  AND2_X1 U70 ( .A1(simpleNot_15_port_z), .A2(rand_reg_1[2]), .ZN(N5) );
  AND2_X1 U71 ( .A1(simpleNot_17_port_z), .A2(rand_reg_1[3]), .ZN(N7) );
  AND2_X1 U72 ( .A1(simpleNot_19_port_z), .A2(rand_reg_1[4]), .ZN(N9) );
  AND2_X1 U73 ( .A1(io_a_0[3]), .A2(cor_port_v_0_1[3]), .ZN(N23) );
  AND2_X1 U74 ( .A1(simpleNot_10_port_z), .A2(rand_reg_0[0]), .ZN(N0) );
  AND2_X1 U75 ( .A1(simpleNot_12_port_z), .A2(rand_reg_0[1]), .ZN(N2) );
  AND2_X1 U76 ( .A1(simpleNot_14_port_z), .A2(rand_reg_0[2]), .ZN(N4) );
  AND2_X1 U77 ( .A1(simpleNot_16_port_z), .A2(rand_reg_0[3]), .ZN(N6) );
  AND2_X1 U78 ( .A1(simpleNot_18_port_z), .A2(rand_reg_0[4]), .ZN(N8) );
  AND2_X1 U79 ( .A1(io_a_1[3]), .A2(cor_port_v_1_0[3]), .ZN(N25) );
  AND2_X1 U80 ( .A1(io_a_0[4]), .A2(cor_port_v_0_1[4]), .ZN(N27) );
  AND2_X1 U81 ( .A1(io_a_1[4]), .A2(cor_port_v_1_0[4]), .ZN(N29) );
  AND2_X1 U82 ( .A1(io_a_0[0]), .A2(cor_port_v_0_1[0]), .ZN(N11) );
  XOR2_X1 U83 ( .A(simpleXor_11_port_z), .B(n_zz_io_c_1_0_), .Z(io_c_1[0]) );
  XOR2_X1 U84 ( .A(simpleXor_13_port_z), .B(n_zz_io_c_1_3_0_), .Z(io_c_1[1])
         );
  XOR2_X1 U85 ( .A(simpleXor_15_port_z), .B(n_zz_io_c_1_6_0_), .Z(io_c_1[2])
         );
  XOR2_X1 U86 ( .A(simpleXor_17_port_z), .B(n_zz_io_c_1_9_0_), .Z(io_c_1[3])
         );
  XOR2_X1 U87 ( .A(simpleXor_19_port_z), .B(n_zz_io_c_1_12_0_), .Z(io_c_1[4])
         );
  XOR2_X1 U88 ( .A(simpleXor_10_port_z), .B(n_zz_io_c_0_0_), .Z(io_c_0[0]) );
  XOR2_X1 U89 ( .A(simpleXor_12_port_z), .B(n_zz_io_c_0_3_0_), .Z(io_c_0[1])
         );
  XOR2_X1 U90 ( .A(simpleXor_14_port_z), .B(n_zz_io_c_0_6_0_), .Z(io_c_0[2])
         );
  XOR2_X1 U91 ( .A(simpleXor_16_port_z), .B(n_zz_io_c_0_9_0_), .Z(io_c_0[3])
         );
  XOR2_X1 U92 ( .A(simpleXor_18_port_z), .B(n_zz_io_c_0_12_0_), .Z(io_c_0[4])
         );
  INV_X1 simpleNot_10_U1 ( .A(io_a_0[0]), .ZN(simpleNot_10_port_z) );
  INV_X1 simpleNot_11_U1 ( .A(io_a_1[0]), .ZN(simpleNot_11_port_z) );
  INV_X1 simpleNot_12_U1 ( .A(io_a_0[1]), .ZN(simpleNot_12_port_z) );
  INV_X1 simpleNot_13_U1 ( .A(io_a_1[1]), .ZN(simpleNot_13_port_z) );
  INV_X1 simpleNot_14_U1 ( .A(io_a_0[2]), .ZN(simpleNot_14_port_z) );
  INV_X1 simpleNot_15_U1 ( .A(io_a_1[2]), .ZN(simpleNot_15_port_z) );
  INV_X1 simpleNot_16_U1 ( .A(io_a_0[3]), .ZN(simpleNot_16_port_z) );
  INV_X1 simpleNot_17_U1 ( .A(io_a_1[3]), .ZN(simpleNot_17_port_z) );
  INV_X1 simpleNot_18_U1 ( .A(io_a_0[4]), .ZN(simpleNot_18_port_z) );
  INV_X1 simpleNot_19_U1 ( .A(io_a_1[4]), .ZN(simpleNot_19_port_z) );
  DFF_X1 cor_m_1_0_reg_0_ ( .D(cor_maj_15_port_o), .CK(clk), .Q(
        cor_port_v_1_0[0]), .QN() );
  DFF_X1 cor_m_1_0_reg_1_ ( .D(cor_maj_16_port_o), .CK(clk), .Q(
        cor_port_v_1_0[1]), .QN() );
  DFF_X1 cor_m_1_0_reg_2_ ( .D(cor_maj_17_port_o), .CK(clk), .Q(
        cor_port_v_1_0[2]), .QN() );
  DFF_X1 cor_m_1_0_reg_3_ ( .D(cor_maj_18_port_o), .CK(clk), .Q(
        cor_port_v_1_0[3]), .QN() );
  DFF_X1 cor_m_1_0_reg_4_ ( .D(cor_maj_19_port_o), .CK(clk), .Q(
        cor_port_v_1_0[4]), .QN() );
  DFF_X1 cor_m_0_1_reg_0_ ( .D(cor_maj_10_port_o), .CK(clk), .Q(
        cor_port_v_0_1[0]), .QN() );
  DFF_X1 cor_m_0_1_reg_1_ ( .D(cor_maj_11_port_o), .CK(clk), .Q(
        cor_port_v_0_1[1]), .QN() );
  DFF_X1 cor_m_0_1_reg_2_ ( .D(cor_maj_12_port_o), .CK(clk), .Q(
        cor_port_v_0_1[2]), .QN() );
  DFF_X1 cor_m_0_1_reg_3_ ( .D(cor_maj_13_port_o), .CK(clk), .Q(
        cor_port_v_0_1[3]), .QN() );
  DFF_X1 cor_m_0_1_reg_4_ ( .D(cor_maj_14_port_o), .CK(clk), .Q(
        cor_port_v_0_1[4]), .QN() );
  NAND2_X1 cor_maj_10_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_10_n9) );
  NAND2_X1 cor_maj_10_U14 ( .A1(cor_maj_10_n6), .A2(cor_maj_10_n5), .ZN(
        cor_maj_10_n10) );
  NAND2_X1 cor_maj_10_U13 ( .A1(cor_maj_10_n9), .A2(cor_maj_10_n10), .ZN(
        cor_maj_10_n8) );
  NAND2_X1 cor_maj_10_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_10_n11), .ZN(
        cor_maj_10_n13) );
  NAND2_X1 cor_maj_10_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_10_n12) );
  NAND2_X1 cor_maj_10_U10 ( .A1(cor_maj_10_n12), .A2(cor_maj_10_n13), .ZN(
        cor_maj_10_n7) );
  XOR2_X1 cor_maj_10_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_10_n5) );
  XOR2_X1 cor_maj_10_U8 ( .A(v_1_0_1[2]), .B(cor_maj_10_n11), .Z(cor_maj_10_n6) );
  XOR2_X1 cor_maj_10_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_10_n11)
         );
  OR2_X1 cor_maj_10_U6 ( .A1(cor_maj_10_n7), .A2(cor_maj_10_n8), .ZN(
        cor_maj_10_n3) );
  NAND2_X1 cor_maj_10_U5 ( .A1(cor_maj_10_n3), .A2(cor_maj_10_n4), .ZN(
        cor_maj_10_n2) );
  NAND2_X1 cor_maj_10_U4 ( .A1(cor_maj_10_n7), .A2(cor_maj_10_n8), .ZN(
        cor_maj_10_n1) );
  NAND2_X1 cor_maj_10_U3 ( .A1(cor_maj_10_n1), .A2(cor_maj_10_n2), .ZN(
        cor_maj_10_port_o) );
  XOR2_X1 cor_maj_10_U2 ( .A(cor_maj_10_n5), .B(cor_maj_10_n6), .Z(
        cor_maj_10_n4) );
  NAND2_X1 cor_maj_11_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_11_n18) );
  NAND2_X1 cor_maj_11_U14 ( .A1(cor_maj_11_n21), .A2(cor_maj_11_n22), .ZN(
        cor_maj_11_n17) );
  NAND2_X1 cor_maj_11_U13 ( .A1(cor_maj_11_n18), .A2(cor_maj_11_n17), .ZN(
        cor_maj_11_n19) );
  NAND2_X1 cor_maj_11_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_11_n16), .ZN(
        cor_maj_11_n14) );
  NAND2_X1 cor_maj_11_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_11_n15) );
  NAND2_X1 cor_maj_11_U10 ( .A1(cor_maj_11_n15), .A2(cor_maj_11_n14), .ZN(
        cor_maj_11_n20) );
  XOR2_X1 cor_maj_11_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_11_n22)
         );
  XOR2_X1 cor_maj_11_U8 ( .A(v_1_0_1[2]), .B(cor_maj_11_n16), .Z(
        cor_maj_11_n21) );
  XOR2_X1 cor_maj_11_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_11_n16)
         );
  OR2_X1 cor_maj_11_U6 ( .A1(cor_maj_11_n20), .A2(cor_maj_11_n19), .ZN(
        cor_maj_11_n24) );
  NAND2_X1 cor_maj_11_U5 ( .A1(cor_maj_11_n24), .A2(cor_maj_11_n23), .ZN(
        cor_maj_11_n25) );
  NAND2_X1 cor_maj_11_U4 ( .A1(cor_maj_11_n20), .A2(cor_maj_11_n19), .ZN(
        cor_maj_11_n26) );
  NAND2_X1 cor_maj_11_U3 ( .A1(cor_maj_11_n26), .A2(cor_maj_11_n25), .ZN(
        cor_maj_11_port_o) );
  XOR2_X1 cor_maj_11_U2 ( .A(cor_maj_11_n22), .B(cor_maj_11_n21), .Z(
        cor_maj_11_n23) );
  NAND2_X1 cor_maj_12_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_12_n18) );
  NAND2_X1 cor_maj_12_U14 ( .A1(cor_maj_12_n21), .A2(cor_maj_12_n22), .ZN(
        cor_maj_12_n17) );
  NAND2_X1 cor_maj_12_U13 ( .A1(cor_maj_12_n18), .A2(cor_maj_12_n17), .ZN(
        cor_maj_12_n19) );
  NAND2_X1 cor_maj_12_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_12_n16), .ZN(
        cor_maj_12_n14) );
  NAND2_X1 cor_maj_12_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_12_n15) );
  NAND2_X1 cor_maj_12_U10 ( .A1(cor_maj_12_n15), .A2(cor_maj_12_n14), .ZN(
        cor_maj_12_n20) );
  XOR2_X1 cor_maj_12_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_12_n22)
         );
  XOR2_X1 cor_maj_12_U8 ( .A(v_1_0_1[2]), .B(cor_maj_12_n16), .Z(
        cor_maj_12_n21) );
  XOR2_X1 cor_maj_12_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_12_n16)
         );
  OR2_X1 cor_maj_12_U6 ( .A1(cor_maj_12_n20), .A2(cor_maj_12_n19), .ZN(
        cor_maj_12_n24) );
  NAND2_X1 cor_maj_12_U5 ( .A1(cor_maj_12_n24), .A2(cor_maj_12_n23), .ZN(
        cor_maj_12_n25) );
  NAND2_X1 cor_maj_12_U4 ( .A1(cor_maj_12_n20), .A2(cor_maj_12_n19), .ZN(
        cor_maj_12_n26) );
  NAND2_X1 cor_maj_12_U3 ( .A1(cor_maj_12_n26), .A2(cor_maj_12_n25), .ZN(
        cor_maj_12_port_o) );
  XOR2_X1 cor_maj_12_U2 ( .A(cor_maj_12_n22), .B(cor_maj_12_n21), .Z(
        cor_maj_12_n23) );
  NAND2_X1 cor_maj_13_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_13_n18) );
  NAND2_X1 cor_maj_13_U14 ( .A1(cor_maj_13_n21), .A2(cor_maj_13_n22), .ZN(
        cor_maj_13_n17) );
  NAND2_X1 cor_maj_13_U13 ( .A1(cor_maj_13_n18), .A2(cor_maj_13_n17), .ZN(
        cor_maj_13_n19) );
  NAND2_X1 cor_maj_13_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_13_n16), .ZN(
        cor_maj_13_n14) );
  NAND2_X1 cor_maj_13_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_13_n15) );
  NAND2_X1 cor_maj_13_U10 ( .A1(cor_maj_13_n15), .A2(cor_maj_13_n14), .ZN(
        cor_maj_13_n20) );
  XOR2_X1 cor_maj_13_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_13_n22)
         );
  XOR2_X1 cor_maj_13_U8 ( .A(v_1_0_1[2]), .B(cor_maj_13_n16), .Z(
        cor_maj_13_n21) );
  XOR2_X1 cor_maj_13_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_13_n16)
         );
  OR2_X1 cor_maj_13_U6 ( .A1(cor_maj_13_n20), .A2(cor_maj_13_n19), .ZN(
        cor_maj_13_n24) );
  NAND2_X1 cor_maj_13_U5 ( .A1(cor_maj_13_n24), .A2(cor_maj_13_n23), .ZN(
        cor_maj_13_n25) );
  NAND2_X1 cor_maj_13_U4 ( .A1(cor_maj_13_n20), .A2(cor_maj_13_n19), .ZN(
        cor_maj_13_n26) );
  NAND2_X1 cor_maj_13_U3 ( .A1(cor_maj_13_n26), .A2(cor_maj_13_n25), .ZN(
        cor_maj_13_port_o) );
  XOR2_X1 cor_maj_13_U2 ( .A(cor_maj_13_n22), .B(cor_maj_13_n21), .Z(
        cor_maj_13_n23) );
  NAND2_X1 cor_maj_14_U15 ( .A1(v_1_0_1[3]), .A2(v_1_0_1[4]), .ZN(
        cor_maj_14_n18) );
  NAND2_X1 cor_maj_14_U14 ( .A1(cor_maj_14_n21), .A2(cor_maj_14_n22), .ZN(
        cor_maj_14_n17) );
  NAND2_X1 cor_maj_14_U13 ( .A1(cor_maj_14_n18), .A2(cor_maj_14_n17), .ZN(
        cor_maj_14_n19) );
  NAND2_X1 cor_maj_14_U12 ( .A1(v_1_0_1[2]), .A2(cor_maj_14_n16), .ZN(
        cor_maj_14_n14) );
  NAND2_X1 cor_maj_14_U11 ( .A1(v_1_0_1[0]), .A2(v_1_0_1[1]), .ZN(
        cor_maj_14_n15) );
  NAND2_X1 cor_maj_14_U10 ( .A1(cor_maj_14_n15), .A2(cor_maj_14_n14), .ZN(
        cor_maj_14_n20) );
  XOR2_X1 cor_maj_14_U9 ( .A(v_1_0_1[3]), .B(v_1_0_1[4]), .Z(cor_maj_14_n22)
         );
  XOR2_X1 cor_maj_14_U8 ( .A(v_1_0_1[2]), .B(cor_maj_14_n16), .Z(
        cor_maj_14_n21) );
  XOR2_X1 cor_maj_14_U7 ( .A(v_1_0_1[0]), .B(v_1_0_1[1]), .Z(cor_maj_14_n16)
         );
  OR2_X1 cor_maj_14_U6 ( .A1(cor_maj_14_n20), .A2(cor_maj_14_n19), .ZN(
        cor_maj_14_n24) );
  NAND2_X1 cor_maj_14_U5 ( .A1(cor_maj_14_n24), .A2(cor_maj_14_n23), .ZN(
        cor_maj_14_n25) );
  NAND2_X1 cor_maj_14_U4 ( .A1(cor_maj_14_n20), .A2(cor_maj_14_n19), .ZN(
        cor_maj_14_n26) );
  NAND2_X1 cor_maj_14_U3 ( .A1(cor_maj_14_n26), .A2(cor_maj_14_n25), .ZN(
        cor_maj_14_port_o) );
  XOR2_X1 cor_maj_14_U2 ( .A(cor_maj_14_n22), .B(cor_maj_14_n21), .Z(
        cor_maj_14_n23) );
  NAND2_X1 cor_maj_15_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_15_n18) );
  NAND2_X1 cor_maj_15_U14 ( .A1(cor_maj_15_n21), .A2(cor_maj_15_n22), .ZN(
        cor_maj_15_n17) );
  NAND2_X1 cor_maj_15_U13 ( .A1(cor_maj_15_n18), .A2(cor_maj_15_n17), .ZN(
        cor_maj_15_n19) );
  NAND2_X1 cor_maj_15_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_15_n16), .ZN(
        cor_maj_15_n14) );
  NAND2_X1 cor_maj_15_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_15_n15) );
  NAND2_X1 cor_maj_15_U10 ( .A1(cor_maj_15_n15), .A2(cor_maj_15_n14), .ZN(
        cor_maj_15_n20) );
  XOR2_X1 cor_maj_15_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_15_n22)
         );
  XOR2_X1 cor_maj_15_U8 ( .A(v_1_1_0[2]), .B(cor_maj_15_n16), .Z(
        cor_maj_15_n21) );
  XOR2_X1 cor_maj_15_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_15_n16)
         );
  OR2_X1 cor_maj_15_U6 ( .A1(cor_maj_15_n20), .A2(cor_maj_15_n19), .ZN(
        cor_maj_15_n24) );
  NAND2_X1 cor_maj_15_U5 ( .A1(cor_maj_15_n24), .A2(cor_maj_15_n23), .ZN(
        cor_maj_15_n25) );
  NAND2_X1 cor_maj_15_U4 ( .A1(cor_maj_15_n20), .A2(cor_maj_15_n19), .ZN(
        cor_maj_15_n26) );
  NAND2_X1 cor_maj_15_U3 ( .A1(cor_maj_15_n26), .A2(cor_maj_15_n25), .ZN(
        cor_maj_15_port_o) );
  XOR2_X1 cor_maj_15_U2 ( .A(cor_maj_15_n22), .B(cor_maj_15_n21), .Z(
        cor_maj_15_n23) );
  NAND2_X1 cor_maj_16_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_16_n18) );
  NAND2_X1 cor_maj_16_U14 ( .A1(cor_maj_16_n21), .A2(cor_maj_16_n22), .ZN(
        cor_maj_16_n17) );
  NAND2_X1 cor_maj_16_U13 ( .A1(cor_maj_16_n18), .A2(cor_maj_16_n17), .ZN(
        cor_maj_16_n19) );
  NAND2_X1 cor_maj_16_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_16_n16), .ZN(
        cor_maj_16_n14) );
  NAND2_X1 cor_maj_16_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_16_n15) );
  NAND2_X1 cor_maj_16_U10 ( .A1(cor_maj_16_n15), .A2(cor_maj_16_n14), .ZN(
        cor_maj_16_n20) );
  XOR2_X1 cor_maj_16_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_16_n22)
         );
  XOR2_X1 cor_maj_16_U8 ( .A(v_1_1_0[2]), .B(cor_maj_16_n16), .Z(
        cor_maj_16_n21) );
  XOR2_X1 cor_maj_16_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_16_n16)
         );
  OR2_X1 cor_maj_16_U6 ( .A1(cor_maj_16_n20), .A2(cor_maj_16_n19), .ZN(
        cor_maj_16_n24) );
  NAND2_X1 cor_maj_16_U5 ( .A1(cor_maj_16_n24), .A2(cor_maj_16_n23), .ZN(
        cor_maj_16_n25) );
  NAND2_X1 cor_maj_16_U4 ( .A1(cor_maj_16_n20), .A2(cor_maj_16_n19), .ZN(
        cor_maj_16_n26) );
  NAND2_X1 cor_maj_16_U3 ( .A1(cor_maj_16_n26), .A2(cor_maj_16_n25), .ZN(
        cor_maj_16_port_o) );
  XOR2_X1 cor_maj_16_U2 ( .A(cor_maj_16_n22), .B(cor_maj_16_n21), .Z(
        cor_maj_16_n23) );
  NAND2_X1 cor_maj_17_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_17_n18) );
  NAND2_X1 cor_maj_17_U14 ( .A1(cor_maj_17_n21), .A2(cor_maj_17_n22), .ZN(
        cor_maj_17_n17) );
  NAND2_X1 cor_maj_17_U13 ( .A1(cor_maj_17_n18), .A2(cor_maj_17_n17), .ZN(
        cor_maj_17_n19) );
  NAND2_X1 cor_maj_17_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_17_n16), .ZN(
        cor_maj_17_n14) );
  NAND2_X1 cor_maj_17_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_17_n15) );
  NAND2_X1 cor_maj_17_U10 ( .A1(cor_maj_17_n15), .A2(cor_maj_17_n14), .ZN(
        cor_maj_17_n20) );
  XOR2_X1 cor_maj_17_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_17_n22)
         );
  XOR2_X1 cor_maj_17_U8 ( .A(v_1_1_0[2]), .B(cor_maj_17_n16), .Z(
        cor_maj_17_n21) );
  XOR2_X1 cor_maj_17_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_17_n16)
         );
  OR2_X1 cor_maj_17_U6 ( .A1(cor_maj_17_n20), .A2(cor_maj_17_n19), .ZN(
        cor_maj_17_n24) );
  NAND2_X1 cor_maj_17_U5 ( .A1(cor_maj_17_n24), .A2(cor_maj_17_n23), .ZN(
        cor_maj_17_n25) );
  NAND2_X1 cor_maj_17_U4 ( .A1(cor_maj_17_n20), .A2(cor_maj_17_n19), .ZN(
        cor_maj_17_n26) );
  NAND2_X1 cor_maj_17_U3 ( .A1(cor_maj_17_n26), .A2(cor_maj_17_n25), .ZN(
        cor_maj_17_port_o) );
  XOR2_X1 cor_maj_17_U2 ( .A(cor_maj_17_n22), .B(cor_maj_17_n21), .Z(
        cor_maj_17_n23) );
  NAND2_X1 cor_maj_18_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_18_n18) );
  NAND2_X1 cor_maj_18_U14 ( .A1(cor_maj_18_n21), .A2(cor_maj_18_n22), .ZN(
        cor_maj_18_n17) );
  NAND2_X1 cor_maj_18_U13 ( .A1(cor_maj_18_n18), .A2(cor_maj_18_n17), .ZN(
        cor_maj_18_n19) );
  NAND2_X1 cor_maj_18_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_18_n16), .ZN(
        cor_maj_18_n14) );
  NAND2_X1 cor_maj_18_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_18_n15) );
  NAND2_X1 cor_maj_18_U10 ( .A1(cor_maj_18_n15), .A2(cor_maj_18_n14), .ZN(
        cor_maj_18_n20) );
  XOR2_X1 cor_maj_18_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_18_n22)
         );
  XOR2_X1 cor_maj_18_U8 ( .A(v_1_1_0[2]), .B(cor_maj_18_n16), .Z(
        cor_maj_18_n21) );
  XOR2_X1 cor_maj_18_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_18_n16)
         );
  OR2_X1 cor_maj_18_U6 ( .A1(cor_maj_18_n20), .A2(cor_maj_18_n19), .ZN(
        cor_maj_18_n24) );
  NAND2_X1 cor_maj_18_U5 ( .A1(cor_maj_18_n24), .A2(cor_maj_18_n23), .ZN(
        cor_maj_18_n25) );
  NAND2_X1 cor_maj_18_U4 ( .A1(cor_maj_18_n20), .A2(cor_maj_18_n19), .ZN(
        cor_maj_18_n26) );
  NAND2_X1 cor_maj_18_U3 ( .A1(cor_maj_18_n26), .A2(cor_maj_18_n25), .ZN(
        cor_maj_18_port_o) );
  XOR2_X1 cor_maj_18_U2 ( .A(cor_maj_18_n22), .B(cor_maj_18_n21), .Z(
        cor_maj_18_n23) );
  NAND2_X1 cor_maj_19_U15 ( .A1(v_1_1_0[3]), .A2(v_1_1_0[4]), .ZN(
        cor_maj_19_n18) );
  NAND2_X1 cor_maj_19_U14 ( .A1(cor_maj_19_n21), .A2(cor_maj_19_n22), .ZN(
        cor_maj_19_n17) );
  NAND2_X1 cor_maj_19_U13 ( .A1(cor_maj_19_n18), .A2(cor_maj_19_n17), .ZN(
        cor_maj_19_n19) );
  NAND2_X1 cor_maj_19_U12 ( .A1(v_1_1_0[2]), .A2(cor_maj_19_n16), .ZN(
        cor_maj_19_n14) );
  NAND2_X1 cor_maj_19_U11 ( .A1(v_1_1_0[0]), .A2(v_1_1_0[1]), .ZN(
        cor_maj_19_n15) );
  NAND2_X1 cor_maj_19_U10 ( .A1(cor_maj_19_n15), .A2(cor_maj_19_n14), .ZN(
        cor_maj_19_n20) );
  XOR2_X1 cor_maj_19_U9 ( .A(v_1_1_0[3]), .B(v_1_1_0[4]), .Z(cor_maj_19_n22)
         );
  XOR2_X1 cor_maj_19_U8 ( .A(v_1_1_0[2]), .B(cor_maj_19_n16), .Z(
        cor_maj_19_n21) );
  XOR2_X1 cor_maj_19_U7 ( .A(v_1_1_0[0]), .B(v_1_1_0[1]), .Z(cor_maj_19_n16)
         );
  OR2_X1 cor_maj_19_U6 ( .A1(cor_maj_19_n20), .A2(cor_maj_19_n19), .ZN(
        cor_maj_19_n24) );
  NAND2_X1 cor_maj_19_U5 ( .A1(cor_maj_19_n24), .A2(cor_maj_19_n23), .ZN(
        cor_maj_19_n25) );
  NAND2_X1 cor_maj_19_U4 ( .A1(cor_maj_19_n20), .A2(cor_maj_19_n19), .ZN(
        cor_maj_19_n26) );
  NAND2_X1 cor_maj_19_U3 ( .A1(cor_maj_19_n26), .A2(cor_maj_19_n25), .ZN(
        cor_maj_19_port_o) );
  XOR2_X1 cor_maj_19_U2 ( .A(cor_maj_19_n22), .B(cor_maj_19_n21), .Z(
        cor_maj_19_n23) );
  XOR2_X1 simpleXor_10_U1 ( .A(n_zz_io_c_0_2_1_), .B(u_0_1[0]), .Z(
        simpleXor_10_port_z) );
  XOR2_X1 simpleXor_11_U1 ( .A(n_zz_io_c_1_2_1_), .B(u_1_0[0]), .Z(
        simpleXor_11_port_z) );
  XOR2_X1 simpleXor_12_U1 ( .A(n_zz_io_c_0_5_1_), .B(u_0_1[1]), .Z(
        simpleXor_12_port_z) );
  XOR2_X1 simpleXor_13_U1 ( .A(n_zz_io_c_1_5_1_), .B(u_1_0[1]), .Z(
        simpleXor_13_port_z) );
  XOR2_X1 simpleXor_14_U1 ( .A(n_zz_io_c_0_8_1_), .B(u_0_1[2]), .Z(
        simpleXor_14_port_z) );
  XOR2_X1 simpleXor_15_U1 ( .A(n_zz_io_c_1_8_1_), .B(u_1_0[2]), .Z(
        simpleXor_15_port_z) );
  XOR2_X1 simpleXor_16_U1 ( .A(n_zz_io_c_0_11_1_), .B(u_0_1[3]), .Z(
        simpleXor_16_port_z) );
  XOR2_X1 simpleXor_17_U1 ( .A(n_zz_io_c_1_11_1_), .B(u_1_0[3]), .Z(
        simpleXor_17_port_z) );
  XOR2_X1 simpleXor_18_U1 ( .A(n_zz_io_c_0_14_1_), .B(u_0_1[4]), .Z(
        simpleXor_18_port_z) );
  XOR2_X1 simpleXor_19_U1 ( .A(n_zz_io_c_1_14_1_), .B(u_1_0[4]), .Z(
        simpleXor_19_port_z) );
endmodule

