
module AesSbox_keyAdd_correction ( clock, reset, io_state, io_key, io_out );
  input [7:0] io_state;
  input [7:0] io_key;
  output [7:0] io_out;
  input clock, reset;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         AesSbox_keyAdd_sbox_io_o7, AesSbox_keyAdd_sbox_io_o6,
         AesSbox_keyAdd_sbox_io_o5, AesSbox_keyAdd_sbox_io_o4,
         AesSbox_keyAdd_sbox_io_o3, AesSbox_keyAdd_sbox_io_o2,
         AesSbox_keyAdd_sbox_io_o1, AesSbox_keyAdd_sbox_io_o0,
         AesSbox_keyAdd_sbox_n128, AesSbox_keyAdd_sbox_n127,
         AesSbox_keyAdd_sbox_n126, AesSbox_keyAdd_sbox_n125,
         AesSbox_keyAdd_sbox_n124, AesSbox_keyAdd_sbox_n123,
         AesSbox_keyAdd_sbox_n122, AesSbox_keyAdd_sbox_n121,
         AesSbox_keyAdd_sbox_n120, AesSbox_keyAdd_sbox_n119,
         AesSbox_keyAdd_sbox_n118, AesSbox_keyAdd_sbox_n117,
         AesSbox_keyAdd_sbox_n116, AesSbox_keyAdd_sbox_n115,
         AesSbox_keyAdd_sbox_n114, AesSbox_keyAdd_sbox_n113,
         AesSbox_keyAdd_sbox_n112, AesSbox_keyAdd_sbox_n111,
         AesSbox_keyAdd_sbox_n110, AesSbox_keyAdd_sbox_n109,
         AesSbox_keyAdd_sbox_n108, AesSbox_keyAdd_sbox_n107,
         AesSbox_keyAdd_sbox_n106, AesSbox_keyAdd_sbox_n105,
         AesSbox_keyAdd_sbox_n104, AesSbox_keyAdd_sbox_n103,
         AesSbox_keyAdd_sbox_n102, AesSbox_keyAdd_sbox_n101,
         AesSbox_keyAdd_sbox_n100, AesSbox_keyAdd_sbox_n99,
         AesSbox_keyAdd_sbox_n98, AesSbox_keyAdd_sbox_n97,
         AesSbox_keyAdd_sbox_n96, AesSbox_keyAdd_sbox_n95,
         AesSbox_keyAdd_sbox_n94, AesSbox_keyAdd_sbox_n93,
         AesSbox_keyAdd_sbox_n92, AesSbox_keyAdd_sbox_n91,
         AesSbox_keyAdd_sbox_n90, AesSbox_keyAdd_sbox_n89,
         AesSbox_keyAdd_sbox_n88, AesSbox_keyAdd_sbox_n87,
         AesSbox_keyAdd_sbox_n86, AesSbox_keyAdd_sbox_n85,
         AesSbox_keyAdd_sbox_n84, AesSbox_keyAdd_sbox_n83,
         AesSbox_keyAdd_sbox_n82, AesSbox_keyAdd_sbox_n81,
         AesSbox_keyAdd_sbox_n80, AesSbox_keyAdd_sbox_n79,
         AesSbox_keyAdd_sbox_n78, AesSbox_keyAdd_sbox_n77,
         AesSbox_keyAdd_sbox_n76, AesSbox_keyAdd_sbox_n75,
         AesSbox_keyAdd_sbox_n74, AesSbox_keyAdd_sbox_n73,
         AesSbox_keyAdd_sbox_n72, AesSbox_keyAdd_sbox_n71,
         AesSbox_keyAdd_sbox_n70, AesSbox_keyAdd_sbox_n69,
         AesSbox_keyAdd_sbox_n68, AesSbox_keyAdd_sbox_n67,
         AesSbox_keyAdd_sbox_n66, AesSbox_keyAdd_sbox_n65,
         AesSbox_keyAdd_sbox_n64, AesSbox_keyAdd_sbox_n63,
         AesSbox_keyAdd_sbox_n62, AesSbox_keyAdd_sbox_n61,
         AesSbox_keyAdd_sbox_n60, AesSbox_keyAdd_sbox_n59,
         AesSbox_keyAdd_sbox_n58, AesSbox_keyAdd_sbox_n57,
         AesSbox_keyAdd_sbox_n56, AesSbox_keyAdd_sbox_n55,
         AesSbox_keyAdd_sbox_n54, AesSbox_keyAdd_sbox_n53,
         AesSbox_keyAdd_sbox_n52, AesSbox_keyAdd_sbox_n51,
         AesSbox_keyAdd_sbox_n50, AesSbox_keyAdd_sbox_n49,
         AesSbox_keyAdd_sbox_n48, AesSbox_keyAdd_sbox_n47,
         AesSbox_keyAdd_sbox_n46, AesSbox_keyAdd_sbox_n45,
         AesSbox_keyAdd_sbox_n44, AesSbox_keyAdd_sbox_n43,
         AesSbox_keyAdd_sbox_n42, AesSbox_keyAdd_sbox_n41,
         AesSbox_keyAdd_sbox_n40, AesSbox_keyAdd_sbox_n39,
         AesSbox_keyAdd_sbox_n38, AesSbox_keyAdd_sbox_n37,
         AesSbox_keyAdd_sbox_n36, AesSbox_keyAdd_sbox_n35,
         AesSbox_keyAdd_sbox_n34, AesSbox_keyAdd_sbox_n33,
         AesSbox_keyAdd_sbox_n32, AesSbox_keyAdd_sbox_n31,
         AesSbox_keyAdd_sbox_n30, AesSbox_keyAdd_sbox_n29,
         AesSbox_keyAdd_sbox_n28, AesSbox_keyAdd_sbox_n27,
         AesSbox_keyAdd_sbox_n26, AesSbox_keyAdd_sbox_n25,
         AesSbox_keyAdd_sbox_n24, AesSbox_keyAdd_sbox_n23,
         AesSbox_keyAdd_sbox_n22, AesSbox_keyAdd_sbox_n21,
         AesSbox_keyAdd_sbox_n20, AesSbox_keyAdd_sbox_n19,
         AesSbox_keyAdd_sbox_n18, AesSbox_keyAdd_sbox_n17,
         AesSbox_keyAdd_sbox_n16, AesSbox_keyAdd_sbox_n15,
         AesSbox_keyAdd_sbox_n14, AesSbox_keyAdd_sbox_n13,
         AesSbox_keyAdd_sbox_n12, AesSbox_keyAdd_sbox_n11,
         AesSbox_keyAdd_sbox_n10, AesSbox_keyAdd_sbox_n9,
         AesSbox_keyAdd_sbox_n8, AesSbox_keyAdd_sbox_n7,
         AesSbox_keyAdd_sbox_n6, AesSbox_keyAdd_sbox_n5,
         AesSbox_keyAdd_sbox_n4, AesSbox_keyAdd_sbox_n3,
         AesSbox_keyAdd_sbox_n2, AesSbox_keyAdd_sbox_n1,
         AesSbox_keyAdd_1_sbox_io_o7, AesSbox_keyAdd_1_sbox_io_o6,
         AesSbox_keyAdd_1_sbox_io_o5, AesSbox_keyAdd_1_sbox_io_o4,
         AesSbox_keyAdd_1_sbox_io_o3, AesSbox_keyAdd_1_sbox_io_o2,
         AesSbox_keyAdd_1_sbox_io_o1, AesSbox_keyAdd_1_sbox_io_o0,
         AesSbox_keyAdd_1_sbox_n128, AesSbox_keyAdd_1_sbox_n127,
         AesSbox_keyAdd_1_sbox_n126, AesSbox_keyAdd_1_sbox_n125,
         AesSbox_keyAdd_1_sbox_n124, AesSbox_keyAdd_1_sbox_n123,
         AesSbox_keyAdd_1_sbox_n122, AesSbox_keyAdd_1_sbox_n121,
         AesSbox_keyAdd_1_sbox_n120, AesSbox_keyAdd_1_sbox_n119,
         AesSbox_keyAdd_1_sbox_n118, AesSbox_keyAdd_1_sbox_n117,
         AesSbox_keyAdd_1_sbox_n116, AesSbox_keyAdd_1_sbox_n115,
         AesSbox_keyAdd_1_sbox_n114, AesSbox_keyAdd_1_sbox_n113,
         AesSbox_keyAdd_1_sbox_n112, AesSbox_keyAdd_1_sbox_n111,
         AesSbox_keyAdd_1_sbox_n110, AesSbox_keyAdd_1_sbox_n109,
         AesSbox_keyAdd_1_sbox_n108, AesSbox_keyAdd_1_sbox_n107,
         AesSbox_keyAdd_1_sbox_n106, AesSbox_keyAdd_1_sbox_n105,
         AesSbox_keyAdd_1_sbox_n104, AesSbox_keyAdd_1_sbox_n103,
         AesSbox_keyAdd_1_sbox_n102, AesSbox_keyAdd_1_sbox_n101,
         AesSbox_keyAdd_1_sbox_n100, AesSbox_keyAdd_1_sbox_n99,
         AesSbox_keyAdd_1_sbox_n98, AesSbox_keyAdd_1_sbox_n97,
         AesSbox_keyAdd_1_sbox_n96, AesSbox_keyAdd_1_sbox_n95,
         AesSbox_keyAdd_1_sbox_n94, AesSbox_keyAdd_1_sbox_n93,
         AesSbox_keyAdd_1_sbox_n92, AesSbox_keyAdd_1_sbox_n91,
         AesSbox_keyAdd_1_sbox_n90, AesSbox_keyAdd_1_sbox_n89,
         AesSbox_keyAdd_1_sbox_n88, AesSbox_keyAdd_1_sbox_n87,
         AesSbox_keyAdd_1_sbox_n86, AesSbox_keyAdd_1_sbox_n85,
         AesSbox_keyAdd_1_sbox_n84, AesSbox_keyAdd_1_sbox_n83,
         AesSbox_keyAdd_1_sbox_n82, AesSbox_keyAdd_1_sbox_n81,
         AesSbox_keyAdd_1_sbox_n80, AesSbox_keyAdd_1_sbox_n79,
         AesSbox_keyAdd_1_sbox_n78, AesSbox_keyAdd_1_sbox_n77,
         AesSbox_keyAdd_1_sbox_n76, AesSbox_keyAdd_1_sbox_n75,
         AesSbox_keyAdd_1_sbox_n74, AesSbox_keyAdd_1_sbox_n73,
         AesSbox_keyAdd_1_sbox_n72, AesSbox_keyAdd_1_sbox_n71,
         AesSbox_keyAdd_1_sbox_n70, AesSbox_keyAdd_1_sbox_n69,
         AesSbox_keyAdd_1_sbox_n68, AesSbox_keyAdd_1_sbox_n67,
         AesSbox_keyAdd_1_sbox_n66, AesSbox_keyAdd_1_sbox_n65,
         AesSbox_keyAdd_1_sbox_n64, AesSbox_keyAdd_1_sbox_n63,
         AesSbox_keyAdd_1_sbox_n62, AesSbox_keyAdd_1_sbox_n61,
         AesSbox_keyAdd_1_sbox_n60, AesSbox_keyAdd_1_sbox_n59,
         AesSbox_keyAdd_1_sbox_n58, AesSbox_keyAdd_1_sbox_n57,
         AesSbox_keyAdd_1_sbox_n56, AesSbox_keyAdd_1_sbox_n55,
         AesSbox_keyAdd_1_sbox_n54, AesSbox_keyAdd_1_sbox_n53,
         AesSbox_keyAdd_1_sbox_n52, AesSbox_keyAdd_1_sbox_n51,
         AesSbox_keyAdd_1_sbox_n50, AesSbox_keyAdd_1_sbox_n49,
         AesSbox_keyAdd_1_sbox_n48, AesSbox_keyAdd_1_sbox_n47,
         AesSbox_keyAdd_1_sbox_n46, AesSbox_keyAdd_1_sbox_n45,
         AesSbox_keyAdd_1_sbox_n44, AesSbox_keyAdd_1_sbox_n43,
         AesSbox_keyAdd_1_sbox_n42, AesSbox_keyAdd_1_sbox_n41,
         AesSbox_keyAdd_1_sbox_n40, AesSbox_keyAdd_1_sbox_n39,
         AesSbox_keyAdd_1_sbox_n38, AesSbox_keyAdd_1_sbox_n37,
         AesSbox_keyAdd_1_sbox_n36, AesSbox_keyAdd_1_sbox_n35,
         AesSbox_keyAdd_1_sbox_n34, AesSbox_keyAdd_1_sbox_n33,
         AesSbox_keyAdd_1_sbox_n32, AesSbox_keyAdd_1_sbox_n31,
         AesSbox_keyAdd_1_sbox_n30, AesSbox_keyAdd_1_sbox_n29,
         AesSbox_keyAdd_1_sbox_n28, AesSbox_keyAdd_1_sbox_n27,
         AesSbox_keyAdd_1_sbox_n26, AesSbox_keyAdd_1_sbox_n25,
         AesSbox_keyAdd_1_sbox_n24, AesSbox_keyAdd_1_sbox_n23,
         AesSbox_keyAdd_1_sbox_n22, AesSbox_keyAdd_1_sbox_n21,
         AesSbox_keyAdd_1_sbox_n20, AesSbox_keyAdd_1_sbox_n19,
         AesSbox_keyAdd_1_sbox_n18, AesSbox_keyAdd_1_sbox_n17,
         AesSbox_keyAdd_1_sbox_n16, AesSbox_keyAdd_1_sbox_n15,
         AesSbox_keyAdd_1_sbox_n14, AesSbox_keyAdd_1_sbox_n13,
         AesSbox_keyAdd_1_sbox_n12, AesSbox_keyAdd_1_sbox_n11,
         AesSbox_keyAdd_1_sbox_n10, AesSbox_keyAdd_1_sbox_n9,
         AesSbox_keyAdd_1_sbox_n8, AesSbox_keyAdd_1_sbox_n7,
         AesSbox_keyAdd_1_sbox_n6, AesSbox_keyAdd_1_sbox_n5,
         AesSbox_keyAdd_1_sbox_n4, AesSbox_keyAdd_1_sbox_n3,
         AesSbox_keyAdd_1_sbox_n2, AesSbox_keyAdd_1_sbox_n1,
         AesSbox_keyAdd_2_sbox_io_o7, AesSbox_keyAdd_2_sbox_io_o6,
         AesSbox_keyAdd_2_sbox_io_o5, AesSbox_keyAdd_2_sbox_io_o4,
         AesSbox_keyAdd_2_sbox_io_o3, AesSbox_keyAdd_2_sbox_io_o2,
         AesSbox_keyAdd_2_sbox_io_o1, AesSbox_keyAdd_2_sbox_io_o0,
         AesSbox_keyAdd_2_sbox_n128, AesSbox_keyAdd_2_sbox_n127,
         AesSbox_keyAdd_2_sbox_n126, AesSbox_keyAdd_2_sbox_n125,
         AesSbox_keyAdd_2_sbox_n124, AesSbox_keyAdd_2_sbox_n123,
         AesSbox_keyAdd_2_sbox_n122, AesSbox_keyAdd_2_sbox_n121,
         AesSbox_keyAdd_2_sbox_n120, AesSbox_keyAdd_2_sbox_n119,
         AesSbox_keyAdd_2_sbox_n118, AesSbox_keyAdd_2_sbox_n117,
         AesSbox_keyAdd_2_sbox_n116, AesSbox_keyAdd_2_sbox_n115,
         AesSbox_keyAdd_2_sbox_n114, AesSbox_keyAdd_2_sbox_n113,
         AesSbox_keyAdd_2_sbox_n112, AesSbox_keyAdd_2_sbox_n111,
         AesSbox_keyAdd_2_sbox_n110, AesSbox_keyAdd_2_sbox_n109,
         AesSbox_keyAdd_2_sbox_n108, AesSbox_keyAdd_2_sbox_n107,
         AesSbox_keyAdd_2_sbox_n106, AesSbox_keyAdd_2_sbox_n105,
         AesSbox_keyAdd_2_sbox_n104, AesSbox_keyAdd_2_sbox_n103,
         AesSbox_keyAdd_2_sbox_n102, AesSbox_keyAdd_2_sbox_n101,
         AesSbox_keyAdd_2_sbox_n100, AesSbox_keyAdd_2_sbox_n99,
         AesSbox_keyAdd_2_sbox_n98, AesSbox_keyAdd_2_sbox_n97,
         AesSbox_keyAdd_2_sbox_n96, AesSbox_keyAdd_2_sbox_n95,
         AesSbox_keyAdd_2_sbox_n94, AesSbox_keyAdd_2_sbox_n93,
         AesSbox_keyAdd_2_sbox_n92, AesSbox_keyAdd_2_sbox_n91,
         AesSbox_keyAdd_2_sbox_n90, AesSbox_keyAdd_2_sbox_n89,
         AesSbox_keyAdd_2_sbox_n88, AesSbox_keyAdd_2_sbox_n87,
         AesSbox_keyAdd_2_sbox_n86, AesSbox_keyAdd_2_sbox_n85,
         AesSbox_keyAdd_2_sbox_n84, AesSbox_keyAdd_2_sbox_n83,
         AesSbox_keyAdd_2_sbox_n82, AesSbox_keyAdd_2_sbox_n81,
         AesSbox_keyAdd_2_sbox_n80, AesSbox_keyAdd_2_sbox_n79,
         AesSbox_keyAdd_2_sbox_n78, AesSbox_keyAdd_2_sbox_n77,
         AesSbox_keyAdd_2_sbox_n76, AesSbox_keyAdd_2_sbox_n75,
         AesSbox_keyAdd_2_sbox_n74, AesSbox_keyAdd_2_sbox_n73,
         AesSbox_keyAdd_2_sbox_n72, AesSbox_keyAdd_2_sbox_n71,
         AesSbox_keyAdd_2_sbox_n70, AesSbox_keyAdd_2_sbox_n69,
         AesSbox_keyAdd_2_sbox_n68, AesSbox_keyAdd_2_sbox_n67,
         AesSbox_keyAdd_2_sbox_n66, AesSbox_keyAdd_2_sbox_n65,
         AesSbox_keyAdd_2_sbox_n64, AesSbox_keyAdd_2_sbox_n63,
         AesSbox_keyAdd_2_sbox_n62, AesSbox_keyAdd_2_sbox_n61,
         AesSbox_keyAdd_2_sbox_n60, AesSbox_keyAdd_2_sbox_n59,
         AesSbox_keyAdd_2_sbox_n58, AesSbox_keyAdd_2_sbox_n57,
         AesSbox_keyAdd_2_sbox_n56, AesSbox_keyAdd_2_sbox_n55,
         AesSbox_keyAdd_2_sbox_n54, AesSbox_keyAdd_2_sbox_n53,
         AesSbox_keyAdd_2_sbox_n52, AesSbox_keyAdd_2_sbox_n51,
         AesSbox_keyAdd_2_sbox_n50, AesSbox_keyAdd_2_sbox_n49,
         AesSbox_keyAdd_2_sbox_n48, AesSbox_keyAdd_2_sbox_n47,
         AesSbox_keyAdd_2_sbox_n46, AesSbox_keyAdd_2_sbox_n45,
         AesSbox_keyAdd_2_sbox_n44, AesSbox_keyAdd_2_sbox_n43,
         AesSbox_keyAdd_2_sbox_n42, AesSbox_keyAdd_2_sbox_n41,
         AesSbox_keyAdd_2_sbox_n40, AesSbox_keyAdd_2_sbox_n39,
         AesSbox_keyAdd_2_sbox_n38, AesSbox_keyAdd_2_sbox_n37,
         AesSbox_keyAdd_2_sbox_n36, AesSbox_keyAdd_2_sbox_n35,
         AesSbox_keyAdd_2_sbox_n34, AesSbox_keyAdd_2_sbox_n33,
         AesSbox_keyAdd_2_sbox_n32, AesSbox_keyAdd_2_sbox_n31,
         AesSbox_keyAdd_2_sbox_n30, AesSbox_keyAdd_2_sbox_n29,
         AesSbox_keyAdd_2_sbox_n28, AesSbox_keyAdd_2_sbox_n27,
         AesSbox_keyAdd_2_sbox_n26, AesSbox_keyAdd_2_sbox_n25,
         AesSbox_keyAdd_2_sbox_n24, AesSbox_keyAdd_2_sbox_n23,
         AesSbox_keyAdd_2_sbox_n22, AesSbox_keyAdd_2_sbox_n21,
         AesSbox_keyAdd_2_sbox_n20, AesSbox_keyAdd_2_sbox_n19,
         AesSbox_keyAdd_2_sbox_n18, AesSbox_keyAdd_2_sbox_n17,
         AesSbox_keyAdd_2_sbox_n16, AesSbox_keyAdd_2_sbox_n15,
         AesSbox_keyAdd_2_sbox_n14, AesSbox_keyAdd_2_sbox_n13,
         AesSbox_keyAdd_2_sbox_n12, AesSbox_keyAdd_2_sbox_n11,
         AesSbox_keyAdd_2_sbox_n10, AesSbox_keyAdd_2_sbox_n9,
         AesSbox_keyAdd_2_sbox_n8, AesSbox_keyAdd_2_sbox_n7,
         AesSbox_keyAdd_2_sbox_n6, AesSbox_keyAdd_2_sbox_n5,
         AesSbox_keyAdd_2_sbox_n4, AesSbox_keyAdd_2_sbox_n3,
         AesSbox_keyAdd_2_sbox_n2, AesSbox_keyAdd_2_sbox_n1;
  wire   [7:0] output_sbox_0;
  wire   [7:0] output_sbox_2;
  wire   [7:0] output_sbox_1;

  NAND2_X1 U33 ( .A1(n25), .A2(n26), .ZN(io_out[7]) );
  NAND2_X1 U34 ( .A1(output_sbox_2[7]), .A2(n27), .ZN(n26) );
  OR2_X1 U35 ( .A1(output_sbox_1[7]), .A2(output_sbox_0[7]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(output_sbox_1[7]), .A2(output_sbox_0[7]), .ZN(n25) );
  NAND2_X1 U37 ( .A1(n28), .A2(n29), .ZN(io_out[6]) );
  NAND2_X1 U38 ( .A1(output_sbox_2[6]), .A2(n30), .ZN(n29) );
  OR2_X1 U39 ( .A1(output_sbox_1[6]), .A2(output_sbox_0[6]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(output_sbox_1[6]), .A2(output_sbox_0[6]), .ZN(n28) );
  NAND2_X1 U41 ( .A1(n31), .A2(n32), .ZN(io_out[5]) );
  NAND2_X1 U42 ( .A1(output_sbox_2[5]), .A2(n33), .ZN(n32) );
  OR2_X1 U43 ( .A1(output_sbox_1[5]), .A2(output_sbox_0[5]), .ZN(n33) );
  NAND2_X1 U44 ( .A1(output_sbox_1[5]), .A2(output_sbox_0[5]), .ZN(n31) );
  NAND2_X1 U45 ( .A1(n34), .A2(n35), .ZN(io_out[4]) );
  NAND2_X1 U46 ( .A1(output_sbox_2[4]), .A2(n36), .ZN(n35) );
  OR2_X1 U47 ( .A1(output_sbox_1[4]), .A2(output_sbox_0[4]), .ZN(n36) );
  NAND2_X1 U48 ( .A1(output_sbox_1[4]), .A2(output_sbox_0[4]), .ZN(n34) );
  NAND2_X1 U49 ( .A1(n37), .A2(n38), .ZN(io_out[3]) );
  NAND2_X1 U50 ( .A1(output_sbox_2[3]), .A2(n39), .ZN(n38) );
  OR2_X1 U51 ( .A1(output_sbox_1[3]), .A2(output_sbox_0[3]), .ZN(n39) );
  NAND2_X1 U52 ( .A1(output_sbox_1[3]), .A2(output_sbox_0[3]), .ZN(n37) );
  NAND2_X1 U53 ( .A1(n40), .A2(n41), .ZN(io_out[2]) );
  NAND2_X1 U54 ( .A1(output_sbox_2[2]), .A2(n42), .ZN(n41) );
  OR2_X1 U55 ( .A1(output_sbox_1[2]), .A2(output_sbox_0[2]), .ZN(n42) );
  NAND2_X1 U56 ( .A1(output_sbox_1[2]), .A2(output_sbox_0[2]), .ZN(n40) );
  NAND2_X1 U57 ( .A1(n43), .A2(n44), .ZN(io_out[1]) );
  NAND2_X1 U58 ( .A1(output_sbox_2[1]), .A2(n45), .ZN(n44) );
  OR2_X1 U59 ( .A1(output_sbox_1[1]), .A2(output_sbox_0[1]), .ZN(n45) );
  NAND2_X1 U60 ( .A1(output_sbox_1[1]), .A2(output_sbox_0[1]), .ZN(n43) );
  NAND2_X1 U61 ( .A1(n46), .A2(n47), .ZN(io_out[0]) );
  NAND2_X1 U62 ( .A1(output_sbox_2[0]), .A2(n48), .ZN(n47) );
  OR2_X1 U63 ( .A1(output_sbox_1[0]), .A2(output_sbox_0[0]), .ZN(n48) );
  NAND2_X1 U64 ( .A1(output_sbox_1[0]), .A2(output_sbox_0[0]), .ZN(n46) );
  XOR2_X1 AesSbox_keyAdd_U8 ( .A(AesSbox_keyAdd_sbox_io_o0), .B(io_key[0]), 
        .Z(output_sbox_0[0]) );
  XOR2_X1 AesSbox_keyAdd_U7 ( .A(AesSbox_keyAdd_sbox_io_o1), .B(io_key[1]), 
        .Z(output_sbox_0[1]) );
  XOR2_X1 AesSbox_keyAdd_U6 ( .A(AesSbox_keyAdd_sbox_io_o2), .B(io_key[2]), 
        .Z(output_sbox_0[2]) );
  XOR2_X1 AesSbox_keyAdd_U5 ( .A(AesSbox_keyAdd_sbox_io_o3), .B(io_key[3]), 
        .Z(output_sbox_0[3]) );
  XOR2_X1 AesSbox_keyAdd_U4 ( .A(AesSbox_keyAdd_sbox_io_o4), .B(io_key[4]), 
        .Z(output_sbox_0[4]) );
  XOR2_X1 AesSbox_keyAdd_U3 ( .A(AesSbox_keyAdd_sbox_io_o5), .B(io_key[5]), 
        .Z(output_sbox_0[5]) );
  XOR2_X1 AesSbox_keyAdd_U2 ( .A(AesSbox_keyAdd_sbox_io_o6), .B(io_key[6]), 
        .Z(output_sbox_0[6]) );
  XOR2_X1 AesSbox_keyAdd_U1 ( .A(AesSbox_keyAdd_sbox_io_o7), .B(io_key[7]), 
        .Z(output_sbox_0[7]) );
  XOR2_X1 AesSbox_keyAdd_sbox_U136 ( .A(io_state[0]), .B(io_state[3]), .Z(
        AesSbox_keyAdd_sbox_n71) );
  XOR2_X1 AesSbox_keyAdd_sbox_U135 ( .A(io_state[2]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_sbox_n107) );
  XOR2_X1 AesSbox_keyAdd_sbox_U134 ( .A(AesSbox_keyAdd_sbox_n71), .B(
        AesSbox_keyAdd_sbox_n107), .Z(AesSbox_keyAdd_sbox_n75) );
  XOR2_X1 AesSbox_keyAdd_sbox_U133 ( .A(io_state[1]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_sbox_n126) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U132 ( .A(io_state[6]), .B(io_state[4]), .ZN(
        AesSbox_keyAdd_sbox_n125) );
  INV_X1 AesSbox_keyAdd_sbox_U131 ( .A(AesSbox_keyAdd_sbox_n125), .ZN(
        AesSbox_keyAdd_sbox_n108) );
  XOR2_X1 AesSbox_keyAdd_sbox_U130 ( .A(AesSbox_keyAdd_sbox_n108), .B(
        AesSbox_keyAdd_sbox_n126), .Z(AesSbox_keyAdd_sbox_n74) );
  NAND2_X1 AesSbox_keyAdd_sbox_U129 ( .A1(AesSbox_keyAdd_sbox_n74), .A2(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n117) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U128 ( .A(io_state[3]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_sbox_n124) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U127 ( .A(AesSbox_keyAdd_sbox_n107), .B(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n128) );
  NOR2_X1 AesSbox_keyAdd_sbox_U126 ( .A1(AesSbox_keyAdd_sbox_n124), .A2(
        AesSbox_keyAdd_sbox_n128), .ZN(AesSbox_keyAdd_sbox_n127) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U125 ( .A(AesSbox_keyAdd_sbox_n117), .B(
        AesSbox_keyAdd_sbox_n127), .ZN(AesSbox_keyAdd_sbox_n100) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U124 ( .A(AesSbox_keyAdd_sbox_n126), .B(
        AesSbox_keyAdd_sbox_n100), .ZN(AesSbox_keyAdd_sbox_n120) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U123 ( .A(AesSbox_keyAdd_sbox_n125), .B(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n61) );
  INV_X1 AesSbox_keyAdd_sbox_U122 ( .A(AesSbox_keyAdd_sbox_n124), .ZN(
        AesSbox_keyAdd_sbox_n73) );
  XOR2_X1 AesSbox_keyAdd_sbox_U121 ( .A(io_state[0]), .B(io_state[6]), .Z(
        AesSbox_keyAdd_sbox_n48) );
  XOR2_X1 AesSbox_keyAdd_sbox_U120 ( .A(AesSbox_keyAdd_sbox_n73), .B(
        AesSbox_keyAdd_sbox_n48), .Z(AesSbox_keyAdd_sbox_n64) );
  NAND2_X1 AesSbox_keyAdd_sbox_U119 ( .A1(AesSbox_keyAdd_sbox_n64), .A2(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n113) );
  XOR2_X1 AesSbox_keyAdd_sbox_U118 ( .A(io_state[1]), .B(io_state[2]), .Z(
        AesSbox_keyAdd_sbox_n119) );
  XOR2_X1 AesSbox_keyAdd_sbox_U117 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_sbox_n119), .Z(AesSbox_keyAdd_sbox_n66) );
  INV_X1 AesSbox_keyAdd_sbox_U116 ( .A(AesSbox_keyAdd_sbox_n66), .ZN(
        AesSbox_keyAdd_sbox_n115) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U115 ( .A(AesSbox_keyAdd_sbox_n115), .B(
        io_state[6]), .ZN(AesSbox_keyAdd_sbox_n14) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U114 ( .A(io_state[0]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_sbox_n116) );
  XOR2_X1 AesSbox_keyAdd_sbox_U113 ( .A(AesSbox_keyAdd_sbox_n14), .B(
        AesSbox_keyAdd_sbox_n116), .Z(AesSbox_keyAdd_sbox_n65) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U112 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n58) );
  NOR2_X1 AesSbox_keyAdd_sbox_U111 ( .A1(AesSbox_keyAdd_sbox_n65), .A2(
        AesSbox_keyAdd_sbox_n58), .ZN(AesSbox_keyAdd_sbox_n123) );
  XOR2_X1 AesSbox_keyAdd_sbox_U110 ( .A(AesSbox_keyAdd_sbox_n113), .B(
        AesSbox_keyAdd_sbox_n123), .Z(AesSbox_keyAdd_sbox_n122) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U109 ( .A(AesSbox_keyAdd_sbox_n61), .B(
        AesSbox_keyAdd_sbox_n122), .ZN(AesSbox_keyAdd_sbox_n121) );
  XOR2_X1 AesSbox_keyAdd_sbox_U108 ( .A(AesSbox_keyAdd_sbox_n120), .B(
        AesSbox_keyAdd_sbox_n121), .Z(AesSbox_keyAdd_sbox_n109) );
  INV_X1 AesSbox_keyAdd_sbox_U107 ( .A(AesSbox_keyAdd_sbox_n109), .ZN(
        AesSbox_keyAdd_sbox_n94) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U106 ( .A(AesSbox_keyAdd_sbox_n119), .B(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n45) );
  NOR2_X1 AesSbox_keyAdd_sbox_U105 ( .A1(AesSbox_keyAdd_sbox_n45), .A2(
        AesSbox_keyAdd_sbox_n116), .ZN(AesSbox_keyAdd_sbox_n118) );
  XOR2_X1 AesSbox_keyAdd_sbox_U104 ( .A(AesSbox_keyAdd_sbox_n117), .B(
        AesSbox_keyAdd_sbox_n118), .Z(AesSbox_keyAdd_sbox_n104) );
  INV_X1 AesSbox_keyAdd_sbox_U103 ( .A(AesSbox_keyAdd_sbox_n116), .ZN(
        AesSbox_keyAdd_sbox_n43) );
  XOR2_X1 AesSbox_keyAdd_sbox_U102 ( .A(AesSbox_keyAdd_sbox_n104), .B(
        AesSbox_keyAdd_sbox_n43), .Z(AesSbox_keyAdd_sbox_n110) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U101 ( .A(AesSbox_keyAdd_sbox_n115), .B(
        io_state[3]), .ZN(AesSbox_keyAdd_sbox_n25) );
  AND2_X1 AesSbox_keyAdd_sbox_U100 ( .A1(AesSbox_keyAdd_sbox_n25), .A2(
        io_state[7]), .ZN(AesSbox_keyAdd_sbox_n114) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U99 ( .A(AesSbox_keyAdd_sbox_n113), .B(
        AesSbox_keyAdd_sbox_n114), .ZN(AesSbox_keyAdd_sbox_n112) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U98 ( .A(AesSbox_keyAdd_sbox_n45), .B(
        AesSbox_keyAdd_sbox_n112), .ZN(AesSbox_keyAdd_sbox_n111) );
  XOR2_X1 AesSbox_keyAdd_sbox_U97 ( .A(AesSbox_keyAdd_sbox_n110), .B(
        AesSbox_keyAdd_sbox_n111), .Z(AesSbox_keyAdd_sbox_n81) );
  XOR2_X1 AesSbox_keyAdd_sbox_U96 ( .A(AesSbox_keyAdd_sbox_n109), .B(
        AesSbox_keyAdd_sbox_n81), .Z(AesSbox_keyAdd_sbox_n84) );
  AND2_X1 AesSbox_keyAdd_sbox_U95 ( .A1(AesSbox_keyAdd_sbox_n94), .A2(
        AesSbox_keyAdd_sbox_n84), .ZN(AesSbox_keyAdd_sbox_n101) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U94 ( .A(AesSbox_keyAdd_sbox_n25), .B(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n50) );
  XOR2_X1 AesSbox_keyAdd_sbox_U93 ( .A(AesSbox_keyAdd_sbox_n107), .B(
        AesSbox_keyAdd_sbox_n108), .Z(AesSbox_keyAdd_sbox_n68) );
  AND2_X1 AesSbox_keyAdd_sbox_U92 ( .A1(AesSbox_keyAdd_sbox_n68), .A2(
        AesSbox_keyAdd_sbox_n48), .ZN(AesSbox_keyAdd_sbox_n98) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U91 ( .A(AesSbox_keyAdd_sbox_n66), .B(
        AesSbox_keyAdd_sbox_n68), .ZN(AesSbox_keyAdd_sbox_n33) );
  NOR2_X1 AesSbox_keyAdd_sbox_U90 ( .A1(AesSbox_keyAdd_sbox_n50), .A2(
        AesSbox_keyAdd_sbox_n33), .ZN(AesSbox_keyAdd_sbox_n106) );
  XOR2_X1 AesSbox_keyAdd_sbox_U89 ( .A(AesSbox_keyAdd_sbox_n98), .B(
        AesSbox_keyAdd_sbox_n106), .Z(AesSbox_keyAdd_sbox_n105) );
  XOR2_X1 AesSbox_keyAdd_sbox_U88 ( .A(AesSbox_keyAdd_sbox_n50), .B(
        AesSbox_keyAdd_sbox_n105), .Z(AesSbox_keyAdd_sbox_n102) );
  XOR2_X1 AesSbox_keyAdd_sbox_U87 ( .A(AesSbox_keyAdd_sbox_n33), .B(
        AesSbox_keyAdd_sbox_n104), .Z(AesSbox_keyAdd_sbox_n103) );
  XOR2_X1 AesSbox_keyAdd_sbox_U86 ( .A(AesSbox_keyAdd_sbox_n102), .B(
        AesSbox_keyAdd_sbox_n103), .Z(AesSbox_keyAdd_sbox_n85) );
  INV_X1 AesSbox_keyAdd_sbox_U85 ( .A(AesSbox_keyAdd_sbox_n85), .ZN(
        AesSbox_keyAdd_sbox_n77) );
  NAND2_X1 AesSbox_keyAdd_sbox_U84 ( .A1(AesSbox_keyAdd_sbox_n101), .A2(
        AesSbox_keyAdd_sbox_n77), .ZN(AesSbox_keyAdd_sbox_n93) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U83 ( .A(AesSbox_keyAdd_sbox_n48), .B(
        AesSbox_keyAdd_sbox_n100), .ZN(AesSbox_keyAdd_sbox_n95) );
  AND2_X1 AesSbox_keyAdd_sbox_U82 ( .A1(AesSbox_keyAdd_sbox_n66), .A2(
        AesSbox_keyAdd_sbox_n14), .ZN(AesSbox_keyAdd_sbox_n99) );
  XOR2_X1 AesSbox_keyAdd_sbox_U81 ( .A(AesSbox_keyAdd_sbox_n98), .B(
        AesSbox_keyAdd_sbox_n99), .Z(AesSbox_keyAdd_sbox_n97) );
  XOR2_X1 AesSbox_keyAdd_sbox_U80 ( .A(AesSbox_keyAdd_sbox_n68), .B(
        AesSbox_keyAdd_sbox_n97), .Z(AesSbox_keyAdd_sbox_n96) );
  XOR2_X1 AesSbox_keyAdd_sbox_U79 ( .A(AesSbox_keyAdd_sbox_n95), .B(
        AesSbox_keyAdd_sbox_n96), .Z(AesSbox_keyAdd_sbox_n91) );
  INV_X1 AesSbox_keyAdd_sbox_U78 ( .A(AesSbox_keyAdd_sbox_n91), .ZN(
        AesSbox_keyAdd_sbox_n90) );
  NAND2_X1 AesSbox_keyAdd_sbox_U77 ( .A1(AesSbox_keyAdd_sbox_n90), .A2(
        AesSbox_keyAdd_sbox_n94), .ZN(AesSbox_keyAdd_sbox_n80) );
  INV_X1 AesSbox_keyAdd_sbox_U76 ( .A(AesSbox_keyAdd_sbox_n80), .ZN(
        AesSbox_keyAdd_sbox_n88) );
  XOR2_X1 AesSbox_keyAdd_sbox_U75 ( .A(AesSbox_keyAdd_sbox_n93), .B(
        AesSbox_keyAdd_sbox_n88), .Z(AesSbox_keyAdd_sbox_n92) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U74 ( .A(AesSbox_keyAdd_sbox_n92), .B(
        AesSbox_keyAdd_sbox_n84), .ZN(AesSbox_keyAdd_sbox_n13) );
  NOR2_X1 AesSbox_keyAdd_sbox_U73 ( .A1(AesSbox_keyAdd_sbox_n81), .A2(
        AesSbox_keyAdd_sbox_n91), .ZN(AesSbox_keyAdd_sbox_n89) );
  XOR2_X1 AesSbox_keyAdd_sbox_U72 ( .A(AesSbox_keyAdd_sbox_n77), .B(
        AesSbox_keyAdd_sbox_n90), .Z(AesSbox_keyAdd_sbox_n79) );
  NAND2_X1 AesSbox_keyAdd_sbox_U71 ( .A1(AesSbox_keyAdd_sbox_n89), .A2(
        AesSbox_keyAdd_sbox_n79), .ZN(AesSbox_keyAdd_sbox_n87) );
  XOR2_X1 AesSbox_keyAdd_sbox_U70 ( .A(AesSbox_keyAdd_sbox_n87), .B(
        AesSbox_keyAdd_sbox_n88), .Z(AesSbox_keyAdd_sbox_n86) );
  XOR2_X1 AesSbox_keyAdd_sbox_U69 ( .A(AesSbox_keyAdd_sbox_n86), .B(
        AesSbox_keyAdd_sbox_n79), .Z(AesSbox_keyAdd_sbox_n59) );
  XOR2_X1 AesSbox_keyAdd_sbox_U68 ( .A(AesSbox_keyAdd_sbox_n13), .B(
        AesSbox_keyAdd_sbox_n59), .Z(AesSbox_keyAdd_sbox_n46) );
  INV_X1 AesSbox_keyAdd_sbox_U67 ( .A(AesSbox_keyAdd_sbox_n46), .ZN(
        AesSbox_keyAdd_sbox_n42) );
  XOR2_X1 AesSbox_keyAdd_sbox_U66 ( .A(AesSbox_keyAdd_sbox_n80), .B(
        AesSbox_keyAdd_sbox_n85), .Z(AesSbox_keyAdd_sbox_n83) );
  NAND2_X1 AesSbox_keyAdd_sbox_U65 ( .A1(AesSbox_keyAdd_sbox_n83), .A2(
        AesSbox_keyAdd_sbox_n84), .ZN(AesSbox_keyAdd_sbox_n82) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U64 ( .A(AesSbox_keyAdd_sbox_n82), .B(
        AesSbox_keyAdd_sbox_n81), .ZN(AesSbox_keyAdd_sbox_n32) );
  XOR2_X1 AesSbox_keyAdd_sbox_U63 ( .A(AesSbox_keyAdd_sbox_n80), .B(
        AesSbox_keyAdd_sbox_n81), .Z(AesSbox_keyAdd_sbox_n78) );
  NAND2_X1 AesSbox_keyAdd_sbox_U62 ( .A1(AesSbox_keyAdd_sbox_n78), .A2(
        AesSbox_keyAdd_sbox_n79), .ZN(AesSbox_keyAdd_sbox_n76) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U61 ( .A(AesSbox_keyAdd_sbox_n76), .B(
        AesSbox_keyAdd_sbox_n77), .ZN(AesSbox_keyAdd_sbox_n24) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U60 ( .A(AesSbox_keyAdd_sbox_n32), .B(
        AesSbox_keyAdd_sbox_n24), .ZN(AesSbox_keyAdd_sbox_n70) );
  XOR2_X1 AesSbox_keyAdd_sbox_U59 ( .A(AesSbox_keyAdd_sbox_n42), .B(
        AesSbox_keyAdd_sbox_n70), .Z(AesSbox_keyAdd_sbox_n72) );
  NAND2_X1 AesSbox_keyAdd_sbox_U58 ( .A1(AesSbox_keyAdd_sbox_n75), .A2(
        AesSbox_keyAdd_sbox_n72), .ZN(AesSbox_keyAdd_sbox_n22) );
  NAND2_X1 AesSbox_keyAdd_sbox_U57 ( .A1(AesSbox_keyAdd_sbox_n74), .A2(
        AesSbox_keyAdd_sbox_n70), .ZN(AesSbox_keyAdd_sbox_n40) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U56 ( .A(AesSbox_keyAdd_sbox_n22), .B(
        AesSbox_keyAdd_sbox_n40), .ZN(AesSbox_keyAdd_sbox_n55) );
  NAND2_X1 AesSbox_keyAdd_sbox_U55 ( .A1(AesSbox_keyAdd_sbox_n72), .A2(
        AesSbox_keyAdd_sbox_n73), .ZN(AesSbox_keyAdd_sbox_n69) );
  AND2_X1 AesSbox_keyAdd_sbox_U54 ( .A1(AesSbox_keyAdd_sbox_n70), .A2(
        AesSbox_keyAdd_sbox_n71), .ZN(AesSbox_keyAdd_sbox_n41) );
  XOR2_X1 AesSbox_keyAdd_sbox_U53 ( .A(AesSbox_keyAdd_sbox_n69), .B(
        AesSbox_keyAdd_sbox_n41), .Z(AesSbox_keyAdd_sbox_n15) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U52 ( .A(AesSbox_keyAdd_sbox_n13), .B(
        AesSbox_keyAdd_sbox_n32), .ZN(AesSbox_keyAdd_sbox_n47) );
  AND2_X1 AesSbox_keyAdd_sbox_U51 ( .A1(AesSbox_keyAdd_sbox_n68), .A2(
        AesSbox_keyAdd_sbox_n47), .ZN(AesSbox_keyAdd_sbox_n67) );
  XOR2_X1 AesSbox_keyAdd_sbox_U50 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n67), .Z(AesSbox_keyAdd_sbox_n4) );
  NAND2_X1 AesSbox_keyAdd_sbox_U49 ( .A1(AesSbox_keyAdd_sbox_n13), .A2(
        AesSbox_keyAdd_sbox_n66), .ZN(AesSbox_keyAdd_sbox_n16) );
  NOR2_X1 AesSbox_keyAdd_sbox_U48 ( .A1(AesSbox_keyAdd_sbox_n59), .A2(
        AesSbox_keyAdd_sbox_n65), .ZN(AesSbox_keyAdd_sbox_n62) );
  XOR2_X1 AesSbox_keyAdd_sbox_U47 ( .A(AesSbox_keyAdd_sbox_n16), .B(
        AesSbox_keyAdd_sbox_n62), .Z(AesSbox_keyAdd_sbox_n28) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U46 ( .A(AesSbox_keyAdd_sbox_n4), .B(
        AesSbox_keyAdd_sbox_n28), .ZN(AesSbox_keyAdd_sbox_n35) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U45 ( .A(AesSbox_keyAdd_sbox_n24), .B(
        AesSbox_keyAdd_sbox_n59), .ZN(AesSbox_keyAdd_sbox_n60) );
  AND2_X1 AesSbox_keyAdd_sbox_U44 ( .A1(AesSbox_keyAdd_sbox_n60), .A2(
        AesSbox_keyAdd_sbox_n64), .ZN(AesSbox_keyAdd_sbox_n56) );
  XOR2_X1 AesSbox_keyAdd_sbox_U43 ( .A(AesSbox_keyAdd_sbox_n35), .B(
        AesSbox_keyAdd_sbox_n56), .Z(AesSbox_keyAdd_sbox_n63) );
  XOR2_X1 AesSbox_keyAdd_sbox_U42 ( .A(AesSbox_keyAdd_sbox_n55), .B(
        AesSbox_keyAdd_sbox_n63), .Z(AesSbox_keyAdd_sbox_io_o0) );
  XOR2_X1 AesSbox_keyAdd_sbox_U41 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n62), .Z(AesSbox_keyAdd_sbox_n52) );
  NAND2_X1 AesSbox_keyAdd_sbox_U40 ( .A1(AesSbox_keyAdd_sbox_n60), .A2(
        AesSbox_keyAdd_sbox_n61), .ZN(AesSbox_keyAdd_sbox_n51) );
  NOR2_X1 AesSbox_keyAdd_sbox_U39 ( .A1(AesSbox_keyAdd_sbox_n58), .A2(
        AesSbox_keyAdd_sbox_n59), .ZN(AesSbox_keyAdd_sbox_n57) );
  XOR2_X1 AesSbox_keyAdd_sbox_U38 ( .A(AesSbox_keyAdd_sbox_n56), .B(
        AesSbox_keyAdd_sbox_n57), .Z(AesSbox_keyAdd_sbox_n29) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U37 ( .A(AesSbox_keyAdd_sbox_n51), .B(
        AesSbox_keyAdd_sbox_n29), .ZN(AesSbox_keyAdd_sbox_n34) );
  INV_X1 AesSbox_keyAdd_sbox_U36 ( .A(AesSbox_keyAdd_sbox_n55), .ZN(
        AesSbox_keyAdd_sbox_n54) );
  XOR2_X1 AesSbox_keyAdd_sbox_U35 ( .A(AesSbox_keyAdd_sbox_n34), .B(
        AesSbox_keyAdd_sbox_n54), .Z(AesSbox_keyAdd_sbox_n53) );
  XOR2_X1 AesSbox_keyAdd_sbox_U34 ( .A(AesSbox_keyAdd_sbox_n52), .B(
        AesSbox_keyAdd_sbox_n53), .Z(AesSbox_keyAdd_sbox_io_o1) );
  NAND2_X1 AesSbox_keyAdd_sbox_U33 ( .A1(io_state[7]), .A2(
        AesSbox_keyAdd_sbox_n24), .ZN(AesSbox_keyAdd_sbox_n31) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U32 ( .A(AesSbox_keyAdd_sbox_n51), .B(
        AesSbox_keyAdd_sbox_n31), .ZN(AesSbox_keyAdd_sbox_n5) );
  NOR2_X1 AesSbox_keyAdd_sbox_U31 ( .A1(AesSbox_keyAdd_sbox_n50), .A2(
        AesSbox_keyAdd_sbox_n32), .ZN(AesSbox_keyAdd_sbox_n49) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U30 ( .A(AesSbox_keyAdd_sbox_n5), .B(
        AesSbox_keyAdd_sbox_n49), .ZN(AesSbox_keyAdd_sbox_n20) );
  NAND2_X1 AesSbox_keyAdd_sbox_U29 ( .A1(AesSbox_keyAdd_sbox_n47), .A2(
        AesSbox_keyAdd_sbox_n48), .ZN(AesSbox_keyAdd_sbox_n3) );
  NOR2_X1 AesSbox_keyAdd_sbox_U28 ( .A1(AesSbox_keyAdd_sbox_n45), .A2(
        AesSbox_keyAdd_sbox_n46), .ZN(AesSbox_keyAdd_sbox_n44) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U27 ( .A(AesSbox_keyAdd_sbox_n3), .B(
        AesSbox_keyAdd_sbox_n44), .ZN(AesSbox_keyAdd_sbox_n23) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U26 ( .A(AesSbox_keyAdd_sbox_n20), .B(
        AesSbox_keyAdd_sbox_n23), .ZN(AesSbox_keyAdd_sbox_n36) );
  NAND2_X1 AesSbox_keyAdd_sbox_U25 ( .A1(AesSbox_keyAdd_sbox_n42), .A2(
        AesSbox_keyAdd_sbox_n43), .ZN(AesSbox_keyAdd_sbox_n38) );
  XOR2_X1 AesSbox_keyAdd_sbox_U24 ( .A(AesSbox_keyAdd_sbox_n40), .B(
        AesSbox_keyAdd_sbox_n41), .Z(AesSbox_keyAdd_sbox_n39) );
  XOR2_X1 AesSbox_keyAdd_sbox_U23 ( .A(AesSbox_keyAdd_sbox_n38), .B(
        AesSbox_keyAdd_sbox_n39), .Z(AesSbox_keyAdd_sbox_n37) );
  XOR2_X1 AesSbox_keyAdd_sbox_U22 ( .A(AesSbox_keyAdd_sbox_n36), .B(
        AesSbox_keyAdd_sbox_n37), .Z(AesSbox_keyAdd_sbox_io_o2) );
  INV_X1 AesSbox_keyAdd_sbox_U21 ( .A(AesSbox_keyAdd_sbox_n35), .ZN(
        AesSbox_keyAdd_sbox_n19) );
  XOR2_X1 AesSbox_keyAdd_sbox_U20 ( .A(AesSbox_keyAdd_sbox_n19), .B(
        AesSbox_keyAdd_sbox_n34), .Z(AesSbox_keyAdd_sbox_io_o3) );
  NOR2_X1 AesSbox_keyAdd_sbox_U19 ( .A1(AesSbox_keyAdd_sbox_n32), .A2(
        AesSbox_keyAdd_sbox_n33), .ZN(AesSbox_keyAdd_sbox_n12) );
  XOR2_X1 AesSbox_keyAdd_sbox_U18 ( .A(AesSbox_keyAdd_sbox_n31), .B(
        AesSbox_keyAdd_sbox_n12), .Z(AesSbox_keyAdd_sbox_n30) );
  XOR2_X1 AesSbox_keyAdd_sbox_U17 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n30), .Z(AesSbox_keyAdd_sbox_n26) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U16 ( .A(AesSbox_keyAdd_sbox_n28), .B(
        AesSbox_keyAdd_sbox_n29), .ZN(AesSbox_keyAdd_sbox_n27) );
  XOR2_X1 AesSbox_keyAdd_sbox_U15 ( .A(AesSbox_keyAdd_sbox_n26), .B(
        AesSbox_keyAdd_sbox_n27), .Z(AesSbox_keyAdd_sbox_io_o4) );
  NAND2_X1 AesSbox_keyAdd_sbox_U14 ( .A1(AesSbox_keyAdd_sbox_n24), .A2(
        AesSbox_keyAdd_sbox_n25), .ZN(AesSbox_keyAdd_sbox_n21) );
  XOR2_X1 AesSbox_keyAdd_sbox_U13 ( .A(AesSbox_keyAdd_sbox_n22), .B(
        AesSbox_keyAdd_sbox_n23), .Z(AesSbox_keyAdd_sbox_n10) );
  XOR2_X1 AesSbox_keyAdd_sbox_U12 ( .A(AesSbox_keyAdd_sbox_n21), .B(
        AesSbox_keyAdd_sbox_n10), .Z(AesSbox_keyAdd_sbox_n17) );
  XOR2_X1 AesSbox_keyAdd_sbox_U11 ( .A(AesSbox_keyAdd_sbox_n19), .B(
        AesSbox_keyAdd_sbox_n20), .Z(AesSbox_keyAdd_sbox_n18) );
  XOR2_X1 AesSbox_keyAdd_sbox_U10 ( .A(AesSbox_keyAdd_sbox_n17), .B(
        AesSbox_keyAdd_sbox_n18), .Z(AesSbox_keyAdd_sbox_io_o5) );
  XNOR2_X1 AesSbox_keyAdd_sbox_U9 ( .A(AesSbox_keyAdd_sbox_n15), .B(
        AesSbox_keyAdd_sbox_n16), .ZN(AesSbox_keyAdd_sbox_n8) );
  NAND2_X1 AesSbox_keyAdd_sbox_U8 ( .A1(AesSbox_keyAdd_sbox_n13), .A2(
        AesSbox_keyAdd_sbox_n14), .ZN(AesSbox_keyAdd_sbox_n11) );
  XOR2_X1 AesSbox_keyAdd_sbox_U7 ( .A(AesSbox_keyAdd_sbox_n11), .B(
        AesSbox_keyAdd_sbox_n12), .Z(AesSbox_keyAdd_sbox_n7) );
  XOR2_X1 AesSbox_keyAdd_sbox_U6 ( .A(AesSbox_keyAdd_sbox_n7), .B(
        AesSbox_keyAdd_sbox_n10), .Z(AesSbox_keyAdd_sbox_n9) );
  XOR2_X1 AesSbox_keyAdd_sbox_U5 ( .A(AesSbox_keyAdd_sbox_n8), .B(
        AesSbox_keyAdd_sbox_n9), .Z(AesSbox_keyAdd_sbox_io_o6) );
  INV_X1 AesSbox_keyAdd_sbox_U4 ( .A(AesSbox_keyAdd_sbox_n7), .ZN(
        AesSbox_keyAdd_sbox_n6) );
  XOR2_X1 AesSbox_keyAdd_sbox_U3 ( .A(AesSbox_keyAdd_sbox_n5), .B(
        AesSbox_keyAdd_sbox_n6), .Z(AesSbox_keyAdd_sbox_n1) );
  XOR2_X1 AesSbox_keyAdd_sbox_U2 ( .A(AesSbox_keyAdd_sbox_n3), .B(
        AesSbox_keyAdd_sbox_n4), .Z(AesSbox_keyAdd_sbox_n2) );
  XOR2_X1 AesSbox_keyAdd_sbox_U1 ( .A(AesSbox_keyAdd_sbox_n1), .B(
        AesSbox_keyAdd_sbox_n2), .Z(AesSbox_keyAdd_sbox_io_o7) );
  XOR2_X1 AesSbox_keyAdd_1_U8 ( .A(AesSbox_keyAdd_1_sbox_io_o0), .B(io_key[0]), 
        .Z(output_sbox_1[0]) );
  XOR2_X1 AesSbox_keyAdd_1_U7 ( .A(AesSbox_keyAdd_1_sbox_io_o1), .B(io_key[1]), 
        .Z(output_sbox_1[1]) );
  XOR2_X1 AesSbox_keyAdd_1_U6 ( .A(AesSbox_keyAdd_1_sbox_io_o2), .B(io_key[2]), 
        .Z(output_sbox_1[2]) );
  XOR2_X1 AesSbox_keyAdd_1_U5 ( .A(AesSbox_keyAdd_1_sbox_io_o3), .B(io_key[3]), 
        .Z(output_sbox_1[3]) );
  XOR2_X1 AesSbox_keyAdd_1_U4 ( .A(AesSbox_keyAdd_1_sbox_io_o4), .B(io_key[4]), 
        .Z(output_sbox_1[4]) );
  XOR2_X1 AesSbox_keyAdd_1_U3 ( .A(AesSbox_keyAdd_1_sbox_io_o5), .B(io_key[5]), 
        .Z(output_sbox_1[5]) );
  XOR2_X1 AesSbox_keyAdd_1_U2 ( .A(AesSbox_keyAdd_1_sbox_io_o6), .B(io_key[6]), 
        .Z(output_sbox_1[6]) );
  XOR2_X1 AesSbox_keyAdd_1_U1 ( .A(AesSbox_keyAdd_1_sbox_io_o7), .B(io_key[7]), 
        .Z(output_sbox_1[7]) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U136 ( .A(io_state[0]), .B(io_state[3]), .Z(
        AesSbox_keyAdd_1_sbox_n71) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U135 ( .A(io_state[2]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_1_sbox_n107) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U134 ( .A(AesSbox_keyAdd_1_sbox_n71), .B(
        AesSbox_keyAdd_1_sbox_n107), .Z(AesSbox_keyAdd_1_sbox_n75) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U133 ( .A(io_state[1]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_1_sbox_n126) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U132 ( .A(io_state[6]), .B(io_state[4]), .ZN(
        AesSbox_keyAdd_1_sbox_n125) );
  INV_X1 AesSbox_keyAdd_1_sbox_U131 ( .A(AesSbox_keyAdd_1_sbox_n125), .ZN(
        AesSbox_keyAdd_1_sbox_n108) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U130 ( .A(AesSbox_keyAdd_1_sbox_n108), .B(
        AesSbox_keyAdd_1_sbox_n126), .Z(AesSbox_keyAdd_1_sbox_n74) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U129 ( .A1(AesSbox_keyAdd_1_sbox_n74), .A2(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n117) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U128 ( .A(io_state[3]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_1_sbox_n124) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U127 ( .A(AesSbox_keyAdd_1_sbox_n107), .B(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n128) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U126 ( .A1(AesSbox_keyAdd_1_sbox_n124), .A2(
        AesSbox_keyAdd_1_sbox_n128), .ZN(AesSbox_keyAdd_1_sbox_n127) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U125 ( .A(AesSbox_keyAdd_1_sbox_n117), .B(
        AesSbox_keyAdd_1_sbox_n127), .ZN(AesSbox_keyAdd_1_sbox_n100) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U124 ( .A(AesSbox_keyAdd_1_sbox_n126), .B(
        AesSbox_keyAdd_1_sbox_n100), .ZN(AesSbox_keyAdd_1_sbox_n120) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U123 ( .A(AesSbox_keyAdd_1_sbox_n125), .B(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n61) );
  INV_X1 AesSbox_keyAdd_1_sbox_U122 ( .A(AesSbox_keyAdd_1_sbox_n124), .ZN(
        AesSbox_keyAdd_1_sbox_n73) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U121 ( .A(io_state[0]), .B(io_state[6]), .Z(
        AesSbox_keyAdd_1_sbox_n48) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U120 ( .A(AesSbox_keyAdd_1_sbox_n73), .B(
        AesSbox_keyAdd_1_sbox_n48), .Z(AesSbox_keyAdd_1_sbox_n64) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U119 ( .A1(AesSbox_keyAdd_1_sbox_n64), .A2(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n113) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U118 ( .A(io_state[1]), .B(io_state[2]), .Z(
        AesSbox_keyAdd_1_sbox_n119) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U117 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_1_sbox_n119), .Z(AesSbox_keyAdd_1_sbox_n66) );
  INV_X1 AesSbox_keyAdd_1_sbox_U116 ( .A(AesSbox_keyAdd_1_sbox_n66), .ZN(
        AesSbox_keyAdd_1_sbox_n115) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U115 ( .A(AesSbox_keyAdd_1_sbox_n115), .B(
        io_state[6]), .ZN(AesSbox_keyAdd_1_sbox_n14) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U114 ( .A(io_state[0]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_1_sbox_n116) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U113 ( .A(AesSbox_keyAdd_1_sbox_n14), .B(
        AesSbox_keyAdd_1_sbox_n116), .Z(AesSbox_keyAdd_1_sbox_n65) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U112 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n58) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U111 ( .A1(AesSbox_keyAdd_1_sbox_n65), .A2(
        AesSbox_keyAdd_1_sbox_n58), .ZN(AesSbox_keyAdd_1_sbox_n123) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U110 ( .A(AesSbox_keyAdd_1_sbox_n113), .B(
        AesSbox_keyAdd_1_sbox_n123), .Z(AesSbox_keyAdd_1_sbox_n122) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U109 ( .A(AesSbox_keyAdd_1_sbox_n61), .B(
        AesSbox_keyAdd_1_sbox_n122), .ZN(AesSbox_keyAdd_1_sbox_n121) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U108 ( .A(AesSbox_keyAdd_1_sbox_n120), .B(
        AesSbox_keyAdd_1_sbox_n121), .Z(AesSbox_keyAdd_1_sbox_n109) );
  INV_X1 AesSbox_keyAdd_1_sbox_U107 ( .A(AesSbox_keyAdd_1_sbox_n109), .ZN(
        AesSbox_keyAdd_1_sbox_n94) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U106 ( .A(AesSbox_keyAdd_1_sbox_n119), .B(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n45) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U105 ( .A1(AesSbox_keyAdd_1_sbox_n45), .A2(
        AesSbox_keyAdd_1_sbox_n116), .ZN(AesSbox_keyAdd_1_sbox_n118) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U104 ( .A(AesSbox_keyAdd_1_sbox_n117), .B(
        AesSbox_keyAdd_1_sbox_n118), .Z(AesSbox_keyAdd_1_sbox_n104) );
  INV_X1 AesSbox_keyAdd_1_sbox_U103 ( .A(AesSbox_keyAdd_1_sbox_n116), .ZN(
        AesSbox_keyAdd_1_sbox_n43) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U102 ( .A(AesSbox_keyAdd_1_sbox_n104), .B(
        AesSbox_keyAdd_1_sbox_n43), .Z(AesSbox_keyAdd_1_sbox_n110) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U101 ( .A(AesSbox_keyAdd_1_sbox_n115), .B(
        io_state[3]), .ZN(AesSbox_keyAdd_1_sbox_n25) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U100 ( .A1(AesSbox_keyAdd_1_sbox_n25), .A2(
        io_state[7]), .ZN(AesSbox_keyAdd_1_sbox_n114) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U99 ( .A(AesSbox_keyAdd_1_sbox_n113), .B(
        AesSbox_keyAdd_1_sbox_n114), .ZN(AesSbox_keyAdd_1_sbox_n112) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U98 ( .A(AesSbox_keyAdd_1_sbox_n45), .B(
        AesSbox_keyAdd_1_sbox_n112), .ZN(AesSbox_keyAdd_1_sbox_n111) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U97 ( .A(AesSbox_keyAdd_1_sbox_n110), .B(
        AesSbox_keyAdd_1_sbox_n111), .Z(AesSbox_keyAdd_1_sbox_n81) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U96 ( .A(AesSbox_keyAdd_1_sbox_n109), .B(
        AesSbox_keyAdd_1_sbox_n81), .Z(AesSbox_keyAdd_1_sbox_n84) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U95 ( .A1(AesSbox_keyAdd_1_sbox_n94), .A2(
        AesSbox_keyAdd_1_sbox_n84), .ZN(AesSbox_keyAdd_1_sbox_n101) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U94 ( .A(AesSbox_keyAdd_1_sbox_n25), .B(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n50) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U93 ( .A(AesSbox_keyAdd_1_sbox_n107), .B(
        AesSbox_keyAdd_1_sbox_n108), .Z(AesSbox_keyAdd_1_sbox_n68) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U92 ( .A1(AesSbox_keyAdd_1_sbox_n68), .A2(
        AesSbox_keyAdd_1_sbox_n48), .ZN(AesSbox_keyAdd_1_sbox_n98) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U91 ( .A(AesSbox_keyAdd_1_sbox_n66), .B(
        AesSbox_keyAdd_1_sbox_n68), .ZN(AesSbox_keyAdd_1_sbox_n33) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U90 ( .A1(AesSbox_keyAdd_1_sbox_n50), .A2(
        AesSbox_keyAdd_1_sbox_n33), .ZN(AesSbox_keyAdd_1_sbox_n106) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U89 ( .A(AesSbox_keyAdd_1_sbox_n98), .B(
        AesSbox_keyAdd_1_sbox_n106), .Z(AesSbox_keyAdd_1_sbox_n105) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U88 ( .A(AesSbox_keyAdd_1_sbox_n50), .B(
        AesSbox_keyAdd_1_sbox_n105), .Z(AesSbox_keyAdd_1_sbox_n102) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U87 ( .A(AesSbox_keyAdd_1_sbox_n33), .B(
        AesSbox_keyAdd_1_sbox_n104), .Z(AesSbox_keyAdd_1_sbox_n103) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U86 ( .A(AesSbox_keyAdd_1_sbox_n102), .B(
        AesSbox_keyAdd_1_sbox_n103), .Z(AesSbox_keyAdd_1_sbox_n85) );
  INV_X1 AesSbox_keyAdd_1_sbox_U85 ( .A(AesSbox_keyAdd_1_sbox_n85), .ZN(
        AesSbox_keyAdd_1_sbox_n77) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U84 ( .A1(AesSbox_keyAdd_1_sbox_n101), .A2(
        AesSbox_keyAdd_1_sbox_n77), .ZN(AesSbox_keyAdd_1_sbox_n93) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U83 ( .A(AesSbox_keyAdd_1_sbox_n48), .B(
        AesSbox_keyAdd_1_sbox_n100), .ZN(AesSbox_keyAdd_1_sbox_n95) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U82 ( .A1(AesSbox_keyAdd_1_sbox_n66), .A2(
        AesSbox_keyAdd_1_sbox_n14), .ZN(AesSbox_keyAdd_1_sbox_n99) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U81 ( .A(AesSbox_keyAdd_1_sbox_n98), .B(
        AesSbox_keyAdd_1_sbox_n99), .Z(AesSbox_keyAdd_1_sbox_n97) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U80 ( .A(AesSbox_keyAdd_1_sbox_n68), .B(
        AesSbox_keyAdd_1_sbox_n97), .Z(AesSbox_keyAdd_1_sbox_n96) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U79 ( .A(AesSbox_keyAdd_1_sbox_n95), .B(
        AesSbox_keyAdd_1_sbox_n96), .Z(AesSbox_keyAdd_1_sbox_n91) );
  INV_X1 AesSbox_keyAdd_1_sbox_U78 ( .A(AesSbox_keyAdd_1_sbox_n91), .ZN(
        AesSbox_keyAdd_1_sbox_n90) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U77 ( .A1(AesSbox_keyAdd_1_sbox_n90), .A2(
        AesSbox_keyAdd_1_sbox_n94), .ZN(AesSbox_keyAdd_1_sbox_n80) );
  INV_X1 AesSbox_keyAdd_1_sbox_U76 ( .A(AesSbox_keyAdd_1_sbox_n80), .ZN(
        AesSbox_keyAdd_1_sbox_n88) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U75 ( .A(AesSbox_keyAdd_1_sbox_n93), .B(
        AesSbox_keyAdd_1_sbox_n88), .Z(AesSbox_keyAdd_1_sbox_n92) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U74 ( .A(AesSbox_keyAdd_1_sbox_n92), .B(
        AesSbox_keyAdd_1_sbox_n84), .ZN(AesSbox_keyAdd_1_sbox_n13) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U73 ( .A1(AesSbox_keyAdd_1_sbox_n81), .A2(
        AesSbox_keyAdd_1_sbox_n91), .ZN(AesSbox_keyAdd_1_sbox_n89) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U72 ( .A(AesSbox_keyAdd_1_sbox_n77), .B(
        AesSbox_keyAdd_1_sbox_n90), .Z(AesSbox_keyAdd_1_sbox_n79) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U71 ( .A1(AesSbox_keyAdd_1_sbox_n89), .A2(
        AesSbox_keyAdd_1_sbox_n79), .ZN(AesSbox_keyAdd_1_sbox_n87) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U70 ( .A(AesSbox_keyAdd_1_sbox_n87), .B(
        AesSbox_keyAdd_1_sbox_n88), .Z(AesSbox_keyAdd_1_sbox_n86) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U69 ( .A(AesSbox_keyAdd_1_sbox_n86), .B(
        AesSbox_keyAdd_1_sbox_n79), .Z(AesSbox_keyAdd_1_sbox_n59) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U68 ( .A(AesSbox_keyAdd_1_sbox_n13), .B(
        AesSbox_keyAdd_1_sbox_n59), .Z(AesSbox_keyAdd_1_sbox_n46) );
  INV_X1 AesSbox_keyAdd_1_sbox_U67 ( .A(AesSbox_keyAdd_1_sbox_n46), .ZN(
        AesSbox_keyAdd_1_sbox_n42) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U66 ( .A(AesSbox_keyAdd_1_sbox_n80), .B(
        AesSbox_keyAdd_1_sbox_n85), .Z(AesSbox_keyAdd_1_sbox_n83) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U65 ( .A1(AesSbox_keyAdd_1_sbox_n83), .A2(
        AesSbox_keyAdd_1_sbox_n84), .ZN(AesSbox_keyAdd_1_sbox_n82) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U64 ( .A(AesSbox_keyAdd_1_sbox_n82), .B(
        AesSbox_keyAdd_1_sbox_n81), .ZN(AesSbox_keyAdd_1_sbox_n32) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U63 ( .A(AesSbox_keyAdd_1_sbox_n80), .B(
        AesSbox_keyAdd_1_sbox_n81), .Z(AesSbox_keyAdd_1_sbox_n78) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U62 ( .A1(AesSbox_keyAdd_1_sbox_n78), .A2(
        AesSbox_keyAdd_1_sbox_n79), .ZN(AesSbox_keyAdd_1_sbox_n76) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U61 ( .A(AesSbox_keyAdd_1_sbox_n76), .B(
        AesSbox_keyAdd_1_sbox_n77), .ZN(AesSbox_keyAdd_1_sbox_n24) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U60 ( .A(AesSbox_keyAdd_1_sbox_n32), .B(
        AesSbox_keyAdd_1_sbox_n24), .ZN(AesSbox_keyAdd_1_sbox_n70) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U59 ( .A(AesSbox_keyAdd_1_sbox_n42), .B(
        AesSbox_keyAdd_1_sbox_n70), .Z(AesSbox_keyAdd_1_sbox_n72) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U58 ( .A1(AesSbox_keyAdd_1_sbox_n75), .A2(
        AesSbox_keyAdd_1_sbox_n72), .ZN(AesSbox_keyAdd_1_sbox_n22) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U57 ( .A1(AesSbox_keyAdd_1_sbox_n74), .A2(
        AesSbox_keyAdd_1_sbox_n70), .ZN(AesSbox_keyAdd_1_sbox_n40) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U56 ( .A(AesSbox_keyAdd_1_sbox_n22), .B(
        AesSbox_keyAdd_1_sbox_n40), .ZN(AesSbox_keyAdd_1_sbox_n55) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U55 ( .A1(AesSbox_keyAdd_1_sbox_n72), .A2(
        AesSbox_keyAdd_1_sbox_n73), .ZN(AesSbox_keyAdd_1_sbox_n69) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U54 ( .A1(AesSbox_keyAdd_1_sbox_n70), .A2(
        AesSbox_keyAdd_1_sbox_n71), .ZN(AesSbox_keyAdd_1_sbox_n41) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U53 ( .A(AesSbox_keyAdd_1_sbox_n69), .B(
        AesSbox_keyAdd_1_sbox_n41), .Z(AesSbox_keyAdd_1_sbox_n15) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U52 ( .A(AesSbox_keyAdd_1_sbox_n13), .B(
        AesSbox_keyAdd_1_sbox_n32), .ZN(AesSbox_keyAdd_1_sbox_n47) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U51 ( .A1(AesSbox_keyAdd_1_sbox_n68), .A2(
        AesSbox_keyAdd_1_sbox_n47), .ZN(AesSbox_keyAdd_1_sbox_n67) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U50 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n67), .Z(AesSbox_keyAdd_1_sbox_n4) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U49 ( .A1(AesSbox_keyAdd_1_sbox_n13), .A2(
        AesSbox_keyAdd_1_sbox_n66), .ZN(AesSbox_keyAdd_1_sbox_n16) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U48 ( .A1(AesSbox_keyAdd_1_sbox_n59), .A2(
        AesSbox_keyAdd_1_sbox_n65), .ZN(AesSbox_keyAdd_1_sbox_n62) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U47 ( .A(AesSbox_keyAdd_1_sbox_n16), .B(
        AesSbox_keyAdd_1_sbox_n62), .Z(AesSbox_keyAdd_1_sbox_n28) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U46 ( .A(AesSbox_keyAdd_1_sbox_n4), .B(
        AesSbox_keyAdd_1_sbox_n28), .ZN(AesSbox_keyAdd_1_sbox_n35) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U45 ( .A(AesSbox_keyAdd_1_sbox_n24), .B(
        AesSbox_keyAdd_1_sbox_n59), .ZN(AesSbox_keyAdd_1_sbox_n60) );
  AND2_X1 AesSbox_keyAdd_1_sbox_U44 ( .A1(AesSbox_keyAdd_1_sbox_n60), .A2(
        AesSbox_keyAdd_1_sbox_n64), .ZN(AesSbox_keyAdd_1_sbox_n56) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U43 ( .A(AesSbox_keyAdd_1_sbox_n35), .B(
        AesSbox_keyAdd_1_sbox_n56), .Z(AesSbox_keyAdd_1_sbox_n63) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U42 ( .A(AesSbox_keyAdd_1_sbox_n55), .B(
        AesSbox_keyAdd_1_sbox_n63), .Z(AesSbox_keyAdd_1_sbox_io_o0) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U41 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n62), .Z(AesSbox_keyAdd_1_sbox_n52) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U40 ( .A1(AesSbox_keyAdd_1_sbox_n60), .A2(
        AesSbox_keyAdd_1_sbox_n61), .ZN(AesSbox_keyAdd_1_sbox_n51) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U39 ( .A1(AesSbox_keyAdd_1_sbox_n58), .A2(
        AesSbox_keyAdd_1_sbox_n59), .ZN(AesSbox_keyAdd_1_sbox_n57) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U38 ( .A(AesSbox_keyAdd_1_sbox_n56), .B(
        AesSbox_keyAdd_1_sbox_n57), .Z(AesSbox_keyAdd_1_sbox_n29) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U37 ( .A(AesSbox_keyAdd_1_sbox_n51), .B(
        AesSbox_keyAdd_1_sbox_n29), .ZN(AesSbox_keyAdd_1_sbox_n34) );
  INV_X1 AesSbox_keyAdd_1_sbox_U36 ( .A(AesSbox_keyAdd_1_sbox_n55), .ZN(
        AesSbox_keyAdd_1_sbox_n54) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U35 ( .A(AesSbox_keyAdd_1_sbox_n34), .B(
        AesSbox_keyAdd_1_sbox_n54), .Z(AesSbox_keyAdd_1_sbox_n53) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U34 ( .A(AesSbox_keyAdd_1_sbox_n52), .B(
        AesSbox_keyAdd_1_sbox_n53), .Z(AesSbox_keyAdd_1_sbox_io_o1) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U33 ( .A1(io_state[7]), .A2(
        AesSbox_keyAdd_1_sbox_n24), .ZN(AesSbox_keyAdd_1_sbox_n31) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U32 ( .A(AesSbox_keyAdd_1_sbox_n51), .B(
        AesSbox_keyAdd_1_sbox_n31), .ZN(AesSbox_keyAdd_1_sbox_n5) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U31 ( .A1(AesSbox_keyAdd_1_sbox_n50), .A2(
        AesSbox_keyAdd_1_sbox_n32), .ZN(AesSbox_keyAdd_1_sbox_n49) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U30 ( .A(AesSbox_keyAdd_1_sbox_n5), .B(
        AesSbox_keyAdd_1_sbox_n49), .ZN(AesSbox_keyAdd_1_sbox_n20) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U29 ( .A1(AesSbox_keyAdd_1_sbox_n47), .A2(
        AesSbox_keyAdd_1_sbox_n48), .ZN(AesSbox_keyAdd_1_sbox_n3) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U28 ( .A1(AesSbox_keyAdd_1_sbox_n45), .A2(
        AesSbox_keyAdd_1_sbox_n46), .ZN(AesSbox_keyAdd_1_sbox_n44) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U27 ( .A(AesSbox_keyAdd_1_sbox_n3), .B(
        AesSbox_keyAdd_1_sbox_n44), .ZN(AesSbox_keyAdd_1_sbox_n23) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U26 ( .A(AesSbox_keyAdd_1_sbox_n20), .B(
        AesSbox_keyAdd_1_sbox_n23), .ZN(AesSbox_keyAdd_1_sbox_n36) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U25 ( .A1(AesSbox_keyAdd_1_sbox_n42), .A2(
        AesSbox_keyAdd_1_sbox_n43), .ZN(AesSbox_keyAdd_1_sbox_n38) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U24 ( .A(AesSbox_keyAdd_1_sbox_n40), .B(
        AesSbox_keyAdd_1_sbox_n41), .Z(AesSbox_keyAdd_1_sbox_n39) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U23 ( .A(AesSbox_keyAdd_1_sbox_n38), .B(
        AesSbox_keyAdd_1_sbox_n39), .Z(AesSbox_keyAdd_1_sbox_n37) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U22 ( .A(AesSbox_keyAdd_1_sbox_n36), .B(
        AesSbox_keyAdd_1_sbox_n37), .Z(AesSbox_keyAdd_1_sbox_io_o2) );
  INV_X1 AesSbox_keyAdd_1_sbox_U21 ( .A(AesSbox_keyAdd_1_sbox_n35), .ZN(
        AesSbox_keyAdd_1_sbox_n19) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U20 ( .A(AesSbox_keyAdd_1_sbox_n19), .B(
        AesSbox_keyAdd_1_sbox_n34), .Z(AesSbox_keyAdd_1_sbox_io_o3) );
  NOR2_X1 AesSbox_keyAdd_1_sbox_U19 ( .A1(AesSbox_keyAdd_1_sbox_n32), .A2(
        AesSbox_keyAdd_1_sbox_n33), .ZN(AesSbox_keyAdd_1_sbox_n12) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U18 ( .A(AesSbox_keyAdd_1_sbox_n31), .B(
        AesSbox_keyAdd_1_sbox_n12), .Z(AesSbox_keyAdd_1_sbox_n30) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U17 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n30), .Z(AesSbox_keyAdd_1_sbox_n26) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U16 ( .A(AesSbox_keyAdd_1_sbox_n28), .B(
        AesSbox_keyAdd_1_sbox_n29), .ZN(AesSbox_keyAdd_1_sbox_n27) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U15 ( .A(AesSbox_keyAdd_1_sbox_n26), .B(
        AesSbox_keyAdd_1_sbox_n27), .Z(AesSbox_keyAdd_1_sbox_io_o4) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U14 ( .A1(AesSbox_keyAdd_1_sbox_n24), .A2(
        AesSbox_keyAdd_1_sbox_n25), .ZN(AesSbox_keyAdd_1_sbox_n21) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U13 ( .A(AesSbox_keyAdd_1_sbox_n22), .B(
        AesSbox_keyAdd_1_sbox_n23), .Z(AesSbox_keyAdd_1_sbox_n10) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U12 ( .A(AesSbox_keyAdd_1_sbox_n21), .B(
        AesSbox_keyAdd_1_sbox_n10), .Z(AesSbox_keyAdd_1_sbox_n17) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U11 ( .A(AesSbox_keyAdd_1_sbox_n19), .B(
        AesSbox_keyAdd_1_sbox_n20), .Z(AesSbox_keyAdd_1_sbox_n18) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U10 ( .A(AesSbox_keyAdd_1_sbox_n17), .B(
        AesSbox_keyAdd_1_sbox_n18), .Z(AesSbox_keyAdd_1_sbox_io_o5) );
  XNOR2_X1 AesSbox_keyAdd_1_sbox_U9 ( .A(AesSbox_keyAdd_1_sbox_n15), .B(
        AesSbox_keyAdd_1_sbox_n16), .ZN(AesSbox_keyAdd_1_sbox_n8) );
  NAND2_X1 AesSbox_keyAdd_1_sbox_U8 ( .A1(AesSbox_keyAdd_1_sbox_n13), .A2(
        AesSbox_keyAdd_1_sbox_n14), .ZN(AesSbox_keyAdd_1_sbox_n11) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U7 ( .A(AesSbox_keyAdd_1_sbox_n11), .B(
        AesSbox_keyAdd_1_sbox_n12), .Z(AesSbox_keyAdd_1_sbox_n7) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U6 ( .A(AesSbox_keyAdd_1_sbox_n7), .B(
        AesSbox_keyAdd_1_sbox_n10), .Z(AesSbox_keyAdd_1_sbox_n9) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U5 ( .A(AesSbox_keyAdd_1_sbox_n8), .B(
        AesSbox_keyAdd_1_sbox_n9), .Z(AesSbox_keyAdd_1_sbox_io_o6) );
  INV_X1 AesSbox_keyAdd_1_sbox_U4 ( .A(AesSbox_keyAdd_1_sbox_n7), .ZN(
        AesSbox_keyAdd_1_sbox_n6) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U3 ( .A(AesSbox_keyAdd_1_sbox_n5), .B(
        AesSbox_keyAdd_1_sbox_n6), .Z(AesSbox_keyAdd_1_sbox_n1) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U2 ( .A(AesSbox_keyAdd_1_sbox_n3), .B(
        AesSbox_keyAdd_1_sbox_n4), .Z(AesSbox_keyAdd_1_sbox_n2) );
  XOR2_X1 AesSbox_keyAdd_1_sbox_U1 ( .A(AesSbox_keyAdd_1_sbox_n1), .B(
        AesSbox_keyAdd_1_sbox_n2), .Z(AesSbox_keyAdd_1_sbox_io_o7) );
  XOR2_X1 AesSbox_keyAdd_2_U8 ( .A(AesSbox_keyAdd_2_sbox_io_o0), .B(io_key[0]), 
        .Z(output_sbox_2[0]) );
  XOR2_X1 AesSbox_keyAdd_2_U7 ( .A(AesSbox_keyAdd_2_sbox_io_o1), .B(io_key[1]), 
        .Z(output_sbox_2[1]) );
  XOR2_X1 AesSbox_keyAdd_2_U6 ( .A(AesSbox_keyAdd_2_sbox_io_o2), .B(io_key[2]), 
        .Z(output_sbox_2[2]) );
  XOR2_X1 AesSbox_keyAdd_2_U5 ( .A(AesSbox_keyAdd_2_sbox_io_o3), .B(io_key[3]), 
        .Z(output_sbox_2[3]) );
  XOR2_X1 AesSbox_keyAdd_2_U4 ( .A(AesSbox_keyAdd_2_sbox_io_o4), .B(io_key[4]), 
        .Z(output_sbox_2[4]) );
  XOR2_X1 AesSbox_keyAdd_2_U3 ( .A(AesSbox_keyAdd_2_sbox_io_o5), .B(io_key[5]), 
        .Z(output_sbox_2[5]) );
  XOR2_X1 AesSbox_keyAdd_2_U2 ( .A(AesSbox_keyAdd_2_sbox_io_o6), .B(io_key[6]), 
        .Z(output_sbox_2[6]) );
  XOR2_X1 AesSbox_keyAdd_2_U1 ( .A(AesSbox_keyAdd_2_sbox_io_o7), .B(io_key[7]), 
        .Z(output_sbox_2[7]) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U136 ( .A(io_state[0]), .B(io_state[3]), .Z(
        AesSbox_keyAdd_2_sbox_n71) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U135 ( .A(io_state[2]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_2_sbox_n107) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U134 ( .A(AesSbox_keyAdd_2_sbox_n71), .B(
        AesSbox_keyAdd_2_sbox_n107), .Z(AesSbox_keyAdd_2_sbox_n75) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U133 ( .A(io_state[1]), .B(io_state[5]), .Z(
        AesSbox_keyAdd_2_sbox_n126) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U132 ( .A(io_state[6]), .B(io_state[4]), .ZN(
        AesSbox_keyAdd_2_sbox_n125) );
  INV_X1 AesSbox_keyAdd_2_sbox_U131 ( .A(AesSbox_keyAdd_2_sbox_n125), .ZN(
        AesSbox_keyAdd_2_sbox_n108) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U130 ( .A(AesSbox_keyAdd_2_sbox_n108), .B(
        AesSbox_keyAdd_2_sbox_n126), .Z(AesSbox_keyAdd_2_sbox_n74) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U129 ( .A1(AesSbox_keyAdd_2_sbox_n74), .A2(
        AesSbox_keyAdd_2_sbox_n71), .ZN(AesSbox_keyAdd_2_sbox_n117) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U128 ( .A(io_state[3]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_2_sbox_n124) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U127 ( .A(AesSbox_keyAdd_2_sbox_n107), .B(
        AesSbox_keyAdd_2_sbox_n71), .ZN(AesSbox_keyAdd_2_sbox_n128) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U126 ( .A1(AesSbox_keyAdd_2_sbox_n124), .A2(
        AesSbox_keyAdd_2_sbox_n128), .ZN(AesSbox_keyAdd_2_sbox_n127) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U125 ( .A(AesSbox_keyAdd_2_sbox_n117), .B(
        AesSbox_keyAdd_2_sbox_n127), .ZN(AesSbox_keyAdd_2_sbox_n100) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U124 ( .A(AesSbox_keyAdd_2_sbox_n126), .B(
        AesSbox_keyAdd_2_sbox_n100), .ZN(AesSbox_keyAdd_2_sbox_n120) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U123 ( .A(AesSbox_keyAdd_2_sbox_n125), .B(
        AesSbox_keyAdd_2_sbox_n71), .ZN(AesSbox_keyAdd_2_sbox_n61) );
  INV_X1 AesSbox_keyAdd_2_sbox_U122 ( .A(AesSbox_keyAdd_2_sbox_n124), .ZN(
        AesSbox_keyAdd_2_sbox_n73) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U121 ( .A(io_state[0]), .B(io_state[6]), .Z(
        AesSbox_keyAdd_2_sbox_n48) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U120 ( .A(AesSbox_keyAdd_2_sbox_n73), .B(
        AesSbox_keyAdd_2_sbox_n48), .Z(AesSbox_keyAdd_2_sbox_n64) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U119 ( .A1(AesSbox_keyAdd_2_sbox_n64), .A2(
        AesSbox_keyAdd_2_sbox_n61), .ZN(AesSbox_keyAdd_2_sbox_n113) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U118 ( .A(io_state[1]), .B(io_state[2]), .Z(
        AesSbox_keyAdd_2_sbox_n119) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U117 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_2_sbox_n119), .Z(AesSbox_keyAdd_2_sbox_n66) );
  INV_X1 AesSbox_keyAdd_2_sbox_U116 ( .A(AesSbox_keyAdd_2_sbox_n66), .ZN(
        AesSbox_keyAdd_2_sbox_n115) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U115 ( .A(AesSbox_keyAdd_2_sbox_n115), .B(
        io_state[6]), .ZN(AesSbox_keyAdd_2_sbox_n14) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U114 ( .A(io_state[0]), .B(io_state[5]), .ZN(
        AesSbox_keyAdd_2_sbox_n116) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U113 ( .A(AesSbox_keyAdd_2_sbox_n14), .B(
        AesSbox_keyAdd_2_sbox_n116), .Z(AesSbox_keyAdd_2_sbox_n65) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U112 ( .A(io_state[7]), .B(
        AesSbox_keyAdd_2_sbox_n61), .ZN(AesSbox_keyAdd_2_sbox_n58) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U111 ( .A1(AesSbox_keyAdd_2_sbox_n65), .A2(
        AesSbox_keyAdd_2_sbox_n58), .ZN(AesSbox_keyAdd_2_sbox_n123) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U110 ( .A(AesSbox_keyAdd_2_sbox_n113), .B(
        AesSbox_keyAdd_2_sbox_n123), .Z(AesSbox_keyAdd_2_sbox_n122) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U109 ( .A(AesSbox_keyAdd_2_sbox_n61), .B(
        AesSbox_keyAdd_2_sbox_n122), .ZN(AesSbox_keyAdd_2_sbox_n121) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U108 ( .A(AesSbox_keyAdd_2_sbox_n120), .B(
        AesSbox_keyAdd_2_sbox_n121), .Z(AesSbox_keyAdd_2_sbox_n109) );
  INV_X1 AesSbox_keyAdd_2_sbox_U107 ( .A(AesSbox_keyAdd_2_sbox_n109), .ZN(
        AesSbox_keyAdd_2_sbox_n94) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U106 ( .A(AesSbox_keyAdd_2_sbox_n119), .B(
        AesSbox_keyAdd_2_sbox_n61), .ZN(AesSbox_keyAdd_2_sbox_n45) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U105 ( .A1(AesSbox_keyAdd_2_sbox_n45), .A2(
        AesSbox_keyAdd_2_sbox_n116), .ZN(AesSbox_keyAdd_2_sbox_n118) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U104 ( .A(AesSbox_keyAdd_2_sbox_n117), .B(
        AesSbox_keyAdd_2_sbox_n118), .Z(AesSbox_keyAdd_2_sbox_n104) );
  INV_X1 AesSbox_keyAdd_2_sbox_U103 ( .A(AesSbox_keyAdd_2_sbox_n116), .ZN(
        AesSbox_keyAdd_2_sbox_n43) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U102 ( .A(AesSbox_keyAdd_2_sbox_n104), .B(
        AesSbox_keyAdd_2_sbox_n43), .Z(AesSbox_keyAdd_2_sbox_n110) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U101 ( .A(AesSbox_keyAdd_2_sbox_n115), .B(
        io_state[3]), .ZN(AesSbox_keyAdd_2_sbox_n25) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U100 ( .A1(AesSbox_keyAdd_2_sbox_n25), .A2(
        io_state[7]), .ZN(AesSbox_keyAdd_2_sbox_n114) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U99 ( .A(AesSbox_keyAdd_2_sbox_n113), .B(
        AesSbox_keyAdd_2_sbox_n114), .ZN(AesSbox_keyAdd_2_sbox_n112) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U98 ( .A(AesSbox_keyAdd_2_sbox_n45), .B(
        AesSbox_keyAdd_2_sbox_n112), .ZN(AesSbox_keyAdd_2_sbox_n111) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U97 ( .A(AesSbox_keyAdd_2_sbox_n110), .B(
        AesSbox_keyAdd_2_sbox_n111), .Z(AesSbox_keyAdd_2_sbox_n81) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U96 ( .A(AesSbox_keyAdd_2_sbox_n109), .B(
        AesSbox_keyAdd_2_sbox_n81), .Z(AesSbox_keyAdd_2_sbox_n84) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U95 ( .A1(AesSbox_keyAdd_2_sbox_n94), .A2(
        AesSbox_keyAdd_2_sbox_n84), .ZN(AesSbox_keyAdd_2_sbox_n101) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U94 ( .A(AesSbox_keyAdd_2_sbox_n25), .B(
        AesSbox_keyAdd_2_sbox_n71), .ZN(AesSbox_keyAdd_2_sbox_n50) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U93 ( .A(AesSbox_keyAdd_2_sbox_n107), .B(
        AesSbox_keyAdd_2_sbox_n108), .Z(AesSbox_keyAdd_2_sbox_n68) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U92 ( .A1(AesSbox_keyAdd_2_sbox_n68), .A2(
        AesSbox_keyAdd_2_sbox_n48), .ZN(AesSbox_keyAdd_2_sbox_n98) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U91 ( .A(AesSbox_keyAdd_2_sbox_n66), .B(
        AesSbox_keyAdd_2_sbox_n68), .ZN(AesSbox_keyAdd_2_sbox_n33) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U90 ( .A1(AesSbox_keyAdd_2_sbox_n50), .A2(
        AesSbox_keyAdd_2_sbox_n33), .ZN(AesSbox_keyAdd_2_sbox_n106) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U89 ( .A(AesSbox_keyAdd_2_sbox_n98), .B(
        AesSbox_keyAdd_2_sbox_n106), .Z(AesSbox_keyAdd_2_sbox_n105) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U88 ( .A(AesSbox_keyAdd_2_sbox_n50), .B(
        AesSbox_keyAdd_2_sbox_n105), .Z(AesSbox_keyAdd_2_sbox_n102) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U87 ( .A(AesSbox_keyAdd_2_sbox_n33), .B(
        AesSbox_keyAdd_2_sbox_n104), .Z(AesSbox_keyAdd_2_sbox_n103) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U86 ( .A(AesSbox_keyAdd_2_sbox_n102), .B(
        AesSbox_keyAdd_2_sbox_n103), .Z(AesSbox_keyAdd_2_sbox_n85) );
  INV_X1 AesSbox_keyAdd_2_sbox_U85 ( .A(AesSbox_keyAdd_2_sbox_n85), .ZN(
        AesSbox_keyAdd_2_sbox_n77) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U84 ( .A1(AesSbox_keyAdd_2_sbox_n101), .A2(
        AesSbox_keyAdd_2_sbox_n77), .ZN(AesSbox_keyAdd_2_sbox_n93) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U83 ( .A(AesSbox_keyAdd_2_sbox_n48), .B(
        AesSbox_keyAdd_2_sbox_n100), .ZN(AesSbox_keyAdd_2_sbox_n95) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U82 ( .A1(AesSbox_keyAdd_2_sbox_n66), .A2(
        AesSbox_keyAdd_2_sbox_n14), .ZN(AesSbox_keyAdd_2_sbox_n99) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U81 ( .A(AesSbox_keyAdd_2_sbox_n98), .B(
        AesSbox_keyAdd_2_sbox_n99), .Z(AesSbox_keyAdd_2_sbox_n97) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U80 ( .A(AesSbox_keyAdd_2_sbox_n68), .B(
        AesSbox_keyAdd_2_sbox_n97), .Z(AesSbox_keyAdd_2_sbox_n96) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U79 ( .A(AesSbox_keyAdd_2_sbox_n95), .B(
        AesSbox_keyAdd_2_sbox_n96), .Z(AesSbox_keyAdd_2_sbox_n91) );
  INV_X1 AesSbox_keyAdd_2_sbox_U78 ( .A(AesSbox_keyAdd_2_sbox_n91), .ZN(
        AesSbox_keyAdd_2_sbox_n90) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U77 ( .A1(AesSbox_keyAdd_2_sbox_n90), .A2(
        AesSbox_keyAdd_2_sbox_n94), .ZN(AesSbox_keyAdd_2_sbox_n80) );
  INV_X1 AesSbox_keyAdd_2_sbox_U76 ( .A(AesSbox_keyAdd_2_sbox_n80), .ZN(
        AesSbox_keyAdd_2_sbox_n88) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U75 ( .A(AesSbox_keyAdd_2_sbox_n93), .B(
        AesSbox_keyAdd_2_sbox_n88), .Z(AesSbox_keyAdd_2_sbox_n92) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U74 ( .A(AesSbox_keyAdd_2_sbox_n92), .B(
        AesSbox_keyAdd_2_sbox_n84), .ZN(AesSbox_keyAdd_2_sbox_n13) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U73 ( .A1(AesSbox_keyAdd_2_sbox_n81), .A2(
        AesSbox_keyAdd_2_sbox_n91), .ZN(AesSbox_keyAdd_2_sbox_n89) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U72 ( .A(AesSbox_keyAdd_2_sbox_n77), .B(
        AesSbox_keyAdd_2_sbox_n90), .Z(AesSbox_keyAdd_2_sbox_n79) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U71 ( .A1(AesSbox_keyAdd_2_sbox_n89), .A2(
        AesSbox_keyAdd_2_sbox_n79), .ZN(AesSbox_keyAdd_2_sbox_n87) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U70 ( .A(AesSbox_keyAdd_2_sbox_n87), .B(
        AesSbox_keyAdd_2_sbox_n88), .Z(AesSbox_keyAdd_2_sbox_n86) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U69 ( .A(AesSbox_keyAdd_2_sbox_n86), .B(
        AesSbox_keyAdd_2_sbox_n79), .Z(AesSbox_keyAdd_2_sbox_n59) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U68 ( .A(AesSbox_keyAdd_2_sbox_n13), .B(
        AesSbox_keyAdd_2_sbox_n59), .Z(AesSbox_keyAdd_2_sbox_n46) );
  INV_X1 AesSbox_keyAdd_2_sbox_U67 ( .A(AesSbox_keyAdd_2_sbox_n46), .ZN(
        AesSbox_keyAdd_2_sbox_n42) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U66 ( .A(AesSbox_keyAdd_2_sbox_n80), .B(
        AesSbox_keyAdd_2_sbox_n85), .Z(AesSbox_keyAdd_2_sbox_n83) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U65 ( .A1(AesSbox_keyAdd_2_sbox_n83), .A2(
        AesSbox_keyAdd_2_sbox_n84), .ZN(AesSbox_keyAdd_2_sbox_n82) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U64 ( .A(AesSbox_keyAdd_2_sbox_n82), .B(
        AesSbox_keyAdd_2_sbox_n81), .ZN(AesSbox_keyAdd_2_sbox_n32) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U63 ( .A(AesSbox_keyAdd_2_sbox_n80), .B(
        AesSbox_keyAdd_2_sbox_n81), .Z(AesSbox_keyAdd_2_sbox_n78) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U62 ( .A1(AesSbox_keyAdd_2_sbox_n78), .A2(
        AesSbox_keyAdd_2_sbox_n79), .ZN(AesSbox_keyAdd_2_sbox_n76) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U61 ( .A(AesSbox_keyAdd_2_sbox_n76), .B(
        AesSbox_keyAdd_2_sbox_n77), .ZN(AesSbox_keyAdd_2_sbox_n24) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U60 ( .A(AesSbox_keyAdd_2_sbox_n32), .B(
        AesSbox_keyAdd_2_sbox_n24), .ZN(AesSbox_keyAdd_2_sbox_n70) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U59 ( .A(AesSbox_keyAdd_2_sbox_n42), .B(
        AesSbox_keyAdd_2_sbox_n70), .Z(AesSbox_keyAdd_2_sbox_n72) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U58 ( .A1(AesSbox_keyAdd_2_sbox_n75), .A2(
        AesSbox_keyAdd_2_sbox_n72), .ZN(AesSbox_keyAdd_2_sbox_n22) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U57 ( .A1(AesSbox_keyAdd_2_sbox_n74), .A2(
        AesSbox_keyAdd_2_sbox_n70), .ZN(AesSbox_keyAdd_2_sbox_n40) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U56 ( .A(AesSbox_keyAdd_2_sbox_n22), .B(
        AesSbox_keyAdd_2_sbox_n40), .ZN(AesSbox_keyAdd_2_sbox_n55) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U55 ( .A1(AesSbox_keyAdd_2_sbox_n72), .A2(
        AesSbox_keyAdd_2_sbox_n73), .ZN(AesSbox_keyAdd_2_sbox_n69) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U54 ( .A1(AesSbox_keyAdd_2_sbox_n70), .A2(
        AesSbox_keyAdd_2_sbox_n71), .ZN(AesSbox_keyAdd_2_sbox_n41) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U53 ( .A(AesSbox_keyAdd_2_sbox_n69), .B(
        AesSbox_keyAdd_2_sbox_n41), .Z(AesSbox_keyAdd_2_sbox_n15) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U52 ( .A(AesSbox_keyAdd_2_sbox_n13), .B(
        AesSbox_keyAdd_2_sbox_n32), .ZN(AesSbox_keyAdd_2_sbox_n47) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U51 ( .A1(AesSbox_keyAdd_2_sbox_n68), .A2(
        AesSbox_keyAdd_2_sbox_n47), .ZN(AesSbox_keyAdd_2_sbox_n67) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U50 ( .A(AesSbox_keyAdd_2_sbox_n15), .B(
        AesSbox_keyAdd_2_sbox_n67), .Z(AesSbox_keyAdd_2_sbox_n4) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U49 ( .A1(AesSbox_keyAdd_2_sbox_n13), .A2(
        AesSbox_keyAdd_2_sbox_n66), .ZN(AesSbox_keyAdd_2_sbox_n16) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U48 ( .A1(AesSbox_keyAdd_2_sbox_n59), .A2(
        AesSbox_keyAdd_2_sbox_n65), .ZN(AesSbox_keyAdd_2_sbox_n62) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U47 ( .A(AesSbox_keyAdd_2_sbox_n16), .B(
        AesSbox_keyAdd_2_sbox_n62), .Z(AesSbox_keyAdd_2_sbox_n28) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U46 ( .A(AesSbox_keyAdd_2_sbox_n4), .B(
        AesSbox_keyAdd_2_sbox_n28), .ZN(AesSbox_keyAdd_2_sbox_n35) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U45 ( .A(AesSbox_keyAdd_2_sbox_n24), .B(
        AesSbox_keyAdd_2_sbox_n59), .ZN(AesSbox_keyAdd_2_sbox_n60) );
  AND2_X1 AesSbox_keyAdd_2_sbox_U44 ( .A1(AesSbox_keyAdd_2_sbox_n60), .A2(
        AesSbox_keyAdd_2_sbox_n64), .ZN(AesSbox_keyAdd_2_sbox_n56) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U43 ( .A(AesSbox_keyAdd_2_sbox_n35), .B(
        AesSbox_keyAdd_2_sbox_n56), .Z(AesSbox_keyAdd_2_sbox_n63) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U42 ( .A(AesSbox_keyAdd_2_sbox_n55), .B(
        AesSbox_keyAdd_2_sbox_n63), .Z(AesSbox_keyAdd_2_sbox_io_o0) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U41 ( .A(AesSbox_keyAdd_2_sbox_n15), .B(
        AesSbox_keyAdd_2_sbox_n62), .Z(AesSbox_keyAdd_2_sbox_n52) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U40 ( .A1(AesSbox_keyAdd_2_sbox_n60), .A2(
        AesSbox_keyAdd_2_sbox_n61), .ZN(AesSbox_keyAdd_2_sbox_n51) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U39 ( .A1(AesSbox_keyAdd_2_sbox_n58), .A2(
        AesSbox_keyAdd_2_sbox_n59), .ZN(AesSbox_keyAdd_2_sbox_n57) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U38 ( .A(AesSbox_keyAdd_2_sbox_n56), .B(
        AesSbox_keyAdd_2_sbox_n57), .Z(AesSbox_keyAdd_2_sbox_n29) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U37 ( .A(AesSbox_keyAdd_2_sbox_n51), .B(
        AesSbox_keyAdd_2_sbox_n29), .ZN(AesSbox_keyAdd_2_sbox_n34) );
  INV_X1 AesSbox_keyAdd_2_sbox_U36 ( .A(AesSbox_keyAdd_2_sbox_n55), .ZN(
        AesSbox_keyAdd_2_sbox_n54) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U35 ( .A(AesSbox_keyAdd_2_sbox_n34), .B(
        AesSbox_keyAdd_2_sbox_n54), .Z(AesSbox_keyAdd_2_sbox_n53) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U34 ( .A(AesSbox_keyAdd_2_sbox_n52), .B(
        AesSbox_keyAdd_2_sbox_n53), .Z(AesSbox_keyAdd_2_sbox_io_o1) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U33 ( .A1(io_state[7]), .A2(
        AesSbox_keyAdd_2_sbox_n24), .ZN(AesSbox_keyAdd_2_sbox_n31) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U32 ( .A(AesSbox_keyAdd_2_sbox_n51), .B(
        AesSbox_keyAdd_2_sbox_n31), .ZN(AesSbox_keyAdd_2_sbox_n5) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U31 ( .A1(AesSbox_keyAdd_2_sbox_n50), .A2(
        AesSbox_keyAdd_2_sbox_n32), .ZN(AesSbox_keyAdd_2_sbox_n49) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U30 ( .A(AesSbox_keyAdd_2_sbox_n5), .B(
        AesSbox_keyAdd_2_sbox_n49), .ZN(AesSbox_keyAdd_2_sbox_n20) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U29 ( .A1(AesSbox_keyAdd_2_sbox_n47), .A2(
        AesSbox_keyAdd_2_sbox_n48), .ZN(AesSbox_keyAdd_2_sbox_n3) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U28 ( .A1(AesSbox_keyAdd_2_sbox_n45), .A2(
        AesSbox_keyAdd_2_sbox_n46), .ZN(AesSbox_keyAdd_2_sbox_n44) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U27 ( .A(AesSbox_keyAdd_2_sbox_n3), .B(
        AesSbox_keyAdd_2_sbox_n44), .ZN(AesSbox_keyAdd_2_sbox_n23) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U26 ( .A(AesSbox_keyAdd_2_sbox_n20), .B(
        AesSbox_keyAdd_2_sbox_n23), .ZN(AesSbox_keyAdd_2_sbox_n36) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U25 ( .A1(AesSbox_keyAdd_2_sbox_n42), .A2(
        AesSbox_keyAdd_2_sbox_n43), .ZN(AesSbox_keyAdd_2_sbox_n38) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U24 ( .A(AesSbox_keyAdd_2_sbox_n40), .B(
        AesSbox_keyAdd_2_sbox_n41), .Z(AesSbox_keyAdd_2_sbox_n39) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U23 ( .A(AesSbox_keyAdd_2_sbox_n38), .B(
        AesSbox_keyAdd_2_sbox_n39), .Z(AesSbox_keyAdd_2_sbox_n37) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U22 ( .A(AesSbox_keyAdd_2_sbox_n36), .B(
        AesSbox_keyAdd_2_sbox_n37), .Z(AesSbox_keyAdd_2_sbox_io_o2) );
  INV_X1 AesSbox_keyAdd_2_sbox_U21 ( .A(AesSbox_keyAdd_2_sbox_n35), .ZN(
        AesSbox_keyAdd_2_sbox_n19) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U20 ( .A(AesSbox_keyAdd_2_sbox_n19), .B(
        AesSbox_keyAdd_2_sbox_n34), .Z(AesSbox_keyAdd_2_sbox_io_o3) );
  NOR2_X1 AesSbox_keyAdd_2_sbox_U19 ( .A1(AesSbox_keyAdd_2_sbox_n32), .A2(
        AesSbox_keyAdd_2_sbox_n33), .ZN(AesSbox_keyAdd_2_sbox_n12) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U18 ( .A(AesSbox_keyAdd_2_sbox_n31), .B(
        AesSbox_keyAdd_2_sbox_n12), .Z(AesSbox_keyAdd_2_sbox_n30) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U17 ( .A(AesSbox_keyAdd_2_sbox_n15), .B(
        AesSbox_keyAdd_2_sbox_n30), .Z(AesSbox_keyAdd_2_sbox_n26) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U16 ( .A(AesSbox_keyAdd_2_sbox_n28), .B(
        AesSbox_keyAdd_2_sbox_n29), .ZN(AesSbox_keyAdd_2_sbox_n27) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U15 ( .A(AesSbox_keyAdd_2_sbox_n26), .B(
        AesSbox_keyAdd_2_sbox_n27), .Z(AesSbox_keyAdd_2_sbox_io_o4) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U14 ( .A1(AesSbox_keyAdd_2_sbox_n24), .A2(
        AesSbox_keyAdd_2_sbox_n25), .ZN(AesSbox_keyAdd_2_sbox_n21) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U13 ( .A(AesSbox_keyAdd_2_sbox_n22), .B(
        AesSbox_keyAdd_2_sbox_n23), .Z(AesSbox_keyAdd_2_sbox_n10) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U12 ( .A(AesSbox_keyAdd_2_sbox_n21), .B(
        AesSbox_keyAdd_2_sbox_n10), .Z(AesSbox_keyAdd_2_sbox_n17) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U11 ( .A(AesSbox_keyAdd_2_sbox_n19), .B(
        AesSbox_keyAdd_2_sbox_n20), .Z(AesSbox_keyAdd_2_sbox_n18) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U10 ( .A(AesSbox_keyAdd_2_sbox_n17), .B(
        AesSbox_keyAdd_2_sbox_n18), .Z(AesSbox_keyAdd_2_sbox_io_o5) );
  XNOR2_X1 AesSbox_keyAdd_2_sbox_U9 ( .A(AesSbox_keyAdd_2_sbox_n15), .B(
        AesSbox_keyAdd_2_sbox_n16), .ZN(AesSbox_keyAdd_2_sbox_n8) );
  NAND2_X1 AesSbox_keyAdd_2_sbox_U8 ( .A1(AesSbox_keyAdd_2_sbox_n13), .A2(
        AesSbox_keyAdd_2_sbox_n14), .ZN(AesSbox_keyAdd_2_sbox_n11) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U7 ( .A(AesSbox_keyAdd_2_sbox_n11), .B(
        AesSbox_keyAdd_2_sbox_n12), .Z(AesSbox_keyAdd_2_sbox_n7) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U6 ( .A(AesSbox_keyAdd_2_sbox_n7), .B(
        AesSbox_keyAdd_2_sbox_n10), .Z(AesSbox_keyAdd_2_sbox_n9) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U5 ( .A(AesSbox_keyAdd_2_sbox_n8), .B(
        AesSbox_keyAdd_2_sbox_n9), .Z(AesSbox_keyAdd_2_sbox_io_o6) );
  INV_X1 AesSbox_keyAdd_2_sbox_U4 ( .A(AesSbox_keyAdd_2_sbox_n7), .ZN(
        AesSbox_keyAdd_2_sbox_n6) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U3 ( .A(AesSbox_keyAdd_2_sbox_n5), .B(
        AesSbox_keyAdd_2_sbox_n6), .Z(AesSbox_keyAdd_2_sbox_n1) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U2 ( .A(AesSbox_keyAdd_2_sbox_n3), .B(
        AesSbox_keyAdd_2_sbox_n4), .Z(AesSbox_keyAdd_2_sbox_n2) );
  XOR2_X1 AesSbox_keyAdd_2_sbox_U1 ( .A(AesSbox_keyAdd_2_sbox_n1), .B(
        AesSbox_keyAdd_2_sbox_n2), .Z(AesSbox_keyAdd_2_sbox_io_o7) );
endmodule

